

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
g7azmhtm6FcP7uNFjuXJjN8Z6yccOPk3SSjzvKB27peFKmnPmQmov5+YTGwYqqN9LpdyiUExk8K6
vPnJqontvQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MFrqn2K0Cr7TmQ5al162oDGiY83d+AkTWOgFyXPYrTNznygR/tx44RAp24ytphNK9p6shs2EFMg/
Qqz0l8DCWiVEoJ/T8vMpnAn7Y+poGVGS1qAR3qE2njrl81VcGBZJeFaWIudhfr/DLTuuf2T/dWDU
YpelM3KbfYNPPiPy8PU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FZca5XZouG+/BYoQ8qrJTmnJanku4IprIWRkO6VciHehE5WehR0wsZJhfKlqLEeY1oTPA4bXaxmY
NjYkrop4EOwW8t47/hj2kFLI1OKUAE/TAhCGg/aNSOViUbB3dUomG/y+TBuDt9L6g0Arj1vb/5Pt
IChc5ZdEfRr1lJMTpFfP+5qmEH6lePPdzgPZATPB4Zrj0P6EyiEsU1FKBuAKd9iYNGiLCxVomaz0
3/RwK2Nl+/l4mc7PJt5Hso+4s1qHb4s2wD+OgbIwdH26ZkEnKVFpaLiuWQKu9uhDLGnsBMPf7XDE
p29f+mrvP9Zi/3nonA2aBKrTwR7XuH+ZYoakxA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jP68OjlYJglq3zpmKrXOhq7Sex8XNW8fQKp4hUNmuw06OOoKhQASNTnjtyVjAIk/VXb64ViBu1ds
cNMJybDSWBhnChfJq4h9PNybShGJXxSm3NDOo5wUHKf10Eti3fSotB9rVks+tNdTEZo4O97kgfdD
G1FNOqlsYcQiShEGLLiEQ2yYtgJBxJ+jc8mFjIEfPhAYy1ElrvtFEpnhkNS2LfE7xdWOQdO/XoKK
ibeY08pgncTI3pvO6TMbXushf0AX2S7hgfk8ysZrT+0gktqFrJnyR6oljS6VVPLtRNW2vo/cC8XQ
Bzvwwt4cpSo5KLS4XxB6qClZipItck2AUEdIbQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o7jAZIoXlFbFtDYmtXhfRBlb07dhBb6Wp03mlT4T0FXtvccSHWhWZgc+VUNwt6TohLihOwvSipPP
XVXpGL4pUVYNdQBCVpFzhMkt6jhyUgsF5t10yI5Of6YEfQrDHigceoBukM3+/zJHPprrPQE6FUvC
wXSGhBCXnHJs1R+n4l0714w8/WftPQhlD9QGQp1qT2VARQXUKBRxcRjxe9TcLfs0P4xnN7uHu0R6
JTmV+MHmhGpetSZGx+B2Wa1MQofUPURqwE70IwBoUhdXH8+39DT5I6x2+wMY6RcVATnhNd2BCgPd
RzAhwfrcqRiU9aB+eNNdFR8ve9M2nGMmV2JxZg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Cl1Dz+fZIDYEIQuUd0pSg+5jknmtX/JERd+yOZ2SRaVra/4pU/eCTjEXMzhz4VFGYB6dgUxMsGBk
nL2WNdn/uaSPpi6mNF0UHQvZik4pUkYPrnRbFveVqW8i1t95SG0RW96uD19206lWrp5U1lqc4fH7
sfKHi8ZpU3MAg0DOO0E=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Qqp76m2aV9ue8Qai7QUavb+lhRYdu/txrnwYLzwTe0vS0S2OD1vxr8VeIT3bF/ZuXlTGm4S/UCSF
bgOPp7VqEOeGNfsSPK+VpQ+foQMENCQYccwKquBDSg/sLjpPK9uuoGLBLxjw2OwsRzplVFXiPcRN
LYK1/FmCP7RJBNgmhh/ti99a+WSl6i2YIIRGocNplQlG8FXq8ZTTHd/x2Gtdf/zGvJOy/fNsos6S
Oq9yJ0rMmbGeWbri5c04gZM08pUmXBsivgOHm2IVEZZFM4SBqrsi0xa52hs2kelc3iKJcWiTvU3X
0fJP9qNFuIjXBPPZvEYwhVtIh6DwiIC2viSscQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967856)
`protect data_block
g4MXYLIO/zzgxWsnFKxy8mK347xma9qlqEn58IDvZo8KzaB5A5YTYVOXKirHzL9/Ky8N75dUpQ7I
kd9Z5ZgaiL/uD7N/v5HKrcB6V4HL2CsoDl8DZV079T53KtQtnsPxSJRfb8aUkPRI9kk+8hip7vwm
q1VcbmmZMqutItV6W1BYIet9wjWtzz/EY/FQLI0Rthw8f1ab9UpQ6frLP2zsYSRthwPwHEj674ko
pY7NdUZ+079cZp1OSzu/78bA8SOzdZrNRK3EtBYQfyXfqyOoK2+j6RXu35QcQBztWT3ZpIs7czU7
iQhyjX3hQgourtaZeWTSmoQgf3MJ6NasjBnrAmZwUYfWxII67fQXJYacrx4W7Atdrz4DT2Fih9wu
Ybd6EAKUdp+LZUipkj7xvF9+9GGexFSkafWP5ueWkaAvqEYlhFQSWlnwpWos/4FBrTf5XBm21jTQ
OynUejSOTk/xunkhAPrFm0przdg082Usy3RTy7HsRSDanpn8OZIyT5ptIIeOnr99CNAr8aiO68Ad
IEkdW6ITZB69gWFa9hDdOQpKFW2I8VtM+qJaufZ4L1HJZnhDcCkZyT3wDq9ezwMTk3UBbHsyRZnk
QDTcolZmQ0AjtBKohPWDl6WR2hSRgfDZzvlCXPRgUIqP5M2W0hIs0zL4K7WJ5kQIrUgwMfvWyIO0
WL5s8bN4hlBGKor2VCzVqJm8yNZkKRJSAqQTfE8MpLUjuH+VnDbeWGI/Fssl1jwraCyflpiXs2OI
WJnIHy1Jma/HSw/QB9tGYBW7Ul5Q9nD0NPqBggYFFGNQ+WKxzPVEGRtEDFr82TQdRnSLfgm8T0D3
0PH0SnnEj10zGgL0EmO9S6X2izeVGH4uBKhWHvi7e3gTBh+BUhlkwKWolYkkhb7CemeA/PIq5uKA
t7hD3nEGFLozON5f7/4O5AybLmjhwXTO29l015kJO5DFCMLjIdv9Av6KgomAIxEHcYXwMkiF9903
YjJ71qE6coMJb4RM3dqqdQoPve4U140xZLpSBCHzY6Bwp8HhpxdzYOrdvP8sSYCV6A+y/LENpZpJ
nAwM9LuqKYchYOhI8U4LVJrPguRXN1F0ti8lrW72IO0NsuyywSNlyrPbGpoHXAgVGMZUQVqQCPVF
hiA2Mmhh5MYdHJQO5W6UlcKB8DIie728Jx9X4sYHxDjiZhzVPp1LOdFzEvT4RakMSQYOQwV5kcV9
094XUBy3QolzOQQCO0W/xt5AcoHN/plWnA+lq0y7Ws09gNl9dZRNSI3A7ryqf6vLvtxV85H+/pwT
/tkU5iiHzUUy/rD9Vdb7WT1VO+uQ4bEJZV0BrBXwdsL9ZFVhL28kBIgL50B9au6uElxksem8FAAA
qB49Gid3XpSEHOwEYEmq5E5vqFFEczLQGeqygxvRJSwb4/nkfro3CZ9GfP+lOc5HxOwt0OvK8lCm
JdiHMA5evdggYvWy1GyEyhe9u1iURjDDKa9coZVf8AFE4QSuriECQZzGmadQy+XyX46aUVuqfkoZ
BdBQaPvnncJsO6Ml5r/Pz8X8XZRpxBDIFfyLiCPurcd9Ft7A9YQT56q3YdkqXypJaWB3ID8Tne72
sEIqGoyeXUxMNVD/QKdnGSG00PJhQJKpbn6mxllN80CPdZhx5smSrbiqUOwQnWgY4oC1NepPmhjS
MKO2QFqHjECSBICtNFPLdkuGvUVcW34SFvyO6RG3eRllZsOfk55SX2p+XHw7UTc/NrdE/0ZEQi99
bqMbeMiMwqUkmdS6Kvdh34sxUApHNGQFhvEKLXI+UbCYkoOzzxwp/xHMYf42Evi+Vso+loqLEQPi
ntcKc4hlphk9h9Vd8zwuzoWza9w6nUj8PE6H+PqO1M0H/UAHW0CV6Njgzy3TnACf+50/pg+F6GLp
aNQW9JH1eSyjHmAIP7bRbSjev6NC0ioKcc3wTXWGEFLqFXsQJs4gUE+SDVfcMuih2Z6O5S7C8wLT
YgeTp+qigXIZUfKooWdyWMLzzGm5Qszm32m9NO6FK4zHKM3s7AR/ubvv0rxGGuPusoeTdtCRyTwx
9LDyLgYYmRW7aaSzCzkUeZodS2FkKStBtiaKxfvbaiB3pNb3SKewvByASUSigeGrLVPNkjA5H8AT
etapZ1cDAhk3T3eusACqhjODiAhFqzMavB9s6HOwQ73i1reDfpbI4FqUxSQ/mS15BDcypELvDxVp
c0ifpN0nbYUaCMGHHAZ9ojaWUjoW4H8lo1WYOwpeKsardCjHJGlu81EviE0leFZKfX2fIQFEfyXS
mL5qPZxBsECzwkiCrlFggBlfueyQqnwGIoE8JqUSlA7Kk0TJhx2tfN9TPUNJ1U2RVLJqgnbK5s21
Nw4puJ8Gvl/z6fG2lljOmeOoA/upxwNqsaZuYRxeTkrJfCbEyfOnN4jdROdoHdPrfjG6C5N8Z3De
y0wVskyDNWbJ5N0xqyM0+m+OppPLOiMq5YIy5XO8AXfYaMtgJ1Y5VO+NU5/9Ko3TF2PPs99LZ8yZ
aH0ILjic9J/Retdhp+qiCLQw5+PnX9Lv7OMV+DPdQPGxzTnjxiKxRJ4fqx0Z84oUv10ttI6TurPP
x//1X/5vmc6xx/IMB2iA4ytuZiM8tVqd+6bSId+MRhj/JjiCVdK4K5p6PEiAkxH+kqzhmdpowruW
MRn0R1LYHB8pnw/odOTsycXBzc+EibXxjdsAe2OGNDLNUMdlJgKSdUTAqUuvLOHvOaxsCrUdCDYT
WizvTJGBCxf76Eh07y068SKGpCOHjsLtDG0xlyZRa1RHhM4fimy32Ftal2vAq1KKmRAhTFaoo7WD
Fm+S7UZKbQWk0Lq5DK5pLFbb0qyJV+ghRDsKLSbBIjWA0Y8XNZLkB2F/c23JMb1D0jed6K6Zj3Eq
etMPrMMyVtScT2L0M+VEHL42OIrJBZ4W3EExQyb/9YJgGwxacwDOdJ/5t4u/sjlJRvnQDkwVYSPZ
F4HM8gABI9n4ii0WlmsEP6qNIWbv9PV8sshl4Kkbrd0VrhXh5nTEzktM4J7Wgbqpi1IHTm2lKid8
WsnjEgiHT0aNzgcIvMPoZw2a4Ts/XBJDeCzxuFjADe1bJNY6fbebu/011fsitUv8YVAnusR47BM1
a5RMA762CFqtzPpa0VE6E5DTevwNPY1U1JVwhbP1IGXE7Ub/e2ROCq4alHnYQZxabVrR6bdO9cW5
hgiREwSe0/IQ61t3nh017QZ9HhbXf9pXUD2T66/fyYujiyafM4g3OALjywPyRpBmOGt+A0ZCo6aT
c62oWZLoiKu5d9YJDMI5MFnSegDGO0IxPdOxc4bA4gSGDdSSvksWfyGhWM1Rb7DlwSJ4cZWExPAb
YUjOxeAwRAuQLBzzaOh12xBdvtEnT+W9TUIqluDbidZ4W3W3JjfLp9rwuS5zm2KJwJZyQwSHcH00
JteQ6bcRGqt5nLD5vwpn7S+kAlEPNyI/c+i0RRb3h7Iqcr2NSOVIPQj5TpAGsf8G/3O+Y5KPi9iC
HGW6UvxJ3ZTJUOWVlw59oXI4fMqHHW6ABwKmFO+Wa7FaNaAnyeRk0sIypwKjV94SFdrpAmfx9Pmm
phEg2DlGsjFQ9MpZn2yjM8M7XMOS/yIQIlZqwtGxhCMHS/ERVyVM+ztxsL3bKbgx7UaOuDzjgHnc
R65vXRSe+UevSCnPwzGRoqAEHegnojfd9bDiaKPQjszTjlVCTNTGMKQutCCHKgo/nJ3+Q+rv/c8S
OmSwEU8oj06ukT65uczI9/PnMByCGCiFCgHB9v7JagnCBqOJx3ThCWLKP6kfdaSKE+bHoAa/DAz4
AGNnBTIESV+EkKsAlPwRTA1PIzXMUJ9vPfrWw4g1lndzhKbwt4doIlXEXH99YmxQvQVr7EGWGLKh
ddKuo4ktpK9KFy5JcRHrc0ShPBg0ZSF7C8NbV/IwuHK5JbJrYIBUkOvW0uJjKOLVMU6uC7aO3L7f
4YrYGNk6DGL5ecgodSSVjkjWtzZ/RQhpENnNagErKu8nl0RazejP2i4PnQKnu8yXg6fO2bqieRUm
rKYJR9/e00mFU2wnbSG4uJCo6ftx8Na3epL32gJWa072cK1jgRfQq5C46gwxkFed2mXxhg5QazN5
yx5zd2ABzPTBoooVWeqsiIEuSW/tQpNoEE6fZ93n9fr2rbwRgYutlS9m3GlML5HezolztTx1pUQl
aYBgocUhcgBTxwfqvl9dVaCXP+yM991BFTPpccVTtT/axZ+by/PAuhY3D1uVQs1L7K2AVDUb7t3p
niYOKbbZAenY6IxKgXrxealsM/VRRLVMwRpmX+4QJ4wI51EPLBVg81FoLwpbp6yQ05OSwWJQFY8V
tpJR5uvQ4+Ejv4gdpFhmKL2XLDBGOi/ZpIxblVMURBggsX2Z2iIxtv3QXxNUiop0Ih6en12TD+YY
ytVAa0bgPGB+lVxOTAResdRhonU/8hu1qW18PO7FdG0KdSrLS36PVqWUq+TAfv3JJgerY2zCjGfs
2jd7L/OQB13zUTDK8+wEbTXqLpP7853TnWIO3x+i5pym0IYCpxjRyC7bvmbdHJLHirdlpxSg6wAS
VrI18iJGS5hXPX8Jk3L0hIoDz9v1fPkkymK1r/qlDTF6naB19Uz2QmL2/NpQn2wT+PlCOOZPldXe
1OnL5/Q3oQyGKF6WExzLp8Pfe9WHph1xulw1lo5FRIegKEuQ2QDUWGQo5DEtnVCiq83AoFU1ezXn
ZDiOTQfv4yyg5g/tgSWB5Grrln519ZvUXVx6ub0OY7BPLW1Eex1IapLT+g1tgxQL2Lw/EchkxeRP
nxbzJOiyZHhCdWbE60QQN/fvqUFGo5xjFSZ9VtxwVJVBKvbX+M3b1TO162EgiMDlkJj2le89x+/+
ltnGS+BHqn5d2w6BIkO85cxPHw7d2WI3s+fI948lpmc+516l32lWgsjCW2SXHJPf99zYulynOxSl
HneKn5XCflt/m9Q/a5oz00EuHMVWh+dMmAsUNs34z7Uj8zTVZRz/BBiOaX7x8AbKRBHJK73nFKLl
otunBN5Ibm81EozA85R2Dt1rAzPjlJw/9xiqsVzQZ4gElSNMyBXtMwCkVF6z4xbRpwCObiZL+p8Z
c3A/4WHHVwzHjXG0G8kq/ejiVcWYq/QplZkt+hFkfG/3EdYiVPrVqREYGHk5+YitsoKBhOu5D/sl
6UqrDrhqAqp0f/q1Dlhg4GH1QEOobUc1xt4+Qu9g2j2uHa4nx9OkmfAyBh9n0VBhNQ+2k4X/eogO
Y5Obfe6OlzHBy0l2UVYviVNc3PLyQXEvGftc4eNYntrKMVtnRbF2G6hcGU65v9J/wLLnUVyaYPpv
eHZEmmjjMlYOD834+E8+cM6tCNgDIbSXO8g0CjvlT/0xhOUKGXQp52vJYCRAUh3qcDSZt2dbxOJ4
M5gcLW9IZxwZAyJEWU5Tj/kXQq6FDT5zJZxyL4Uiyp1iZtrWt8cAeO5YaXIWgd0ifYaeO/9Utw31
KJE0Ddd05+cRU4+FuTkiOROIfn9ZhPFods2JzC6kkiE61nSuX5Z1wEI1S4GrrEDQQJjoqr/Y2qsf
9EZFUNG5ZwWRU6n1cwutLpe2Rpma9owFiswjLBizbl/kLn+ZqqK4X8nV4bHNw3oYiv/LnSq8I/cF
XzP1tZUeP8/9fvIL1PQZ1fceRqne0vC6cWxpEJCOk+aCL/QBbA9iIGhmcPew8xbKgS++U9UUaBI6
C1C3yKT472SDjKZh5GWyokrkoYhyFN1WB/npLusV+wEF/ZPngbATZDaOb5q8dWOhkmhy8xRo6qE6
rGHVXiRwn3zWLdygXe/PqhuEjgxQmP6oaocDqtNC4CIhhJFofxXdWXMIUOz0lhUfLVa+7xhKSuza
5+0wF8hhTmmJP67oUW+tDKJCWE0a87ogjtqkiw0JQYMVcR8ATD7apl6RupscUz8xDfkwFVfH47OF
U1hM3HHP+dLl2rQReEATHgvtxp2ZGFg+YhHorh73l0sOgiHWbMYEzoq4jw07AJEpEnISh50rqc5D
H6iPvPC/eSOzc8xt/jTT0OS4sjX4j2BHVhVuO2ZL0/5IprKc02d3CbemEbnj9a+I0JFh59J6CIAB
cXK3F1I0bfM4fv/Qe7JaXURGArDXeiO/R/C8GON6aPgGCiQ6hN12D3Fzn2NQA73TkyNHIInqBJ6B
RFUdiZSa8aGntVD3Lwy5DVNi0oC7EewbGlkbOkm7gLscdZLH7Z1fvnujDqnBxRQF7xN4e3wexgAg
vV5gf/jnM3SBUaDdelHtmArgg879ecaOpDWhKd6Om+h3fg8+3YPcpsK+uA1R0Mnb0+eomX3B/jyi
1LWqSMklXLgA1iXLQFg9SUcbSkcGj3EyA+Wu5K86C2jYi4xb5as7aSClGdRnd1akimiCw1gCFGDD
ywAF/1ckQxFbEWaLrwO3XmqBh81HPxF7IpE09pP2KPmpjBepOQu1YYfe9kteUTjTRkuoloFJwxcW
A1wjZiBovnfbr+DaSuijebuNOuoa6s1CFH+ZwADjBnoA+KrYR5JrmxMt4hFl7dCswKyKELdZtZp7
VdB4jpSPITctpxysgvepvGxI5qXv4V0k2NxUItHR+qa7XBeuCZhOpCEdRIeDoK83+mhv1SW9uQkR
rT4kVi5IpPndFc+X7gYv4tEq5OWqpjtBlSE/10CtQvF9aUTKZ+eMmin+CnzYI1+4AJ2OR6aHJr+H
4cqOySLRB+QwcnM+jftMi5BYbY5SvLwIx+n44vl+dDtDNn5x/VWE4ixX4tkNWxC6hVOvp66xgAJP
GCCe1oANl4wcIzlj8ume77BhD15BDGxz9xbEKeZxAInWkezafoy4jy5Y+PoIKmHJUZYzxNWhMDDb
rF/gbs0n6moyZRkW2sGfTE+ob2C5UFwriq6I1h17wZpOjervM+Tx949cH5A7rw/MOyTC/6OML25H
GuUt7UjkYlCqMkxXTUQEXJhgXWpk6OumOvm1nADLe0rehpa1Lk7Z6QWilZ/XPgStr0N6GIB1KsB3
SFNnf8FXS7Rs0SefG7tUti5IFlQFYGHLnvF6ftvtaHFOgOmydoe1SS3ZxxZ3moNyYINOBdUXUoKg
1SEhAMdauvf/4Lhq1Rwhq2sck8mfZGGtRoqFVDDo67kEbFAE5gBqtkz74cqCueyWSwKjLjoM03XM
e9GrMh4Yx0EU8MsaUc6qTeH0oywEbke7Wc+h4e+Knkybuh7NP5fkDQHwRUADu8s2E2TJtWbh/Zsc
pZVoO7D3h8ZHJD4hcN5apNgQ1umeb9kmDPahHXt/n7d8XnmDr5npYKVd3FKOUC6dMDuIe7VKWzPA
9SiVUsA/AZCL8q6LXVXpPyB6lMNeR3IhdTxeYKANi8jgpJupM7Fz/mfo2PBYhPX4yqJ1ZStgeUb4
ayReNQl11eqZSoi9t/MA549SdTDkJ+xMHtFaqeQHTt5aD5eQdkc8YMVwfeLOFHyYu7Y5GUY8jxmi
m1V0b2R/rzTlEFfLTeAUZ3Iq8vXPRb/E4FaUtsQlnss0fFZhKD3wUmERYxUfV8y+OEwIKWijTUvp
6X25pkJS+jSozxjOmcZcz8PLnA1q2K/XCxxJZrtwDxA50XsNZaD7EaS+VE/AUYQ2uGfDkOMfNAVi
AFmBkjTaOWi4zRNKfXabMGBzpJiTKsXQ5pxiobkh2tM22IEC+xQOi4uWiwMdAC7MXXdjOyjmSZus
+YzyesSGtJppc6Nx8HCpc984hJgUq9lLwvFC+OmBHOCjWVGMiJYx1D91rKZRp8Dooax6Cdy57+9i
b6DxCV4EqGcyVHXkrMcB4Um67oRuZ4CI5BekxtjcmIb7r62o1AGBYLOWfNKhoI9iKQnjEwKrI17t
TlJ+nVa4fxM22Dr9/Zyulbaot44LIpyR/NKJbGvSJWAsh8EUvAwOJUGTBAVJTOBQm4rxtJBtE0hJ
w4QI6zfYoATFVgzYzg+7mMYWGcdewJtbggiduLheQax0dwFd7TpAon9kZrQBA27fILyRlVcNIjsh
rzKPsAMXcipSJCaK3AzDRRsFqfwNBfdFXr58D4JMdoyoitpMn5osOCETXG8hCK501Yk3fks8jrlL
/KPjCABJNnt4x/G0htEsMeNsqvDMUaHAj9mrnEtFQ0XTCbIDI/7hd4AA9y/zJFFJKL2aaqcsWL+T
Sx1B7o/gbIuKSUiUmDAI3J78LnRXcYgoD7un9iz3J0ZdEPEEAKyMLpfdf2RahMx092ulZg/X4NKk
hlWZ0RSUJbBMDek/oZ0n19A693u06L08ZFvYgqDrhlkeenCrwCTRKXEm8wGNXFyhu8UWVwuqtfMU
JBPfOAVsj4gB8ualb41LR192rdJrd5e0uJPlAXuJlGRqrdW+X5rRcfSs/McjslwBqrWIl6WZtT9p
gKnXSGlJc+HEWV4vRjcvQGj6XGOytZkb1UoUCkyyZRfIBkCmEUG4eCNHIsochrGplUBscGa/S0G8
hKzr1kYPsnwSIfo09tapfwSsA9SOJ9cQ80t9R8UgJ/7p15bRD1w6zhQRSr9rkDzXgavPGOX0kTMo
CnYEkUINumUWMwpS6v20zRBHmzdg/3GTNbhH40ota2fhGGJQiHNdlYAdTaxXF6WAMl+pPb1cDnPF
+gaSEobVkqJsyjdhc0Euvy1Z/wkZvGHOYbgr82G0HpEZSJUiS7075HYdd8XxZM9i+ukeAZ5/eOwN
a5xf8m9Z1JD7E0fnlbnBB13fUEBpMbdErHTkFi/AWNrIDqP244NDwpX/dx5qXGOmgmPC0wG7Iq0w
TwLba1ou7J1Sl1nfzo7zc2rj8Dg6hysd0XNIoXcqleduNq7pnYFNwRuM4SmGEdBhBMa6Es2y0bCT
uTtE7LyJUx9iJkHoM4X6pGCoJyQB9987FGXvNI5X1VqnK+dVEU5WjOYsCqisPWKxKVPKfv8NY/9W
ZUJ/ZpmkNPUkZOGpw3aZHr2TfJQV88mLlzdm3VmnF++BrVSK4CzbRTLbexZYTTEwVHppM/YMGCrC
jzJesjSSMI3FdaXOgWgZLmdilx+jPHlU+mw6t43+RDrazh5lS4zZmMrdWb5JXm/9tlmTVmoJgOk5
oeoP3IQdiYs8LKGYYRO1PYGE9mjzTPTTzZ7FOPAQe+Dw1ptCS+fHuIWiNBFeLrArbSjqNm8IsBHV
gyvwamja8P1MQecZU5ey1I1fPrewk4Lyq41xiums2j9iIQDRmnFN93CAhQhzdko1mAVSk2ClViDr
zQqGVlv9dK8/+Cg/1tRbF8MA1nSwe89eWmNTxwS4Z01w18LvW8IauHYz+XqogCs5smgNBrthjYVN
JD4uTBaQhprplbTGgt9uxwp/eNaS3ul1betejkncOzlouJ1g/7mTmd8wxtfAuxdX1CR5I2PS+VLw
djeyu9ChIZ8kwybaYzxvDSrpObHl5a7j67jd5hlsauuDWKO5QOcmgFFgCEx+r4+ZHBv5RnJwmVqA
S/0qfeNGQeGnpnsfLjBpGA9ePCAcfUjVCj/wS//uJdlqcbtHc1WX4NXOaGvqAVmPQWE1oUmEeI48
/VAPxjRCbM3U7cBegFuTpiAUiVpUu369TTOR5ZJeGulTrSd3w+lL7EA8A9v1UdBimOepqPz1sJnQ
MdhtR2b+9muv+/bd8hCux51nwVhY3YTWjvRTqgoIAaWf0HAwHTd8NALrlRQwnC8haCJhGVpW33zq
7aTNCJZHP4nWB63/7sXxvVHGq/cb2Yvj1896DhIzzzDmlEBiho3WuUZ9AExexE+itURoknBsm131
C+ARIo8quDekAzuDLpKrDjFvzMthxNWKeEFxXRdfdjrGY3oS8FKzMV4Kwbheg5xoIUUJufk6ahcv
I/njaKKgquhc1ZxYWhtZdRaJbQCS7QarThbWvKP5kMj9aRT/zgtepF8/uUYXE6MkQoqE6yWU7ntM
nkcBGFmL4rX2xGIqSywQyQ7+Yt/maTPCJN7x0xCcWmtTMKIFBgnzpQ3NlALJeAYy0/SLJDkaMgU3
zstwiY5ALccs/7+IJwW1bODtZswXsbaVqjsn/qKOSfj8QXFr8TOTu3LZdqiAxuL0Hum6feY+6rpQ
zPcCia7B8yutxDsgrA9nI3rrokSmEznC5UuzRTchsHtg3RxkCXU9o0yE/GK7a+6VIQ3Oq7mPsYNb
y+AiKJFVuQaWQSgUr8IU3nJlOvBzVjgFKKNllDTtxP5cHY+9nS2sgEufR5Ec/+a+xj9pMiTiisYB
GRpu62EEWqPMnCV5D96FWajtDTLVB0+Y2bO0PLKReyXvEgbvzXq/7eqj8GentYKQ9UtOfYaUOYqE
28gNALSfzfveXvh7d+IC8CG4R3QUzhy4KdL9hZcSdnuiUAkkLSGyWqBJflzI7rb8klmM9/UfpHrv
vY8SUNCqN1GJFAlHQKft8D0A5/ehhjFJvVtBOQx3m+7jQ25DN1kEYTDfH//3bcIu3B/1XwFXhtvk
4ezF3FnMQnLEKl0rWNDt7254RrknAvgZamklRXfPX4S+pKtoF0v1vrbaPjv0OajUSqJ5Cdv6RqQJ
iEVhHpTc5yeUZFOqVgyJ8ggfxhGfmg0E8U8G1EE6f9pnwniPalKhaBSv13sSueqKP/ac4uPDg7cS
MvbcRRum8kI2yP/zOQcm5H/3mEV7jTEIsMGdGotCVnZp3AM+fN14ZaBbb7POjpQDhNdjM3L3/q2J
Ng61ETUREFH0UwAJnC+v/O+ecJ3MKrmatzsBi6Q1/Fd/Fghvj+9Uz59K/5ZxLEtI5SGVnPctPlXc
WFIg5dk/uZKyiigosa0jtB/B3/0J4rzsajbbMGL00WlDeYTcROhNDRTlr1i8buEK9NS/dEhZ/qIR
CE6XUMDYxGwRMit4L/wBnPhCOMQqLb1TlHSHrrC7DO66USHvJ8kYdicyJxGNeXJx46rfMFHV5gLh
79AlX9ek0bXQ0gM9h4TMu21ZPlIJ71rdwOgPGaVq41AInVrOpqtkq/U6+/MQ2K8YjsaoFmN6uAUJ
jV4KeG0wNgPXdgatPH/Gc/R7inMsvY41SxS+vvYv5jgIkfxP+J8Vq2gqUpVFWd0iP2qCh29/lhmV
jbAgCRz4CSJXssivUcP8nvJ8U/UX60+QMq9u+Er/oo7x6Fn6rucetT6Tb7ECxdMhrgklkcMJwlOy
EAErAJzTk9Pl2bzKugwFRr23bvZ9rdoen7tfWB88hHlEVuApsvvwyowrx/qUBP9B0egzk7eIvHdR
MICPkpi7kAlTbTMREr9sPp0wKQSVAUQWegqY33sW5F+8FqKRCpOAbjvYP1z5wPaoO7gumZSiccw5
z6n+CX8odmooIUpbg9XXy0K7L9s3fbUVU2totY/nmteLOqlNz2gRrsIUt8jGAXMac8QgNRrHfXw0
QnJwYno8M3y5dkVlvTgm31FKNLcZ3+I0xrn7DJ2tdyd37Z26c2ByXxQOQ8CkPCqL6ogPeQigBCRk
fPTuA2mpC+ZxZ4a7Sugx2SCzdsp3L66rFi4kEZwJ7KVQNbUyt6XuFJxKxy2h1qv3nI0/Dk2zt7nN
r3FMqHjXP4vvfwjBdtsybCqJbkmlsrAljVwCEKrNdhVzn9/oiIyZVr1YC+nq3v/JPjhNJQ3hmdWi
qr5PtBRDD5sNe69R51J9Puk77q5cUD9fiy78eVjYkAfXg1GgI+zYjDhbDg0PAXHQL2gJ/sO7Ygvi
Z8dTmeDv1idKeiaTkBmZNFGScCJdxBJJJiKM+efsvwYGefFxBQ+V8WC4hvtAe6F2g/jsQbJYHzp0
uAwRTqnXPqyHKs/7vFF0ErutsP/XS2p57iavh9gIQ7Qi1wB49/5C47NthQald5STFWG5CG4UzeAD
LwMm3K8iBcDy0TWK8JYBzLAQM1imdXYU9DBfVdgRh22b0iZMCffUlPe0VWl0n5lpKA/ZUDfYuHtx
HbF5uKDSKzBIgSSDZvP2VT9c7OT3+shxRgojTOVLyWzVMjLMfYrwkenGEA/9VerFoBRw9T2zZiw2
a9a1fNJQOeQ9f2m5AqlDLvXHnJmyDxIBcIMaZMyWrwOROXMnu1ZyeG+Bkuz+SDlrYTrNS1DxNd5K
YjS7gf7YhSe+aTqe1Gxo11WHDy9ckgun46rTCtOvo007iBH4F5WlX6hGFfMPUqTbHN7RQCKApRkD
F6s1Tev0IEdiw4U1fD36i1VDUPgdHAA2mecn1b5b2dU0Xqyu8FqPZZGQVDTQ4PR/qoxOLekStRTR
XjDJS1Sc+JjF7+Cea0jdoh6VL1T3XYK1hN9PRg/ccsQ+k7lG41Bh1Kq2Q708P+Lfq7RdG/Q7upWw
Ce0Emqw5wiDPdvF7DVvuC1D3V9FLHQRxqYcI4keozdDWoNl9Vz+9Wn7G9YUECMl/SUprU2ALrA6S
jNwO/q5K1xuQAfmHhsgtpZShTeo344BoW0ls5kcr2Fw16Bd3ZBYzImKRUxG18QGOPkOFLUARtN9x
Sg6hl9vxyZ+3zKZPYmKFExXcWQf1aXQ6myAtpu5AV6EDb4pk/S7bv9jlEDh8kBr5jAoLYWAMguWi
59C+pV/gNbdE46gtmpmFsvvXQO44JzphxRX6iKfPg7hiJ7E5wc+EMdKfjEq+tjfJ0NkBWAmBvO48
ryLHJGpLRC83wkWI+GLBlD/3Kwhk3E3oAw7WI7cMwxK3qahbJUDR5gtrwP1nYjnaLSpiQE7yFwGf
xlKRDOp7GvJL5hgbuaBEuXVdBFCLmd+RbBUQ54a7ZR2zjxX5kDYvI5UWV75NGWArqDaShj6/sB0x
KCheCOm0CWVb3TO6fcH4qRad26ZSGLeB4KtKmPGDPr7FPEN/cx0o0agkzET8qwC65DHbiuRYqKfW
UnZnK5jXhifiplVaBcINs1dnr3yHPjBBJJfmBkilN7INlVrIw6ZRiVWUIvjUC+aCGmlVIuqEAeSM
popzVIo9RZ6s4VMLjUmAmFpbsHxbR3bO2kuvBKGbmLbg3lDJ9ZYNt27xsIie5Yh5fskVYPwTqKqw
nOepLi/ItkYFomuQY57cI66tt35D7clKy2BRvSOBHMNOMKE0yxc7dj42kamWLZ7XfHJmQ0JU5Il3
oLd3UoXljn1RbgHG/ilBgq4byENQE0PfCgrjsPyhTr0Q3H12DxRL5oQmmDIK981AsltcmdDc2D10
qQvK4r0KdfBoljRoGAF0zhbRWH7t+/R3R0fuDCsOKfNkbRfcbLAgmRPE+/xyiqoduHg0vquHMswA
B+HQXidt8H6ji/+KAXpqW2BfHx6kd0LK04yYXBCgcHb2In9SA8PGggQGTFI9cuh9Nv2ZIIbdUFCA
k3Nt8Ai3Bhk4CPe1DOexZAWLsUxtMosK9y2r6SnNpuxV70tyZIqHZ1FTkeIQ66ya+kO+f7xiYGWc
AMSXqSchfC1fzj4dQWoUd+T81h9r5BhIs+Q0vDSLWZt5Hgc7d4XVISbxiEtYiAIBKeDxATgILXpZ
tegx4jSX2xPO0fUs936TsxVleZpZXzsFkAyxTPQThShWgFVhal4MzuDQEoSkByIQSKlQq20hB6Qr
3OCcCSsmCggmO/gNCGX8aIcdg2FZGJMsIwad8XYmpmSAEoYtUD8R/J5N6K/ILbn4X4eDyJbTiKQg
VLbZEK70kHHTagbMwebBnMYWciE43dDED3zz+lpixNSkQnQd1WLA3GyNxK+xc0Th3SISm0Bz4qjd
ocQGW0LQfZPoAwlHb86/WzU06Er0cgOZC1aZMufcyJRV+WaGgVyeHgw44mEnbfS/uQlMe298HABR
Ol6WbXolRJK9/SQu2BEddoXvr2SmZDEB5LF861aqmW9mTsBiPwLWpt9cOCB7vXvPyIJsEEXpzYVY
p2G3l76R7lVzQZe+Ih+l3ogZ6jA8vHcf+PcCnVeYfFfqLcDdKuZtvLsL30CoWCBj4vK5CxfpiF9/
velxxkgl82+G+VLkQLD1upOFp5zPl2bThtAkPGRnqCJ6bjMrMCROkyH6DPIy7uX6EYAX1quAsIMO
54bQxNdhixWaos5w3D6zVQyHTSB3rgsf3ajpYV0GcgfUQu1EUkBQrOMoH5xCppBy5eVKBCYDZB+H
jcABgb0CJBIc57nHuMDXdh7LVw9EztXBuS39HBTsl58sblB/7KcY6GQlXED2OTImEJ/D/4yPgwcU
EFXh3wXZ7x5lhV0qTKYk/TCeAhDTWfMFjS4XvEiTguIoNRRf+XmBSYtcLnZ+okJOHI5ze0Xcro/O
bNZSF0N1OpLjm4H6rjJPAc1LZcM/X6UwcNs5YN30NeoCGVnrGOk0RG5by/84rOPQ9Q8xItEzGYOZ
YFPnxmnhPMpihr8yAPGMxeeCAC83H4D4OpvwX+DQ/ubgut3Qezc+hatDy5Su4UxYhW1Y5AuVox7S
Les1kHvL/NPrrygiRXfhgZRNqDWER3fvuKTrKjprmRpOmx5aQpCgkN1JHreTGZSY6AD1axBbz1kZ
gVQF5kemBQQfscN1fwt4peJ02+n/7LMtU8Hi9cr2lHlTnP9nKZleCZR7ZYyrkqy0uO6ffDpQo2OX
f+l/2nyPhr7p9I66W5dqtnCSxL5wUxUTbeCH7J8ldSA6MaBhAQnjRbxk85puOn+GOZuhYCYH0SnL
feZvVFw6/NCnMRDTvE9x32zBc1AoW+G2XeHnlb+HZJmWdbROSd1yMEvKMYQCATGLxsD6sw8NkeDy
3yNUX0q1m/vDwTPJ1iUOooEgsO/cdVevseCaznBQlwgs0/r0+41iVNv7Ti/uhSEJYPj9kgIzcll4
+4Qgui5x7MJLQatzoG3JlBWidm+1rdEY3b3teyzI2siEgEPFPrIVa1HrhnJSZaJp1l+Mrj67U6KY
GoWl23KAK5NceYoq9Bgczx41o4FDFMzVlYxwDCc6c376RKHMRc8Tt+uWDhna0n5S+sMQ2WDqlwVd
wPeosJ9fLTqZciX5rsSrrc6Fz981oCYoE3TJd+9Fcdh3Amn+9CUzJKXPgu/XxTgZ0RZQudxYR9ti
GxqrOFI+lBTzVq3u/9upg+rD2C+HObPTdYgkAA0OYZziq8gL26re5v12HwKFrl5iHNIiVNfZQNey
A6+4Vb8fe1wgtxdIo4ShWX1rEBGPdrqQjm+6/QUQtlp0aXw5h9iRLf2Y11meXOyZJVqBj1a4zHDB
Av42dGQ7/lqdTVxXaX0q1+fMV9M3pYHAlnNeN+5wtyEyZqljV+U8bMDuX+H2ADBzwSSAvud8r8gh
Jxu9CLQNGUDeADeIiU9StE9/PC5ie+nayvYwFsVvjmnXMVSZ6apU3+NQGQgBKqaNKSxua70i3+qp
sMpR68xBE1sbWyQEUVFzOt+rYvUbSLKedChayUzprfO/3aU8MLc+mT2FYpL0p/noM2fmLB4cWUXU
wdYSomfgTwAeRZ99faY6dX9+OajLG4hxlDj8vL0fRHpb5LxoCUrqXoWtzfHpFLJUKtRNh6uzaoVR
C5GITplOtA+60sL23VOYIf8Dk+FMo0ucRFCBpLv1o3ZA8NfyJ9twJ7fVdZyL4Odey4VL5dIH7aCq
5C/INiwonW3C6Hs2dvk+/AGkGejbLIFBFXfTU23aBTXUDWqXxTbP8MDaV6Z2lwyVw9sc4nUSAZoM
iIlNMZASZ0l3WlF+WCGWL3CWp3+FRT9n7Kbb0zFrb5NxttUT8x3X50Gcv4ACaQeyzRwVJJGOh19A
xcfYKBYH0uRbvKymspEMgVbZcVcdC1FDqdIruzgntlfR9L6fiaDD6JoDzgnlvS7/NW3y/+s+EwMj
+hOpiruPUMpPBr0Sl3mmK9KX1L7nqs7OSpEADs0m6FERwmxo1IwR7fSPeSttMtBGeikSZ25RjKJ4
AtinZ2xLzWngZuPc8fQp0w8DKYEg+NFwCsSkl7r8sBiD1bEd0R5xRHP3fnl5KY/4lL8gzCo+Gran
xoVMX8jCA1BESRVfoNb++wgGRpfsx/8H6zk1Nf1R5m/LxmSyJqyh1w95cRoTDegVJIZUAy1qufFs
ZNgL5GrZe1EoBjOrmEPB5jeDJXlHe90veYP+il3XCG0b/p413GLrkeTqhtK6lefMn8+TENqCZQA8
qYR8jFR3ussCtsp4MN+MjhmKCg78iLVa0gsnxaeM4hbRDHfvoEXO0K3p0xFH83oeyXw/DDsHRlhu
TCYE0COyNdImABRsQG5IbMkOOswdr4ajnZemdgYxOLfcC6N2UaOJzKU4U7GY33sCjiunUe/AVxsR
8LTY7SJWlBA22yC5KGvChPG9cjDO6cbG3y5ujO931QMmmz3j39fwyYxwspqdLAudShaN3pSwGegT
plxbzYhX8J1+cFmEXZHHnmlmTE2yCdsAY/w26fIW4h8DbmwkjhMHyDKaHbpxeDkTadWxKwOMfWLl
mEH1/1wvsTANhOOFxX+Em1wyJNFi1bumyPn06jizl9/rwzUQtAp968WKMn+MKEJYB20eNFEbGHF1
lCvEBB4cmeS00GNX6bh6OU7LqRFO8wLLVCuGLjl0O8u8Nw7g2mt9lNB9zk8ZG8ZInVwAgpxA1scY
vRMkWtGQlqmIa4ZjeihrwGYYsIur/gIKyN/aXnmsKT8xroVgar+J+1cbXxGOBA0MqYWNH9a0UJTy
ElvJNWpIay3hNyAtcTKMl+ja2NhSuZjN+yoNLdgAs4A1K4JA8wXqn3acGCjJyz3IJVmPnaghSu8G
ixNfIJ3pEIdkk38FMne5jtQL01c8LPF8JS7N2WKHUpp4AWmSulL7bsF7cWqLy+lbwyoF4x5t/LeW
ptqm1XfvzSxBzMySrlL4qLYSUsaCCyq8iCYgDSqN68uynv4dvU+rJ5NKgl9fOoh/FeA7WOAWPU9Y
85YytbdsSe0pZ3i82G5veL13pFMhmzZ/NStiYBZvVUivJrb7uHwEiMuy4mIMa9stYuNlhbDQAuTw
z0k+wLX/ZVMwgFIz1CNr8yhG9U6DPrysEsCTclpORnVw16aEb3Lf42AcmgLSUpEII5x8UucmPcKU
nnly1+jcCePPEiCnGjSmqvT0+5EqvbvB9PhuXBV2J9c3XDYIPZkJoujZCUNNvFvW5Mq/vXZJrILS
NFSN1illC7IJAvLSzEGym7jqLZ1mkMZIRPCg/A2nKyl29dREDlPhf09/uECp5aw2O8oEJoqBk9Or
6aZTAocOJt0F1bVKXTXnCCE3fT0HzejOS1eSwmMRppYHIzKwjWtTg3GCxuSgODckNRpO7WHc8l6Q
jJkioqksL4ZxtiBTO+9QTyJ7tIpdr1gs5FghT8uDyeDLaIO/HwPo8OTiYFmO7CC7XsuNQPMby/k6
tctnOeKoYVU4C1QA5hHh973WGokIL7Kb2f+pU7+fz5MM1qk3Cgs836rb8SGHEcA+xHGMTGcLA3PV
zDCt2Kcwg8NIEJNkA8j8/NHlP/4AE9q9RAxPmv6R3Pa2uqFUzaJgyYjOBYqQXtl5ahs41brf7UQe
aXx9b9dpVKsh7ljTV1JRK4I+uEJpzISWXE3ueKiYzvYVcKk6DSa67iYGcogtuQyAKWzSZJZTAiu8
9ojnmWc59Ic1/0vbGwE8Yvmg0LL4OqeIoNw6BqUhbmwTHtP/pQUlQ24BPZBXnA61I5ReEy5yic2T
OVhEZSNLUZgg8HvphLPCmbB7xtDH2nQqU4i4zd6ibWjrA/PJ3YYY2PaHQ64E+DAYwYtFMWHs01sa
AN7esL63k7NnUyqURFcyka5V6UF0m1SnQey05hrvj8yhWFcBZmaXEhLDs7PphbF05oUBdpNgsKjm
kVMAlu2ehwXSfCOtXHHM265lb6yofkVM0e8Q3puIet2Xlh3t+k6iuwm9UzH1txNJC7ZnntrVYoPB
m5Lkn9zcK2IdTYFDm6Bs4lBvkvPAruCBwKzy93nUNWLofnNd4H8xKNnVZFTqhaoTnrgOLNJ9JgPz
ifAs1rnZLpfQprcK3gbP2If0xnqdb8ZXzlqDF8xHRE5E86UxY0zj4RGMrIQ4t/CLP/dXwhGu0azB
9oTAa+rTqbgMHWScn7Dc6GmF/De4iYPcNk+y1w2Qbm6jtUcks07+rj57Pa8zwwcX2fCAb/yuMzf/
iglNJ6kWGjk2UtWpiUJ3xat/h1NhC9+pXmZdeTth+WRISF333hARrDyN6BvmJYG1WDh1UURS3/RB
5b+ClIGwp+/hZBSyf3f3MgTOc12rFNwRHFqri5OullPawLAVPufhdxT7H8ztx4rg49n0dUKZesu+
1EQOiJ1ehZJbVphwj1un64ESBQ5WzaVtmeB/NRpB58UAb86qCjOWK94XW8eqlcTRkgF4hAzHiVJz
mGGF8fj9Zi7IVdPsLN28pB/HoSSPvaFJzwNDP4VjNmnEbKTe+hcPbz5GjU3kJ3toEv5XIs0qOnZs
7tpFlgI+jg/VEco+K9K9/USQayAOwj++n4CxL38o8Xlwq4vXf6DgFGePemHm3MP2ndH44jspgd9m
twLfxeB57eTYzL1ikAe3sN513xSnlaT30UWgYKIc3EGIC6AlseOhvcrb98zojTaN8tyiNyTCzc1e
TqKZL0kXXBaJOMqHR3LI3nA5gTDp12C4Lf2eQrCw8gt43oorGHewmwynAP5AzbXLl/JaeSnDrr+j
b88ZmeqfzHm6SzzRuHAVWgSQq4lVqETwSATxr/eL6TVd+9tg7Z80VXhLe2tW1KTbFtnx4SiUhQva
uqVpX9EGWT9+PB+YP1rPc1xxMz8TBr4RxTrGur5s3yRjAR/13NnU68r4rst1GRJBcUnXq2ghxh2W
HJdzHnaspJDkbRB2EBBTaEaekhVTHycJs7PSRxNt24BYlo4znrO8C32Ja8cvJA/xjo+7XVNkQMPo
niRsdXcX64GDYyQR2BRSKCinlXZrLZHYMp0181qkttEUA21BWXLOaJu7Bk6G5DuPZ1OCHlowBF4j
F85LH+0Fpqqj2QTsnJvYcC7NKPpVcZ/NeQ6+6axtQAbBIPhHuN5yM3y2Ml2N11XBkQTD4foENuCY
p4XYoTO4PPX6AEMx4cexHAwAp0QRtYJvsYpZaOzavf3k3OeOzzM5oZlhrRYMkYO7ih3jj5mH+nYZ
0RADCEKViDmrPppP134u+vnrffxW2oLOHETtyowM9TcDYbsHa5X30PCWaRydsZMXTgF1y/Mr2UCJ
aE8jvuwHwlsNr8ZmY8O7GOGZJ2d0btPUrsFU8cx7tiHFRrw7miXlXJXk+3QsZTR61cjOrOG3lG5s
IOYZsNbyhTooHTHVHSoGAqJ6p8zIH9SMx+7yhUrGNslSTBOuSw7bwCRdS6LiYO1RaeXd8nlBsyeK
yCy5mYuqLaIEztHkENQpijB7qhNu6SzH1WWiBYk3MaiBt8acoRdr5UemhC2WToKrRwfBS9RSfrGp
1S5/pfb8jSpoRzHn2x6ez3IXBNHn//GuG/G3dViqwrRJHvDwj2401LIXphIVz6I3a64q9FYdotB/
8T/5eUZ6pRUkcNAhVHddZ37EBX5Kf3+izr9iJhkqmMi73MClxICAYF7E15vX7Onzx2ikzwYfYUZc
GeMJjAlOzUlKbOIl/tM7KxiAdVFzS3FjBlGy7GZGRYTJ7XdbioOWjnIJOZCdiwpDpQ/uphQASRZ+
sOpOqG/E31WiGgEu6HUx0hPvATGXCu+k7rlPpLTmBM8uRcdXApzEtbnBqiz61XrKXmis4OH35UUD
7QyluXiBJhP4DYQzKrVH2/ESvG40wJp2E/8lolaIlQ/itfOxH52WRAMl4PWZcREPyovErwNiTjWX
RmjnWiUsPC9l+GOJxb2xKzoWATma8oRclp/i/iS4F94sii86khCS08YUs07a/J4g1Cod3ZhMzypL
C/yl5jh2dXLPItqiQ0f4IgULsfDNn5gAsp4PxQn5pA8GbSyqqoUygHDAX9H2LECZVob26el0mbEu
tcPNAquKQ7DfOpzWCcYM1GdzUVWxKTB4PgLHvyIZffN+KlbllO4hOir3lM/faRs6IYuxft2lAaAi
wAwIVT+VVrHBQfV2LszR15Zhmub6hQ+QcoI4tcaysOcpLp5s3JgMV6JOaHTobufj/e/LTHFbxTth
r97+eZEeOeSFLmonXEblQN40Ee1jgsRyYHiv9KXIkCGSKNH9y5N3N72yBJYM4oJsRWb4EKyK/qiO
l6XbJS9zv+Jss2SnZ7oYhGArQCsIA2FmwsLekQyoS5NC8fkjTWyKzxRcPOpSmL81mcKvrSsZEphC
BxWMgQ4iY+pFiwNGXC4LOa4BsNZsZGOD4AqljGDrVYA13jxixIN53uYqa8IAi/yLRD6X2YdnA5ev
9PPdOCJYD9eAszr1LNHrk6FUTiHb393EkPsBcFd8LWOO+iA6otSrL5pDCVIBCilf6DIjMhLpM7c2
VfYj4qp5VEml1m3FQIAo4UX5+wMN2QlsWcDQkEMN5Lnt0rvqDqdRuhhwwyhOjwoG5/VrrmIJ0eyt
feEwFdGd9By0N5UMVSjj7RZg0J6gofuCqIW2tZZLAugXX5fZKji1pbnIr91+QaWi6twoj9AEgSVA
XS6Yt/NhCOAr5Zg5Gg39ugJy/rJP66ugUVaztR0qu/i5/JNcTOgXo1sT871aiKtTm/6zan5Zf8tA
euOBFxgrgCe7pDZGVu7u51FFibGbrNU7RJFalK4rCR9KcdiuxT+5NQexWFM8CJhHy/rA7X6497y1
WkB4UYYXyxu84ArCCGqQJxYqWs/rlpTtRk4p9qcb3tSD7VuYj82QFDoCr3e0MpyBaDbhiwQpGgED
hreVvHMnYf6xAmKLko0XlkvLhCCUbrkBPlJueYpIFPdGtfkAx/d3Qyg/oqA6s9iutcPav8BwpWRB
Jnl7dZ7h+UKeqR1aRk4MkfKwjFVBV5PmYd5rKL/GF7defRPgjRr2ST7z9x6/w3yt+4LfJSD1i38l
vA4jRpJUb4ChWS3F1vRu7/B3kLa209uchRX+N6SR7RibKixQtcx+ra0haAN6CPLmjmAY1L4A94uo
4mm6iNp30TlJ/ayfrEA+SOg2rlp/IXF7mkAJvSQBb0YkiDRL4xdvJf1T46yeUZXTV35eVMRonfQg
fZ3Um/f88yodIlsV3WLaDfr7zNah8yXUkqhmEN4OCxAgPtUf7R6WdD0mbqG6uUo6/TxbHt6iqCDj
SWOA/uUw5I6l6jr6vIZMjjVGp9GAKMXV3w8K3MWdDAgfCcCW97F09OhMDZpafo7CIVqo0y13VmN0
ESqRwf2Tmet2AagRiI7AGd75umgSheJqijDcUD+7a1QT9t/d19HMOhsjXtCeDoM9zWn0vVlMJ+ga
Sl5c+of0mB/VHUO0pN3OGwq/rtE6UYRZVDG1pS2iUeZhY/4D0uNdELwgf1+Uy4q/CQRPZR09R/Rk
nXvJ2PwMHCxTOfQes1qabB61vQIssX/POiTBAYoEeoJD2S7NuXF9whiG9qC+M5kbDMXBXUSJ98ir
/hPh/NU8+Wpmcq0/TM9fpFI67ww9PoTt07zUNdd20QBqwOjmjCfqxW+7CpNkGymyiHli/lUo4cl0
OJ4Kvs8wwZ4olY1e4rnBc5phcYcu6xnPR1hNh5aL8ImnAMCVOWx0iObM9SJaecdlAS7LNZ7XcPO3
iPuclSf7VflsFGYXbXd8UIS9JCWzdHndJa8WkpbIawSMqMQ/hbGwx62hCdAX1SN7pXGYACudu0a2
FfKS0hHhCEKA0qI7N1eLf5LMaxzOOdrCHCKfBm86SsLLRsWQGmMLJTzZluyweavu3YzgmOvMI1on
hp9gtrCKzBpbtKLbBQF8ft/O6r+6KCNKeoaIh32yuzqThKqc1KD4ql+5eGRwwMp07aOvnM50XS7R
HYmfgcGTDN0F8InZEaNU6qKDT5Pzs4StPwjgaFfF1OCnqxXoJp5LkNCgHanFfAs9Dty5tVHtML8L
RdJ24G642SR8Ir4Q3R1+6w+t+g3M6ffzKIOuGM3N/Hem5tFGDMCFirqYehlQw/1fBuYzZKbRcxbS
VrWiJSrV3TbRbkM+XtzNy2h7WymDhKBMpObzxYJN+0TOmDXvWpQZ1eYIKsj8HHr/ml+vhsOQC24Z
d2Az/+DyPtvp1wOdpRcN91QNSm4JOUo5VM4vpRIki4OBliizwaEtZtyZvI6U7GjHuJOya1Ka2cT2
hFxniK4uSRAa3p7hAWE8abY81AwuocJy+Vnn50SRQ3pYANjvuWzKuMTTKjFe9QN9zjeE/eYOVcRY
+62UoJ3tA0ogI+me9ZoTJijveQtimejCFVwIMBrEAVi125xVg7kKYnTU98bimEcjSKeCGrCVFl1G
cyyjI7ug1hiwDFE1sg7ayORRTSA/ixCwrlS4GwUxN9NaoXyi+WSgR9BYl8lSJZQ8hcq72aVuB4hA
V3YGNmKK2Id7utqFr4SSLoHbr1xjbWZZczoe9T3c2jxByy5f5/Mf/aAbdA9kUABxmrPKDpzTvuQd
dLWBkcYmI09+26DzhWI+RkRdgB+KNWwT0VcOzoreuhB6RX6FajYj2v1RY9l9cYkHdG/2Wfz+xyM1
n3g8/XabF+eRsUn2LMaEQInLFUpj7pMMzSFz1wdX2nNYQdBCGm3zXCMLzAnEzNXlY2+49jbLK2jl
EnkN2osDC4le+ekOJef0C3+KKHciXWD13/ri5v1AdIkuvxtK+Exihqs62Q590ZLIX680zxc/UIye
oQyiu4WDsOSMdgBvERF9qMIFfgxQI6kW6E0/xPZDlkqSs9p/3lRVgCl9oM1rhNx04MAFVwupjgDF
5gQ3LAFTZQY8jo0/UNeQU4uGq40oA/2w/v5DNHvtUQuLmdQfdD2JgUnaKmPfjSqBr3NW+490yQzF
10QPvt0O1TxK4ZfVHWsztYmfU4TOzyTACUPVNUeXs74vje8iigRIibMour/f6LgmyTdjf4wh/vmT
x99+3W3y2dXTmFxyORO1/v9MXsFzyiKlzq/2TBPU3AVsYSIvsA2kU7wqCYA08Us8hkKLW/3S+hKM
ziiJzG7H1C6WlmAmXAmjG5FXEKcrkRyXu2J0OKe9BVoH48fEXGFCVH1GaEk4g50Xls3uOKnxAog1
F5SkBO98AFDs1oVpJBgna5heLMjJD3fUGRMjZHuU2p+QldU8CxRMhcG3oKF2sdcTZ93sddsGnLPR
XdBTLbJ2gikQrWkBUYqdvmZpJ7lPX5/UWIbsrHlAMiF/MrXBF9RRGellvNATxZRoe0vqd0v/3wyN
owM9wC97E7OHZW7q7GF6qMrTrPvKiK1dQ76EvFjqNVpX37VZKQ60cQfMGdg1v2HU5Z5LDuD17ABX
BQuQdQSANy6WjNIv3DHZ28egUTvKPKda0UkKTfjpwr/rxLB+QNJMLnJ20baW7AY9kBVzXXLxu2Hj
EQOy4DiE8x01c9k/N3BFc5QqPDpfLgar9AQ82htNAE4m1CBovbh2sQ0TswoNNUa0rwzU/5MZrDIr
/UHAT4Aq8zAT2453jVoTjjfizWSEwgA1hXq4ASIC22pw1JXzTUY2y+OKJPj6ufwQIXFot9rAzomx
VUL6uo0hHp+GSyms5Zp53Xn4CkQOVHgbtCH9XP2CpFGIDGLDCKrgFUb+i5mO0RnlR9uh23b6uuTj
QRO5WAfgAS9OmoN4Qdl/wKcYs1bL09iaB676liIEPxFwzKvxYPD6PtG1CLtU8nAUas3nQBOXtvtt
+eN8fk7m+mv7f25KGC4pN+AR0SOFyD+IqyMt0g1nUA3rUsiTn/ABcdMadzeBFOz/rk2CDgRlSXKh
qkj5GVoXLK1lcTgGC+tUugIFX3v/ADF8/HxtFpIvEjGcEGqyf997l6JwMGpjbI97aB9h6Emn8qki
OZA2m6dOYUuyCpgfY7QlApBd8rT65sNprdDOXmwQ63Uxy/KTgWmI5g7Nw3WecHDiZ2yz8HTqlovx
m+GrPKKz9cWv/uGG1RsdJ3ypKJoSZvMLJhjpM7kXBIYeiii6fsfwKwqi9DaKWjvCMa1H1DCFzRgJ
nPPtrsZ7IspcN4u2SLa+6S4PTSpJd0xZC133s0Xk89qAFUbu98n43FQXydg4HFeIx2ErSyUvsn6k
MWKwIGthdb/vHGe8hk4CLXBnhDAYIbI+xS+IhhnwwC/q+kpn81uU9bbpEoetnYSKKDYc4g4eqH/L
4p7KZP+NTUG7QbLrhFEehBcD2HQJffRskzCS4Q/dkqPRUfw4SPvIwy8cCdeI95jW/VangAKseyvi
FIoQt7M83Za44WD6LgqxhkadaA/unlR9hBncYWT6b5e5sc5taWKgV6Iab3pg/Nh3Sd2XsBIKeehU
jXTkQzLuOkfgrdAeGWLYUhycZDlkoz+NKBxUkJqCljha6HNFL6mgAFP7CLUdJCw/oxB+w26tLOzH
bCkJ7X4oRXw9czOQjigeX9PALXUvcB3BQmqbnnWnPHi3x6aPInPF8etzWYTCmfkWmUPOAClV4Ghi
/TU7gFDYvVQqMMmviO1l0RwXTE4AB8wXk/SaPiqaoyqhJo5EISLcEhzj1puSlSqykWAjJFoYZBoC
4DeTwIucqXN0CXS0S5348Re5zuDJqxxECuAur9lYYcmzR6nxqUvj4HzIWDuo66G8YtUUJMbcdU2r
k4WU8z+ZksOd5bUglOMMLarG9GAMf+W6Q6aYyh5oyH+6SwM1OOh8JWl4iBX5NyMcdXJ9QIM6ZE8x
V+HJ3TZCkw/ZIK+0pRPCYqAkfsZZ+IO/hluBnY5kO0Wndm2spNIBP4dadJbAOFnxbY150aGWMptv
uuD/3By50jyVl377frtp5/DoXp4EbCUnn24e2VqUCAwvsrjugJ2TFJwUg17+/PdAA/AT5kvRGgMz
84xLMq26LgJx8W3f7tzmpjzRqNGR2RXVyxNu6miAtWIgPtkWQuvpyhBcUUVT4zpYCv7tmxSH4EbI
NVtbVXJn4Ctt/V5j3Z77+X21TRYlo6pzMWCP36Jn/sJCTBJjKgWySSEBGSG6O698V8/ltXjmKE7b
sOOPigWNVZZtJykFztnboIhxkl/ZnTGHW8LFSygiKXv7sytSvXWD0g9Phwkh0VcfZqZ8ycw9Ih2Y
vwMufJoldnzpH6gvlE74v7t2DGj7Ibrl0LHkI81RlF6BHt2bnlTlodGq5juc2h/jeilJl5dLx9/C
ZjummzcQ8F1qZMg3HlsSQ2hqkyfq5zW6TBoV1t1eFr8pX3QzUhAEgOHYPAavaAySZGLy4YJoq/OD
OXZFOFkBoufk8/S6AfT4DD3Q2Qhu5VA6uLcJ+Edv/ayTBiH+gc82QTrnMCQPNtbvojwqph+m1pwA
gbyP9r1X3z5YsjO/CF/oLtOTIeJERINlbhNHEjnA0IzrhIWD6o/Vlbbcp9wNiZZ0H61BTEdejfrd
9RXRbSxGJZI7Lxn3k3t04nLRm6kR0PTUVB4x4g4AzDuiAZm2dDlUX6syjy33B3/FvIt9okzBW4Hj
in3RbTw2nu6AgtGv31zZYH8SNGPVVL9kQXAR5Nh48ro/XsoTyAf3ugUeeSPfx1lfQP9SRk62Z2dQ
D4inec8sUk56nCSDc9pRwS99GJEAveJQoBM7PovFgPoCvGpAPLkCIcs1vgHkGOUg0WlFlK6+xm5x
uSJ2s4QOp6Uei6bqcfqOpUDChfehsO5np61xnC+sBxoa1pc7Yj/rOTRZk4viV+l46eBqoBhQMZsM
dRDT1DbeXpvX/xk400oc96b4UsmrcBKmHxb8rGai+1UultVkDcqB1wVEfN8BLbWCGmxReUPD0yhK
7LHZJnwvrxkofxHpS2MnYIqD0jfMQu47anjrdDxJtpGZVujv7mWtyIGu2OHV7fc1Jybik16ODlEj
3G5i7Hd9U8gGvXyeuGP5MMM8KINWG80DbslMLGISNfhCxClVzG4dedTTzl41ueJJ4WgWaozj6rNA
LDW9mdAlIIyHwrOO1lnBNJuCqS2AEx/z00iVNrUsTTWixc5Nm6BjyGojoQWBUSFbOjs0bGmD6ylM
I7WDOmGmM0ykRxaFHvAcFuq9MdzHR0MQAm4lC5GZ1yLosELotI8ZruOFaqAEm73CMj276uv+A7l3
J0bSX1XeoSrG+D+08WX5d0o9NtQYylKAtZ3cABF/Dd/1i4kdKYCYDS67ruoCvXVtraaPDuUm3kBC
lFkhTZX5nkdEgMz6IY5vThYFp5UWmHWj5JUmj+T0nZBbNa3W/1xibgRKcnJKlux5ofN8V8appH1u
DyXVfNz1eQXi6EPt1ELvwC+dp7tV6qoGHPHGVbXM84GYFp60cgrBdn0GtukXhzolsocAwjivcC4W
vbITjO3JqVj0QlXRausxuiK/P6UXwoojljatxEDeJ/vNmsNDGnGcCE+B4MPbU45EqDj9Ui6PHC3/
+w+QfZe/F6qlyIls0/gKasHa0fW75qsOS+PfqPi6ZLYSnWHkgdLmRIybe8IueERKPePXekcyWYCx
ki09xEet+SnpArprOYlxteMSr8VuGs3qFpzB39tH0dlAG6QgnBDRWATBTV5Bjxuc6wIWivkNezuR
bymAM2VdwP+TrdQE1HeBpex9YZVvuMrxeiCsXwvqTX+Xx2q/DCzATWogR5A0P3oU9LTqgmQ0z3YB
zbtYS6WBH2nrRgqSYUkakQ+/Qs5vX3p8/lyezAlChDcsZwjgFuaxdwRlV14rWL+iUGvfzp0nf6vU
JbOg0I/6SRCEEvgKVlmrq2AsCmTtZVaKuF9hIZF/vT3iNdSbcryIwPqfyZwmfQJ9pAVDx7jnT0DK
8/w2N6IgoqOJi4xc7+VQVi0ksO3gtd+54pcIg2puFbku/+9lVM3SwJjnEbhVmxAII1l3c1J6tmDE
8RC5Sel7rPOkUhzED/WzdyKZU0w9kSQYGHUtA5PSs1hKglSoMGqEbZFgXnD2RfuVpE/M5ze5fzTR
U4KmTymxR/panzez8WKjYQtJd/WsiTMLKxbVucpaYgLEMVr6m38aZ8oublXb3+O/iX9mco5H0D1/
6HWIR7PwJs3WG30SEBzuwoKg4J68/ft9LajvRpiuNkhDxR2IMGwaRQr0KIIds6pmDV4/pfveboMg
0yJ6eUQf0S6RbCO1MjB+0Hm4qcFjIde8U4A8jI5BLmT+YZFQeun2PMLM6Q2dj0z3mmm4iV5NR8M7
PQBlMXXv0WMtlKippSXsyl157TNniLfnrq7NYB3ZxTykf0lt20VuZzDM2CIA3c1SVb7HjRNmNnhz
omWxV2tm7fA3dGs5g4rfZxLbyRYkkJEznp39thNp84DidQOan2/4K3/VDdEqRKjIGXfIPz2R3tMN
VUzafrIg3rdtcF86d+BL6ClWVa29QGn1vOny6DmLquxgxW2j2Bm2DWAVpeubOTO3GihGpGHlNFaU
mYiR0t5pH3EeecPruj7nZGf1IrRw/U5PHkuOd/1wTd0JqZTnhJMKQCSMK5L9uAE5708FQG13UNjC
wPtd8M1oKCDQIsLvD4Xm0XEUnFRsLcQMAeM3/BZsZMER6GHR8eRq+VGK+p3tYDLypExNZCv9QVCv
1cb66m/PnIQe4Olw5QA8zfVsD4LpU8EWYmgC3zHoGqNkF6fECvuzh6FTLybk5m5nt/Hs43fOeltB
XwGR/rilVxJo2lr/8eMDm5MuisJPJsvb0IdI8MwYKqDnmuvmyUtjBNIAJdAiZfk7qFHHoRYp7Lxq
8t/WqcHjPe1BU+tXx7/BeREgSv33NO/HFGw3chFU7Fj0LEyeOVEVSVxaoMB0//Aw8e+mgFpinOb0
fYLqQjI0mX/NWPnEqr0HbEtT03ps/ujdb2IutCM5ki5NPdJHkZzD2Gsglr0AxawbSXmGc0f24/wj
/xIBCxctNBp02+TjAq+cNZCy140O37o9iMfvZ3bV5+pOOPLZDyd5ln/mYudLxBulPxZ5A11Ld4se
QmUAW8sOfAIyu33HQ9+mwiW34htk4uAZf0JZuBBXc82S+L1wLoU/9Cnbrxsp0spyzW4Z02koxknn
ADQHBDBXqDZd6D0/+sofAWVOulpO/aHYYWNIPSl8/JpO5Kvyde27yKrpKhLVl5+DRISUdWQLBEST
EkdKS+ImTi6KRNAihYUuXq9PmaoWJvsrkwyx6C1qo5pvA8RLLrwbWuKcoYPzTvE0IqLvpcDvBRp/
quSQYfqjt8eU4oFaZ6M8CbgxZuxZ2g1gHQT9+ZGG3BfI9UPbOmyNZ8+CYApQzRbSHGdCRCKpysJc
+VnxoKFx0sixl4ZubyiyBzxd4wRLtITDuma34ZJg8Dp2olObsQ0aTXGcG8VIuRBzVlJGcApj3p5o
GN7ZN2UcI3nt/uDut6LPVqWqTPWDIV5hhPaQu8tvle+TkRdDClDwJOyGZwaa/j2F42LxVsD/FxMD
bwFWlhbTAE3DOhV8u0WL2rDqB8W6rHK8B6uj3TPDl0tgyHLXjdbvb4BIJIv7KkCltfbkCGw9g51V
7FK0rZtE5dmC0s8ChhwmIXF5VvlNBhg2mWjbRhvca+lYUzRhM1NDSI0WyLKZR+Ul+Vot04D+zQK9
TYzoIOvzjKzmkoQo5LFsJoaoV9qBazs6f4O/xwjzaY284bMx17ZK8OJJ4vuY1TV2Zn5MTO77RGME
tsIPJOwjtme5UinO0j2xwHC9AZMz7A0JE1El9pDmPoIhheiuE10GWxVVZ4yJJ4LpXB9tJIYhcklB
HznIgaA+7tc42taRb6fRMB2U1EgrF3lPRbtGrQkysMLCaKBHUsJPUjQrkwOH1Hyxs9vWmeKBxAYn
wLIE6GKo3DjgcmPHf9vZlV/UjGIC/jOYWyD5o0G/cZwZcLW70t9VBG1xfbtiKINXTtw0BazvXYko
DoZPHdxPZy+ZhYEdtQS47EJZaFpr2HDndfHtheD1UM0xAb5yiVeEpvueYSWlEg5+/VEjXkdBtktY
XSQBoK9UbfbVD//636O3PEA2wDKziUcNedseJPOslFiGyopekpkBUMtuH+HZ8ckmMC+j/GYoifYN
IoEFo2SLuSQusd/S1fujBIZaHXYh2ad3cODpCOD2iCQRxv/998alNC0m/8BpNpfYiNg7ljrWOnh2
9LNypFdrak65b66R3rgL+30l7n4ySGdlOHLzFptiU9MuvAIfW6YnCk/E1ppD81x0Sm57HhZPp+xy
zYjqYrLPGW2CPhNkrE1q9xG3DxE26j+kmjOQOSvAY5BUz1X9MLEXeox8nm5rFzSSpqmbYXcWL1ky
l378+YABwkcYutcbkDg3R3BOxrijIIXj7yc0jTl9dCb2u7imSgSQsMk92IcMjQ59/7/t1BXCv0uV
tKlb2H6to6nPAt8c5L3hGjFf642sWBCfw8hxP2w/ZZUZqwYMVY9xdJIImM/sZ+LNyefxH5dyd8Ni
CHjBQ9nt+61jGlxV9HuJt0+ETI4sndIQTSS+ZJ5d7RQ6t8VGsv0skHZhYm1ahZk3jcNFHSz2Iwk+
FewVXr3L5t3a7KrnOoPi3weFr9tRVM28E0NNxXsoMNNQESLnyuOQGo7b9Z+RoYk3A4g3y/JacpKa
ZZOgzflVescfmIztcpUi904PL8ppT7Uo+x7VxfFEyECloOFTBjM6WGQpWGZf4tfJt1nZUA+SsC4g
q60plNpgX8bs6O9zxz6CPYvMZiJhy0V7u1jGrFSXv0IajQDG2Nk//eTe0UxfekeWDOInOamO+o4D
uE0PwpwpOH0vRAGoziqCx1ZzZbkKTG9ZWpowVzI7tzTCBsM86+eMGRlwr1Ur6Mxip7h6UH9CGhfJ
qQRRRzvPZYJD4TZAOJ4filsfc2GGRe4ANrmbeEeJEsOI8KRnfBRxfmxDYyjEqLEAJgEl4e3HE5Bq
yRYI+0SRovb2h+N2Bqkn3shZDTjM54pp9FArFsgPa3JKVROSj3cPRn3Dp0ELgVCxQreXly6GabGm
tu4EBdzGgXU5zrPurpmC3HkXT9iSY6ippPjbYvJp2hnW2IcQMRljs9or1T1t9cWhEPvmtwongL4S
ood7zSnEMEFYyX+CHNgE2EHNGu7ng17KX7oZxbpAiQnEpCk+YhDBDisbpVb2uLmpnZ8vFJDfg8RW
RrT1fVySmGe+q6LFnXoD6O5hoDRUhNoTWpQ+sFn3MLcFH07xr8r8C2+1GUybJ8m9o0GH9/thDNZo
iGYy5FWnj4R0M99wQ7T7RGxFxOYAv0F5WDdRH5TCRveGvKQ8j6Ei4gGlp0FDDidxtmfkgZa0SxP+
QM7VYNIsfZZUwQD5KZw+iXRCg9tBNOxhqxYO2+GNhBAIewj/wkkht0ZPzrNs1fFOhfvd+A6F89nW
DD9BXDZpSXfPD4D+Rc53pHafp8b8HUhUS+qqf1rKaLUxYYWyJ+ZvbCDLwANPddbB38bLjPxfpRq8
52IUn0uLPzlx6yUbVRwdMra6EBMEQUb9HKITyUgQUZvplsIrzmUMOlg5L2ACGSQ0A685jQy+RDZN
7rshkea353dmBOeok+beILrxtlRyPfgtWK1j1Jp44mXpOPklRMa/aylKe4I0ncO806wBDg/Nw8Ie
zAaVpeWu5uSVBHakY9jtVfqahKd39j9iGXEmvwY6a3XzHTrgqttz4dwWXsfdfdWi7WmXbpdDvl2x
9103I1wG+QNJtjdH6RKvXo9VsuSn3MYbdQP0YnZGM+uGHWX0JqoPngUwZmulK4+feDgO+tDLkgQB
Vt2c08rBwnw9mgIGY6dpOBIeoCpw+age0BSKmSr1h3iaz0hL23hEFPBYs4lUhLIPizRYQZkqbwjX
uS68HfJ0bT+3OtkXH8GC9yW5WQcdRS+g88a1qZin9QzXkFIxt6vnhkUEqVBvM5rFv5CL5M0BQioq
2cviNZ1XwcJHPlxoJ7ZjV+rUZVchUiLgzUlz5yEbbd405cKqrmtFnq6QQGkLPSlaZ0Isbt+K2HOH
JnKpQhvcBTVmbZaagwupvtAMPfU6uO0+aOgN087WV7s9+YfmdCTTqIwVVE/DQo2WgenSY+vjthp4
Do0oEEN7f6Q2YynTb/CQKHRnDgWYc8yPtOPbmBlg5cPjlPLOUc08fzO6Yerj1kUVivl8dDVolf2l
vos8eyWN+oXAbjoZ6vSHa5D7Oy4VrTQCF4KbuifvKars7O8mQvnMC39AgshcERrLHXm8X39iM5W1
A+5SmmJ4+J3eCFOst/4vYa+PBWwIoVfFYzrfvCJuKnQBj7MYoEUAsSjvFwc/JcpAhhIFkseBucDM
vxXc2qTqnwTJ6d8HLLQ7UatQNM6QKqAIzIhyxVUhzj3LTBM45JZ3p+zO/HjljqaTIgBjxzk5U6j0
HXn+EWXviHbU3eMsjd7mRdiMxcc7ZnY/LWRAXQKGi2v2pPxNhtAECUBWnCGCv6vMEh4pJzKkg0wl
vuNUUAUPmuHfxdvG3qX9I2yF8RDEXuwfV3FhwVb2M3r2OFjkGZZsIdJWuVNspoGnFhRLoK0o04RZ
HGjjrZd1i1rxXT7uG2zDIP4rP6q8GytaB34VcokUUKQr/4EukzJAsioU6ArPE0EoM5wcWBj4KveR
81fomDdrFw7ABotCEw0IDGQZpwBx4vk7lc3iK3WMs+aBR5WLxpVFtoNzzsj3oa8EHSMW95W8jBhn
RHQgFRqlRBeS1jvT0Q5T++suiA2W0/RjDfDIhJizUjA+L3JbHum901TEX2b8PNIIUEqmY547nbFT
XV5UlfhLWcV9R0H6F7y4CDPe7xsuyRSS40LOPpA+KoPPt99ShkA2EftHztXIjbCRzaPaNNxZSWJO
Y3eW+Wp8R2S1aZJpm2sYNUCyn95XIuVM5u9RpzyQkEWa+LjU4IfI2MUhB+iaQ9PiHl5T1znCL5d7
s7AMnIiQP/afK9++cE91OHGtnAQZksSnV9/WaeV6tOjkiM+DEcdsiXHJUXjLsnDudny2/G9/CSSI
ydUTcTHcrnQLweaNjJw/3lmSEV1ekvAdTWR7doq2oVHKZX6EKx9JobVL0rxr0tCAf9aKdNz5naum
bGBZLd3QsNDxGE5GJ3HbsOhtW3rfDQzy0rH0/rSVGJTEHCsdUZc2HD6xtHlz83Jm55yJMvuKCYDs
ulmLUrpY9v4OhQBU6JG90UylQFfUc2Fge4dfPYQWCawzqBs4HS/lsTt+UupCXg1IFZxyLPbsPoUL
vWwpYua8daloix1IJLnK3M13M6BJXNuB0mc3T93vMz2x9pM8qk2IOvnHnO0ARfJsbjCKrDYIzZRq
p0PyR14iNW4Mdf36n7AthaKZ7BrvXx3rBXHXzqO4rf8EAOaGY+9lfkPdMAcQWMcEkaLOFv7CE4Qp
EcyHXuRdLobaAxcxWO+iPvK7xRwYy1dz/hl1a7OkNIkMuyQuZv22yR2DY0n813RctcaoZkOMz7X7
nFrHp10uTpm3M6PM9/nns7NAnwEB8JoJD79bvxgHaZXuTTG84kD7AW5fmb3l9VCd9hPciUx+j46J
Upkxgm9hENytbf+62raaLOvwdlaGth0SQS9btEEeMs+Njg3HVTvCpw3iC2AknIrPRM70o2UZp4CS
M1G9NqR//t/cEUH6aorcbQ/RaAoWahqLmYJcS77BtE3MNgVv689JzXAxaEzcLX3T8Fd6zCTOU054
/kERkYZFeRIhtu5t0O1DrxV1SRfQiwCXy+jFHLFFXLObcpLl2QzIPbavncRg9g9HVGIo9GOLZ125
B3PeQpwP/R/hFKJyCZwfwJZIhrOrdYjZ7w6lheG9oRHfhhtOet6hdk7OosPwvRUl895/1NAoW4r/
7AIbb7eSGFBQfakFfsAiLHTham6WoJwkaW2MsTayW1VmHl8H0Eo24i4Jr6V4Zl+dKz67T1ZQLO+1
eI7IMShr2wVeARoXfkKgovh2erLs2ZZonBxjK2OoX4xm2uAiWMiNFqbE/PCk9+O/H7g/Z3CyD3FD
facynCi/HhQa9GEwoLjGU6mKCqx/Cg2qR1DVUW2qr98n1Z+cxDQXJcMLnimz1XqHnMOZsTj6bBs8
cZlEzfKh2b3DneUESMD5769hRL8bZX6bibRsu/zeAz395O7RoEPexyX70ucMgMcRpP3H4SY++QEZ
7ACJV4jtBD4fbmr9ZH6koXdGKqiI3HD4S2sigyskaQvpEgmH/bLk0mZZma9ArescVefJx20n6GBm
UbYW2l4sHCBU2Rj1PPT6wCFYn3QwUSCVrnez+B5wP/IO2mY7pDCxbHHT/d5iNbcx792+Bcr+io7Y
xqMRt9KVUW/2qhrY2NCeTnYYpeQIBux/CI56IvgtPwFtiwD8xkPOb/OjOh4kJliEfIjJL2YkkeYC
usZYLOcG7GbSXFXi1D72V1TnEdvhud8RCM9MhQZ3184c5m8iyx4AM/01BdVm0IiNTm3Xig0cMZwy
h/rRcvqrYn4ZaZcXAnm2tagEHAFKzGGEKBUkZPtyFEhBIZU6Ir+4ZzD6e+4NcVShbX30QN0yI9OR
6KgXV48pByPGECIxIrd8VOSmGnESFEwTmin3AivM4SDoyIjCq+n1inhaxjFHA/5measeDZ6o6xAQ
/mPJ+KnXMYC+Yv3xx5/iEMvty0a1IO7hNNgPovKYaw8DhTcX9etSmLpiPjuIwlLvo8y/YC6Zucoc
1vCP5ii2Vr8LbifEEwUgOZXYQOh/svx+SqiUmTgiPaY8OgZXHBdSqZYj3n2SKUHn4eR1CFJU9A/s
AcA+TWM/XJX0HdTsuQXdL3lNpAOwzQvB9FCKOoxYt8g3bPj0UfbyaZRWsvS8alOQGCBJaKCXiKkH
QmaJm7u7mfAkiql9BDjjfu3zf+SAXmqEBe79e1awJupgSubk5RkhgbySMtscaLa8yIdrtWWzixut
rDZtrCiMmTEC5oCehvbr/EOMeowHqm1dlM1+K+xRSghS4iTPMiCkWR+OYv7oAYNmoLF5wymn61E1
QtnAnq+sUKmV8WD4Hc8zDm6WyBgilDqfP+tkF3X0ygdWrYTkoVKT+e5Dlv7gHzQvdsu3zLGGAgYH
oc2DvxStHy6kqV3mrb5Zffn0dWc/AQJ0pwJgnHpHCRNBOewDeJt705za65AUlwogAX2bfs+rFd90
+Xy0AdaNqBx0AnNDcTc9L2GlzUIeat8WeM64IbQOOOZGxyvatLZLFECpPWKGdXPMbcyrIRhUigcP
xWVdxe9HQfBiBXf61NwdcOgVewWLrNCjIMJ49sdDA09pSxl3IaPd+ROTdQgxO5i5sQ02BtGb2spF
YM2Hxi7eDK3/uuQ0HXttpcvt+NbOGdTMo9jEE8DhabFQLlhZEWy/OntzuFVV/fpRmaRkY1FKXfKH
mINWWY1N56xxNZSsvTPnw3tBGJqJXZmQQ4p1DF5WWNuybGhJ5OpofebEeNVEzWVbtJGSQSIcQPSf
NAfiV560XrzyLQWdpP6mDC0wd+UBL2BAoQDgUArFisb1zhxhLUbHylwxL/yoDmldSyrTtkdmGMEF
R6HFoGYemlfvKVRb58khqQgC2F/4I5pWNWn9YJM13DScv4spz55vPovPtNUGGOZc8P7Ajk+sPIDG
R7ohVB4o9GZQbIpCEY8EQs46h5BQQWssYsZnimBfV3j8+udWjOV6WNsf8pMvDx6LUS7Uxx1BkQeG
3szrPyjuB4uiLNdku5gr3qEtOOwNbBU3OhW1MB5+tStP9QVrNh5y37KeF40fux8DenjToBMepa22
APucmsxLbB5ghjOsOCgnEInna56KjGtTsGr1QV2Coe3ODBn+QTNtrV8IzDMdAqqzO0BV6UMfZw+V
K55re9vJ9OoELQKjHV7M4i7ZgaxAa5Dk63LTpvZFFfi7Q8TmGa+1YYW9HC20Yyf0CdbDlS/vGBza
rFasVlpFgNcIF77g72nmwzlCux6sMT5r08MYHr87z/TGbaGfyIQ3jxvLY4RN3cYFwNnlPWl5Sm9H
60n7/UOFqCxEWx/Pv3oy4GViAKjcGKWVOssdcCjHrS3izN5J6dvndh+/1OKqi9uMS8s88oaNsI+Z
VPi7BXfcu2fMo5TH/NajYYtuXttjGYoeSzHEz8o8eW4oBDNZPkV/P4tFzBBImQzoSJPTnhJUB05X
g/bHR8diTKEkIGe1Iti9pHZQZ7qWS1G+t1z8398FiTPnp64lujUShr/3ZMpoeueTu6BHSRlKF6G5
WU6Bn3cPR4VuwSLJq2DW2ctfU0u2UIaN3jlkKwqDIsFezUlTkUvrO+sp+6lFS7mMMRA5GxG97VCo
eORxXaKWcEF2JLcGrJQ8vcFS1V0ZCm0MT/EMMBQoLBzv2z42t6NUqxK++WXrhJlg+AN7lQM1sVnB
V3zpqndi9XWvnKsh4lgWgfZV1N8bjx9/eeY5DPA2ocLCTQicI+YwMtrZZkWd9n0jTJZwl/6sXryA
RcvqedxYLw4NM79365oD0JfvESu2XbLrQOYxttBq59Q6LhvwnuZgrETv/WmxH1t/nu3pdb1x2wgU
Wp5/r5KPwLutTwFFrK0zUUuIOV8zjP6TQQtexkrEHqncM6Ayb21Q9MDMJOAqW0Al+CN//yM/v8ho
oVXMG4KNbyjaIR8xR1pds1he8Osc47wrTx9fpToSEhYPx7CDAy/asMI3QOTsRmuSOYXWlbmuY4mD
tJoDPihB44RMqapN1+q+sLA7qIVMIhrOF9QumbxJqlkXI+wt25bd9A8DgNjlY81L8r88aE1VDsCC
047khyPyaIilhoNU9mtin0OrtU7Edy9MEORYhHgnPjsohhwj1B7tt6ylI1ugBUBRxZ1VgsY06+wm
wvAMMT3Eef3DRB2VLxTSB/AOXT2KoMMHeswo4ePI8WuwS0zDjJZUZ1Yrb72cAieUI7fL7UKrtwWv
Oyn0aMHn8tg+tvVojfWYIzpKivhkGejfBgjT4oO8RUUx0HmALzPBalPgB8VdgGCatZUBVPLF0VDN
o25XvbmgwUhEpCVIXk4E4P51KX7FtTd/SrW2g+dPA+A5tgqnA2UthuUYsqame1S+Cx9NE+G6ec6n
sqr7lWBEduorKUndHnLixeLej6KyzmaJJEmMbT2MBxao/RfdRResHaPcFQY7gKx987RAZTkwBePO
dW4M+Y4H/mta91d1F59Rknd9yzo48nrWxg0OCGVh+V9nwbvvyHsx6NbjTSHDUBxjTiPG6fn3mI6O
vhqhrUks8O8GEy+xl/l5lg5lSm3jUTYthBoVlRq+BI7T78bX42VbEjCry0VjZG4H91+Q3zBcNKat
7t3lKSXhSnA9izMGI8I8/J6eijTOJVWx4zLiH0CU56d05JqocC6qrrqACX3dJrPbsIzd9DbHAnWH
OGaCrTblxx0senMZJiTE8A7sYMNvJ/QJ/Q7EW2k8vRmK/M43QmX7ZwzsSxKjN+Y7OM/CwS4/1ddF
Sil9nT/FM0ilcNdY91y1+nWyVk2uYwUDkEm2F6ZozVSxSWftRsm+f8Jpb/YJibYJ+RdhOG1dYVHc
Eip1W/m+JWOuTNnswCyZaMfpFxJS2twj1SRNvleikoDiDdoVs/qzwJPqNQhV3FvDvVTvIsz0LXR+
vZDYUe5XbLKgLq9Fol/cQUPYrwDy+FpBBr3g18OEAduolyR4h6XSlsWgZlCfR6oWuVgCCqOjJnZY
TCurqSq9tjbdUY1n8Yu0Lr9NCyigktC3KcuIiC3ACGybqhtGXWdRoW9xWkNw1/z+jMyUt+YKEb/I
w0aH3CKFhQHXtTUQd0NWJx9ToX4epEdXNxagVyAijuhmbyP1zeXC7S5EZRBp0J9nhHwpnV+qo5ep
N9e9R96vIv/ouRU2OrqCz8NUvNJmCosk8+/tcHn+00AtGd8hxQqu+mh3lsUZH+3xLj0k1jyNr5XL
GvcG6NU+38Y2UOZtKmErJ9Ilrin1HYEfArESJckfg9cmrxxbVK5ZwemgH+Jv8NT131GSAysjNLRe
2Ie3e+FFOJw++mLesDutPdHbWdkD/sNv9GIHRKQRpY7M5y1j6Mq5wUnn2Wznc0aer9O2RLcBkGZB
Qvoq8VNnWgsxyQAnD5JfOUGMAadYcrMlhsiBZfkPe5B4urWqBOng2OSnccTddmdIh8tJYl0lP+dT
3rwllOo5AmBJvI7SNA53w7XpPJTjCqnE1Sq3GW69aBpbVP0Oi0NFr5vgfMz17iK9n/OOFaQmdMiX
hMH3hlO9BlDMomaaBgTtKJJutWF/lyITH/ltoWsDvBpUp+DRf4ILiRDfaZM5CX1EI/uP1xvMbchm
E9fYUro6Af99Kvz9P7A0Q4yA1NF2IYs0I25OLveIuzMTkamRHrIDaQ+T5G3jw8/vIbNMFVbuaeUT
ITRCwgnSiDUXGWWpe5raEzWwt+gPPbbvCvtw6uGJRycA0Y8kIlLgg0MxsXf+w1aKrQlCD6SpJT3n
yy8BwsrPoMvF41oaDPfIPMHSSxCayv3TzlnPIel6YVLO3aL5+CGQ+cNwmVxFsNcU4W09VK/0ajyK
ejVZ483R129UpvEHbT+kT8v6Vlrir0gIw//jLJo7iCpLoUBZwWFykC+Gw4L2LN1ug0LhEN0ML0cE
RKr7cL0w6KWJq8TDUPDcPQrCA2MHgTIV1a2oa3dDZnh7nxuJTrxXoTFtI2IRVkwchLDL0PhsevBf
ONvxvp5jYYcD8fkwoa2Q6xEq9lYefOG9+QBZY6FGUqO8b0B/dgTKI3uKKfqlStnky2HlWqaXGy2x
KpKhrL2iHt7aBWsJNtVua/T3pdn/z6nddP9q1uU/u9q4cbCSLbA8/4nRxPamm/XwYZWVqLyGawTb
HTI8a7HA50mBY2/pov90jfXUXSl/duyigg2IWAEdU8nfmoXJxho2cbC/aD7OY7Dg523E9+P5pGoM
6dJIX+2Wb4tog0JAgbLxCtGsxk4w0c0TeTsGuN6TK28RLzgECtrJdbnD5M9oZ1GJpVMGdwxQuh0U
/otpBSWtco5FOqwDyVni/PzVNM5d3sQc90SjNtl2NoSFtJ/SHnO7TXRw7Mq26x5SQEEsU4joHgUs
LY6mdB75DTxEm1D3iHEXhKOBz14a3Qv6Ibe25JufxpzwI85X9VsM6KVl7HF3PS7mw/+b8P1Xg4LV
s4zjHfveYzMmRG+lCZ1vY6Ho+f1iWPwOhF7NMGLkaau4nH0y8Y516uTMkKldR774tr+Ljsg2jUc7
WHVppcYAemBqFhqBD+fdCgvyy0d6Fg+EvNcNIZGaQ/fRBppAgXZZZW9g0Aa5deRADos7luUq4J5T
14RcmUyvUZpGpHT1iOoFdp7SGlGkE4yw4tnStBj0ywAmbJGnwx72xEBZFW2dioX9hOLIuOy6wtDK
meh06rAdojFcKiu/n3iWU4mfMU8KuyGXkCuBUxDdcgHL6Bo1ZVI930TA10XPocqPFKuvUV1ouQCl
QAa9cf6Hrfha938VdH4qCqiSgTBsTIu4421KbVlr5piMxYUp2rDBHv7Ih+o1Hj+GnaO7+oRTt3dc
BLrx8tDXIS2WEVJWWnV3aqc1BTIaFmIPe8CivImMOXBmJvWfygxokttivlQYjbPhvNvqsKSvQo2n
Dde0enxw8vi9hAYQRhU900GPzfcmAAWJ7EJf4cSO3iyq4rnkKamES0BT3CRzpdGaj9YpqrqG9Kvq
xfkHfvEXnQv5wD1E6fMmepus9Mtph2eAuLGtqtwNaI4qGf329YtlP45agiCUSX63v3/+SeM4gLe8
MQUOy0CFhaTCYCq3eaYBv6ognxqcQXYV5q608rKKSJcnhhEuh94OvOOMJg+pXC731gKyk/1iP3XS
CGUfqYuQjNooIGIF0DvA/CLgqyh+LtZ99b5E6ATSFyFiOaVXa5ITH4nhpnBvTyyKtIvL6/f07TGU
O/90Ph8etFGOis5WonZ1K1GqqJW1kqMaZF+gv5jD1aLjjUvjeQeuM/FWMTY1t/t5+O2RwcRWnmQf
1XdNWCcg2dN/9A5PGcFvM3jloXkBpbdvh8iyTDQuFTsS0cDILf2EFZwIqMu38i1LO0iaTLB6ZREn
+5IdtAVfgofPF2OWEx4zx8kl4pdRr7xJ/5jFc/hGhrdLpyLYiNgjGsUICxdKPbSzgUIpHCZOtlC4
liC6L+BlYtpCUf4TIHST6kXwt+zJFlGdJdZaAfZ0RO7Fdzxb0fAvdlk8imVOCwzeabsa12jDctPc
nUR5icKQsd1JBTvRY6HV1wRO4WTByT8i7q+3SZRqMAySC8wZ96rRaHcUheziIS9vqHQWGqnCR1tj
rzpjOSq26LwrQ4zmUtHA8dgsnysbyALLen6btum3N1TfqLt06Xoy3gK1iJEaW7qdJ39hTjbMv0qK
lnl8GOVxFnQfdWxjlIy6VSPJyfwiQ9id+PKlwNdlCWFWBeHWwmVM7olGR2EAIpU3EZ2cwkwbYINS
X5xuHZeGeElCdwr40awevQFaf3kg0DQTJLf+C9f/+b+ex78303Zzhertyb7ZFD5IiL4QtlsQ8JX7
jmyxzSbLyJ8JdlxKvAdCqTcmfgNN+bKND6dvTA4SmExdiI/Bk02WW8XmlTBDtbJWf4CwPuY2Zv6I
m1/PExkMyDZJqrFqqBSEgHeXuLHFvJjQrEMYhVjKkgQ6LqrGrdmekKWoa6rgwfXyhELZ1lvtgu0r
5QKeNqSrWnsS7ESbwfaD5S3YYdIj76Ro7HQRgHFoGQU9Vz3DHIXAsoLAeCaM+EOYBeGNfNnsi/7Q
0VL0OVHSZlUEuxUccQk+nhHguWGIQJT6AXwgbPWU1ZBb9CWeZ39K0zpQKZEJi1xtFyPt+JBcdsof
ngtCOTIK1fzRuEMtXLW0QYMjvLLKtuAgZQNffxjmLZ8pSYM9+3acBgfDJqTsl1kFpTRllNeTDBOc
oqwKt/53/h9EesuWGiQ5Vc+gi4dZKbGeWb+vMrMOm8XTCTD/LmvLWoAcUuw9vvcsWSgOPjCKeGWT
iqfZTZdMyibyKrKn7fhoiI4w8YMxcafTI+B/TotEVTj49GrYIgQb17SX8qRZxhWgQ0ASiuS4Ttbm
pt5EtcEOFVLC6TqqzMuyIPJJ0biIstz2nmkz6HvBBZSDQ9QGSseaJ8dwJNFks7V69YAzip8K7gdy
NknMNb9Sn6hLEyaVb2rKHvavRlrC3GwQwxN8bcIVqBIZPIxrftRXAEJyEKJHgtMvJcop4VzkBXyX
f7gneNkZvzNot9ooHGLM424yCoe1OmY5qwXDLswanNyeDqRRmZXJI4FvEb2E4AxCjG7DNxUL3H+e
6ziRVmjlyZ0lAsnYf2TV7f5C8f5yr8SK/PuPkM4FeBLjoh0nv/zouB8OrjyCHnLGfvoziIpM46yE
pdXSteFq+bc6qR0T+FkI6KjbMtl+WQoBiTf0l+VHgx7gF3WQIb+cXjfz9YWClMeWDX3tSR+iDJSm
rjKS2Jcu+nfj65AYtu6hXKPBzlJYf2cTb0+jHjzdBK1VK5HkVloGELAURpCkjZe3bAJJlF3K1Bt2
L9NzjmMbZKhp0G/+jQnq5OUmi0IbBtGm+NInGejQaXoSjM78X1adUSKiLkmLvYYOnwbiuUoSeOq2
ZZ1jeN45ldGaOH4rXHP5YyKuG0r22kbdUBLqUYG1eEDytp5S9fS5EMPy0JQgNsk0wiOLgie639V8
34fh6rYL1QEhkG8HifhuNZwM6hzZ2ycra6R1rwpB5q8qv4LZTrdnTle8DYDFXM6rq3YTRt+EWEJc
RowNRqGBmEqhOKvuvT5JXMbWNUC83HE8R5iZ4B1AA1yHfPQlj4qv/COa+57Mqky9CZmZGB/kIJJP
PnQM3vOl6CzulkvycOkwNRnSahuDXL8csRiUcqfzie1yNbAY9b/sKBpjvPwYTyz4m4S/1BFyhGuq
9QybCrs3lgT3Mcr5mhS0X1+e8qw5ZfJ5xztsF9L7lFkkt2msIC4mRdJYCxpt0slvLQHQjc1TcxH5
L03W6lSXmNu5Eau7mgrT7PRj7AVj8aQU95oU7r/oR6/QsjuSbImtI1gzidZuy6jXyjo/wLhmSlPh
RWhPJy50Yo6ykjvgfn5yBOpmQySwp/iyRsytavPZDanVvUzFbrqLgNKTpr78aFZYY3ar3nFGkPRc
HwxdjZFjJjAjAHbmHht1TcxyfKn0wb0JQGeKBZOx7APp6xGIPACalA3nYwi6F4WetabAapkC4tV1
JpqTMdtnUTJMflljM3GIj2+/QRX2rpTkeMVlGWBhHEmSDo0M6VBwZaV7WuHoiky+f1gCvAUKN9+D
z3D/5fTRI2EryTgJSG4TvbDq4qTXsXp9k2t2dTEzPypqYwhfIbNM8BbOLLlM5bWl7A2Dm2EH2wZZ
kNS6OH3lJtO2TUSSA3nWwU58dqoWxuPHU6vYDAKmbY8jkGdMbtiH0ABgI779qr34b7O3IdRzIviT
4Zpq+yMuY4F/cMurjvM8W6p78kuuWQh4zraDGtOIP5Yzyqv2R2jffDXfJPes7gOW8IXf100BeSyH
psJOeQaGg/dQTTP3TE2IdjR23Clq3mYQ1OGsg9FhsaBfqAETZ3AmC674/jDOqEpwG/rTN85EzSMq
+n/cYoNdgAdj02VKKZ2CE+3IYEWMvY94aBEuv+5nIWaDhLiINl6EHRs12CvubQvC5XUHK3yD98an
JtLznxVcr8NLlA/nF6AFu2vIV3F/pCNc2fv+ygSBhywYgdWjdX3RSCM9mIoOXPM2mVHMedoqolY+
fvNOzCVnXDtfJU2fXZYhwOs+MhPO3mGxPbzIwLw0M4Wvbn6bspSLJ2cjIiKcGGn24GIayQSz5KLU
iBKMng6xLVCsdsod5qq+js+oU4xznGoAIaX0rNP0usLACov39sTTZBDKIh7Bajpw86I9OZV3OSYY
sQ826rVUooESohN+ETfM0DeOvhUThSDN9saBjCWhkvGyOc2TK4BXHXBY84xSyjSAsfQH1Z7lei6w
s08tnpYlV09CHTh+LRb0SmUmHsD0Tz2eIoP5DGfmgSylHTwSOCo8T3G9qW7dPo2GJlCbgdPZKBFT
Ka5x65RzObmpt4O2AOcWTQcaQLmkdX3acXQhrFZBCK1fvAX+7W9UI92QzlktdWJcU+2UIj2Tknaz
5nFwEew0YMehUlUBZAg5TKoLwYEi1KnzvGyK/WofN3oRco/WTxysBLecORUgzvSCmpEcOrRzTdMq
Vn6gOEqVFceIzHlSG1x4XE2PunWdeOfAo5fnfZKlRvubdxSCKISq33cpt5+SGMIqlm5rLWEgdM9m
nq8F7HiutphQBUuV78/fDdATxEkH/lqZ/8zTlFk+71T+4QG24b3jURk27CE/RucdlnB215t7oAHQ
+cVGHu73ukF/nb4eXpwBcENLN09PalvFdSJQbb9QPJhClpP0WzFK1DBkNE4Muomsb/39OnjKdasA
zHPZLXypTEsuGwz6bD8CF4T7ZyEGMS0p/ga9u4gsh2U2paq+ml0javAG4VMkSRkprs0Q6Pvk1lvf
n3VPHHjTjBhEOgmPBcd7YUF4NwQKFnoCsx053PoDWkKEnAjGFOeC3LJjQjb3lREMPrWBbd1uNnen
eDvQprKLi+teYAoiVEiaghMTQ6j+V4a3aARDG/1h2jcyQ+iqdQwr3cqPA3WF/jdJGJJvusIx/OfL
hLhVTPx8mI0fw+PvuDCOkYW/JcKvbHxiLjJvu9oirhX1s4ecOdGTQri6gMrRynw6p4v9oicO9IwF
E+vu+8hirnn1Er2r3K4TP1ZePRWfIgk4q0/OBZw1PBlRPZno33S+LJKvgAyph1GmEjHDGpvuYkEn
zhVw8wACzMFgblDJNzhz4SxBpQt1jKbhLl8zN2oofgiQG9G7hzE7k8eDAr6FuG4Jk54IJPvSVp28
ssAJH8pdlcuZIpxQKYWRScwSrHiHebvnVuvJ0RS5AI+61xaO6fu/cM2CBvCpHKV0NhpyWtTIuP3w
zwUfPZEzrZdeApzgYY7uBCuVEwPWuCdTmopipFvsoJZcwOOjLkeMp0K9JHS1vKtORdY4wrL+zkbK
2hxOmZ5xIf49xhwRTnrB3C/epbx2lrBlo4Th011E/uDW/cwI6cvY2IKTBpLaRqqMgbS1u3GMUbsm
v84P6T3tPQVzTG8/xvJmHxV7x0rWiEYmFewMWTa63dHRnkwypeKOxUMUeUFZD1VzJ3SjspTbm4L8
G79JxeJ//oeZrqNVpxNmCS1MFGJ/ERFX68Blf1xADh3GfPLxFYePE+DDMmjuvyytqE/4PbmvL9hx
ACMOM/FZzUQqOxNAsdOxizBhPe/EGTqFAlzP5U2QVmqhYoUpLgGILCtY04FFGidIMPLEuQR9E2tW
CUU3Tc3m1iFgPbdA8pxR3RCGyUSX/3ttKKI6YDym2k798mjXOhFvdQT9MIVaKKxTUqAbeeH24wrI
7PVBi+XKw1JVPWO5oSDZXEAQJ8Nb6vgFbQtHfRLNlN8Dy+snPLGGbz6qH6JwkJ9/uVxuiZc8Rf81
GMj+eWKS8Bl20NIxHCX51LwnzwWWwaa2IloVnmYO2wp0fyPGFtAssbd2EWDfIAId41TB6ohXEQGJ
RUe/g6qMa1YA1+1CP4WXe86ZVo3HZVm15k3BBAuA5qzg7d0QxGK+Zwj1RADJjGMQ8PqNSlsH878M
zOUgqaONyX8IJy8qx8BGRxR7EEu25Scp1Z8QOIA9eJyTpn0lclmkItZttduoLBybZkqp5pcyfrU4
MrMfnwXeedAzOfmPohqPh64PsiPnp1EoBIs1YuZLGwJokYW7cnGBdI4Lbuzyi730UfCteoVhJqjO
Re8vcjpZJg/ClFvr1SACl0a435g6QUr5mf1oCs/r1heAFmHodgvJJBkOypqvxLg7W+P5f4TSzFXR
9xzhpz+MJ1WFOpRoVOXCsTQS64eoxJGZG8R2EiXJKDfyO3PYVsFOoG1I3E0PL+ofCs6xQViLYRYj
DeIp+0wd62hbQVcODBPvkTCy5flQ+3xAWcVQyKBUYNIKFRami3sFI8ukDsWs/JuTe46/Q8T3nxcS
QETXO0Vb6vXA+AGZ2JzCO8cW+KT3vnPix9G0ljh0IihQGA7yzLMYGIdYFAJUD6FNv6jxT2qtC0dE
IwUgn19IbjWbKwvXhL2rsNwKgwsfvbchKWn5AB8rb0murR8AVdhvfFsD9fiYEBNPZq8ogXgZftEf
S+3yT3rfZyfSMUv34TlIGYZtau3fVOhxE9D9w7luLRQy9PZa2RL207SyNuu0Peq8NjB+ygGsmQgH
iBEh1P1GbQqggH238vLbbDujomUjnfBoFlBw22TcFN0sMm3noa4JrcykyY2MGnG/CILfFm0mtdzg
/8HXx/vwKfxOAu02SPn2iScsa2LjuYkA1Rwj/hYzLsofO5FBlSJJCBw0b/TPGJRF90rnMbc6BetZ
6Q/iEdCyHU4tIejQ500zL8AkTtz9/CVvB65aozv0aQ68n+gL3pHjvRuD2EOLrxzDM6JtG6cFkj3n
0jsblyf3tUC4FA0EArRbT3BmFzI/PpPGme8Dnh7JsQuc7XJOtY7g0Rp2SipTg6p/D290wvIgW0pZ
v1lYJAo3IWkwlcfYWefHkYnc40UFK9qh9oCQkJduN1vswnVUsnLr4WuZpX50uXpprJn0IBj1PEwp
DLNE18R0jCJrNHdj0Ax7kpX8POnUjgoGAjGW1C+aV7Zd22EuXdUd9QCeRUQZmP635DRqfbzZjLOH
GcAvjL+jlxe9hU9kHI1q8xDQYxKpe75SOUhNVIS3AAhG6UAfve+XItkbljMPqIrkB6aUxq84jtm/
ZggPbfD06s2kQ+PsUmuf5yoYEqeumeNJwKttSo/ZeRPNj4qeI7eZ2H6B3R17gbENsGZt5hejmpkv
T+eBuwBKS4Z3fm/WgFbjTZTq4qLMYmz8FYyPXKHDSUkoGKUmP1r6nZbYrcoTOqw7GPt9ZZip8WzB
EyC3US9o8N1YeSoCDGGMi0vsBHtnRxOSaXrjoFSMmEFIBk4yavjx5bZ4DjvwdN7ZesqaH85o6PtD
Cd7QmzsyadPYaicym8TOmu97a8+R//S64k4cs7RxOaMSMQfUZh/3yUTiaOxrx+3BkQecTvJnxGHy
6fHTUk4MAbVc1/aVysYmBJzBj9VCfjjwdm6NtlADCA/1PIH576B0Iw56SxqmoHCCCB7az+xlYKk9
Xew/IQdFCjkrhR2XQ6oHZNEETv6kkvuehcPhuSz9Yf0Ax9cBMOIKns6tX4RK9sae8yAhojUb3nSK
fv2tT1JYQ9sp93ZWKwAO4fnvrT5ImPRMYtPOyQuchIEFfH/M0ZpC3yxP6bAg1G1QuKTKnlO47xLl
X0gSmEYxkHG85YA9e/c/oIElBWq5qbXKpVHIIuBZVg9ebsVrFC8FToUvRQTL5A3y44FcF/Khjgo/
OTa/K4WevWoW0LG+yh3dOfYz6YKYGJyAT8q1vN1DGEXEwl6sHw/W07t89mTHBpqdyNWXy0Q0lhw6
ZSR3XYYCs57tl7zYbt6oiNAl+IJm5lPd6H+kImDsutcJZc/a46OAY4h8aox+hswGu40MRH1o0OjF
0GPlQSE7zKbJRxEHHtv+2AencxMXkbHCxkRitgg03v5AEY9lrywrSBCdW1kYveXoMUjPch0QhtLP
iiOAU5N05nTXNxlbw5iDs3DKf/xMIif0BO/RvApcOnSPf+GH+QG/r7A4FyzXxB9xxdVmb7PHEw5V
6TgXL1S39QvJSnNP9hG311aUiwWe5z0NZ9AyeP2zPvq4QFyUzhD2CrSutljt6gtUrXjz43/R4uzS
p8OiLe0jhOIpNMISNuxztOmPydYaa+2PbZ6Oqdsv/GXcoFtZTK2pq0eLYh1holm52sUwFhOjQlTN
X9i5nyDOlnq2FxjOZNsNc4L4kzD+5f5oUzi8SArTd83Yo35ea2JDo54sqEEDdlqjPjvr73+K/pyu
Owjbnn5yuyteanL8z4go7fl+LXIJIeV0/TNFzpmUWFiStmuf97wrqa2KvSFWQuMYrDI3PTIFrH1v
RagvVZqLxJUw8Qf7//gtSwa77LE42n3bldVkqqjPuoHBb4fL0FFgqaU+IxShJ4mT0AxcyJITu0uQ
r2thqYe/TAZ1BNksMIBhsHl5at6qk+4fN0IZQSZ3EmAx33/laPQ3Itu1XziD7XK6EpWFrvOsxbGF
IHZtMBt6dh4FVH6FBcCwDKqEyT6RqoPHtZjlbXvISgUls2zjotdHSNbI4gc1PgVwxfjfF/JKr4ai
yp7SgmELq97x/5zEdxTXbqocpKe8mEi68cuf8loWT8rlKdQZ7TnEuyiRZeid9P/PzqWgwHNa7ee1
rEjnMbazgtTPnaCGaLIzWMZ7o40GutmOSd3omjVPYcLmQhKNJ278318YFBNA+UOTtA0ipWV3CDtp
CUqcTaTTlbqyqDpN1dLeHKQJY7Y2H/Lakgxzsg8QvxLd846sRdHpJjR6hZCYSGRR29USUXS6hHtR
QKdt8ag+fH8M6jyxQlDiZAXbXD8fLJ6Ptdn5Yw2FIHULA63Kzi4sqLLWdgQ31IZfLmwPrhdVzCYr
rz7mABu1b77MhebaKYl9xuFblh6eh5wh1Or1eBOmbNBhDPkC8EKGbAUB+eiXRZ0cePuxrIOWCeop
y2LTKmge//EsoViraWYANZwjpB6sNpYZBCNjF9ftKL2VP/x7njaD6g+C5jzfcOkvTLdvHbCz+AFU
t/00TF7MVs4yPvrf7ogiX8AHxmOID4YOul+QEPFUVEzeInU3qAkMZNLYOyKLQlg+d8/+LXkCceNs
n1D0y/Y5GarS+TPLfRGbOad+Q1rUZRYTeG/ceZJLrnbI4kh4wTFfS36XW+mszn7M/WE66gN1i5Na
knLmdrWnyhTcFdzRLXI7fiJRPwojTvhZf84+P+QxJzEgAV8c8Sx/jijbk2cthdXePA/QvS/gGe/x
peJWrA+hHvzCPJCNXeP0hHUtjCeW0vvPlnRtWybcyKW6gqb8h9bx8v4mLYSKSFm+b9G0SmIczXtt
DTwV9JClmAk2ZLLkJs0UwITeCIHe133wpSwVjXceGT+2+QYjjRxpnkwV2AP18AnZtPLVqD6njOq2
BxWKDPY8soEMriK0bFYQsrCtVzCgxLP1w28gVApDkXSjhgw4TAWNaYjtaQ2DdFJIKr22d+2471qs
1pasF5chbur9KuMzqYPbpLiqII+VIYwbcjstga7mkP210MbPtpK7R/iPbDVsH9AU7ZM0Mu2OaQm/
+rTm5GwudexFc7iR5//L/rbhSuTt61EOhw9ZtMFbrSW8RxHxTtrIp0b0xOg9p47yRMfG32839kbL
raK+zJa0YZsBXTK+gSZC1xZrANUevRnrlzTYFOKLMtueklg2E5FZqsbH5+PhVRZR+522mIjH8ewN
oXwjJRE1UQoy20dh4JGyDLviETiA21C3hLXtpcOjQlpEaY8roIRSfT2p0KD+i7BxlYnVmeIib1Ii
qfIEKo3W+uCTNJqFSJeh+lVxzgAtAXepulFQzuEvOfNdq//8D7LGKapsRJqKNcXYhdzBc3RBz69Z
h99UJ4wSW/hsQRr1shUYD8+LAZhLNDEy6kqR+pNZoOvYLHVGMtI9SNOz8FiB8nqJGEiKX4XSi9LU
GEHvV1AivjYzsFMt6TdBIMAxqpg0uxsHfiI6d/PQL84yi8RxyaE85GrZ0aIF9lLrYiGPG96TKS1d
VW2bC4lb21Z50I442Lm7rtqIYbjd8KMkJSS3DhlDMaXiTp04L+fvNaqVNluEIhlgGRQwCosnz4kM
LjVSZHlI5jTMhg99Y8OoVw9cUUqaXc0nLpW61JGaSsLiKrP9Od73s13//5Sgl0CiHgbWXbkE320u
bf3hutx9H/7QINLyW0kHfSPCAQ9WA+ZkTvPms7BzP77CPVe2OaBIG02SrD5Ec3ES4xhng5IFVuUT
L2DkMr7TREEk1LzcFyNRMKf5XirqBLmuW0zNUC8X7LHjK/I/TjAbcYb30z/ZtdpFgKKnNUTvM8zN
/D+lmtvpXBt9/LltJ+/nfJE9Kci9Lghp4PCq/h7PJgbBEyoSkz1ACbcEupgbrS0YLSPLUnEtCrff
u0jIMoV0u78mb57sBd0cICfqJRJct5+omER4tHSv04sbUzHNP6Z+1RxJ/qSomzBu6X9YXG486QK3
iq0UGQcsQSW4ExMqd7aFbwH3pWleXFskLC2uiqTukBYJrU7RXEZvxDs+OytZdmDyzhiI6hWEjNKB
Sp5wCRtuEcTGlEpy3WH8EwRio3/HsnlUCgHLbMNvKUpuLKu/SpJIc3rt0f8u15BND1xXiSLqHjvy
6Tlcf2RwYYbHnt/WrpSywGeoIRNWw6RWLza8zgMaNMkAWiFju4tCsYj9/hGbPh4Q6rvbMHqFMxaR
lEv/4Ih44l9iN+jFXW6/gkZ3ALJZqwyMENoSsiet+9ToVAYNve3enUHIym1MzQ0MMa45qvB/ZyM1
CjV79TEKKFFk/0iFzk8IdaWELL9TZW77B6nfaXZ3QnotHpE2HlZhTnHV46ndTbd/8Lh+P16JqAqW
+iKUWB3gc2rC6FNfq/1NenIBw/V4OthBYO0Hb9Zv8yFhKPKYgoDIjqFOKUl90lEXuwBK85aLu/aY
Zn3z3v+YhjrK3cv37WfIDfSbj96htO8at75RBpzv2HNv7f3GL/pYGHv9177/hTNzgbr1VdBfgHc+
TiTBd1w+2nQpwmO9qzG1oEwvg4bMjO8IjajH99ahczck/jFRFArFZYFglPr4PkkKg1T0y8Kb4E1W
5kUs22ebfWzr0UBYERPAbcSOcrxbTlOzq66k78lSo5X0e9dQBp+31p7SskMWLuRqgTobcezAHvJO
3j8nGxxF2Y7c2aP/5lVkRBp96MCqvm1mm219C1RrNHNqvcxdpZdWGRN9M0ImQroquLjwRax5V9a+
vEI1D177g6CNdsxLk7ynPRMaxvu/231SZTzvbcj8hguRlZwN1RDRwF1scdbBb4u3/OtjO/OP44on
05qgqrSGBxkuVcTt+Z0U7zXHBPa7QITTG6LA93mhK1uBi+MPrXiK12puUk6v0gIDsL/g4u4zlw9A
TOu/5KXXDV0mlIRZbWD8J961rIULmVc01Z6gqp748AHN8abjT5PRzV87u4VlUj7dSDPGn5tY4Fak
tsjh6Pj+psoeMt5xqBHzVUPJhKPLhJQCcdAQ97el4wS4CRujEGem5XxxX58Afv5VecQ6bn3333az
r7E6z/MlW7CePUU9ypQjA92Z5buHKvGhDZNJNGM5zNVxslGCkGYswlh+rpZAcwxPWoiYgW/mC2xx
AIu0BCZiGbjI4CPiogvjCrknn4Xgr0pffCJaiSJ7dmksR2kkGGN0reM0nvfIWGaFHGjkWyIqi7We
msvIQLjm4cF7z4Unohfup5kizGh1pk5LJNw95GlbYAFWvMbF5DZkN1pbW5pJcU9r4287STQZShDa
ZCr/RB+agKnDJqsIdvFmQEaBQinCElkhFl350TVVeGBOFMiPVCdnXoQ2L3Cj8MW5rhvujtBvFVIp
hw67YckYpXHwsR/tKObTAYmfrvMMhNt2UbkMn6MijQ3KN8cUHghZcoLgnwXe7vJ/dJdAikkdFmRC
pmGpDsXVoWRHHVMExFIdQzh1lHKJ86WACChSVMYaCPuCSWioSIzR+3t7ZwHM59CQDsPEXrhVwSov
/JWVM9OYvFoX8+vpO+pfE2Uap/wu0xnYNwP7nhWn6Zzp2IKzcoQl8DkKI2NLrGgPjQ/DhZchxjOT
NQLFy5UW0Set+VY42MsjjuX2Kpy86BsTJpEAHXugOBEoQXIt9EbpFkM3+na1yRNOOTbLtIgPfmpR
XfpnI17trbuZMWfYkpzNSz7vzAzeLZ60KMXYJ9Qm3w0v3ga8EoHZPGkgNLDq36haGYIEL3SLiYLs
/kGbPRUGjxKuUmmruYRGs91We2yW0hZB49TPE8fDr+0D+UOncmKnQhzv6aseR6UEzAFJRALZoaac
stEOF+6Cra7C1EFQ3BBqPCeZSJQ7M0abAPSz4i6ld/GvW7NFMR6FfFCai9lU9ek7PCkCn3KOIUet
d4aUMTxgjcalm4wlsBtLMmeSdAH5xYCBx8bFRSpaY3PS4WFVx06Vphcdmo+WB4zw6lR4cCrGTkmB
N+fD9FwTUnDUjkIgLI7XhrXZB/nMAJvGZt2PWDod9tF9MGuHuHd/QFgpyTP1qNk6XgrDTzNjVF6y
dRhMkuEajb4Y3VPzcXS9cGZC7bGPNOGU4F1iJhbaS5DvzjjVzH6lTMT+SvJbcBowt/A8i1+LoczD
ItdnXvOxOyB36xms2z8LHs4FQ8licPGtWaVfQn4kFdeufpLWj3QIanuARMBJl4xItnTUPG5SZDsS
JWF43VXFnUYzRtdB4lPJBG2VEpApzogNstOetuw1qlZ8YKdhJsV4FQcb8FPLfgdQHoN302r2WKIt
3J9l0+W1PikIcjcIHtasTg4bnX/R0ANOX+BacTYlTexP4DOOgdvi/NBu2u0WOzOXnbkKWX7nJ0hF
bLSGfTn7UBQiUqA45f0B8DXYxBa7Mj0a4QWNDRFHaj1ksIoThE4JCEZbqWwpI21J5fnBCWzniSvm
OjPgvt3jEIyVLyVJ2kwLPTlMlNUIGKTLjVJhSCuc/Cpn/pWK+T6G8q7+as51v7FZULb8IRjxqtli
biS6c4Vb+FF/YyxkNmf0whJohHLTXkj7TTYqMAP03hff3d5TQbu38gpeyyHcR44/A7aAGKffx+Zs
694+XO18o1MTAroaJkR86q82XM66C4K0P7Dq6aHAv6GhkAJYU5v6AtlavJ7OHbetuTPkbRWEaWOl
DnY8H4KKYmQhHThiksSl+2MR4CpaJ9hKLBh28JKLqocxxZsNlFpnx9xi4S90wMjAcF50rPCiW6Zj
YAlzxfFd/hIgMedogoxjlZiNs9mM4tkvTSF1KWdiq4yu0xGLRmM+XuMLWH4FpzQPa4/fFzTnhKMV
68K2gaSFtcMVz/qJgcys1Qe05/fthPK/TGtcCUc2SeC3bEZYEnorSAliA05SE5ZyVep9YZ4J+H7c
uhHalC0hvAgfUXdBz0JrKJ6/Mwj1OYrkonv1f82u7oKz5ta4o3na5I0I/KRmBtm1X3jelT3djt6z
hGkiHIxzQEpGZVCuBTTV4IhDWaJnvxng1SMtfs1WHMHVBw7iWB9xOI8r5fdmrTSBuHE54K8RTr8T
DfzZbRfQm7CgcCf/oy9tGq7VsLyPxrbcMMQB1tvZBlHESPZQ+5Ldp+5c4EwtsIwe0ClwUFljE92n
ZSUXDRpy1G4lF/q3XSthnVGr62UIYZIAyuI1eKHbLCilG20puOhml4C5jVQpmvrb3z2DxMGd50gC
14BbghB3wG204dEZZO0ZjFMoNjjHiwEkkigDStNSKvlOtpCkWH1UVwcYMy4XeZabfZiEFGqnwzfZ
KZEMUNevH65ruB07LXUSF3JcworA7yXL60f+dT2dNo8AF7+C+eEhhfYEnx+2NjXDZOPapK8NIhXP
QkVxTKQrrZlOBff2uny3HPZtYpMs8HbwsCRIBhqvfKPbnhDXDHpe4fwuy7WYPE+S1qk886gyjsIF
i58nd0HSQAhxhmp+FIrCTgBGg+sQ814PKhQa7sg9AzsnYwwWge58WhzuTlAjji0x67fRTuFStGe8
76uftpjBWil+zf3L1Uzv4FLuOvv852TXKE5QlUDwz/46/c5WQBN0ddRoxffUdEE7G5ymjVMvSFAB
SKbZ/hlEHge4kRVohNw9v1rX/F5xIE+LePUInNo0YYQHx9Y7AeZpUrFb3g6C8wW304cDHe21KWvV
8+4TQBH1qcKkjE4z0gZdUrF9sCQTUuvh3XwXzK+F76oGLdgimU2FYe4U2jBSk+rwqSugK+eYYtmM
DG+BlLwf377Ky4C72v6ec7+ZxXrsI8KmbiBVuYVdlNFRtpVcjTvFOPROwNM3vu0ji/O8DGDXzyt7
Zodj0Rep+Lhtf3A/ygQ8e9yxgJAMGCQvABska9hfVUFxcZ5Q04NJRPp2GgklBwdvuvivnnC6s1G2
e94DH9TgN3dc/HT+R2OXuPGdmzrUAoVc6VuYnI6YrTIFctrNlMUWjaZCPRiWLnT8Vc7iXJAJQD8s
owS4rhBN+Caw0uPgy3A6UzBmXNRTZ8Uwc3CBatwZA8ZzWYJdODZw1ZBlrDta5ZLl27O5XCoclHJk
R6OAx6aW6hWoQOdX2CXjgnL9uHmhXuYVmJxoMKee1vL4vZqtOULuqX4CZIDhjBU3yAJNeBw5MQ74
+f/BGduQDX1RjZYgT4M+ogVsEcfCKE5vi4qGt5o8ipYXCf5FbvelCst+J2pG5UlRpDfmZ1DOXdkM
o73ZQU23mMZVqZT1wx3Rw4hNud6JY3yJQ9u2zeVy2m02HVqdB5cpdnEJ9c6JY2x99fBkYWYzqpg8
For5Xga5C8E223M9SxgV/tzRE+D/qmPa/61wKsE1HMl0Q32/qWg7lMVtcRD21ke6gnYHaRHJyIKM
ttswWm+iKtQlar5/6MZMzwxh80eJ++9PDIOvTLtpsIvuVb7N2bOQNshjsJC7XbXtOJOBoLYXwQO4
GMI7tQ/csexL/cHkjxq8JiE62ex9LK8wA/19n1e9cbiYr5LeaGzTSkTx0tuKoWKbRaFkcQGypTJ+
b3QXqzFFGSYQ840JqCDFIdn8N4zpdRr1C/KpC2K/FUEoCGYeP/q/JGDvjYpdvyzUcasXrp1g3jDG
l6f4Uo2UMgBQ7Nvf3kBaqtUhMhAbSIjhi6K4XrQdRTV1endo5WRNfzQz/xSS9vie4Mf2rWCCd5Lo
adz2Cs5sKmTvJNaE5xBakezAsQopwZaqGBaZwI7SUKaw66oWTLn0Djz0qNvU0w/bNHQPALibygD0
gB7uevDNHALUgWaQnYnGcKD1gNxp+GzyX6BXWkDqCPLMAkwrR6DIv9z5U9kDA8wgT1TptLqYA99O
/URg4dxpSACbEnnkf6mrjgCYkcv6/4b2cmbwXb7gaz9dTSKgcodp8fxp2sbvXsrro8/4G1qu5mJ4
6Kc7aMMU7R4hhFwK6zy92Gy2Uzb6Qv2i8wg9BygHievr3QbXPiRoV3NHzEs8oIACLz1lZTtOq20c
5avPdbXoYFd4D0Xjq2SBYAlyDB/wYayskTQflwoNP1BxfS7ny7WLd6Vb9ASDqmjQjg5WsIPo6KoK
Rbcwvvf27a7MDRZcga9G/gzVtg2K6Ewcaoae6uGTzrdwQqdf5So2kvA5/uWmOvxmyoms66/oZ3qf
5tPo9Khne9Rhwxi5aUIMF40VOZyiaETUtsDcvR7AZFkTrPkMUkDEXDnipYRGlDMsP0W8ilLxOQj6
nS4XquNe4T7dmv59CZvejl9xjqcswAAml6hxuMYGGMlK3ICiYe0CtqSg+3B/sHbPBG54wNSvtmhg
AgyiPESIerFG+fgaiSos0Xei3jvncNG3AZgI3OatmKmtO0gLpwJ3FxITguaYErxSJFGzE/0Qb/3D
sMj3+K3VSJG+vCIS8h6dItsFH9A71MRL+01YNT6pdGL1X+bd1ktmeQuli9TsH4Pm6REe0o4JwwZt
nDfrHHIrOyPwNCQZPUgnUxE89N7DmEH8Kej01s1F6HKJLUo9Y0uie5vgZF24RHvhsR335oRVCXDC
vOiv6OFAQ1hFd6Q5xUywZ/ObcOVCZoqJGcTZgvjfc0mgYjNmpKRyJ1iGXbwfa/sWe2qO4EKCSExV
w1C0VjWVGHkgUh1ddzq4Emmac8xtWyASaBGdz2enYeBHn9CU0EursfLNrwk+GtnFp02D2s+DcA0Z
3R/KzIkhg1nrKvFhUi1ylJOgiAbB12Bxz56Czxm9kvwJ20zPYhWbcpwtMfmoMrp7vXOtLpNcbh3N
InLoa5lW2pE8lj8ckQJHUf8D5o6MYOVcFB5JqXWH2F+Nbgl/9n/2z9LO6ucDUG7HvqYSMKyyRIhH
tTRVAdPqfgy3WIFFa9tBy0XNemS42jwHqPbMSvW0aoClJUpO2Vji1AJuY5CLp46sEEL4yzjlIEPS
H6L58XrDhg+KTHEkgRdvbiT6StZYi/oRqxFHlpM1FEC8ycsxUoNDFc4q7Hivk9fZu/LbaFd3GF+X
HnZySWfncf6fpgiMnv73T3SDZruIlu+KjUVvGrSi1a8UexAalijHzdFWkAMebhxllVGMUb4ZItu2
Qm22MvWgUaB0qkBFJ6KhBcoSmHj5jrscP8A9qdPp/5kz/Up267k+czrntelJCNFA+xBECgecItUo
Eusj2qc4ToMvcNXvBW+jqTK/Zu5fG7wl1vlVcEhN5ru32UE2/+yz+AA/CxkiWk2/2dvgPSaQ6Nul
na5fsK+bd4MecwNVAsWDGG0GqGIE+iaK2kBM225eZCbbNSjS+P+KLcmrbJpbR2kTI9JZv7wZXgUN
n4BwUjaCRObsYWaicYs71W+3RlFV+qxIjaA3kG9TPZNm/CT8Fda17Pkgrjanb1tzOFaPTEsRWlIY
VDEkBumgFhbWjt9Koal9+ze2Hegvtnxr5cVmRWEtjzouXNRoXIm8bzmcAjAVg4eUbQeJWQuxwSf9
rRv/oKWKZ2lzcvRcKVjkcXze7Hfae7g6BrRV9iNaUAW5g48QS+SVzktAFB/sS8KO3WujI6uXxgCv
Kw13CtOJg2J9ntKXhkf+hOXLyBRJ1tOCqckGKDhSAvXUoxBK89UI9QPnPdNcDCVEx7zeCrs0tJrI
n4IA1mzp+mZqvWxpC7IcbG949B+MF8e2lDvzsI2jZhLXO08UN7SpGoD9chEaLEPxcW6NV+BR1Ge3
qktkVGaCAjJousBOnu2/oRa6dnxgzAssodSGuQwuN2/jdpyLaYnmdSJT8DsZIeOFeldjDNj8ksP2
oWet3kUNjFqRfjXqC5qX7+NjQKIwK+TM9/rwqUzKDd5Bjd62lbIpnr1SA4nSmKsETJL5dzElVHLg
oH5suwx8torebLbM59scwOWSN/zjZoS8yq3Io3CyNi7c5bxMP88fvUdgfcw2edEGOk5hu6aJEbVl
6b0KTk1fGu8qdmZkxa97z9i8ITxc5UlHMBh9Oj9XdLQUqj5C2kvPMbRCBgTW3rUIpczSbrwmb1eR
GJTPgkWEX0vxJdmpepLSyeJIKwZcqyG8lugJpEUcCxMKuTxwEmlHguiMfhpGx2BC1sXL7E0314rL
L8nqHri9cH5wRi7K41z0uZ9sqnSJTygYBvCA2nOwy9oZiDDaFO43ju9IdNsx46NNjaKtoXP01ofJ
Anl8L8jxy6kZSTuiM4yyV+sKsW4X1fo40SwVsG1C3cpVYzHq86OTW2VpHjMlc+Fuoid8DTGhqJw5
DrXcIZetlgO61CNpfQ82M2xfCI1ay7/etwtYl/HRONaIkNupEk4GUmh22Xj+8urabKgCjiFtS5Ej
X271ws+EjBWv7MunMBFvlwhSvjw9UQGfhTJ8sZH9AeWgnGKcnXKY5vJMp7j4LPDEKxmV4PRLzRjt
z8kxWHKd00oIuZcowhf9bItq0vt7NuhjSVZEmKIg5YP75oikVDMtmBcDRDwKK6fipkI8dj9ABcml
UP3NnynL8Xvw1Sj9IYUdTvdyMe6FKs8SwZtxWYtlsMYKKLelHxMOE+hWRudUAMW1OAsa4RpMQPs5
o1FFLYJX2/sqgGiGUEQBwijmyeEbTfWV9x52O+YuZQFay5/oBXuDbx32CMhnPhu721AmY9Dc77ct
Pjn60SFUqKQN9tl8fCkGixbbz7kPErI80WL9vNmlNNo1UNYo9YIbo8V2vbB7VOZU3VYHeKrXON8W
NguaddYaC+3jrEsuva+kmO8D0q0t8Xc7OlnbZ4hmDdRbqvq2cOa2gkGbfpa82dOsYruOdj4eoAK9
d0ZaP0NKlAFy521C18UzV1g08s0Jr88ia2Y2gsGtzuPJbyq8Qnsa0cHQ7NtOEFIoY9qiF7DmmbQO
RBs5phdn3/KgxCtgArAJRyrL69E6yw0j9Psq+sC5RQeYmpLm4umG60ISEJxvjnGNU9fyDrNuZsCG
sRXlq+wb2WNRHeLmNhceSxeGFWbF1bY1hioFeh+dCFMnRy80onyEfCeBL55MiD/XGVUvJUp4vLlY
VVEfBHRjU+CCrXVaXPVf/d1CF2ROghjB+8937DfYkq/zFjvNyOdm7bHKM/XO7CNIN7iOPJoTJ7Vi
noaU9Rcy0Oj7liEX5X/MBruaYHxvmirv5HpE3EohxzcW3pNE3g6BLZXylf/JJmQo3sdpR2c9i671
3PqpsxDyNENvxwCbCkRkD1i2EbXJtL9aDa0CHxxl6QQIO8A+TWdixfkyTVXaBWfA+kgQbP6nm+Ta
p/DpLdkL8TPPcjyTOaEqCljzorsKZcfR2r0Bv/W7HMAuKOl+RsMpOHQLI3b1tecD0KSVUs7ADVi6
oZ7UIUaT8cKLeoYjoO3e+dQFFv1tf5PQvjSNP9PDfN/gPxg5JknhHCzC3a+NiljECEreZHMSfw3l
lTnjkHYno/YdDJKJVflm0IFCkxXGU7oaQK7bmKX+ZpgpzmrYPGDVtsDyr8bleozZ7umGxBjLUlTM
whB1gaWIv/qwj6a0kP6BIqTpeB5BTWVPWrCZgK35DFlJHyTNgCn4FH/lWnTYsDJTnUhsWATC3sEw
qqb2Z54RC2xUILwKalN9/wzo78yo0KjN4+Lg0XTTi2MXraXwV88Vd7Z1REEN60kYpYdxYtUJ7FMT
McCjbIpXFY/FVEuxc0mUTY3VLsp9QHePoh4jorGlKf/q+qAMdj5hh6fmw3ZA7VuR0FzwBoQtWNRh
iFvtmNwLpQvD2pyaYn4lk50lr/2CwF/mtn8cfTXq7nN1rssGFQv6L/tKw6VyO/fuMO7gkS9RwRUD
Evviv0R7jFWtDeCVPJdwnm/XuAHFBNFmooEclwnYp081xV3DPPALCL7LCMrC+AUcnPN9/P8bgt7k
ALEzlgOYoAVe4kGs3UiNk9AefEJW6LQPAfw+nIESG/7FVpAbY0H0KgMuI+wWMNvsHcx7JFnpmh/v
w+HQ4QO357Ih2XuJEcg0jMovdz/TbKJpHzbsK5c0RsqVXZ++g+eQUtXFRe1D0T3l5Q5uZ6CMYn/m
nYDbyxpStndGvIyoO+hMsGs1CTurE1ISjznh0h0Kwb9EHrHQcpcgA6GxrD5ED7+sqhEaG7a52UmS
zBz/GfS89dHWDbxMw02SQO6aad/CNIyuh1llk0PkgIErbO3K8aO8gJZFYDCWG4jg3W3tEq/asDU3
brLHfEP14j69aQZDsM//o95FUZg3RoUOh2yj+4ZM7AR1MOgm/HHq5E83vwK4A0KGL7U140iIHvzO
zctLTtrmdvkIuhNxq6z08do8fbq2G11nXGxyUPupOzfdssyyGIwGxXld6NuhJjdNcx8GXCXYNiwG
26fJND/ltkO8Fh5P7dPp7lteYN1tNHDhXFGfuUtL2hNajSTgZMcWUPgdvnZcQnEoGXtO1VYK6rvv
4cqpWSPuix6T7r+iaDFVK1qOKL92sLiuo0iec4f/e+WLO1fFuJDm3GAzemf0wU9lMGwWpebKRxk/
VfkveZphI1maU9F4C8jgIToplh7dwIqrABLBi1D8MCDy8BXP2gTorcAsSTJ+2V0IeaRsICQwvsiL
EOrFrS+m5fY3b/lBrkyMPV4Nmd0h5sCH65Ruosb3Yf6v37H6qgVhdQA1ATbJSFBKOgMZQTe9ZsI0
JMNsReo5Y1GfppVxwXCKpEL0mV7D6qli1LJe468WyGzXvd3aUOWbIaknNR1STXtzpTjgVVQCJ6Pz
2i/4sNUR35igiZDSkFiED3fvQ02Cb1tII3xhl6lfTbvMWhDQ+T/PRCB+J3IcqqMzjedzK/nKUuL0
4GC7fHvzoKSyclX38G6qN0tBLTz8cAmD79D3HaUiTfAZII93dKsUG11081txcl5JHcCZwN3m/6u9
zkifYQPsqEldA9l2T0H71u5YOnN58/Sdg3fXdi8gAbzsbsJ8m3WHcuL0cdH4uItjN6FWaWFb/N2r
UbKvPN74d5wRdNjoJ0WEKPsSVz8uQD98B3/YeGGccY9R1ILqLL1oJMFI0RN50tCpKwNbfWv1N8+x
zOALDllypyd0aPnMW8pKKQ/9XpPf++NjLc1BhswoiqT3F+XXDG8CE5wFld/3t6p+2uMBhAzoiPWC
XeZo+B+mV1LQu4c2GYPYC58HqTr118HzwL+hwmVvrxsujf6nL2bI6kLlEZ4an5QMKNcYoV45pUE8
q9clxDQywDmnLeX1vEZSyBQz0kFXwyZPXf4Jh3hyh02hLxWUEecTGLkp+S2JlPTyjegv2vrSAwG/
wY/pWlmQ38DXJZHgv3udojKoHqnj33Lsiq1dthnVtrejuxPLXpMqL0i5IxWyyAvmWPp/mH03vQlg
J0aoAZ/nVM1hvFNt1aYWkTEtKRiP0Dum9lJRt2mTT/Nl+3a6RIk+7RLNRft7Z71/akkS9/lYNsFc
YY3mxPvJiv5ovyZ+01PIW3ibOG5tzwHErFajlpe736STooxicPxhH3uiBZHdp1isVa1dBATA6FtF
1cgDXvf7DH2PSBazYShT7KckZpImZ+GQ3/8R5KTbJnR3aTUR39knWJylNjgDd/3NdBX3xvZCoR9c
wjVzuQhP8kcyDbjALzMRpzJsKl1sTXLgdewCSHK8pdbMftTsmgY6nrDTelBi03WhLjER+HC2bkm3
P2/iThicGgQGlUlZLo/9xcN6z90v1tLlR6RDdJaSp826oso2y9rwOKQiqaKf/01S/pUR9YDzTVTf
MeOwhnLvUoYx52E3Uvp8SD38hTyr4JWFYbi4x5KEY4MegD9X+/DfRl3W+MhKMpS3aN5EE92pdWC6
ASD5qyDueQ7MahF0F49CvXX8k+5dPd+QygVQDs7W0CvPvzjphKSNggMnnfF5702owuyhUMdIWERY
xc0d9E7b+oMI5PVOjOwzzcAX2G8+9MvG4Nqohyw8an8s3S7bTAX8uM0FJemvVLY3HXbmJReCTQ1m
UBswtLMtks/sWATfM8iUYPPD3XBWb646QNjP9ojDNTa11SA0O44AxnjNeX/SwCv/spGDx4J5p7rh
L8LjDuZI1pyLNFLNzlmkK6fwdYOn2XsvgmyWuza9WImME0ahEJmk6mi0Am/z0x3ueiBzKDwjfum7
DvcTFHtM9My5wruCCJwIQSRBKRhUpYLfowShvQHxsBRNQeQ8f2EmRvPGpc+vckwDY1Q2jp2hsBFY
6+FRSEMKTdWDvqTZpuTK/nAJpICQECmvH86qmB16FrH5iVWPiW1/dNeHmNKvmBZcmvu3pFe/NZEp
vsHXn/erS8g1gHFahucN+joGpvn5OCsD/DCCGx96bY/R8I01zD9rXXlX11oIQ0S4tq9f/1iCBy5K
G2/aWydNNS143LM7ZjalTW4+WYYntF0jbAzBz+asOk8Ms/AX40VCex711ktx4Gu/PfpEIhlWnm7M
iB8kIgoW0Cq+ZH0kdQgtzYETfH3K4FcouyMiL9+8MFSxNbTblfYhE6wO6OCQSpdRl0h7htfyrom/
8F0RLftmEfNXm3snWBz3Vh2WkA41YEVd1dgRPk6MLBDdBfNIi4U4qJ0xY0TJ3xBg4QRiWnO+5p3r
lmGKpw15tQcAPCzhFBPRrTlwFDT96vtIz/gt+GFqgTW0SS6WsGreJAcv6llnkIPmtmOY5nZTBipj
QZMcClCXFjlupRJy8GHiRN3CZeb1iXw6rvTyukhIY7GmVhQPlVndHAW12Yt3laKoUmzPgMTewY+z
S6m8sbIpvtIuUIn2wOpqCz/Ff3nwiqZB4aKcQ6cxAuRoVTXOwJpmihJyf4Pcdoo6dlH4brsN651O
aDngM3sJ/7gE7KC+j0QDirWPkdZ2hBbL0csBbPW227ZzAYuCBWTr74G1ttQUoSrsp2VKm7z9izMU
iyqNS3skSj7sB1piqCBrI3l3H7J90uasEBTaLQk8S3P8IvgS+pjqY+w8RxXbPvFIqRBwl7bgQmPo
JEfxf8JCosE4jL6N78TFaF7rei6K4GriJnMJ50IIIh3OVgalGe07hXJUckW2MqP1uvAMo/xBXmOd
MxL+h/BmzxGfAwOimlYsphcs4hXtPYmhn8jy1wfIJSRnvFyl8Xv5w9Dnd7itQazMNz5f9YayZNcf
32mfd4MhzwdpptoEY1nsWcupQo2dVZb+5JZEgMvmpYOe81/B15XVHiCz8wEudLPLCXXQZ8/kfDuB
obkP/E1YwTlJ9Q7IfriHHe8/eg+MMuQz7TXL7d+vc/OINdw9DIisRW011TSwdCUbtagNggv0up2X
YG389yLoSnEA+V4Jv6QRHeQx9sOeaX3p9FLVWDntXYB8BxOOVCSobUXD+0qf2pCXmOspCWIkBm6b
oV74IhXilt6lxG3U4MBXJu19cz65jcNd+Xt2ijJC3EHU7U2eea2jjH3rx8BvLhjZPXYSBmOLATLO
T7MHEkf+o1SkWD25ThzEsUZ3T1KLMQlEZaRAToOzLWpkB8AU58kiZTiEVOw+RmE5Fmx5kQVx4M9I
Akd1b9lq/eMmO11tbWfYUdZfbDVhK5wX8pjVJYxA9FMe9OWcXwQeYGqKrvXGpN8oFLAhVJRiucMS
y6ylWPWu1cgUs9+X7zo3dvbOGgaBvHyDu4c5MmddaM5AF0MF776AvFt9LCo+/BXBnjbMfAwEKgsx
ZHC8B214conZTYkRLZsdQIUtWj1yDP1nwdjaZMnS+WPx7K+0my9KLSsWdEA81r7cV1XjsmqDC44R
Jw5Qe0os9mwB2EcfRRatQggEgF5vD3H9huHDcEuQmxHr2QOluOiHOLu2uijt/6UQjCvOzAiUbIE+
B9W5UmDRAqFtSPieX7DeAaaM11xTlMEFMWjo5IB6fMXMvUFjqIZuSRk5hZFN6qrWsIs52IEm4QwU
Sr07Qg60wGzSK34bpmbz6j/ME3rAF0oIeIR3P/4M9EYUrEB5P4yBiRCMHn3XVkz+ftCYhCJxasdq
omm5JfYBHOb6Sn42U9FydmvKD06ZgL4DbcjCGWsUNjx7MI3azeKJj/dip3CPZtU/G1I/r8j7HtkP
Q0oprileC66X8nkP9ec6YPXQlthu/0QwhOanuO007ly2Cb8jeQDfLUg3lmEczNoGEcmE4VjXaPFU
gJBi2+uRVwO0JzGNpJ/5CNQAVK65tkF/cUaCEAKxQZd9IlMTLNfy4yeAdV1ELq0IHbA5nLK1aSW6
dprEBJ+jH6GLOPcc7aDrUwCzslIXDGGCeAPiif7WvRhzHK6wOSL0Pu8KnCCaTR0U43os3CC2fG5K
Gl04D3g0/sr/hbPNl1/4/rrpSLSM6wEp5KDKyLKRpPCIXm0p7xVLml0DaTniKdbMxvK59yBHFzS+
rSlBngZ2fqVec/UJUXXIeJtTDVEbBjk/1q3UuT3NtitGr38c55ZAuqJuf60P1pI4o/kHBE4YcWhS
nDmE+PZS9dXoLxn2qj7gN5atn66ljTpkTPEK2AV0aroU+qacsTw4Ycn00akd4Sc/O3Ud4IoVfEHU
Q77eo7ImxpYN4F2i2tbc4Fallqp/meeMewd5+41p7O4w++ZmaGyF7BaYx0WR3paN7CkO15ijYnEX
qN/C2ZIUAxJCOBiQLXHzacxbeXcLuDWuh1saWnlgmtYpGmddon7Dn1zyS5iMZAPNywed0mXY6wrE
y7wIH6jkgnG7wjBKAwH8RJoAHkFz5dcyy/s03FGMsW+FOppOAwpCv1HW5z5aKv8cr5MRZgMQiSxu
HjBKRGZba1zF9j4NvNvKdVDcDQTMzn42GDpDHCB9IaN8C7RhMs9797iy+OiC3AZ1EG+ql1CO1UKK
mX2RK4w/rvp+dRaemk2+yd8rNV7CAMu9cIct9SvEjrcflnGy7/VVGiBD7PeBb2yXdmHIUGgDlpEB
ovwkaeeVdHJd+gBgVnf5Dg/3VNpJ28HtmW7BpBEwZNn3OZ4oRrb0Mwy7OH4DMW2zSDBisjY8zpNl
TxxPvUv/9gxnIQujfnU35GfELB+BwhbgviPV2XB6ZeNDYGoFXNCho35Vzh85UyD1UzcXDEep11zq
rthyYGm1WL354p5O2u4dz/Ew5SoAmRxZl75s2v6EmWuFBhltjT+M7pyTcyHhUBzDw4qVe8RG/K2h
StiuHQkP+UCqn1Qqx31UslsqhVYMLtd5dbGP8vRUziqUwcpbCTZwUd9WAPS6FU8b8eB/Z3StghQf
52vo7xgL4LZ6VH9fhz/Eck8B+n0BsVby4m1jSIlTdmhNoJUWngd+JE3WuobqbnkQEokppQCN7Ifw
KF0w9G4KXIOctLVoYPmWKAYphOyrh3tITwz1vSNyxmKHaaiRwjMrCAD462mv5XDdPneGfjkj/TRn
1Qq+CllJXUyEYez1+vGMwvJGSC0xHXPiilTe9mQFFnxOd6rmMU3LUHDliRLMs1I4RYFipEhT3xzd
Bq84oWbQCJiDizC70EX8kApQt2nfcyA2KSYPLqumKAa4fK526lb/YZGpG16gxP0fKFV/0e6EvYIa
EBFHFE/WhakBmspJBLOarqieTnidy3I/sLY3OSzZCHIbkyKPVdURfCd+acXs+4HBy5nuIQyvpHKU
tKymLktGL4l7GAF5mubHgGMqr48/DVcxE1dgs5YaZuYpAyX+Ic8gMgPvXsuKbTHWZYqVU6+iOHA3
RceGjEKDA6RZMRHlquln85MspHqKqIysxwlETgxSLAbT7Lg941HsTvBSLsFee6EaQ+C8vmOHnll3
Q24kHC3Xp/OWhihc47v9CdyER9NXrf8XAwiJdB8bXlr+HSCUm5OoCMvS140Tn6LZX0XILcEy0doj
FaYthmMRKNc/KCXsQabHeB1GoMxt+L+pSVFXtEGJN2pLeVWrNlYfpKTczXGneT5/mpB2FQPp1klC
yNZHI9ajRMpH2I+F4wuSGv0FWeOX8tGPH2745gUxVCPsNLFP3afgTUs8Zx2dNBlwfPkEOhj4c8jc
HruH6ZW21UXK9TjabM/o+WSRzdgUvCI/EAD+Ir2SQxRx5nmIo354ojVDmRzlj/c4mFbZ4lLrrXbW
GetCbv5Ukn0YmDTqhjd0QO/5s99EqjO82AL+JmsfOqR2yIVsYJSiEYVpnWnCeaDu6MDVRov+s7Wq
ALNnkhJLWz8vJbNVvO2LH8ohe+q/oiXC//ep6meOyr50AIRpqtnje1CiJOR1cr89zl0UHFn6dzEx
cnIwSlQTqF/Ql2Mr+tr1KhzXE0wsvtlQCfu/H+BO0r3bcHEO+q9XSwBw+n/CBW0Aj8v6VdqTAjNa
Xy7Q5q2I6koiOA4FVGS570REI6k0agQysHlfOJyKXBVTjmfHU10S+whmJQKznj59i4Qz4Ebv548d
hhDQzN8jL1zWnmF5R/LkfECPF4okxb8nIixSWyizunX2qiwcOnts3nA6YQE2paQK5OyebF1mulY1
WucwoUWaX7aEJuvJWqMp3BNlNhGbwwtbYHxcLiPltOcSZjVmB5KhKiq+iaGIPiC617CZB1VzkvWe
rT0RZ2mY4ZiObgPbGJaWtApcKbaIBSkHRsLc9X5IsIO4M8Z93w41ZrNbx2rf0w7fFWIPCreAjWq5
iEYGYn9xTvIFGkn7wpoADh9961PdZYu9ueQTkcKIK/2CmI6JT28VXjfPoxChxo4qTbOgZXGOvozZ
zOPFiDek+v1Z233Hd3kQ2LSPWIDv4EZGV2be4XOlT2k6vVCegnPOEDt3k81BJJ7BIE1hpJVC10An
uy2eykanoibE2WrRf4JJrVxC7mjNBrgOnwk1mnEtbV16yKkMN0ZHSiBhJBPVIzz58f0sfGclfazv
5mVus5/p/Tk6lQl0gZvczgjLo/OVocjDMDAsUi1Z2XvPNNkWxC2OUDAzAjslZptiDDe7H2nzwYU6
5w1Ynp+4u5Md462k4Tx2KxGSk7HXg57m6U1OMhULpnPCtdsYBi4O1fUZ/JltjPTa1yRlfXJ+8xTR
z+awn9GuVSupBZ1LmRlzm+9kb1QYdA6hTd8INhdQXLrbuUD6ymbtANyITZdlqFq1do+Y77o5MrTd
mXXifz6wgf9ieq7m6oWiG24IQedYYBGauB9tPn/+bGiU3QW/2kQntHibLjUuJ39U41Qr2HJQszLJ
0n3EbqGrqR0dP4xK0O6+iZFsp/bwzVmxg+A02KE2clKH6hfL9t0c8k30BuOYFMLE8eHXpTj2cY7Q
r6iF5kg0O4xKSGwLt2rx/c5vVCgBWxFg62KVL/WY1kM1cidA0mbgEQABKKEsTNa8EaaESUR+6Zm+
HGuabBg5z1lOM6hxFLH4hwV60Rp2khNrcn/qvi//CKkneCJb8McL0StHQVITwCTmN8mFQnHcbzne
ZJKxp6sXHZvOHtagIWI4MVIuMyROG+9oHI9T7iYTOO39CtSVaJ5mGCqEyhN9rg89PU4PuOKgmXwm
OwGhdUNaeVEDOKFm0acvLbCbfffTVoazFdQOTRwES1a5PFMDGkSI/Jsyp6v13WBzgLUgn4znEufi
vv3YK7QmrWTzkhkwG4HWPxn/JpQoPAGs4Nxgv8lyVhwPidToTbFyr8wCiYlbKCjbhrei3lGH7IVc
XbT6Cpd5gZ6bFBsECdcfAadMP5O1hBU+JJ+8/bB089cnN4IcGVICkYIKvg5uBjyD97ZzY+qq1wXd
XjFAbwKFZix9G2Z/o/wdWkB2miiGS2Fz8xYX8KB9fGRN6ZXEWqPg/bgD5CeMFObetDRjRK6S+kbZ
dpMMfnIgyHeof2UdjGJw+L8b/0MjEGIqYPEREDFIacw4ZC+MK3W7WSoWOzqCTzQsc66/gFtlGmx0
gFzwa9ubY2kmM1SHBSSA1xN1e4y9vsUPCSk+5Zhjr0mpRHoanY5sfHpo6kamDYeOzSn+1uquEw2L
tiXrYg4mXQJUXCiYXI0nB/779J/dwdTp6mvfB7z///2e4Mt0+OO4tD7U9na1X6BDoiPX+E7l+Jt6
xWazMCiqgF5CWqhc4g1ZCJTHXHAZQiGWfDSPlrW+G+AkDffEXMuIwXRzCQRDOfiJ0O7XxD4DIJaG
7mFijGKdhd9BuiukC4YNMksbIpLz5oeS0wB3CTOUxhH8FNOAi2AStMVQgSLExLFuj06f9uPhWbOb
F0zWvO4nnScfTaj+ja4xQ1mFaSm4r7q/WU6hGo4iZhsdpu+m964SYg+QZZw3Wp47VHlcPfb1f+q3
5ZOUhmT8J6oAeeQZwJcRFQyXsOG0DLwzKDsmjMmYD9roBmNxsIJeMy8s97clJVGNEpXfLahaDuBE
/u40j4/YxNljnXWbtmTYY8X01LUxdL17p5Nu6GU2L662aacXZ8Vx4S09i8FMbWM1EEwCLyZfFsce
dYs7skoD4C6sJCmU7zj8xB8X6A213PB27VNekfSK2AVDViOJ4Ry9k/Lnbfwa+N2RwRddFp3c43fu
B6Zx01U1Sej4FVIi/yAqfFfmWRGEPQ1yBftsnMxQyZtE0a8ANYF+oUlVIOQPCPR2u/F/s0oBev/K
kNZWmvtuAAgQt26d/BcxySSIMJ8Sc5NRG6OrFOXhA2WSWhTBeHRWG8fWVacwk18s00GOABnhn7HP
Z5603bkyR0WMvKm8VY+Br2K2uV/Qr3ddIRFaJS6CMXj4gsKiD9uHrhSSINhDLF/72oLEdHc/7f61
ulpgPJDDJGcIZw5Ii2rABIrA8Tydp65QDKDuJUewAO9F+eSbioVJvZ7RPbzM3YUu5vEUL+xzehqO
dYti6RhyrOvXOKz7U4FmfGYDZ5xCcV0OOq/F/tp9szIM0xS0FW7/OximnlEiEY2OjdnJ5E0nQbPQ
ccOHZXOaa6U7D/ZbPoQZr4vQIIgIx4Lhsxt8l69Ik3FyQRtwjf468HOM3yQm4ZVaY11vVFOzYnRA
pR60ZrTUWXQcfQt0Bks/xphQabV2QhstPMrUOJvkpFCrfp00q9byaDhINaLIldVqfAfYZnEb/Eyj
+Ypss+GGHAqJcCduDoNVfoUK3FYQc5IqF1EKLeVGIu2QcSdARp9d7efs9AV0Urz7bttQLca93UpV
Uv04VDobWMCyUuZTQ8nfQcy6QQEUsRoIg8k9eyKkB3YRfPClPIk7hMOw+Km/Nd4hsayMWklpSVKe
SrIgZ654fMv7pvAvTC4NqngG6hPltno+jr7CtMFElxn6MbWtWTJVyN+prHRTn0l61qXxRI/FBbxA
Pq1oCqGhNopAUjBgGIVhwoNGtRBE7fntnSizTEXi375GG6hPvxV8BC3l3y1AoUfI7wOi9oGN1+N8
4w6GkrBHh1tROX4ub7QyHpjoBGAZU8YXrQJEdR0ijm7Bi/NaFMqzdvB/2+8syVpW/SDBf5czLKh9
NCHWNGXuADw+6OAfUzApa+4S0HHKCpUCpRnQzk6cW+hwMeLooUe7LhApmbUu+BbC63twNdjgVrO7
HhToJVw4ewSQ1ga7WyD63cD3LrVB8rNC3b0h7uNteycFMjwSd3nGTbk4hKRgDwqoWfjGOku7hjnE
r6Kd9mCcJreDkZJ7A9GxS8iPbn8HwWN6VQsEOQWaWyeXaEsxXwlfLHAL/qv9iKJ9KnTcmtrJ/NjX
rjEzuHgPdW/NTh5p6oKOTyc2qrRSE+fVmE7sOl2pJscdAq/y5sm/TlfKn0feg7gJb72GzfVQ/G/k
zjsR2pMLrMwpC1BCvYZVoDj6+CSMF/qH4ntpKr9Y1NdMa1Lwe7d/kfsVOG5+SbIO9YWNh+bntV80
92HLXPTI0Hc36T5Q4m93ft6zYs/IM5fRA68zW2+aJtWhDdBfxxSfzIKAlxDWMnVtRyhYcMaJlfSs
kSKphDfyNFshXH+9eUAzar/G8drt0hJnQWAv5luQUR9ve8GfYQldyQv64qJwqXkjeTMEI2wpz9MH
p1Cwd5NZcG7yYEPRKPuEkek1xFFbm7LbXQ2USoldcbodlwZ503k4PiCgCZN1H6amAe2a0IGVHYLT
pg7bn99QqvV/Ic9o0Q/cfllp82Jx/zreJFTsw7F5Hk23HQDYBV60viaM8x1gEXCRsZpYjNeFLN4c
xnjTQ8Rus7bWW6462gt2I9nrMg+jBBeZ71aiivrv+WpJM2fUTuyfo4WNzHnprD6/QXMx+4JB3IHw
g3Tj1eAyrTQrqyUk1POaNLYjrI5rwvviiJUcvCsm00kO7ABaLHZCRJNw9YQtuLHZB4Q6NyedNCBH
UkFYUTRgAEnyExo2FD4oAiUhIRkJN4RNens3JmeM7vnBuQifbQbVS3GRjwUsVczVVLt3Az+C6iZZ
R5gfTI4PcUX56clUrc+rnii9x97eELijsuEhDCaS5+kKzSEHWjDr1cSx1354VAR/GTcXloZRCx5o
u6xeClguFq2JxzkXGjqwM6G4hHJHn2XubIKrCc2nbwzOr5Xg6C3FOvYTVcPvp75Y9PZUWFFha7Ak
5eeMJiYNJwYdsC6ZEkU98i9DExVMA9bZq+s0QCceSK4ci1Hj/CEpzr8htAihDCD84WWCGekUWDx0
d+ClrW26DV2NIXlOK9/KkrERze2QRUcvb+2mN6mWogvK/pIlAT9i/jStx/NRJb4s5qNvC+GLDbUM
KOiO/IndVOarl3kq5dxsPUduO95znuG1TYteD4NVAeiyPbgq+mZB8IwGgU+QdP3GwMEneqgahx5g
J2Ba+k3A7mmEOGFc3l/H8MYQJtpEaiABKg8ve0A86k5xPBnzthV48oF1u3WcFAfck+S4TCjYfq06
MnXx0THec1+uDLBem1IlFs21sHqKqUEasxFVm/pq1y/QasWvapO4Y2rCtOhHziSnweKEzJy/hNcF
e2KuT3AA2ouykPHCgwrw51ACWxWO7nPfy6PohCJaoZTifa0o3vbjPoZUKduNpn7WsajYssT+0ybE
oMyj59bHD7DXhH/FD3eDX77xLlmB+7bPjvYmMz423kZ8eIEKlqy5yLB7Rq8sy1p44Em1vXhao7JQ
o5BCxXGv/Gnrya5RSNitl6pcBMQ71j66qJbh7jpkMORsh5gd1f0ivQC/KfjNhGKKgeParesrSfGW
lP3NJ38zJbaPn42gVqY1bWJsBNFC0ZwQ4sw1lfflDTPBA5GhW8sUFhWVQQ3wzKLwALrfVc8iIomf
1ZpTrl8l/kTeU9Wk4pajq48JNBHpJUw3cH4lAV+HCxLrQv9oBtenSan5ScbS/kDxzX3xhz5/IgM8
ixB804pXSC7BoPo4i/0HNDEC8OTyM6rLQUFOFnB68l7CoZsfYWINePzOOKktFtQcoXDvL77Cti2V
bcGUpf3K9MU5Jzl8eXmMqUMJGnorOAqHdY7965om394YsmU1L9WVVhR5ZEj1SO+hHjsiSAAa0eRE
pDwlj7ixaOI/tLPqj8kYbfr2fvpZub8C0A6XnH99cvg7aWei/cawrh2orTUDGAnc8HRTCT9pfVSW
cNTaL/9NM1t4Ne1t8xpqSQB5dvRUJ8/yZ2CS68SUal+GJi2H0lzqTRshXmnr3Th4Lhe5IzCS0pxx
7XmmuL66IKOkRQkUmbc3+DKolt1cmOKA+r/vxj/hdyUjq0H5DmE4uhf24mGjdVCUS+XsSEWvcX8O
yYiA1/sesDccFtdQdUfqAMyHViU6t8SO9fjKjN4tCmWjbCVgt9N0VzXNMHb3ZATI3lKygaUwPpf0
YAy/gjjHfmuU+Udpq/mAlVEfMSAL4rTdtEb/Fsfo+ep63/n0Q/gs3vwMWk+uuOfxxoKgWBcgtP1A
Ddc4mHQ8EHaBIhnKATUWD2YTJDibwF+Gm6aKXdJTdKP2RVnqmLg+0hTXFpkw73tBgrulF3RQmFgy
YWc9oYzN4+5uQMZMMzU7zme2+DUpC2lb7TGTRNGW5vJuEIJrlhkC/PETcK/14PDDk/IGvkYeD9f9
BHhMPKgLuYmufAb/Tnmho2SLiBCvVCsqwLIg6Q25XbelER7Xdwv2CN8s6HLUqJJsD+KecPbkMWeR
Kz6D/icA5B5zi8nUj/nUslCr2tVn3VriSqOEVqeQt82NeA95eIqfgtyF7d5/4WvlraeHxpqFQiKc
eBySTq6wXne6Ritt2NO8e0Jn3RLKdqk9D2mW7rEv9wGUDIXx8umHXQf6lYgPvh9aPHVsboIyZlkO
/Fc9b2PqumuvjKoLhRM0yJKfPTcu8qwW8xK3vXUehFCfVfy1zqCH5+i7Ae3PkXNayZKdqH+KVG30
jAVh2GrARpMmS6odSSBwNR0QkLsEfM6vlaTAVVe0d6oI+IITye/9ivF2bRWMEz2TrEy7PBS4A4nE
nDtZwh6QdcrxvVUUPswofwAhpG6LxnUjwn27SGumW9A1OfSVwa9k3AIbNR211I0e886s/9UXBEnK
XcxN7y7ipPLZJSCSlDkFsxKoq2fgFxxrmSD3VXkzCeRjAqm0dogOOXJc8dDgQ7SjAMEDJzxVxUlU
5y4RegLYd7aqj7ooMoncy3wcvUj24FczKfcU4WvT//OvjWOfNo1Q03Uk/a/eE4RQ3S1MQndfw3N/
eVv5hH1wr+hLyMRdUPSIXJ91qkb3qYeVQ3BJRpjNu8VaFSWuqdAZnx4a9UA1tG12NNi0xWiIhTtI
6yvEzIklnTMPeOPp9DSJl02nWJBoUuibQSq2rF68Q/J2YVtkyatWl7oK6A3mAM4arxGoM0fiP4Eb
FL0fgdT66CoJEhWvZu2U8F+MadkxHtK5Kt5vFntIPaydrrbpWPtEDElhMVcUpjAgfWqRofCYtvjY
WqTu7YqUyBPtyLHTUbKqpSG1Q5hx38eDnuA/gL8QzdkQWLQwEXB1RKM7K8dbvNQtVLmS7tBn+s8A
stLyesG8jKdNtAOXOQepeVjoG0Fz0NwalMu8EN4AZAJsc4Ug6oYwgjasnRHGNQs/UPd13rfqpq+2
2ambfhJElTSsj1/IMy78v2ZvTKoV06/V40uXql9lPnmLKrqC/SMJMCs4bWeZxSl0/P97KSBNoDKb
nGfUnLCklqUp8FwYm5k/pBNgTHimy4v5PBR9t422Ohbkxw+qCfu60fp14AHPdtFIbGdAcSUaiyq3
RXdQQDlqw46H09LFhAeWd0pCe/EigYFYQgYkTXAVl9AaL9NTHRA82qZgkYuL+zYC4RVVyL61gy7L
dNMSkOq51E7O2uCW7XYS5T15iR2B0H2pEJTgSGB0W8VkSr28PeQ972uioKrRYeYKjCVQx/dZMarO
otX2qSxXQMDxYiASDWJaTANsMjO2bXlrslLzbGfvv8te0cbxbi4Mkk6TbGhZ+r0z9ME0LAIWaMck
G3/Nmxv6etXkLpBWmPQmQeeTZ43FQlNuFDxiwLdBViXbvbrqPrbRMaOi45lk9vGmRP5+OQil8TzW
HCIsDQ6CBDA9ssSxJPwSB0AIhXYg68FHW8xaZueqSLOBGbdAtLoA/VrW6FWinJZAGDFi6LlY3FI1
Rol40DorvTERT/YhIWnDwVQ+/TFHurWNccrKMgqL5L3N2b0kEyvTIWTR6Jn9IxTr4+ljgntPUutD
kDASmmD8HgOnlZakHDuhMsHX0VLw0fRMnwgHZGRegT2+b7/50HPXo2oWdeTgNhmNiooZnqMqALwF
fLo6x0B+2QYVgpQcjtyc0Ww7bHrVgF6Vl1Qxn+ZRonOSUtkas3YKFVmdGT8ayQtOuzBWkvh2/o/n
H03Iir8qg5V9D5m8DTZbLjLsG/7XsOf/tYMWTmzvjhmAJTwSaP0NcxAvWsJS1PK0lob3DZ1FvRBM
w8GfGGId3S3F3uX2bpKIbmdtASkw2H29wHCWDiNmXJd5BJWC1MFTmXuCNxfKa0s0jsDvT9XGx+79
HCS1jmWj1D8BayiGvLiXU5aNFQhmv5c7h+/dOv9W/CP9wv+xOHx9Yvqvo9gDbZwnf0n9yU2/OhHu
zJcBmitAJR09Ot3+Wot+iQAN8rI2v3aDoazKIzmOyFaqns9QOvMA8sq7C93FvPNTESHWC3gn8F4K
ZRZZU74+9ZL1VuzVhegRCqREGzwvRVRXRQ9Xv6at3C9SJbo3GXXSVtaDdqrLg2JOxPzQZMYGqMFP
wKh0EpybYeiU4gQ+GEGR5LZZYaPTpxmqmXCAcdxJK9v/23CHwYOrwUHd/kj3odPG3b4z4w5pQXAl
gVyYnC97DVfQ1sLripAfzA2xTjnoUoAmJzGvj3fobta+oAyC2PAH5/zMKemuhSNen6FdvNWzvdUW
Y2g0PmGg/r3/FsHeNACNjfiTifl2oRLNWPyO6HUjNcnW/kz/SZa7TuVzBAbFrBuM1k3JZmH77uct
5gMb2y4HTRfqy6DxqDVUv2ZnMwWrdYveoJI8bfzxwau6rSLUAxo6n/Wctmxc6AptuFAJYibrLMpa
23vOBT1buY2fSDoBiY5HYZu9Dq2et8EgkuPA6WRMhBal6B+ZtT8xdMv2x1n2m2+4tMLfK/tCiy3F
D9aGrNaik29CNSO3xk2kbzSq24Z846fTNpDeUHT6w3xnx8R7E1ju1QH3q+KXAzFdxEc5vgxC5TNH
o6Wl9pehwg0hz8+Hb3B2tCBnM9Ubo7ZaG0/KJPpBbaP+WJz0hkg6/rP4sel2GKA5k1dK3JcMQQf6
srRwwzz4bKdXdK5X/gMyXBeZ0CRuece5e7fNAS6DhWPJUJrM7ZC40sSPr5ryyiow06EA9olFFsSJ
jNq+ixgQX+OeEdpTZthQwZIo/ABmp/sW1vEL9S15MvlNVuiiCwq59JhdfAU5JHot/46zA4bqULHe
x6Vz/j+coc4cKl+oxST1G2n0XaydVIcM7L0m52oS9tbMvtM2mD9H+bepPJ4ju8R6eyweuJ77uNcA
DqiKBIZuLGXKszgnkAt4vMYgzGdKG4u1uPURmNhZIa/3+B32Hh6LkqJ0ZsAJWobOhMEBV+mSNmuK
V5h2hGiwCBgTnVY/rl5j7uGWJ1KrVWJnu9ckyHAaxhRJjLgwfcSGofUVfFSpLENpgHcxyKMlN1BO
C5lwN8fFyASE7TWlT6/7LWqd2TYfA8xAH3Gp65dh+snBrsym8+w1t4DGriqXeWOmV98wojIjhz7O
4S6VKbTK5Ihif9n44Oi6hmomfAksvv9vWl83hOUIS6rHzYU5u8MjQ7VHSlAj5FKe8F96z+gdnZi/
JOC7u3H+uvhWSleL/hBwl9qfzwxkvleMcwv+a9z3N0Sa9XXja7PiETZoDlJSOrRyrmXEn963QiC+
JlQr/6CV4cEnV6edcrOwBJyaLlhyrt/W2RJWtj6zp+w9FEdUFea2igAUtceRfNGZncsb11FCchJe
Gb8vsS0MHN16uosfkfjmvw4X5lQW3bGs1gjaomoFffPXBCRq1MEaoOL/cs6ENaCuGiz8Z2NgAjtb
T3m7/OFI5KJ8hSob++NVUE8y5UlLzUPW12OT6YhVYHmQui/s0YHjCuaFTKE+T7z2vlYgm8+eTT6N
SFwWOBWTVq2Fh1xgpN1m1N58u6XGMUZALzjJ2quzs8mqDop3UshjTemTK8WGf+ualgKvVcv0hsYS
0YNrpx6+7Rpf1rPnOMcXKdn1XxK8Q8MXoBFzjIzantrYtWxPwkDuSErxrhhMWVLgK0nCah9M0HsP
huXt2J7pEwrmIRPfhABA6QrFqEiOx1bJzXCwq+na9Kap/i45aG5/TuyD2FWqXY3abIlxGO55tSsL
L4155mVrJVb23hYxFEwCAClIbUcI2kmlmU/SD3S8FRwoPbvo9awkw4+Vao90n7SdmngzUhKSWV4s
1yIgY+6nmlaJ7yAinFNG+j+75Ez0/8dlx9je8Yj6n9OGeGcLxvrBnvcdEGn+CqykN9N1CQgF++Yh
mt//px3yRtwCNWjyM8k6VNEQroR00cAkHVOMXngneoNSYt1UElMCL5+cYoDVuzqBCfm8ruY0qZpX
vPG4Z8R+1wC4qZfrvXrrnzqMXSnpBlyayh6HTMavpzDj+SaLsX0gc0I42i/b96VzSz8i2Ic/W1YY
Ua6LBq36GYG+UwXsT5SQMuWdyk1r/hRElLXWZSHDXK4VA0ZZi/v7A1JeojEG6NpHO6ULExBo3TpP
zy9Z5i2xnrGu4rzxxmLID/6M9EtqrXKDqGo658tEE4dqaUbTsIapzgSMHhvLldBXXBgGMXyH1ld+
2SoWMDB5wGOUQY6yKliV/KT2qELz+ks0l0ivVTVUSARgbAoLbPKXJ7SWkMortexiSuBrwjB0YhyV
eU9MnGiFE9Dln5dzSald3TbIRwNpvLPONlVfOCpRgTFoFsw4NRHxlBfcnGaSmzx/Z/JJXv83x5by
qf8ziPCXftt58u/vzAU+QifzVBZYPgXCLJPqwaSTh8isrKReI5iLJTldE1sK9ld+biUqjfYQdura
ACJcuqAsQ2R3U9juKD1JyYoy5svEJLHLc2JP09v0T+Ihd7UP3Cj2adwd1ttzi2SC0rWH54vy791b
h/9hY7EKBHUIYR0TXaHkAvUmpJoTv3VSarUMvyFoFKP1HCbaEmcekdaB6Klc/hNcCZklVVO+zS7N
vmOME4y/JgGFA77rSTPeohX45GvjE1OYLiwbpuR7aaH35oAIKQzHNw7zS8nmFhmPdI3oeUsCLeRV
9JPrl21JY45WZuJpz/NyGnc3jhtAb2HADvojeGsNMknQTivrtIQMDc5Qkf4n2CRzrlUnapiMzSPG
e+CaM778CWwax+i/t/CilpitcR4PDYtCXs0N2gvf6lbxb+w9eT2fFaCyUUTCQfrbnaYeGhf9yQM8
FsN9slGcrAmdUyl3XJyrqUCtp2Qbs47kXUIZE3lOlAERA0bm61IGmj4QEhntj8EWKHS/i0xe7z+R
JwtTiHFj/Z1N5BPbYpx1a1vFc0YU4H4NVlOqpiQKuNxvbCHIwWPd3WXgpx3Dn+tc2QJRpDYzwsxA
NI5qNTnkWOqVeLU0btWGBOStZro5D7NMnMmiOmQ55m9b8A50D4b9sto/vyx5U6d0jvQwU5+vethL
reFgGhUeeEVsEQfRkW3Si0Gk6b3PfBlZ485CIm6yfaDd/zO0/9L5cNMNZECxp3X0hcUfLmEQzVKW
5HvXANqYj9q9C6O4T9SW72ZYKNjJskyNwKu00Xg4LmXuObTqIS87BtUfHAmtDaEn23CSyB1Jb4O7
oYctK3dedeH1Yfuka1jhM7AUpp6o6T++qLVBk6XyALc92RGKiFaE/FWPlLNt/EMYRpkpMql9R0pJ
RujeomSfASERArJtkK4TqpO8yRZHwsuAR8qQvHldECNmdb90SVkmZmGzvvCtekPVnjFZjMNzwYaF
kHWfCaV3EEN9J0TX8eiwnA4GGZznfbiM+VFYIUiKhmO+jDsdFxGC6CXyWd0+qL7t/1FRI8DjsdrH
v8ZE4sXmjFtUoTjZqIZBPapbIC/Pd99Rk4wcrVY4nJakeAEIYsIO/+84IDe/ZI3n9U3GUiQ5RVgI
WsYg2P3H2EMl0e/YU1xT7cbyxUYXAqmIanr12CFkvF79jCRl+wWcfnmycdY3WaOk7V/FkY8oUEY9
3JrAWwRjvoAkwVuhTZarvUK5Q4sffyHtHBjHAhjqRZFBepquQPkyr9DMkSKbyxlxNiyL9OBL2HTL
4xtP68VUiErBZ3brv06g7K7I7Zq/fb3rmi9OtujhMb/41oztqAmqbCeizLzQb8dV/Z5FnWCeGmKb
mmwy0D2YUG2gP4G90hEef51OM1XHTUe6+6JIqPnRw9Hu8uK5SgQrRtC2axa/glS51N0dl15OoIkm
8yCCEoCWIG+QcHEOhGj/t9D7m4JCBerlVeZKyJcVvUmjkuxZ1ITew6pBmxlhE/QCuZszRpVpviNX
GAns8UI1Zmrbx0//ipkr6VMXb/6okF0mtxJCgerl14kGRbTt51Y55toA4VNwjept1WUDrFo6gAd2
2yjXKfxQmkE1hS9VZtO5shKEkMJwTW1puiRD1zMktHWS9tC1Tj/Rw8p/OS93u2Etgm+7wrlk2jgI
3XxZI4QLCMs9vFU57GhaU3YdtMTBr9d0mooO/F0v/H8OEWk3HqnZSufZU/0pMcZuwCsGN2se7UcW
iR1EuRqcvfxRDLToez6NXTN/7KZmeVo+Hvrd5mm8v97u6hHWXdeFFRqbUM4166RJrQ9jiIRZ2xFO
b5obgfUZz3Shh2tWYGuS2LR+NbYa4EVi87cJYAUt9YvrcGK66o5GBjukjRD02uvY5FKDDlv/H1I0
yaw+gYBKW8y42Qrpx1tUDXd9IL3ZMLGgxy0wcPK5dUofBpttjmzFme7Z/r1LjeT4nl2Dqo8wIq3H
vfqU2t4g6g4Edf5iH1Xj6BPFuCNyn5jN6nA0CvLe6dF28EBtT7tQEwcKIuXt4MhYb7f+49VM1anh
vVDYtrglxhlrM0kevkn8ihOHCWRTAxhbLzl+/NsbY2rC4RDjch55PIyC/LSU4WQQlfYFjfrzVgvT
6tDzs/WVrYGjBTt01kF5BcqD5lVh7XxqwRJ9cGY1y7qns1wZJeT9HSZzd88/m5hQf5MTTQn/Nlq0
wK29TUL1gQb1LCbkrHlurwMgX3xDhsHY1eckR4LfbHZfOKAfd3ntdpwWENE7dhQSspnAWBfyVOmg
5gC1gDCDRhkCzeEZ/UwTdbifGPvGkGnTRcwzOloglZc0r7Q5bBsERCQsDZumn+12OzgybtlEZbpD
6icYRpuvepNTSpR4AcRCJ49gXf0CrFb8ClZux0kkkgB9x2PxVetdIW7GkrCH3jxEcfI2Dd2CLv9T
vkvpK6Os7Nf2gaYa8DaR9L3hFDTpZL6Q9HD1nwYsrAHExX+Fr8fHHaU+I8K0bUIBvAiYp/TXdBjy
bQBn4Fx2wTn8NCMzcd6aNBYvOoqdtEoEvsEAV390a1WS9DEjNvkQOhDlDfeVt1GEZ3rb2sPTTjqo
Y8oLm7ProuudBCS8LCvEmtxWtvSZ/Sj0S6GMsiQoAXSCVVuxvzLLhrOiMvOrD8Q8szdVYuOeBbIu
WFDjpcuAMqWibx0ndQiSGvVIFpfPg/TDY6qUQI+dy6eXj9XxiRN1UHgTejqN2hVHQEhPZnUkQSJF
3/fCFYpba+zxaGZhOvslyhhqrUjFbraKSOV75iAJS9MRzA7+8Sy1Dg42f/uhGVS3ZCfPB+JaRQve
QYP4ykcaX+Cf6UYspUfsC52H7hzU+/uOOHhXz91BLYCpZiODerHjZCkp2G0UmbU7i/FpWoA/SDfQ
jRjyaVZ+xTEFvI8EtHMU2PCaH4OC0ncMXlWRj3vUvLyj4ALLZSgrQP7M1OxRxXQW9ueB6z2j0i2z
B4nmtkIyS2/fqsYAmhPnfWvnwN+qmeoPC7Fx3FGRkpAtcqrmqkQV56OQgjd5UYG+SIJEXOjywwrM
e1lFPSj/oWO59/kkiudo1CU02rUhsa+KVZwbMZ59A8WhZtxhLciuwQ4bKXtWo1mVhrCgryqIiErA
3o9TG901kHUKUSmZlOA54dIUuO3Hq83rHz+9tdcbNSDyjKoVNJgtDtiCZsi3ZIcK9vCUmaV6hoDm
qJXu0FTWyECPZJJA2EXjwOgulfyHjFaoKv4AGDlLzX3WaQ5GiQ+8Zqf7oqZfNZURXj0oiKJVNvv5
M0V/4qyGq7UlMDLguErcr04wbn/CPzFk9UwtDPJcyJ/ES6hlK7zPR4lc/YB2ju1ZkokATkQ591Bl
+jA2rLJAVzALiVrbWKTOUt6fvb9zoyanEcMOkZpe5YKvowmHlVos25mm01KYpcsFqDeBttYX9ypb
Yr7FXiRxkpkXNBl2kSanNksTqpE9+ta3m3Th6T4tlQHkMGy+P+T5b+l0AY+k0pFBYtdQuO2GnTbY
z9dkp7/4PXiC1VgtO03wVICGlrNVhE7PrO2h3pho8SYLf2PpM/Mfqzkq/uh4LFheWeDjIlsZ3NFG
T8Z0RpNvRvBHudMtxc8bTsnBKq3B0D20ttAM3gZzCi6QCZxJbDXJkYUw95eGLnkiAe+lnhaY9ER+
i+zcc/CMrVAHcTfkE64+xbo5mvfX1E9rQ1o6m0q7XFZDx+ySL8lWUHE5vCrnhThhcE1qDjTa0Dbo
Kw6WT4nnPcXM1CtSyEsOF5GEvhBVe62cUpkOzapm1ch+iUyQqXOEMzQPbfV5Eq9Yg4GpZKCzXg09
wHC6W/otMT2hJsp8HMTNc8EqVnm2OiDGviAtPbevyRA3SsMri0pefmgne3qhiYBe99Hem44WFIbE
JnnMOn+98l6D/SkokObGPOfsd6kWmyYX9XXY/BEVatTa3eGl6p1DR+T5Ea1I44jc2yKsbhiEyJOe
24pdXSoi534pMEd1LKjNGVymR1ivEQgcLgXGBrry+qYFPxuts1PW1wC35pdKKsxag/Vk5VDeTR3Q
RVBe5EGlJ50g7ATiwGpmBYs1hQLPk3tm+M+q86JV7USJnMeccAieVoi5N/isPDxbn+VB7sl2liu1
mg+balW1wYleQVyfZ9m3SfmeL+MU/CFLohZ9eEATCcAWBtKfIiSoqVLOzmQfSB+tAe3cdNxyIGCd
+Xo0gM4zNaGGr8CEo1YpMnRdSy5mRVD9f0rq5PppWboeJt98+XAcLlj5K2kxl2+hSlISETJrknA/
tRDtqTyvXnJydXNpSdBtTccao4NuGJPZykZRa9R2oS2ko5LBQC9J/LMqQ5wOHnu8Lssw0AqFmg+J
Xt3rfpOoWHUzdgJd5f1Kac7ygIZQH0aEMhWwi4A5hOLVUTlP3RyxgFlPdQwrZ8guScCN5A/8P1uD
pRfqqpY/mVlyoFgIMJML4jm6Nzn2pZLlQedcQ4ndm3oCPECFeJvHa5K6cTuFcpmie4Lt/V6MyBeg
Thn/g0CHX9UZd4gZZWHnwmba5Hrxqb0+81Y8L+KL0VvwQgRZpFPHm4ZA7jRlHF5OPzKCH+3A7ra2
WK4EsiMc/OCdoqeh5XnmsV2rcfM9Uj5ZxYAa4ZGcUtAXOTQ4YXYhwtzVBSlg60gbGmm09FD2fYJr
UxJxVKryF4wKnoyr54lU1xFFMvPpC7LWlS6PczdXIclC+bLslwL9k5gOt12sL5vJ682bOfzE9gLt
kiz/R++5fq6wMLE8kZaPaQLumngSH7tsjXiMjnGgSgcOqRRtohj1IRsZaoSiPj1GCl0F1ZcgfeCU
jcI9kREBYFBSNyjHtXAwQSqMxBtklhOyRjxVFuI52QS/82H35qF/iluFPW1EpY9AFL3I9BGvZqNL
/zvWUzJJlz7RvQr9zGUhCaQ4NlB2AT1okAsQM456tgfj4FquCHB5Ps+mea8IopA7hMV7bOKZ3m3P
zoU+Xh6OnZJpoZfLcIDGFwCDu4hjzjeb/S+BUjkq25R6w3u6r3Kw7BQ20RxS2slFdkDcC9EcJh+z
vYVXLbMeuZuub41x9+WJ+Kl6TxQcaODZ5ymetNa+/GwWOXtOpXR20lKh7v9jSV7J32lp/L2v/+Ot
rYnPOYgK4Bmf45nCsgRsAtHQ5DpinDFDC0XJ3muJePYYIWY/qvqkvJssnH2hsEGB3+Fo9oV23oFO
/Wy33BjX30WiAQiHZrhZ5hYvv7i4UC8T4GKLYq6KhBLY3G17aMjh80obvY5s2EJvKTpBY/lJazIH
N/PM0d6FRRORdAFzAkwNkPD3W1YJutI6zUC3YorMgjkoFXyHoYQIvTDA8AoXrArQG236SxjyuV8A
kKMPSdP++iimryzayWP90rBPtCRyA5RRXDePJ4H2OJLoeKEZXpgRJdbBFSIYlFazBe4wCIccnFg7
D+DZZXYaUcGX8egK0P8cEN3rcXOwmM9FUkKqsaXTqmypd0JBdbeyKZQ0eMYRkn35NcHkLEKANqzw
JkqRPJpJkRDNBI4+wF8h5Qb4Z3nXIpD1BZMzC3Dk+2noMuSZBgmxWtnYOlPgMoNQDwSk3VHGkicV
WukSbvISor8Edzys6aCKHIsmg0TP8wlwqKCRw1VgeBFZBXMwG1NX2DWTz2uKIth6W7yAGHhkFCAO
M2DBPTUqVfQWymWj8X35e9FtEXnomQGC9Qdt3Jmb31JE+XzrQrBExUN+Od8u4dz3CY6OjHS1/OnS
+1Ejb902UgjhThivPEnjjJOEPwR4RqkwxBCF6Hp28zMhmBWnfXET0jMsSgbNk+C7bqxt7q9oUmZD
aCNS+pkuTC/wXksnT2I4K/2zpRFhOayaessF+Uplfq5ETdwtUpS4KFgc8TsXcVULuuH7MnP2Z5NV
xlMlA1SGw5lkrgNdhGsW3TpisSvvs2RMmaMLe+nxIuJOgn3DoHxeUvt76O3PLI7IvBT7kOoB4G8h
7rFrdBgULX8KEEqJKTAKWANkLVJkz5hibVXrRbFxjQd+9xat99Fa/VIoWEea23+R899T+I94pjsY
1ofIdIjFVB/T/1V/KradCJZ5BKdq5+70PgULrtS3itQ1afRbs4g6WRdhoFQ31KPJLZbBoiWySxGa
oTpuNAiPQ+MYZwn2utYSrV5+Kj+LRQWoEdGr0tWF4jU7DJTCjoo192sAoGOAGy8MZlbwk7a9LKF3
TA53Hu7ni0tmBMQYqNOPVNxSeaE58FhRMdjfOaAKmoGadEDqVQOCD4sA4KYbAaPP4YgpVk5HORz9
e6Qj62eo/z+Qxu0anF8lyXraX79z6W/NRG5yU4r+oTGmOofYMlYsngAft6WV35+nkePpkIIq5bS2
BlWCaDUdwhyxCI4DkA8z6ay9o7SDuWWu8PlZy0gZ8uAJhLl5qkDXV4Xy+cXjNEXIMPibqUJ5VZ0n
8sA7SO2Nb85DsIZBz92UxfrDH5/G5nS5t3Iya4dEXJQsPQmGse0vSMIUKDRcaBNiWKJKZe/eeqEQ
TMJk5lGHrHT12dlAzF75IXnsBJdNVhsw+orfGCGqfPfUY3BrhUNA6lJapNM3WzImTzZ3Z6vFPZ24
Sc//F1CNUYaEXVzhaOiuJFs22Qt927inopI4NXGEeqKsYlnrpu5Hd5JnBH4w7rw6aj1VcQFZNFHu
u9eQbTq0JlB65c1REC9Z14SZtZlwJ8DdQ7feOYSOwM10jwr3H2zQC8QztKtC7dasUrD790SQS8nS
b4cguAu5gH3FtOsXPXjIsIYlSMbkQKOxGimawCMxP5qGtEl3xlHd/AoNZsFV6vtvHl0CRYVw4xwa
BgW5g4V9o7E46UhzYm7EgCBMOlC1SeuRMMnOu4VWsSGMHN5LuYS5Lw5lxtYW45bQQn9idkpQ5SJj
Q3GLyWZoZVRh8MU3QPWf3C2XQxBZEoHmPQ3ix6wVaa+M4rDFTM8YUqTJFAJP6OTSBZ2gD/qFkmZR
D/UMcbEGezw4TQ2wsL6frdCkntYw47K1zM1SjJu6QY8ck0IEM8IISG13Nw0NjdhBBDgTb20z7QOb
wKIg+n2b8IaXl+Orsuhz0R1fGtwg4uxzWvEaNbr2bufZW1bvfbDFz2iCQHb6ixo7YpTydtW/F8v1
u9Wpa2wzsKJM9p4IFPmXxTyGab5GkCmy+8YTyEovyoiHPgY3S2PBoZf5cZ7ISTGlpIZebDaOttFW
Jq83igQaddzm510LWphM3nRfeuTjQ6wAEoV3wKrBUMZxqWumlvlRVh9INVJDjCeoozPHJgiDN9bP
lwrtFQf63kucrmoUrSOTfr3wH14IPdLfnW3UwvAV9YIqfGNKp6LeoSQ+MsXyGI3stDjoJIuOBjX2
bc1+3MB5IYYl2AmMKuLsbFuktcM+FjCUMiHid3p4PxVpNEUB5n0XsEGW/eNwmGw9fkA2FYS/Zqaj
SZb45BL2RTNBMZv2zZK7H9F7rIoMGgqjivQLssCEdz3lFShq581JDZBz3xGw2cwYJBtFllCvLHWw
kfFonnskXZdD4zGMQPvJHqM27KO4D2XbbvWEnIR9EXt1ZFzk3w9s37DZ9aCjoQ+N0uSNo7CcOfRp
xlD//alBaZ82KDOUhOq+LF+XE6vw3Ud5WwFSK6iXvXzolAeH2N57ShDSo/z+ikxZwCm4u4w7Cp6R
PzfmKRRL4udZrTt/fVHDQyVKvvW/BKp6AsAHVxDwfLrcqr02uO1koIqloQ2bObfB6EypH00c7DhU
3coW8ZiBEFnFefdUhnvl5ybe4jMDNl/HXBFDihgQBG3Bm0R8nDz3K5/Vr+OBvyVj5GnuYSDga+FI
z9U4azRsRM9ODCoIOx7XA1yyyp/E62d0FgKKoavcSe+TX58QnAbJisZ7ODkN6palhbNGUH8ivmAn
wlz4FS2hDptSy27PHtrNZ2ZSDy0wYuVAjfVrKsme918SVWKSXl8Oq0/ayZ4J7Fw0/+wtiwo/G/Vz
gG8W5rjEJLhNEfzDX9YZYKsnn1Ym4DNYTh2+2KtzTxgJ2luWem2RNGddQJjgLV06BCzzivxo2g5E
fzdQ2f5m8WGvBl2cCEGKGcLoR3L7UNcVqFSYuiyum4KiQvoBy5U+T0dWwGSfmX846+H+nDugMhvC
Y/3XaD5dQp9vB7uHFtB6TTLxfnDytUcTih9TGBoGhHla688MqoZpLwgD+F9zs4pS7S+y33DPSDbn
ED0JY/IS/jJiUnKUmNLP6NXtnEPpbxhTKK0yi950Pvhsc0EluEJMjgwvZdX+WJGAUw5oOomVwCFz
hhG0NOvlVmQKQ0/G8c6ltoXaniQQGgnVfTWuqy+ZJM3cyGsgN+ZgfGqEoeSpqtSmMcunYiQFlp9a
5ax/TA6csf9JdF5NxTWVWa0lxkBkjWZXjx7zT0zblCjfWyErQrdRZrPS9nnF6l2rkqBR/JZ2STBJ
DaAim3/1d5DDGG7P5DKAW421/uzOYvJQ6x49z8lGz6eBMu+E/in9CphV2D0hdTjmXFtZWkD3eqde
07EJoxa9wGgvhLUR4/MFjQwC/00SYZqvV1CF3lM3Dv9LaU5kK4IYA4iUoKkpfIOsXhdSdISeWr0N
hiyR396+vf+s26as9p8E5yYtWCuhPX2RZ9LrfLxXkdR7MT86z3CsKUcFv+XY2KqeTgfff5QH82rL
tLTu1HiZzuSCPlO9R5wbn/LWANVQrIGXYarNaWEUEZDiMhdIJCcPBPYP7VP1LFwBeMyEADElGsfc
35+UdQNZirxmRNo/0t7EbR+zatid6aPp/B2MmAZZAySGT4OgMRhqHEAtN/Cgip0F4BpkAgGAXQPS
PGonPvX97P0OgED0bdCV9IEe0GNAtpWO2vEefV6coNKK2TVwkec8GaSGvbzH98jvNy/cgS8D3nlr
ZS8pHOCoNRJvbdP9xiCxL2tRjnAdyjRmMuRsRP5pZ2skyrqHbwRB09WNuQaq13gtlMxS349Hln3S
Bqvy5yrVTwjTlbRyt97eOY94t7YwtJVv0RdhTyhy6q5RH4OO5IgI++dQqE6YW8zoY4CPzjH6naVL
y4b4NsIGi/zUAywHjmn5Chp+ts6dQyvr46HXcbETnKm0j+Ttm0kK8Kkidn/OfYyyH3riV2JG0yeh
8Bce380YccUY7iTFEm8DyHKfn3W6wIBDPVWlPFcxSg8slXY5klsMRJmQu1Ko7CN0SaGs30WLWTdC
zIs0znpxqYGNPMTqoabP12u9BYfrvP3yzK3l7IkQrnGjxfa+9FmlRJimrSuxADyxEr1JkMOxbi/0
m3ZGQn2Qk51j65RvgQUfMPESUZEEstlu+oV1AXDwBiXdd0nTos2829XBuT5qvWsl4N2FnCSzqyJZ
uaxIdzuyQ+ejSKSaiGBT1M+2w6zd+Vck5CTXNE2KgcQ0LVk+1UHDfLEV9PmC9ujSklLiruMPAhG+
/csHmx0BCUBRsba27ooZkOO/CQuyuBP94t6jMXvTU5VyY/LAXOWyXkr+kdHpHnNpapsjFvOUpHf7
DoMQLbcWFwu0keH6pc2Ub7sxeWCj6ivSvlpAmViwPZlEYbqx1I6GbvA5JNtAOB+PfIBEvslzZnuN
Ds9sgW47IoZf6dgb8lUsnwPLf5Ww1q/iQ5YMCUAARuXGvXdeleaqnsHh0R9wgbThmUwnRhWiOz/A
ag7rufRHFGP9Cb3lHBuvfYly1m8/VorZNXGpDCiNAQyaXqqQKorSxhTcTAHg+qXizfAZw9xdXfcf
9Pic85YREfvRx/NJYk3ktBgqxIi8uX21we1uYNTyfaoAsb3GUIOJw6pkDxNUtyksmQplnu3vbXTR
niEA3VptruipK8r8n7KZK5QiNAcZLTD593u+5canCK01s62mKB9rrArsZtG0sXs0aS7t0pWJpVNs
QzHwXmWzZCLcxDb4Gq57FEudDjI49R+pDq0qtnSroAYW444F7oAm034JqZJq/G/pbYAw/wP6gKJH
lgwQ0lGSMfV0WCGHxWSiBKmBBcQhbAl1Q/IzyvhUyuChUtQIdAg96daQAVVRHO5M//VVqh4hGBKu
mcSDkXBEu8t/dXdgIW0lWSyQLE3GtAmNzEYU4ln9KfYp+e4lz5i9qPxx54+/oqN87LIfjcs6WWRc
SLiOg58+rUtmR6kzSji+U/qq94xHrham8ndhO+1YGqum2A9OrCQ/WX6VUTcM/w/4pSRpwlYfhLiO
uJ7vcfne/F/Sn9zut+o3zzJHX9f9d7IbapWTqQr++sjcVyjDRHqaB0FYuwLK3LgYvF/+in3GgFYp
/LGmt1VXugjKeS6rLhIOY4HBu6pxnrVZXz50fMGTlv/cLFziaeygRO+14mVINm5G17VOg91VkHwQ
mM2CywZ3vBxFHgiiJ7gzdzq55RWi2DpRwd1I7ZZ2yd+3Tj+8K43iPpmQ9oFepXyOw6W14hzuO5/b
q+Jx1EnYcdcdsb2vfR2+GRZDInY3hPLBXJMdoOICldioF1txMPrFpplrAK2m9hQbiVPXWCx8fQV2
A7oD3cNzuvG41Z1vnMKNinzSPUYOmds0tmsFoehCtaP4sIxC9pmpipqkHKdPjMy1hW5WwgUrX1rH
NtPrONwlRBwace2ZXhrXyaB0XnJiYq8MSCv4jKNQ8+/L5qJ5HD7BwxMS4lN8lbyjQGgL5lO5CeOq
Ufs/4LdfxgQwLurRTX6y3mWlk4sJ6cLa7zIYtosEHXKqoexk70jjSg1MV7bUl2T4l4tI7B+5lwvZ
xLaVAooyOHdRgQOgfZ0BDmCqmqqgCwvb+TxeJpCH8BpZ8xShD9apun71Qu2SSFsKhNLDP/QplBMp
KzJKG8gPefY3nULJLS/o+I3848K4GMt/VDi2gx+WhYFOfkHwmdHqtMO4fE3UEVBcHZjm9dfmP+td
HNgUJ2hz5uFB9v2bDNbHHxeiq5HXH5gbRo36VrWHsei4NNZQHZtFDXRDjTIv01ER7sBXTyOZnV+3
Q+DVXnfby/mWrn0xp+kPQex1rpwl+V5wn7kHyU64InLbQgJo8PV/bJDUDuzfJoKKwMo3qdiOiOM1
/zf/ZXdxqY1FVqBpiqgWyxvRsB489xICLkj+A1dER1M942+14SLnSGIW/l1mTDl0JEOKx7sl3gIc
pDK7OKxdwd77+dICRK1Jnu0sjVCt9/wTSSwbZKrfm46wTfBS5KkJk/MaSQKzkprSFhQuM3pobgJO
gSjspTrb2VFHtbkfawPOMA1rai1aqFocxVr1odzvAiR+/x6Zo1SPvDvdYy24EIXzdZLlEaGivO0e
XbpwGjhCtQOnWoZeSg45akzsMKZP5dB92bzR1bO35vONJFZsVksFXjjWduyrBMy/5ha9xICyxLlE
1IRTgPeWhih3MLdh/ovQ+GMlxMRH0ZCQdgNr+GY0ocof1Z2RgehqH3R9Sr5zMn97ZzB3KKddrHrh
jyElZnYCIGVyBF9qYgrPqzru5ObpKhmapM3Q7Xco17wtjLCjhcC8KAdBUG7bqTlgSVAoacpcNMUO
4KJk2AqERo0XWvUIeUXDRRB3MhJ6QANa80V+AWivOAHnhtuzCVPEVCpINXB9KPKe5Qs8dvhshGkA
p/U5F69nC+5j8xx4AAr9UFDPSfL9gxFLeLNI1Gp6rMM6M6HMlUsC6+1Y3Eqn66KacqyBUwjNJXuE
nsdf4KtVbQF13P6eQ4sFvCF7uS9f9iAZ+abfm+BW1t68Lmh11bpVgEPwe3gip611BjvQZp6g6RIv
ElpRkVzlsCJ1URp54J3kYf7M7XC3QneeiCG4Q+KJFgjhy54D9CX22W7PfIBXKAMVrgCi2/+1zSmQ
VNyfZpEmVK7TUpgW52Xisig+xqZZqJM2fUbSePnRCwTcsputFo/2Htwx9vI2SsQu0Hk6KB36NM+h
D6OmOT+9uDAh+S5eBXgjT4e8rIcpmrcqINi+VzdBFie8oduf2h3yDHTK9WFh3W+ZJt9R2z6roT88
dWIP5l8NXThgiKXq1rmChbglOP5S7KoLSp4+osYKbb2vKDcvp5Vl/XLYWUYmpKh2BVfn7v7WP/vo
wMSlcIkewJF20yRC5FDcKTnqgAVWQsla75SkQM826K+YNefWiJhguSlyAI9/76USO+qnf2J0VuHQ
SrzDPCTZSxzdcfuWWZ9EepLKMgTYKdIVkkt150nSIVkzPi4Jx5m/wtZEerzLhVdDTnqMfW5I8MmL
R5wGi+fL3cgIOjhpUrT/uwKgxFWD5pJcY9L20T39HCSMsPuk/V3jzE5TjvDoZcksYzrwuDXuJXIL
J3RhwLuNY5VKtRQQ1lmf3rX+FY5Nv42ixLRzdw9pqmwh8+tjCIKwbupSoca4Ch9U5cv0QgrpXsvN
RbcQrfNwSJkx8zdKcAg5/Vgl1quvwVTwgNRSaoLSd9dGzuMzeJb0qw0HbOosHZwxvyfNssZTfYmE
ThfvkVHi0a8PPk2+UJRCuTe9soSaoWzF00//4GURlK+6PXCSy+C+Fhjv+nJ/yphu/BucKcBP6z+g
7DsCIWw6ZH1zOHV8PhLdFfabC4kYiPhgP8CcB4M/jOwdf0F4iimL6F5mDDH8cqceJkaLJaRWRI4C
3pOlLMwlob6YQYWA+CMPQmsnIOnfqEAEHc6n9Y6DmhXFryPO7E6fgpLNKobOMTlr5RAEWb7Moh5c
q6DjQfvzmsAqiD/vLzxltHdiFmYYyny6vpGxNmXbSaOTEXbiuoX8VuFxQOulQqNnCpnu9QmWDhKW
9/DqfFj7lyCn48FZaOaNPdn5qSMKjy2ZZJ1Rlc9LugkQmtB3GgSPuOl2j71ozMtLiY0+WuuL0dLf
bdA/HUjygP8Yoo58MgiW/fLuSHWhDNVJCSEvyG5C/H/P17tkPtWHdyL2AYnaEf8wdhZiHiRH09ju
tdrqlsjM/9JLpS8hxs0p4MgCQ3O1QJ25+uv6ooC6lPI+2rR+1NP2E73Q1IYUOW9bexH3KcCeDp9d
ezvVnHCRkqzt7fbwfxrRN6ZSljMOzRjF8/42rV5jeiyhKhTmAiReR4G7bmB8WdwTC5TO/h7ioTj9
UmvR6uJpJwVusGHaAA6oS6XiaRolv7RZm9cUsJUF8bYovPDJQGhjIIz5zQua0zsfjjXgFe+162AV
RBUfn/DDirqfnmmwxPs69g0TF/dl3Dk/xoni0ZCXxiWAT0KwhImSGOAcFvppgXQmdsfnNUSEHvC0
q210OLv1FdtwS5t0QojrkCxK5OoM6poLQ5yqciBRs0X54bq2fScBK+U/RVjRD3MEhazMXQ3SO3cq
fodrzw97SXiiwbiZMsZP68m7Fj7Rt4gEI+yGp9y6g08RrbykxsIOKXlHaqOZTxpBMi9s9A+jXHHV
szoJgtC0oGKlLRfIPlfPB01624Kg0cRdzJumXGbc6YQhdB1GrR/1Qn8wEzLsM108VgZSRHgNtB4J
atRYzCSPz6txDoCrURSsWGx09J5MavvMNpKbNY/ETdlXqOAypToOAJvrcTuxg1v57Q2Zg+PfvBJR
d2J1q0heyuYprxRBhzn3p7h8JgDoWT4I2yvNsYXRru4pwn+fsWU+AvdzidY7KjB4paoHn0JrnnjI
PnurCV3SHrSeiZUqlzTfjenKz4a7RavuV1ZjzEMVuksSluZcUZBv4fNmFtPLho2DHZPejfzBq8lS
+aQY9kedwaUqHrfHgfuamvXb0vp5kkIUeKXUNhwSS7RMXVQUYVy8aWIQLiCGX2/dMuCyiPcfva0k
Y+kH4bJTyyZ2Zjtc3icvjXzEDuuRDgElCA+iUjtEHnbU9QZdxhoIDAU+UNRDRsW6k3DG8UdonPcw
AgxctESp3ftHtGzR5AtTWZwxLQRnff9LLatKwXIr4LzWYfq4+VkVnh4Yot0ba0eQpmG6/W4Cd7+p
Z1ohnzkpUIa9FKBOB7EuK0jz/DBfAnW0YTRQgt/ClbaLWMgnsxht6MMQeLO5t701OvD9UuKhTaKg
m1lSyKP4h7DUkd8UcZNp5auu8YLR/Z2iB0PSsBxs230NLz3ojfj0ik7CtVfRkcPTGboXb2vLzlww
0BXXKqVStrvM3ca5KLBinIR1GUOfOXGREc0MZThe6715EfXMTDgu3Xh8Cy9xaQbU4FBWVwCNO2Xm
DcA/9h0XgsgcQvOARPWOESqNJgL0XPa5jFA5lwQSkHN9iVjz29wWy4rd7P2qdMPEci88oPxvRFgm
7D+SPxzIFQk94KpAHDptDNVnHb+WVqDkxn3iZUrPe5XcxuPd4/6eL6mkZZq79mKweEvVMsOtADgV
wCwNNpJF29qgVnOVEki/K9ZWn8E4MeSCNLJ1vHpKkLQMWjy/EjqgYJSpns5gb76kqenHixhW+o+i
jVv9DJOkcgqFOIU8EkB5otdg9yaM7x0nBYSoXKjm+43vmvVy++Ko30ZccNCLnNchSbNq9L6ujEaJ
NcqlDuAegHBugk/tAamCKhOjfLqJ7A7TQ6h0gGHGqSPGbvO/z0OXyhSsKikeTzdbwttgZrHXzhFY
GrUr9wuJ8YP+TrbrlhXbFujAFV1gW364TrEg0GZYvdCM9jzJf+n5H5PgdO25s5F5mnK3o6ZMsgA0
7bwzQrO2seoU/IIuuVYqhM3+piXkII8Aw2S39ouApKJfhrJETJ7OwR1kQthogi9Nke8rUy8sKSX2
2f6WDYrDoSYfS1vkcHT19cOll9gRJqX7QSU8OUz5MyteuITQNWbJysGfZy8rvbcpaeUykJJt1+r/
EeyacPczMR2bckBDILArm8Bi49r/HrvYQuCXsP0VeJ5S3XCUlVvHyVJW0rwAstdrOY1vD/MPEDEX
8BT3frHTVuQJXKkH2GFMzzviXM6iBuVCjIxu80QCd/COQPKctaZ1GU/MbLDVZHs2hVNKkBAu3ZMD
as498hEFAnl6sj0udEdwVkVnS+MCICVor248v3HbkoUu9+BKb6HOuV3nB+gv6qmuOsgeBkp/9Mer
v+6susEmtmRaXRxWUiPbtfZcb8Ty5gZU4gvbmzuwrd2cIdmdCAFrBXZGZFDQYU7FLWouBfm4zUwW
4v1rf+VR9u9+jMADyCxTd1VUkhjcpe0SaX8JLgOX+Kd14fRL+VV6j5rk9jSdiP8vP0HjkRumkDk0
IEHTYDXS1+1nZsCBFBFSyOB2PQeQn3yHUpQasA8wcLjuBng6iT+m8Wu4lxIudj8CkKMmpE7LhIo3
cDU4R8pIBQyrv+wyD2k7wNKMy7+iepzHbs1tfn8B42WdkNBkwGiFD2cCBtrOcWqQ3ACmVLnrCOtr
e66NFqUkN6IH3wrDf1xIOHQzSXqpqq95Ivq+/y7UuhJPGdWt9UVcJjet47xZJKhjFvjZqsCGWH6U
trRT3FurT1sS2C1e33k7L3GvdKnlRZp2GufCLxjVu9f7eqmlGAh9cVWe6r/a7EAQQMtQQvO4dkdt
lyfa9aczU+7a7zfROuso2EHN1+KVMzCVTy8IFr8Rsu6cWiRpWr8tLn6/g8nOANgF9bkKu5T6njV9
6sELvunH47ozm36WGBYBGD77/JEWMuCu/9aNpw9oKIKVXQgAftnfs8HxJTxQ5ITA7+2OFHN++/8T
fAtS0ghQHJXo0MSV8KdIH4TTQKsZ6WPXne6c92mfp9pjfxtmdgOZ1uziLu+ZOwZ3mdFTrVsLJ7oJ
vOQ12GJ4PM3fl+3m2KSkh8zI2UPauwEO2AqHpZvQtqTZS4Pm3T9AGcmvhxyLUeajNyH2dcqGT2QB
gb1j6WJe/fEEcfmE7ec1v76sSPFAuM8cuVgwk94tA2kV+lopHTAal4FnXCHV7Nu8+ITmcvxdUj3S
S/fR/VfQsYQOifcbRLPSfEbVUCqvZyiK4tdIhHWEWZ7IKd2l4hyuWmtXoKEm07NamRe/wx5yPJjI
9SOf4xOC7P38w9F1RRCq5CLLy3Xr6ndIacUd0w2IEje65Q7o0fcHGmYO9tmgYsj3BwSnygX0giOv
3s/hVU5vir7P8EfV17xsfirkx13H7ODKo0Tpn5nprnOHYu3RAOPnayVW6fSh94DEVi33xp7FmVQH
D3gixcNRZ0CyRDWu1D16Z/xXee1cJGFnEk094LYlqleVKIasN/v2cEebZcSj310s8GfizBYSdw5n
kwWwQYi+gvQb3X/gfxGgtjsR1h9kgC40m28MlwMjIRxtXWWSZaoZqCXFzr45lN+bu4xlSRVhAv1c
BPPCI/RMp6f/nmQHoTKRkAHfezhVfGio2vAo6RP1wUq4po4euxCYndSU8c2EULhh7UEwrFDzDfHb
+MiV1VLcjy4V1V2toWGqIkin1VTl8nzCYtJu71bfq0wzYl0ACRl5NuZUNHhpxJViBTvsewwp8UAk
+oDMKwrQvIung0/WEJgqTwZm+OUeZFjnp24RecIEEsIC/NwlSS+NDmG0p6qpdMzkIh66hoOEs8uD
3bMdCfr/btjP6TV1QhlxLvRZRCNj6t5ws+nqvm/LwXoD5c3QYmrXmB0PMISRNS5fd40dqEBj8ISE
XEL8WtXytE6pO3q/h9mB8QXBo/6t/cNJ0MokNy9P8SMGJCCAQtvNWgKTsske6Upu5e14jAE3Dwu4
KxxtfqXA9GAtcrZAMsW1rXmDJcbPLn5UpO0NsSU1/EcgvEIrSL5PT+lTx4Mz9p51Woh8gJftnSIa
TINz24FUSg9fhy0MWx/bDSxk4pBQmtBPfejE5e74KoAfvzHILdjar/cYeM+pOXi/9lDLa2ZwU3nR
0ZyK4PdobaVH1wTNiFkgJjx4QjGWhqe8f8ML1WIPbyaznJR82wPF5xWy9nfkir61CiO9eLgJeZT5
o2r7p0EIRaQPyaMI7jGB/7kD0YRHgbjowNtqhGPUyUeINSapw4ISod8uqe5zde8di2B3W3NPeFrO
LGE+ZQh09/rGZmdC8mzWA852xUxit1WXvaKFkUXhHBxAbT+xrnhrIOPS2+yJWEgk5cIVvnRtiYjT
y4+6gRUVI/bcj36S7V5dnpjtWr+QSQb7vDUgqeg99P1p+ENTsZRPsspYGxQDjZi6Rf/ybaiGFuDP
Qfj8ydneuhPG3eH0R+J9fiGRR21V/RRH41xrLosvFX2sf79ICOjtf+Mgv37cMEEG3fFH0WpuO8Pi
2s4wF+9Dc+Gym9xOLRtrvALIJBnwgNmzZDP38eXXPMKUwTYqWj2ZuMtfhy6/fYpq/SHPENc2nEqg
M443FW/lTZqnwHlUIsUkZhlouyNybSBonbNB4RY41Mv4fSXxabWf4tfgQ1jw4gkKgsU/HvMScsq6
NZw114lSMFQLERqF6JFlB/MAkhJfIPaUf8dixS6kupilUWhuldeY5o4wqOMWPZ3X/q51CrylKwoP
K9UhYKnwWtu8rTKfaP9e8Xhh/H75mRxpCC5sysLU+5wrDvY6C4mj7rrhB2p+kp9sLaGsu4RGEsiD
3meSzmeReK0DjpYpgK3lV464Hz/9HCLL32EVqp8PrfyizB5mdOWZ+vJ+y4RTJIg/AiRm2vqsTOj0
3+zWZjUwXxso8gASAKj+qoMTKATjmt2rjwi9WZCDUwHryRlU10QCbp7hYUY0VdhIijRC5NUK0ttm
UkGQG3Psd7pKRcZK8DxSkAuXlrH0aVaptMQ8cO0gghaLwwmggYYnnS219o0enpgjsJvHImng4n2O
/cBUmv3On4eZ/hBWDaLvfKHtTNag+pzymPxRY+mzP+z2e0un83siFr+kpPVMOaYutBs1wISaRH0y
NPs57WzoxFEyCQ8SvRKDiqkFN0gPCyCFidSjJLIw7uOliSZ9FV46uOw86oUGf0BY0cQbFaeYPerm
Axjnw4A/lsEu5apqsWKtzvRBcP4CGwJQtWKE9fQSqdhNCbs2k99LgTCI4xZjU4/Ze1vWz6LixjAO
5jj5OssRus8tjZUDT8RTjGP3JfLyUdGN/1GSi50RLWIJV58pDcixXQpfTrECi3GVkeNNdbexzAnX
DiyoorgomDFDy7E/uBCEEmgpjwiTVaTt/1SaJNb1aRI0DNqdBJr7h6PkROUTsvGkKJ72raoNIqXw
b12q0pdmRIZ+FuH47/uma/s/r6goVHsIvHOaQENV+5H8L7zCsHQhBlbl22uLsemp7DoylQgEqnt1
I64hBNeu8D4s+Zr6fxKa5JuVsQ9DvbIr5oi9KaIbzZ8hpRHbm+TLUCRLjpFSyfGGYqisn+QfN0Bn
jVGPi40qt+ndBswAKGXQS9DFWdgahvyjq2QMGqo4BoL4GskACZowCPcyPgvQOmcbv/9XcCHPdocz
5uFEl6guZxGcBk0NtmB2YmDgyKzGNKKl0m6dEWhGqChI69nsWk3b1rZVXruPP0uBNHRChkQfAXVs
M7WujZS79MQUgBzkfBhVjmvino6B8TMBzJ1zj7CHkwfb+znRRPVXGX2i4yUHd6kNelPcEDfX5uHp
FpCw3Q20SRQEdzf/rqcaRuc90CJ7mZ3qVJoB+oswk/6lSWQUye0n6689COZsdehqLgzddgB3hHN/
03C3zTHDZKFAbN61fEoW4CXUMaA3vttLmyiilIPvh27IthxGvPgiRQLSi6ar/KNeCoQBo3QL6OYf
EnWr4ppJ2WGOmdIyA86Kawi/ca+jdcd+FPy12yaIIccdMm8T9Iyfe76hY032rTEzFR6QRNW6utr6
6loU8egmmhUdE+8muEe/bDU+JctxsvwxAAsb1O83YCV1sF/kjVRQSPe1n+jt/+hEee+cMzBn2mtw
zvHDxTxoD5tnGGI9mXYOR+bI7qXV4x/MSIL3GLKHIv5/g3fO+95FW7wmXOWw1J2DdIWlRTHfqvBK
ANnBfD+DlaPFDiCBzePFDJmVYZXUqLf0MbJbwa7v05sKQqLRe5INDtb2JMMmO3o8zDgI7w7Uf6GQ
7yyGwtiEomUhrtQdFw67tVzCleFtkTfLd7diPPiHMFhok+MSt68Jvd7hDSmMJ/sMNE9RgLLeB98W
Gy0+K+LPsm8zofOqpO0FGcJjA/ANaXOolHIHTICgrTBa51DNQyA784HT5c1X8Wf09vZACNUhb72B
8c1ylAYLP1fccF8GdZf/zDyNiIa0gotqEacJuLvc/OaL3wPeMo/jg/h+uqVQ7QBpP1VqQubJjrj9
+gYHEkqWd35nmOegvupHUigYuzPZ30lryRQUgLOoW94Bd8DlzmrFXHvZfOXrPZuNnrSC1EjXc5kB
HZ1UuJVpH16xS1z+5yW9Ub1+jziL/nQyIVSrzkmjypyA+4p9kGjislSXrTQLY2FcQd9J8d4HnPB5
SbvP2Vdifo4PCN6xy7gezlUWJh3ZzO7O7ImfcIWF3RP/9Xo8FlpF2+TyvxJS8wNXbFtgbIBNUOCD
lbSsX8wZP0YwnkrywxZvJOyZKdeXeAwyV+rnwIbvsOkCldnVpkpBi+WoMwOI3I4zVSXeZmUPpZGP
0uSgT2j0JJpff/MjRdEi961kQT1mDsM/e6/7D0GTTthxtJbQA5RljWWOqbpg00v43ey7JjpfqLJr
zKt9baUMrxcn6+CYxE9Ez7Ey5v2649gRg/nyHOmfzrLkbtzeJg8jHwsw1LSNQoTRMWDSSEren9xF
2LiyLXsPWNefUp380mAvhAZPaxXZuMxk6TdWbuW7B+R+t8XEbBQZwgPem8lJyELYKjXue2hkhmjC
q58896yiXzr26cH/iCJpcj2iIqGBnsy1Lg2cuM8ZqPWXvaUHidw22RhwvP0aVuJR7CDmdpSxCb/s
uSgs4QnIVaBYbRWGWvb9ZxkFTu0jsklbwUv/YZNd6BdWbrvjytNDH2W4hGq+XfcAmKEL0RGgAJTX
u/ktrvtp+r+oRjbmCi706YtQpvF5ahVjLg9fNGU1z1dAZ4A92bCNOFgUj+gIW4FxTPhJ4yIXN245
+R0kUhH5a3i+fg0s8BQrlLKt9PTk3LR1QMYvc6JylK1Mo1OZ/5CYOdTJpDxTmQYbBMljQT2wSify
PvXhqmhq8OLH/PBEP8FNC/TpytOgkgwtslaUEAwOy3uIWzljZA1L6S+04zqI9F+mFAg6Vdj1jeZT
4xQZbWW5AQHuonhZhaPrmEuAlZJY4cE5doPqYIvBU0q4r61LVQtk3ibSKxnNByY6tUM6c4F9M1X3
WTo1XrYNLha3dLpL8KjdcDmr+1UkzRHHahsXmTSOL3QCAYuUe4iJBB0JWjLWDBX15uiQF4NDD4IO
JAipKNDj6kT5muWuDbTrubpwIqBEvUjGiipMe31HZUiefqh6COowsWLaH+T9/FD55TLtSJ5o0E90
bkQ99dgCYuhYhKN4wZjEAJ97dfoGhGdz0YQFuGhnlZPJUsqzjyPUy2yswqy5SBrKFncWz3zxS4YG
xKt7lb1UgyHG4ZyrOseXvhmuzW8usGQqO7xKweaXIpC4mPI6s8REKCB0pppj5HXI5IkVVFMjhgSI
apC2jhETdb9rwkKwybLUHCExasyAbdHiHoPy8wEK5LdgKoGPbz4knoMfGApa4RW8UlwjhaWk7TM/
AneRP8VTzBUdevEfDUqUdkKwMZMQ6TZx69xADRhUY1MTBYlQSDe1B6MHJVXu05AmEldgpETGw1Qz
OePT/p81RnVc9VL90BRCTq4iMO4/BD5BEBQaPm2kpZfhgtWi3+v1NeugVsWKs1D8PJbFduTib0Od
WS9Lh+jYc6XOjlEjycfTOPYdYDgWWL5rvsibujW46OwQqLo4CSXFyLvgLeJmWK+QmcgQXVW02lc4
Dv2IGOh4p64NPlOVGm4J+rsxHPXPdrp0CFLgbXyMmoK/5Tkg7gu4VQRGFykqyACBQabVwfA7Ppkg
s70RglxdzTYzSoqNgjQRthuJ7ssjLP7ghS3t1erI6Mw/AIsuBCwOydnpSffc81SRxL8bJduKgcEZ
qaOE6Djfc3Ohu1YAU0uuhIx/IdQSsGnYWrxbxjkitckmcLLYD65DN53RXnP73bDy7O6u5tp2KBky
Y5fhYovJxPJ2RLReOKVDIPEaAcHRRDA8spMiweUSkWCiyKhAz6XJ9u6ZWLSfYre8b+IPnucqDFh1
Q9xJy6eCYQCEBmidjxiSxAfkmgsK5YZaoLBz8J+gQyOPzIPFDAmabcp5B5lF++eSaTue8L1RdhXm
YRrgkRAqYmNSXgF8Bjx8yUwsorHkx8dS15rg/4uUWgE/MRRik5N77wVYe3ZKWlqXmj5cPgxCY9SK
z0r6t+ca15rBWplsCdsn4f3z5BTcchD4g5VxLZ7Qw4/KfEcbX/AMywTXQ7dtCjQeUJB75m8FXquY
UgWjpYe2OYpzGTPPK26Y57YgYzndsNi+jf4XU5C21i+Xbj/IHgSfBfZlgO3Dgy1TpIuw1A5PHzRD
tQPRiqxHdpboiWqIn3+8laE4OquA/92HbNHUyUfjdDSyNAFlu4ujZKAAubeaVLVKyrjPFf20yeAZ
zmXu6+wRYCypJVAuUvVlSTsBx/aYTYyy9LhUX/1JSJJon1/LMcDI98JQcv1615KPN/HrtmhmrA+e
37uYCn3eJUwFkO70bex9IYQmLprmNxDNW+T3H+x0znwHsS0cJBIgcZnVOkzsQdswzPUpz1GMF7lS
W2Womf9hIZA1JnAuUbJTIdzS9+lF6FtDXi23P19KhXxj7EkdD1QwZxxclEiuki77NjD8MHK+cVgL
9yd0qHwPBed0UX8tO4GwiNXDJxWhLyR3QVa6ALw8Mle33DdvuPP3yAhe8A2FPfVvvY+6GSXu1nZa
qULVL4YSyL4kkApD2H5mrplKws1LhOKnMBkS/S+dnvDY39EzCk1N9QLUc8z0+Na+lSpbsYXHXuV+
A3/LlkRA3X6eCH2wtWWXrS0C+B3IGltkAqBbOK/vFd6I6qsUEX89hg46PK7kqHZD5pT//Xufbdwa
fFxlCsbfavrR87Pz5iRjq2R327MaLN8dZZ2ItsqM8WM7nZBSbwFxF4ClvX0FXwNN/+L4e3oTCyKl
LaGBDtW3knNrdsh9TzIsnNDfq4MjFxm/u0WLbJkbyWQxaXhEJgfIeXU1XcnIysKNihnVL0tS33bV
/fUYGbEKl+edFOAR5D80WXCYPCNeUFVzUu6d2rN+ExODW0+2/EAF5AT87wUPego6IsKetERRrnIq
vQd6U0pk3Jaxw/asYqUqeHSqx2iIxeWCe/46T87ySoA+pxWV2kz1IprHTE8gVP8dSg2+6f1gK03T
RT3pHkcg7+B0a84LGXXf3SzoJBc+kdE1HGqDHYzvb0GB/Ka4r/7l6PKKL8hLP64nxKNw28Ah3HXL
JXdg6C1FLKK4wzon/iPOR0VJOPP2HXmI6vZh10Wbp8E1nlj0n4SulTbIaBn6yxILdoPP6D/5YVRI
kj50Ydv+G5FJZI5wqA5NDLtvbjRfWAlOlmoiHq4vNqKuSwFwyr9Hz9m57gSJqFkkA1xnFR1wO9WP
3sb8+UP55anz+xVHlbbD4Q7VK90Y3VgCiclmLewID/7cHtU0M6OHg4emY3N5lAwjzRS5fenC6ALF
26v+WT4cjb90VK+/wTmo+g54ByMqlkSC/BgiAFsdfbuzr4cjQP1G0Qv7NzDgVVqD9Ay8ccd73jKU
WNY2hws5IPe/e4/DSVaA0ffVMb0V3ygESgsQJVtudvqnrjEKfgSnE15PyNPT2AU9qNcfHeGmX6GZ
rHrrgs8FqohBUWUfgzQYsVDT1pFWiXtm/MPpFFgoYFhzrkg+gDwHfeaXBGMGzJARPdJ4UA4iz1AE
B7Jl00gxACettqgAZMmLjVXdau/FlB3anTW78+m9Ui2omLdmNy1iimtPgDS14zZprnnnc3B1w7F7
LkzIKl5prHcd2RxkG673cIA51vnBiH/hGK4+5rw8uqXXesIT+WRIqbe2RGT7KtlWzu7j0rEGgPJp
Ip2tnv46+fv7CQkTpQjxKmUuusmxdjmr5063FUzUs0mgtbA/nIJOHemC6iZh/7JvnF2g2N3wZoFB
n4NhNxbyyCYxf9uJBzDx+va1XHXvIj6dDJFiYwK1nVeRoXNVISp3uh0L+qIjyfffSZBxllF0bP/+
jjTsLfiTDAEpwXTWaHSQ+dx0sVhjDY4tkSzL406eC479FTUuHwzoucY3E89JeZ5FwM0XeRCLGqUv
ZcUnkJHB5uxRWrmmD8H3WjVkOI+qoyY17s59yzcvRu/VjCcI6WZTavcyTUDp5eJHeFNyPsHDW9T/
Rj7rw73HXpcKlmFd2wdqyJirqz+SAUUKYD9Pj0YfrbEzuQzmLYLxsUu4YMacFKceAqD6q0mf6xC0
ZWz8RbMkYSU8alpjwWzXOiUpbisgoCyuJrAzBlwhBcMpmdkhIXXNJxUoH1oaWUw2urE/Dh6cda60
n2kd5oOQSgqLpy+I9fjCGjvHVk8ycBpXbLnLXY56iSkUsKOhJSrSOHzdCYqPdzQbcg1DxemEUxEY
Zh5b6e0jmdqEuEoiNSqOVAXftaZo81/nUydrOCC1aMeXi9hk51NQo7F879fj5T0ZWRSdgI+YTJaq
ALvckyv1SyYPzGEq06lkPRDc4XykdxNex38gfXzT416CgRui7oxMi8DvzgHJm0jXME9hj4wE0OoW
EV+V0Ic8X7XotXO2RPgd4J1qVqkeaW3FQcn214A8TFTTe/HlBnJa+7NYmSlnVLlOJVo95QqLP/p3
tVbEXLkyJx49o06k9dGaybnxfZ0wWfArYJf3Jc68BqhW8z+4mMcKksu0PebPdTU9zETikeV6lQ/P
k+WyzCDgPqwUaXuGAh4icNfO5TTu4GM+gAyyhnfI4gKwD7CKW0OX5t8DDl7pk9FaSJNiWLy018eN
wKcFjTAiraKw0onmNh3iJ9yHKKUaFQdTVlO+4AGexS5RtEz1pQDf1eAETkTfgFDpEYR+A+10YRLr
HUK8KH93hB5ahp9viWt5Ht+iLaF8LLtHItEcD5WDFss4w0mZiuboP4u0KiKdvcMsHjpfn6WDtRDJ
jeMF5VYQzmSSEZr/OZzbg0HwT2Ma/Wy4qAWmLmtlDtfjz2JACf6ntnUPo87iGuo5VhQMmMBZiffI
NShwylm9PiIKVfsvWRtwuhsMTR6tMxyxc/WLz57OkEQcUlMHUV/1c+qNiwrGeKiH4risM5v595W/
De3N5T0oADbZ3xIu9xYjx/dmNT/BHrBKfWPNZalLZ218AKyflmnnDuG/zbQpwWUIoaCWMOWqtDXx
/M16eivBP9FPPfTv97oGWDHCoUIRNkzCDCx1obCcImB+ZLWRl0S16kco+Tc//Rmo5JIcqGdGS0Ec
ElRfX796DA7uCrQYz2wKr7DARhzifqjxLlIeD5d1wOSuVX9UA2KcEdessu+KzOlDbpzKxaMSOOwY
7BESrhZSnLaxbMA29qKYeho8ptr4mtBRlOTpO058o0Htv8GvLcnErWojLZ7OJ8rLcR5HcHs66STJ
yWGACwKyIvNzr6te2d5U48gTjJHZvFeYABwMd04cQHUiyCskTNRW5CT7EMnFPmAJEg+91TjFklhf
mknhNLftcv50LgLwQxckha4YKtAaNmb2j/MrYCt00gmJcRKWP2oFtSqh/wHDUmACQuYM3wUZ8lIG
YB+U1mu8ABMScJ/To/RZRnD4Up5wjRLKY+0PZAiKfESJw7/efOLJnez/VZwmO0TRpI8VvNdW3q6C
xJBwsRiXjGvlAgYgpIL7kRspwcTm2X0TVFqiYQ6yDLRY6XSKxbpZQF5DbQNcz62mS8LFu8IG+T7y
NvnGenowi0wUtw9vGWKDyQxkYvZGEsrxs7mZN2yw6fVCxuQBiIj2MMQF06ev9ylPttYf5qUBGaBr
OyFnCM7+XVcK9iSteD8T9+a9v6G9KTLeR9ViNfkAZ29q24ThA1Pm/5Xx+6VwfHESGqIKffykrRT3
VV8MykglXWEVxZY9/WFzHQ7KuR9u3HdOp4H2nB5A4WOdQH8PVMFL8Eeq99Ni1b3ApwDAbuL2Udr4
mCDTF0lR/GZRSwb4ZI6KF2rAsMJwVuHhwRaOf2zFOx5XBLCSEyZ202SebmbRj/SJEmIipSA20eA7
t6C7jwTw29I3q+/o59B54k1dO39bPtA4xQwsAqIOfYYiq5/SyyM2QsHb7SBUkuY2zj+qGqphYyCK
VrDEsUcCR0x1MeB4UravJGmOZX0HLibyv7V4ImpBgWXc1B84HHixlbJYpq4EzzzTSR2Z/ctpOBJg
U3E2RLVI3jmQhbpT3rbjYk4Ie2I9Bh+nZVyH6ZqcfEO9l4DfOIKDB+pH+/Xit9FUDpDgkhk7ucGr
HVEStLCyRRCG5/z1hkR9u3+rQikt7mSEpZAO9FbdmLSFt2ae5oB18LtxJ50jGuh6RA2V89wdB/Fo
ZrAmSAp8KGFSyI4FFZbLAzLY/0VhtnTE3V6hKJ5fd2DFSQeS7Bm4N96wP7Y3fZV0Ka1bT4Hwmuv0
ktypzM9zTLmXn1F0hDLNog+2bB85LKcUD4Id3r2K8V9QdFgHqP3HLevqQh/U8RTK1C1RGGCZ+RBB
RVyMpLjESuIULlveQulQwpFAGQ1vs2XQnekYJERqlZveb3363cV3g9lkIWOJhlfewo13l9tjGJhu
hxGr1+yzWxyJHxWAJlL4UIM0u3411gJruqgEnEBxQaC3SPwK873PAy2PWvkK0sUYmeSLIQ17q0P2
rqv7z39IO11iTkTNg7zmplS+o46F02WMb9v5+TqYGboMoCoxokYWzVrou8/Sx38CP4WDVVK/oLLO
9ZKf+OICeLSl0x+63WcsD+l8hjQK6x4/5OIBDpUw78ILEQDbvk954D8i7ci+FQhKx9aJkTuQlEgO
IjqtlXXQXH1JGL6QdKVT+zYzgGYQR+KFSkEjophiLwLdHrwMKGhyDYGeIR+jZlOs5qgX0wmZAVMD
yV3e+DFI1CoBXWQwb+wdU1d/aF4RVud+89/6+UY/hdRntJkVZ2huhei7urPg2Ta9iMfpCKV/0AJF
5wwrRj+xdCh46K4YUTpydpKl9DBVJCdZXnOw+OAk1tQIRXQDA0ywdIisrSYnsrV1DP6jBNv7ocBb
m9XZr6Tps9FDuXy+BGVlOKE2xPAL0h3Hpe3ANlVv0D83n3uT2QIZVqr7GGsYXha0KVtpPHtDJ2dS
00tp7M0F2oDkv55MXSbeE5w+6zcXN6uJx+wF4lBNRqexBXdlISdrA7CwSRRVMEwi02RJAi/F7Y1n
fF6DS8pHmAJ5ZAiXy3LV0B4Puw19zFrfz2daYZgAMY7gSvrwo+oFmwrRe+7DXUqnDXfkMaQa/Skt
kZr+qZoH9+6UxfMZCFYqZRD0Qzv0haAPsub5Bqwk5QzSOqPOsgXc0ms9eNYp+W/NDjvpvgpgVfXl
uhHEK/aI7heQYtuv9MHB1zuJCCG3ssf6QChMcIigZ7foR7xzsP69LelTTGJrtdge9SlvT/WFbatr
4I46qA0pj/zxCb+L/tLY5bDqwU7BkoYSf0RrN5MDknCyMxhI7OqM9luRz9uR8WoutMx/hhMJFdiO
i6zESqCp6dXgxKdFgEILmei1Asx0eR7VtScz7rc4ZyKPK3nwwEYdy6ygwPK2ajyqK2MD3ah8KePQ
6U+v6lLnpKeaG1ClSc1E8ZV++P8HpNOtSETFDYsFYx0I4SHw6aLD4j2XI1PseQRQxUme5WLqSyva
a9IUZ7hx0yYiIz9IcOtEJzEIs5hq8zmkWdNST9HIMhdcU8WBhlMehI8xdJzJ3Q/Gm1sfnPi+IW5g
0HQqQQzVG1/K/ZejFYAqnQR2PifZDSDeMqnhny1c/+h84mitKB9yEqnj2ZTlx0+vhYQ7bM9wE93H
2YaRDaLMLksyxsNEhaAcke1L2UNMuclojM8guqZmKjXTR1YO8BFwSzsMPOWySWTdS1igDKrn24u+
+wgs5uY7PyR1fznrKPQvYcxVA9cBIcdwXGsd1+lKMsPSV+y/ARv2O+wxuwLElyLWCkAkPMlRZRf5
yFnFu25e6WgfUpMSVnvaDCQDR7i64guQ+4zHvWbGqsRTcbeH5R+CYmS0F32Hm4D2JqiWzXZ58ixr
XIZldQbABOhnz6H0xps1Z09ElXVk00zCMm/aA8+CkoXU2xMKuCeWsqLvr/AslAXBCnyMCsFUNO/4
+9zptpYmGUhKY29sJ3amBpm598vI6x3Mbryvqd2bD9hQEGCcHp+BoMNFG+n6KzN9QEcL5ANXm0Mg
xDmwsVp1y7DZSozxBLcvkzBdl1MMZ+6m7toCK8Xjb/ngPhHo4S2+zklk1lfZrHn8JszSKBqkvZPZ
dTwkYGGzgdGHcwIu2cK7tLC+Ddv3TR8WxOd+g+bPtABYar0rPtkOn7DNDnVSdNVAvN+dAUNgMdYg
gZxJ8g+gO2Kan43uP3TSBfMM57DfntFQadm4jUKBv2JR7BZl6D3UpUDQV/YJl3tnUV0fL3AFg+5H
hW43K1EBHmrHgSYqv71nkkknYu6FsUwsChg3sajHTJkuBRKj6wZxz36AZgxVaINqKEQik5zN79y5
gPqNbkOcQy/jvN1f205qQRTPsRmWb4ol33kfoJTJt1GxeLDb7mCNoKEINEsbxj7L53lOPx61kuFR
gkgjEAH8lu2HKMXBemxItS0Gottaq1AILHEANOO2/cqIREEFtc1OzEyXftiKKDI7yrPfRJiPLFzN
YBN7m8A6fiyVZGPHezK5bzmZ8DltP7btW1KOim4Q4W3JdIkVTxhEhiTTXfQBkViV190eVN/tYw6M
1t+9Pdfbqgmga6VzwhyqWj8jBM0DkUh07xT0+R7blJAqSN6WTy8ymxBuSiEuHEqiDZgaMNlqcy6p
COvS45/NlsvOvi6SKPvrt0dSThmA+7U8MIb+l8ZDArw+tdzkH01KFs+E6sZFuZuF1dN8Pv5fr/dK
4ZY8E/q7vuECgJJjvmb1T8QjihYiB7TPiUdBw1OVWNZGCl/jQQki/+MOrQNXgr/8GLCBfDl5ZWiy
QKZ6PQOTLvFRtcvB3cRijkCCuUjfP+9yXLcY9eICJ5VThyCIphYCWS68aTZqFXSxyKbpriNjO+vw
ExdRrGlEP+c6YBijUW+CMlzKGEFlf4v0igtnEx8XnpILB0G6wxQzzpaUzHg69YYHEvl6fEb4Fc2b
K8GOpyJUbrJewhJFhLZgMuhe8xBu1drc5VPo1M8rB9W0nmZhAmjY3zQ8LLqeIL+416PyIjvAkJB7
b8x7UwlC29BOqOz/3hrNtCnZoS5EsR0l4XBVPqZYOGJOGbbjuBMfkTBNEtCGDqo+GL0A0ozALXG8
lBWlugPllsP8TYQMvopPHpX4LhStNssO0hGk0AjvDLdL7/IgM/Z03fU2UcAhDGbzjLRmX2Oweq9S
lW6Dgoeph7eVUd6AfsHm5f6uIBP67HPXayAqRmdumJWOo7FyphosjOHdBTbJeGJwdeO2+8sQv3Sv
UJ75QFxW7WCDWZ/XIDXcF1Vp32RWvCbgTFFvErmfdkhRhzOVXcUEDpiwdJVYFJM4U1boSE6xj9v3
N2DcjOq8Gt+Yg1yfMKLs89F4zOztVrTl4pcdWPRMPbAFHW2LfLrXOAk9eW9tM9lLXJCKH/caTWSi
9t/Hur3xzEMy8cmzP8aBj3pZH8k1QdkG2V5dR7jOrXjbkcSGxWk6pf6HsoZjPRPrLbwY54199RFn
mybtcGNyRVfwF1/oXHBTz1uJiM4W25ahT4TxYCdIiYsbjj+PthhX5EazQOTu7XMQcSmpn+Mr8Sga
/iAo3s6BdosURweLaAgAbYbVpDqjrjsKU2ST1YofHcUlW+gH0cYam73tAS/LdjsGVlaemCwFJdFV
QmSDyzisr0K0OD+xcxKz8mB76/EnaJJg3F7oY6cVKYFp5yYfywPYquDd4j2o9R0qM4d9rQFBZYXU
PKdXpUeGwZ0QtvZ+AwkqZTWLO/9AIN/MRAYBdOVsG5ze/SydQtCSAvEJbX65wwxV6wxe0po7sJ+C
WEg63PhDhNfsGqW+UG6Kg81yRGYIMbmEikOzehYS7Mf0i2HXKzv8acXNowrid4GWVtl5ru9t+ydr
R34yAqyDxHo8nGuxV5rg0A8KJ61h8IWmVlqSXpfCrH5afWBsf9bS6F/jkXipoqk/fFUoNsjt/gwD
gfrM1/i7vLxz6vU8bCWj5IHlCIq4ZaNWUsYiCy3+c8LfJpGwnjGjKJV7xVRMNsoFO1dZv56YMHSO
u5vdq7f447NeaLEPNZreeghj/i4llhwMleGMqIlTdX33mcX4XvhCQiLtXHd/Y1KfG1Q7NuQNk8Jh
3IjBmM0BE77YARLNNOrT91ZpgTgVtazBBjt8vB6i7hv/BzLkM/7MGViAzNOi//M2K9+t9pV1cAcG
cFUZ16ijdJ11HNtFP4L6Dgo/Ifmxx9c+K1/a18JLj+pCKuFStcKWjmKT6khN6aGtsfntazmrw/vI
vfAlHz4t1ECU7kPThDrWp28sWhpLphrCxCU9KsSympL1u3FSdUAtyFiSB8ROFLUl4wJH5VXEDP8A
LvBvDjcT5Gv4elBIHSnWuOPYpb1SJPQ+6IsQWqIJa5Xr0Hhfue0F7j8yKr3QovgF+lJCLVeb/FT6
YogOrppHQLc6Id/sF0l14cyDIVH1o967b7AEVtlClP5Fv2ZQtQ4lfP4Duizn124UK9qfYBeO25uN
pWyHDUtRDmmTMD200cyMmUmE4vbp7gXzEFuRqJCug/4zJeSIFtwQsPmbSvb6aizPTRdF6Jfob6ok
FvwBk2ZFxD1XTDNo/JLkgSPpbaI5kkJGpHliqP7XbuS1IskDQ2mawo+c/5JSbrCxHkvufV+RpWJS
/tD1cCPQL4/WczLFnHGd+u50C3RS4K10Bo4UWHUZFZmunVEqkCiy+lOkg+LZiEMXiQpfiH2staX1
M3JNI4yQLCWqsSeJ6co5kiVsqEo8aStWCwqMCyJ8MVj2fUB34n+d+LihW0Uxwmo2vEnF5RZr7/LJ
ZlcuO8dGGYjKWbkeWLFxpPU/WA8rU+ptEgoOLP6Tn6qZcb+klNt/zKUHkuCa6nP3u1/sMmOvDF7A
zSCmes/m2kLxBCb8y27VOCIG1dkHOHhtxoVGOon2A97PqoxW6UwGSvIBnFy3zFfR90/wbQ8Gtln8
JzNyGtvkdrayeFx2+SoNQs+saXvWHXMVDqRHj/WS4d/Uh+Htek0rQcyFgoL0wVQD0eGwTlTz/2wh
nfqyck9XFzMqP+6d4GtVVrKjeeLojLzr0Q6hHPAvWjfhlfy91uLP1srwtgNxuT67dmd6D8wu16TM
xK9U2j1bFfsOoNwIXJq5bVP6955XcnI/Y9evBGka4AabdC7dWCE6bLXnu9983LhUNajgXxyYzrzY
FhrmsqqK+xYqJBNo6esvEEY5lajgJ1DvlEtojmIbuvmt28DkYNlx2VfJXKP0wW9NDamVxLIXoguN
iViVfpBZA2RxWvGPl/EOb12sPqRA/utvekXbgvSmuL1Oes98Pve+LMxo8LAcUl2J2lCX5YY1n5FY
38FUrBldJu8Qpi2HTZT+TmzlQXVM2RaPLXCwY6Xvy5g7Dn5mg5qp3s2q/bqGmVQDJ6yClLUogo1L
4nRwdfogflqkA5uOQAr6XAbjzCy93S9CX2ybMDUCjZLAerAK745iGOS4zYgcjAp9PxK6M9aisza2
KSjs+TQX3LnIhono2EYSQU0G/ZouFoN/ZBnOjgXMvu2gQHxdQ1ZIfloKz+guKxbav4T6odMlj0f4
ripd2CH0GITP8zYD3iOBKEZS8AVaC+qbVfgfoFqtDdt83g0TrZWZjuXZL4NEbXcPCznWeA+bpNAo
eioUc7mLHl0BJnLltwiLGjgLczLetNoBqtVfU+PdQQPElVo70yCAw+cNTduBbssos2MiGo4I1O6h
lNDcx5X53uQp6jU6RFfD74FxBAJblizQFLWBIqQ19bPNZAjNf4JnG2492yMvlIYDaXiuByF+LExK
dusFHGu1cOv7hLTG93mLkBfDI4/BsVI3SeoAyKpzgHjGUPMQdTGMUDozQUUcCcPPp2prF4W2fHWo
0H07LOTe0mr+2XZQgMmsSuTJu7XH0dtoSCmCOAiMDzFNmGgQ0vH3OB3yUi72vPJcmDrKhb4k7jkO
xKHKnKDoHMSdF7Fs3PVLo5R6bYfUwGks4LXSphRrT3XcqPBb/HxjtnDF365cqOIXggv6Yn9BcN7Q
Jk8xhNpsAl7zZZFaK/omZ7tE+zGTlVGGOf5QruBpzljWrg0NPFbGSWNyPsXe4ZO1L3JymO29fdsJ
0lW5jst0Hlm+zR8+GAayhbDSpJow5qzMthCy8yJlT16aV3FrddDGOOt51NA2clpnI/qJX5pGfhb0
aLiz+x0AQPlR2u5aCdCvwLrcNozKZyJB3mMTBMrnmsCSeN2vkoM0ttPnU8HBzmrwg1SZV5mJQWGi
xtMRO7a4FRfgbyMOv4juxYIrOQ498qw7PEU4u2LNDfA2gOVCmwGY0ZP60vHvIhoUPwNOXyUTBEeQ
yKnwUkY+iLD//OBg+BRS1qbWvb+WjbF4bHvWItGn/oWWZ0gQn3lIZE7LzfVmhgiF3KAPsTGk3wvW
SIDV0gHvjgXx9ooXZm5N+K6QQteqAel3Uzh+VG+prTfQr79nRVMbyBHVv69N1to/1T37RNBQwPDx
8KNpVhXm3bOCUKzccJHM/ZmsDfP5y0Ed1WDYrAoDBxkrYoSu7ad9PBROzV5Js9yzJLFZj61vZCWl
L1U0zP6zL/z6XGEv15jYvaS/yJ/Yge4HBZsVPGijOQ7TnI2bkvfTiGgmHERNQOXfUZqX2f56q3/8
gMoewPAVVuIahmyfNB6N3m0+zzP5ArVyaB5e+0AoQy53LSdI9ZTowu16c/JV/K3fuTIrZlBQguy7
i197AM053Uh7EPnNmPiEq8yGnnE+IL9C8WctmXu3xKRcL/Hozpq6m+pMX+xWscU0TuJjXmf662gA
bjuTjegQ/9A0opSNx5wbYG9CnaWZRlbbmXGfr3WQGdS7HgrjzGzgG/MYbqoILxmnsUPqWz8hXXYW
gTCKvsfqYpgRkiigxxXgjilEfEDwxFiwnqus9XkDhU5Z+eDhgt1RLej3vgPJZEIhL/t/D3As+sB1
3hjznJCTmEuGRyW7HW6zueawH89iGkAkaYKCpe3y5417py6xae6hji+TLMLkYhvL8WuVWSLILSq3
CKTaUylhPeckasRdPcQtkxCVcnnpEBfbGsYcmfEEv/ayEXt2mX5Oj2sAwXuXs5Vd3J/UI4DThknQ
PSccWWMO2MFs/Ic3ScfDvAfdzARV0YBjMBdcw4g1eRGRcFJ0Zb6m6eZJ253V9/cFEBzgxjvJAywb
EzjZtY0po0pUSFANMOkpOHjKm46iJ8/O18wGc1CAoYT5VTaJ+QyxbOY9zZe0Daak6OhpN7RyTXne
ibEAKr2Vs5nsmLNbH2S+GJ2YzdtEWoll3IKsTpPhH3jzLTXEm7b3ixx82efFOFtauhbeb1NCwyrz
FJqxldvzluNg9PKzbGh0JBn3o1VlPfIm4Q6+rW4jACuFE4olkHRlaStYbEMcDh+S8NzwQnbRACaB
Zw7k5RxV5+zhmPp4RO+Q0gFt7pnJ5xDExKMYhOfJ5h/2N7wBam+ntQWtm9bqDDfOIUu7A0PEcBQ1
U1t/yAwKEYUMj2kLFU6mON9hPsfgnLzTztRXiH/rV89cebfQ40364cPOw9PZzRZNw9tSlAh81768
ofhGfvgDyPYb0+Of+J51/GCDq5lh4bWeUetWj1OexIJqm4rOkz9cetrIolj1RDU59iHJyLnRc/nN
G7esT2GcA/RxYcJFV2xPKPJ7dNwov6uYr7yVap6h7w1OMSHa4nsgCD6pq7spU0gXk/kIKUgpiIJj
9j4QiM1Mn/Skb+sKAWSF42ZlfnAUv0r8MqBg9s80QqWP1JYSuJSZhf1wc6l9JmsWqzCI65ZZVty6
iSLMi4U/LWJS44MFi6WTNb1Em1WiVgXA5bftyP/06KKZiLrpBHbFND4PIwV07cPBCrUD2HkPNsiB
xCOuZSR869ozMZGME2Ll24jR/PqZZ42nisEz/c7w1RLHUY5htgcUaNnhv/V7ToxKDhK6k1S49jks
mwFop90qtTq5HcUPYTv7FUYs+GLeI1dldaKrKu/FD9vCs6033pFnRfIttzS6WDQqN/QodOC7KqDo
jfV2CDEx1g8O2aAdxwuN/6O1cIEMZRiBx4ILcBxZ+Zuo8IzsKdP9979AQ4TmIh0KBYwZGdUCdRR0
W1ZV7HhvbWNXGR3v+1/5XHo9vwSE2UJsMbzbrUgHidLOttKPStTlW3QvXonz2IcQYox32Cqf6JKp
mgHEOOLXWzbOrHlTPjB39iiwk+6BcYMbzrMLjQsdVLbnD+Nw/AGC1p8sRwnh2QzCpYK30ANvr2ca
ELaOfVO/SLqEBXXYw3bYf04UeNcp3v3cxMwsfTauDlbuUKz9ZwAaT5jdqI0XZlFpTqbSEsncwTEp
YiqxMcN9zJ4OhwR8EVrxI0J8TWujieSnumTYMkkA/eyXWeBRu8AxK2fhDF/qEzKfKmBvc8VTmuED
46EqZcKoM4XdXI/Rte0Jzpkb+hNIBiwyI2Yur5FU1ZY82OEry4yjaCS9TYbUqfEFKZFnHX12KpKW
IKctp6ehy8rIJ4AIaegLAzT9iEHCl7nJZkKPQ5ojQ1+MAtrgt23p5gstXHCI4AiZIW7IDLlC2LcI
D2xStEBEQQB27W7f6885RaIHOpYWIVf0hvJHnmtuQ2NP1SIUeZYK3G3kIhjDk9BJd4YoKn8kTrgS
3e73jdkKsWjTTLcqttMWYJA8YSNlvVdUGYIfFBBRdVPg6VIdLP/8h/cppQS/vCEzx1sX4X5RoImB
fnZqPHk8BQ9SaRIRjjZAERTxB9AtjB4yfEFnEAtI1ZBOvvh9UZm5RWvCH1qBXfi1/hjekqW/28ol
BXlu7ssN5tdHmy6o2Dm/lJdEtYo4HCMKlmQ9o8ihknq6yJGAf2rvl+rISe9mzJtrcoRqQS1nF7Dp
WpXi94dnSfBi2B28SacYQzHn71tITQ26rnFH5lbE937bZH3dvyjdVwIK5ilF3eGpKdYk4XAqgafb
kb6M4qR8IEiQmhAGwO89zHedI7r4UDlLhGrzU6hHKN+6zzJKfMEVQR7V+0EwF0gS0cUktZW6LQ9v
MZHF0Cs+bGUWBGV7EH9Q2PAUq/2KroAGt/txAwP3V4IR18t8nPq8q4b5wuDTeh7LgAq/bIJa4/w2
TWpvDiMQ1dghYBEWWDEWigpp6H+tDQJ093D49qUYlaMdw9WrqjKK1GnW2/ymgPStkgjPmImhCP2n
Ba0wCpTpvpGNQXTSh4TACiX/DtOJ8sQJdQjku5sjpn3WWlkGIzPnxnFtdpXKscd7E44wQM0XU7lh
5OHfcLn27Gg1YxnTCL3ddGoyv9V6OOGLrUm7Od6AOOU3M71GXtExkevNAM6GsPlwCGiGtQuNAuG5
lMH6Jl/5S0SZM1kGZYbEd9Svyy4BPBLVYckknfp+gNV1f5kkx/EHrjnmptrRb1o9P/WbxSmeD5qN
Xi41uDz8Lw3jhxqtyjJhEe+zIfXtWxRcsUsTgJ5x71da0ZYR2AiAE480AAjuQUzv9gHbmssPYxZM
CzTzBq86Svai3yAI3gQNqNhEgvue2R7qdW6PPCEgxEzrRX3l15fT9on0OGyJaSHbfAyOhr7BfIp5
WUWdNjkfHAmHcPtKRVqi/J6z/RZjZOZEtQS9u7GppII9Nyh1W+Y3oPLHbPtQqaHNLPN4ar2WNowa
78PuK2EuG5VR8xw8FxmBLUuLeqj4jVws+LIqcccD5LvakC9pA8PtN1ZZAMdNT7Tshxv+Li0SwbRq
p/WGdvv8tbZv9hpXj0z93vdL2QDlGMFiHsLBt80D84D4LvOE9tQgcJHksc+CZltoEInHblZxOzGf
Py+eLuVTUyni9j/K171F0a9N8piT+TS1UeD2PIQrQBD6hHKx2WY3msj6N3YzKVZgzQob/pEnqNsX
8CMJCdL3GHVy1BnSkmxYeoSS7TFsaLybpYJY/T02GDTj1jcpOoiSDPEHXffZ6/+wL42+DiKuyZ5A
h77iz8ni8iCWizN4qyVGwf7p4Q9OiLPRYw6VYFFDRxsDTjfKNRtp5cP9j8MoKzuh7J+Q6KVNOD4d
RB19ehI5hWEuFMc0iG6HOmNCY69wrvZagiwkHaDDtTnjr7F1a8z1pNjecsF7ShN4qaM75GlCJ/cO
vKMBN5E2BtDoozMQf4ArRbKwVhK2BeCCG+/xvjFxVssHZsVqPgvrkWvdgS6ujwUzBRz5rNfgeB2+
CSsOJQOFC63P2zIPBIErvaTirnXdXKTWAvLDrISbzlN3jthM+sxP664mVEeY8kzV12sf2hm56PVI
+C2DLtpEhx//xul64qXh1JnqHqn5s3BwcjhSsvlZUWeUzEf89Kf2rtpAtF/fv90l+9Semwn1yVfI
q19jb/xV1Vyk8H/IhCrFTVV/Ow/I7qNRL7Q06aNHRFb2r23gPq+Lv/PYIOO2YACYF5gCIRar1+pI
xCeiNqy6wP37zdKu19gdqMMCniO8PaGphTXI6regS+MxAF9bOcMOSDdVqNrnvBuPsoMFnq4xNK39
S4vLw2UPLuffBtq6xOvVZrHilcPxLozXQeyAMA//g0OrOtOCST/iVq7Sq7If+qMntb/mLTjs+PFe
MOaavAzfO5I3hFjR0KP1OGB38lpn1if/X+UAktlPVd3hkXuf8zwA9sVISyMufjynXy0ZEu68RUvF
3NqtGspLwCVZrucTYDVuC4d1e2qhrw9zqgmQZXiON0NK/h8tS2SuUojRV+AFLBpgvdbIcRGCn50j
O9VI1IvjubYI5836Nrflga4Vxvp4nAuBDbl7KGasol/iQpDekgPbO5cErlSPED01oMrHrbmlpFfH
UmcTiz/5qzF6VW8GYwuNUD/+OJdwyN61LglacqleN4aREHN8Ur6gY6xe+AKp0wTGG8BQEKCncDN0
908CAwLktWDEhMluZ79cNAf0ddgOYgwX276RRiIVc5XqtMrv0mEYE1oTeIq/qKsBwtjWN+Qx0waK
ieP8lW1f33SoR5nO0M2Pvz3JuP5lPXfz+HIvp+dAfkKFzQjqPj1W1AxqTSEX5LlMXvZ69BiMWOuI
vm36/XufPbnjop/416s6FZ5FU52rFj0AhBGXbcjWnpiw59+kSd5EkGKxyjWZZb3KI3XUca4krkd3
qeSSVebmr+NYjXa+Zk+sKFpDCXZn5mm6MwaijRdhgGYhG3riTCdy23COEDPaQSc+zg++QCV/TKjq
vuHyaAXlBlvCts+xlc7dprqPXg0bqm62hIn8QPrFOQvfI60B2GU+uEUl3nWfCdhpBeo7HDJEhu/q
EqHBftuvwF2vNTGBTvr/GSPIeiiyET2OMm135BXDMBDjo+4N5Lw8oXHN6NZuPXsl/GF5m2JPAEt4
quy8hITJ1w3E7ynFKFyVruT9USa/D+0p1DeA3y8qtJecruJu8RQOV65l01qpCjz4+ySgLo5nB1dQ
FnE17E6cY/ueoaP73tLysqY80j3CcLHgHAf2Utk5JywMDI+p44YcnfPlpCkrqQRTi9u2jMwx8hQG
Ua8U77Nx9jZnVQtDhVO2OnDsXFDXw1jmS6WiOiJIL2J8cEAq+75Eu5lspbz+Mr1I5Y0DBw8X61Pd
+1fT99j/KMcHycUxnmwEblBgHh/MJfmmX88d6UowwZLEdOSVrdHxiGjLgig7vFrnOyWw1EwabuYM
j39P5/vNhJkw8wtcWv23lpIU2gNrTQvJvE8Chph098u/JsK/JQGJmro2hGTESqaoi1Bxp+XA+m0v
NLzsc2j7MmcfMznC9+5tW+BvLvpkzW2ChEyAheeE/cpKng5B24Ak4Wrk1BV2GhWz5HLdiFai4Mr3
wsUCGyUU5HZX8MEHpXEWlCFWmePKQYz9t1pewLBgtZzARVH+xeEBqwjr1xQz9s1oynxOOnQ4gcoW
hdjpCRv1tk5dGWoXjcOiKwVINVZybKG/rSS+PenpsDSugo531dopS+4Mhqo5GtXxVeKEX8OE9eNW
UZZCVL7tR9pBz2/sX+TGqmuLLAYrk5qlmKaS6wFzO+llRRZ7rMCCVaNClC3tcPo4ZLRS7VduHv6W
KCS7qXExxm2Dfu2SNgbsqaqVzOWjyodfT1fKB2BfGB8grwX0RqZhm4mAy79S2mrkka1k3IxP12HM
8xopW+jMQzKoP3sqaRIfJiqwfvR5ZpvNWJftVEuFx814x6xLR04h2L5tUshJbtttFb7+JXbhrfnF
elLO70r2TH90LwuOeKeuqgGxrLc+bWcXABn5oqQA1+he4sbSESwSd2ScavvhdZ3/V3xhtC3LZvT2
EwoYV83y6GgiclxbIHiSxB72EJld6FDsoLu1rLcY9IkWIAqcsMMj33ADxzuRF0Hqs9s6gyv9Mkn8
84xeDPl0KkXj02mG2ZgEUqcStLg5DsCJMe/wwHq2nTiqiZtZxEqT0IPCGZz7L6bNpNhwuETe298g
+DFslq/RBjPP7+Md3vSN/s1K5Ea27qELfWdE1YRPH6ytKeS7SBifwmOWBGl3UzOJDiYiAtkhc0Vp
2zNKXd91JHIeHlVMzXhIJ/HUUapDREPktTEAMbTsViWJJXHC1eesCs5Iig9JlX2yXf3RdPIWTLsM
1TBOC46sZgFYgutLwFVcGVcRfkm/H5twU9xzPFL0wfB2CjEwrc6Pk7mvgFU1A1Z5TLfCwI5cCJCK
SOj+kTTANRqqnLAXzr3TlaWZcSj9zLfbASVAxY7z2P5TNGilTZ+QMNkzbQzB1K7eiuBq/qmZxQMm
+agYAqGOreDZdwJ4tRaGeJt/UKWx6I6i59Qhuqb4dquT5xOUqZ9f1w9tCkGc0DnGEqS3Y5rZkiZ/
qYgyuNHU8MexBIICHJx6hkZQ6FsnsEySa61VbZnk/kzEcgxM/sdidaLNWGNjd+GDF0kbMFlpOQvj
ENZb1hA8TiJxn/y9/t4TaWuc8sYMb3xMDPCxuk1od1eLJJVQTcDoNk5FYSyDMuvOQ9+bCUFAQhur
xrBG/ena3wuRKxFaddcBIk0xWLurOp3Ze6i1luLkLl2edB1fgWj7Z7YFQK3TjWPP7jpf+pT3BCRa
OCc+ZhJZ0FIJcQz7KJ7W28aIDuamy9r3loSXP5lJ9KnzqP01tZEUnK6DPvsZ4uoDUMtdfPspsBlC
TJkzzrTlcJ0y7ivk9JI3CqqM6+Vvj+8xeuNJ+ABEidwW2MjcqoIeZHo2iKWkMMDBEQntguiajTuH
whN9kTrrAEgNkQXvnDASt7cGkvqElscn2hlofkv2kLUaLpypWx/0Kilvo/CJhiLI6VHV/jD5F8cS
o2JQxcX7GYeMgZMXbcmvGmu9iPXtg0v928G2pzhGWL3FbTpVzdzDcjVtkyWbc/4JSFRp6afl4seJ
sNhxqZdwRF3+n62nCq0fqutv0tIUmOeGPYnATcv/XWASAQNbd93TbHc7DrbQY+FoqZsmmNUVD/Z+
DAA5fch5EC+CtTG/6iRmsCYp4cY4CO+xkWDw6cz+ureX1/DBYHXC7+ZU4QyV4ROEI2YbbMQWJ9h/
aX1Kp1OWknFepLgiO8QHt1fBE7zEyO7Rp8Ia+r7qe0DMsyS1xMehou4F9p0Jbww26UZtHd1baZ+m
wjEt18NCaGa1c+R90un1ltijMUokkUpCxX+uRAFbN0XHiZNCmKKe8rwWsDdwmapc5EX9W817oZKe
QxXHvAWjVNNWUozlYSfc9XiqVZ6qx+akQWzQtuhLdMG4Hx4JrHP7W1yvjPCaWOldILppW8xUvdLk
I7ofz/E8rSZkig17/rr+1p+tUf/p9N/WQxJvgAltojJy+RHpNg+MQ1HVLh0JwNFyWZ8N8w+RHTwE
9fSOoDHshoML6eipFukZvIimv3Pwk045cVJxFgfLLp09Tg3coOfCemWbyo6aPXogiVgTDWg0Va3U
Ci/WCKPUoDNOm2tEkrRW5meZpFcldcd94yt5vIND1Q6RB7Ni6FL6zyMi+D6qG70Wh7RsEE+8lW9b
qLmp6xaupKy/0MtXsz/eXpTxSww41lZG2OgfW1iR6XdQ/BlQJ7OwTCuEMt0mwmmgEYQxxwE33Uxz
0Pf+Jfvk0U8wtcZ6Cb8xkgHuypge8f5jxHa36aD3sKZPusU1Wi8FtMM2ka29o09Np3nwYPnpGzsJ
rBQbnHaUEcYFrxr3WkpqrMR/3e5GAPo2irFTHJMPd8aC9Ky2+s2XjLL3YW9GnHalTSFfQylSbUO1
swoPm1mtyJuFUpGlFOoHs4axWQzkEKIlZipSW4vnFsLYAeaMmydXDRfNpy9ZXbDGJDqWYiV2jcuy
wUnMmMuqJ9KxNPOrJBUnbEvNrHSQO6/lpHQB/TMShX172bhtNVaCJBsseu37dq08LFVkVQIE6CYd
lZPXvDiYndvctpc/D/duroHE/1HS3GOvn/SNaeQ+l6IhV39qaHfe8n0RzelnVRryObtHeOhLWUGK
x4pgKcj8Ci5YC6ylNxIXjbxpCm76J4Pc+qUBxy6ZgCVXctaLVtoawH5hw/mBzAll5i4tugIGiER9
TL/wBZp7nU1J9R5gZ6NpIeQJkEG2+pULG/wwwDEQ0ynmRmBqAB4jpKNa5ioQxpGTpWLHUihvhS7D
5V/dp08/Y+NSVaYmS9mQeAFXkRu9SrbqQNcbuzRfa1T+a4veLJEiocPGBRb9q1Y+z8VshvNoDj+4
ndW0gh2xRgTtpgdDnfizrXWF2FsGLVmtGd8VsVN4xrCyFEo/R7uWfMZgTWQTBbr7gbbGT3kvh3ek
dEcy/SXW560FQTzW//rg1CqA8ikKArePrGcqQwZUmg/RjZ7XyoaaZmNt/SzuF7CMfzTyIolGlbxd
fLAs7WbSXjvSrxlm9b8NXaGP4XcgMmDRseek99Tla6MDFR/dtm/gQYcTtiFB6fiGnf3hA3d5+LpL
QxM21W94RJW2kR81Yus/LUptJqqRPx+kEMBGcR4fu3rCsQz4/hGa6xia8aGqs7HklUT/0BwydQxv
DkXA7tWxUOeHG6bXGcIo92540dHyWaYK7+j39HwlUksxV9jO2HzuIlST1M87ccYJ0x0+D+qYAlwO
0Kbb8HlBAZcKGegc+VPSwiFEZssRz6MsgvVslgNZVvcVLe1elrFnPQgtdDrImOpAf5xTiUE7Kamx
f4L9SnHVqsosIu0qMTMDOx0rkrvyaOIetlu2X6tLTwqsXquyYVovXW/vz3CXCFphOrnR/ZeWNBq6
xj5YgXrOdFBovxPAJKv4Fb+jFIX635JJS4rD3UDo0QM4DRsSxnaEbjDfiRFZcjiyIM3Z4cPMSh1y
wtvOVR9TF8LTw2iexx6EMnrHLvUIGCSch1FM3qkdsMz3ueoALOmKzM//uAks0zBEJsRWxz/w0z+I
V8xHBEwnliVkY4AGaITNbh2ec7UvvitEIosBRTccrt55ptdlp77/JCNpoht+RBse48hSte3LKtd2
8Mdm9cDOV90rYf2W+NOJOSIyBw03BX8ZRMVifui7dHWrG6jXVcEUdwEELsxZnP3j5wuM0g7i1I/p
VJGyERdGPsYXMN2LM11EwIcwbTp0zN4+5mwg/3FhB3U0JpA7vQ6LVlgKXR64karzeOFwZFi70kbl
mPIDwhRzPK1mXOuMG+xHXRnFO4yHSD5g5tiHcjQ/GuzxCBgIPGXIxqJcONwiVjAiA7SpF6ziAPfL
DudzKK6kqnEKlm/Af3UVmCya1m243CPWhZAFaCFJWBk3/2zZ7Uqmmzk9CuCsXso2KmCvOruurd1p
IcuF/7TU8PVLHxPhCAfb1G5kvdeqOqxvFomaQbzmkdkjfM5ERPe3vkhxcqX3hBAv7Wr+ujyMrgNX
J7Vbd4dAl8KBw/2YBmf1uXowFSjnw+ydZHzFu59xKZU8wrMAMRZ7FkovkVZEzw8YOXwH6Kim58Ir
8Zvuyks/BbKjzZ50My71dqfkCHe+DjdXttO38WW2IvQsYV+1Kjh0OTtuymnv+Mi7jYo9JIiWW7Do
O2HZDvN2eMwPeixowNAnnxWBNCxhFTb3Bduq03sXnlP3h3mdLRaf1AWka+qv9azWgQjxrA3056bw
t1lkNMWytKTuTou4BLG16D1Iu6XYVCGogKog++ha/0qDi6fUyOMA3tEWdGQNxHeNiVmPa+NcNPSX
o99a14MqJx7pwQRJTnOC5EU7Ta2MBPspCdbtu+suOiHg83REacsSIso9FDpt8lc1O3KsLP4iWnVo
hDus0uSjpPAgNin325Pzk++3rVk9G18MZWMBnpKINti9n8R5tBi6rdbQJaMM/tE38qlize+/BArA
0afgWoLNuKRHXbT4wESw6n1rgNd8v/vr80JqgZKRWF8/MDJoad16btk+fgA2eQR7tL4ayaKI5ddE
wiyCPjsKIo1Bl5PKmc1i45qpu8WEM1MEMQc+CU6jBz2ge+sRaz6jmEKJS9ACtOsgMB2ktA/fR3/X
r9OpnQWccF8/FSqe9950dAff/Qz/ky14xsso70I3XPbSAx5yzEiPi/eqoDN+GmFS9ryBu2re8SIu
4r2bjH77rdpixN4MbH8wp4olmAhR0RWEiQCsl/+wS2Z39DnLHbsbKZ0l22B1R6SDK6L9Bhhp3qie
DTGf/PK45sDDd0Adm5+3/zZKeD2dOozgPVbqMi0KrpcS6aqlDzly2SvzyML5A5qHC0QBhvzFD03m
KF2/qoRdpHGqsR4F3zB7ba/iPBPdGgJOkTJspTUg8rRDAOD7wcWQOXqg3B5enoz2sQn/ZUC+gJNI
w0/1VQHtjAcNFAT6flIwPniXJIr5R0tot7WMqsPtkw9npEkiQwRtRHDts1+S5lMbpUbAIhMTxkwC
aeml7+PqJYrTyoWyCkmR1jTOKe/BWtXfRmiKJdY9GA+p9G44w+VcKxnpXXGwdO0DysBAXY2n9eTI
YdU5rot4BoNqW5vPZ7wI0boZRTTIR9qewboqUK+uSGXyqppuCNwSrSWcLBYH1IFcdnaS2M0HkXhR
Q3OH3tOp/Pm7g2Qh9adzabDckG7FtB7eI6J777zbciMCoZF0QAvKGXkpIP3ssUu2bGSl/M5frlaT
+QqyWSxkPETGyo4vnTidjVIrt1dTqprG8SI7jjgVbqisVtqZmDxW0cZ7EVL7bNhjI5w5yI28sbwU
T9t+iReaXRAM+QTAftiJjEf0Wc2tcFMlaOOF4pNz1C6yz6/b5c+Hkr6z8h1PN4wLULp5keq24zFn
RG87l0UGu2SSVPho/eQVYsh6aBe+n5dnEkqamfwZLGOaS+INHJzhAoL9FW76ZZt6k9xyKi64fIHd
IV4k4B/7+HMg16bx1iJZ90JLwgGxZOVD26aJY2VNfqTy2yiR2hRwFeV4opBxZfzi4vHgw6Voue4R
h+mYzDU+tZXdBUM3+v3N+FozGSeUSUH2qkMXtuuLZpjVzuFDICNubFO976KYhVmde/Xvh+1OtuuQ
aocO0OY/uNuK5IYMSYCnC2PfALxEItrfVz4uPmSbkq5YgWiaGCo19mA75Nl6q/trhuarvra87bgg
Vj91ouCH95WwKMIcuDt5L5gLuu9Itpy+rogKyNsbbA59i98gfu5RPzQOJc64s/gvxoyC+35Xh1LZ
sdtp4NpVUHVMen86UN0/5gM8goWNr6YkB7ocA3gLv3nk6KR0Fikz4AhPKAVp0ahijX8VKgRmHrkr
fdaBtQye/JoNo8D3Pt3czzZ1AaMR8/V4GNGGHeIK0dMk9UFBEJUKHqeHwiP/bG7lpYUZ8tYus44F
Wz/x4xYd2OMj56CBXc7Bng7J/HzOwkJ4f7TmnYZRwbeZ632UznB8RBJCAUenCbV5feFcqesRb/kD
csWCvCm0Du9BaktXXSay82uGUeslfNjY4luNOYrETnrLwcz6CKDhz4oxzpAplqQ5Nwx5tnQG9PXK
z2ZfcIPq8w36tx0HUeVPnvwYtpTXCEDaSlgIZZoOsVs7HYnjqWM8nsYRbhM8TUsGymIoWuP0aBX7
dAeGn/dBKeVJ+A8ASuIcFru7eGQl0f/pihccgKu560I/0Wgql2gAnXVBizfOjHIL+5cJmwkmAB0i
XCrAM1S6q7Gwr94rFHr6pXBDWdUjmlG31PgkpAvZkeMboGJhvRJxAht/29CI4tQBBQbgIzp8if91
U3vV3Bjd4hvTqVt1Zfj0b3q1sDypAyt3g3Cl02osDDLm/zXS4e8JdIAPia2N7rlhHcx1PjgzO9oi
n71rTCIWLnemtwPlOQhNMEHq+q1veEnOsgMwdkRipngcI0mT/TA/5qTYSYu1uNESULnIK68jVsfq
FHNzhXY5fwikU+URsQYP3Rw7IOR35MOaPKr40KNRrbWN50B7zC9IDtElZA6fXtxNZpf+Zx8xmhQT
MU+6HBI+BNsqwk/BTmMAVUrUp9Ujdne0JtOs1tmNhWtNsCiF2dyK4ebqQqhsUgtIOIGThwIkbqpT
B4wN849uaIrscA9na5YsiWvWlyfTohsmfycB9WyPTyb5A7xvnEDuqx37lchlFp0Y8seaJ9IceOnH
jRAnsNmwY3r1icrYn0IIAVwmOl/zTm0nFQjN52ibXEqpaH1Ug4YX8sUaZ+SS1UDEdI1T5z5kf4gw
CwsoMVrfteckMkZPBgAzCgYssPJzgy/bKgBMVfWNUHaaJMmHHxvs1KkuSHMBlDMe1rPw3rL0o4sB
52gv1iDv8Km3P2iwIfvsYAkRXDeZGLTr6z2jMT6zJvXycgJMP/xJvy4RgXRa4U3MI+X3HKj6uQFn
j3IDuHkfHzQoivYXufaafbFFSIaaukkJr+GfjBztdwKkxBt1eLuYDVFhM38Qj2zD1BWPyax+MJzf
qs4f6aTaKY5qWHzidk6nPErZfmkV/ZlnsMISGeYJhyBoLB12L1r18gHPSPsJaT2Iw9GCYnNTg78Z
3hukhLfbbUlfy0NINS9GejJAPp89uw786C/2PDIzKf6hut63SyZxQ87/iGQLvDAAihDvw97/T0Lm
02MqJ4ux5fHqGGbcbv/hfArPhe5nxg4AC1E7w8c1qIOZDciKyAuN3TZqPUEvTsJj6zXvH1n9xKI/
DvQuNebZGE6ZvtVLgNUUeBc11K8CTWdhwp2F+G/JvWmmyOXDtjb/C8MS1EQivEQbcFwvzoszQO/l
PfHKdD6LPLwx8X7xwTboofX1aGBb5PSUq0GGoY2gduIZELdPERjuwdGRwVYZrhXvx29LSviAKypu
qGKkh2vsrn05qwpiLw8xqAaSwrZUpTPHI9XwbpcTDATXxU7rJRCCEJqfJcL1shyfb4PP9/uKl3CW
1EU8yZvmqzBJuQGsziW09oL1+mrbt6iNAwAXBquo8ble9gMNHyzqvelVrfi3lomiwZ/BYA3Axcs/
F/1qRNn7Bsf3emXmz0cmHbFAiOCqX9NEoPRit86rm332DhSbOLhfCXLoQtk6+QueAn04xmK8ZLSM
qUvjbdWns5Q78+xGvALhRoqJ5xCeR2E4shrNQixUBmrZHgYPHpMten7Sa1Qrr26bPzpLZdiR5UBT
mz8U7kmspMqcFRqDZipxt4QR9luGPgzq5PQHfu0fMNbZDqI5S12cgsRn11uUff+laLqSwgg/Cm9K
a+80YmomCMsqH90e4WSTM/lcpDz/tdE5EA70eMGbiSHp1VxjyduxtExRJSntKuICijBuleUQLRlM
tbFocbRa3yXpBPNdhbXjekY/GQ3OjhK3goqoaPNGUjgsyFJA5+TLr8Nn+FCIQj1PPjwXCJTlqHmZ
FlZGZcMHBjqSses2OSMss/vmBFZ8We8J1ZZriAtebIvcJ8eLQU0RwwgBpLNWwmyYjHHoqDzvAUDO
NxYON2lvq4qurYrICdF0D/66251x64z1CqqJHXqpRck9ZXxuf8eZ/EviDxu23G2FJmOSIZImexV1
5PwFvkpNnehhtijHHWHWa3Z6RbX/dH/dToihnuFHELr25BEhvLlNpqmj4AeVVPJMUdsdRJV4kNVP
gXlJuguoHgVNLkAJbHKycBAcYjuPA6F/AGhzPiO9Tvj9esJ/ERMe8BkFjrVC5RlILQAbX3RNgQ9f
lsK+5fUqbeiTCDZnVm9LHcD3DtT7b+hZJ3FjrNcPsdz1iJn9QoWdVUeMbJUMluTHG1NYxbxGDhBT
lWRTofgcmyw3XuXwfZKiZzfLU06UwFWZYTZEfxM43fqdCfKvRsc2Be+ZdNtC0+/6wPn1jZtkbdVj
u6DupMKZEXmbbn1ddU9f89Z4bTiopfYmAYKm5vmVVkYaMScRf62NAvALGlWUiPISuChpeJ827Bjh
5BlW5NBtvqV1hcyaOKnx4trn71hv4knkiRpdoK/dmAdAVwJSjkXrzCAjJx/T6z0tHWoBDhUMJm0w
cdtIfmdHlcuIMDy81b0iOm3eE3OHZtB9kvJGb1jCQ5wolqTOMU2bSBIwTwV+DsPGFGCyzJphjlDB
Fcf+pK+HXo3V39ugsTGQVp7noina19jpMoTRXcvgqE6pl2+Os9d5/OgzlWtPpooOPdREYZmkI4Zl
nFY5VGwDUh1/B4GG7YtXn/tg8tK8YX/+9DO4TJGkDk8lKH9eljyO5oa1Ysci0774LzYsvPETyicv
2ozU22ZtzxQuN8P4iRQl9RRcLV9DJ+PUDmdQoeTaBpc+flI11oc8BRioAUE5b49K3r2fJYSnkdcA
Kd8EY7WpQSRmsIUqyLsp3nVd4w6w3z6j/+8kG8LrDPZhrnnJ//cNKS8ZCEg0q7rvwrKzGSNZPKNW
uGLOpz0V2egQ2EONe+/qZp4QIW0LAzwpQWb29hoYhPZubhr7Y5qGesHXZm4mNyynbgWCD3CRv5L0
vr63251N4r1nT9Ze244xbQ6QDWodswi9T97vuV7iL2cHPw6rYSSMWV8jF0KmNsoWKBmnwVwabEJN
PpffZd39paXAg7z0ToP7KZtPmD8ynn8IsvsHWQa0l+bHRXcu6sSLZLXSJ8T3cHz1GWpZO8NH4M9k
+oGt8XxzJdPksc/IQ2bqLgobkB8DjmGbn5IuUWKjElRDJKAyr/HY6v2a3mqudsoh+2GWwAhF26ux
uvrwYfqlTfGd+RsG8+34xdp4E/i2q8S8sWClLGDIbmRs2Y0+15K3a20HZ8ahFIkEk9vUbM0wcEEC
VneH9GmD4IcYbDs0VQHmO3mquS0CPXwJS+eEv+6At55p3NnkPrG8fjuvPQgyGbnA52E7plqh97pi
jqgzlczKYiSLltxNx/RWTnPu5wMIkfyabEghrzMln8hNcHml8rsNx5TmBX691jGYJZ9d2GDQz/4l
1rROvnZT/Ce5BgJjItPI/9bzjyudWgSHFIVtIiv26qbI+z4ETeZ60RI13A1/e1og2L5yBw2YihNa
7WDmGRzmi2Y0DgneEYvxjMfFL38lkoK0MV9egSWWdCGerXuO0G1gbN+IcSQ0zt3XqmAJLTkqYd4+
5xEGJSWmVysvNNULh0jQ0UklluV/AzY6Q7vco3KQKS+ownBbrSd+rnLQpcvKOjLLcBNF+XAtASUp
22uYN4ipcMjhgAsKHQ2MIJb/DHy1wkZcNU8gNh4VJ/q+kdEoqH9U1pnWJvb3fIGVfurN55y9MMMJ
aL4MEFxVKqWSsJEZQnz2Xo6rMKA4Q58ighc8fHJPRZF0wkKeGhfSvLdQ/TWbpFPM4ZGdQsA5VTY/
Nk0QxMoSxLx4HH3bFIBr892+rtLOIhPzzpz/nzZ0cm3TrMgRx5piil9U4n0zOADQiqrv+ayIIo0f
iN43/1olD12wJ009JK+8xB6Attnsc2QjG3FiRDDrcMxs3Sg33WTWQyIEw2E1vDwc/ca+Kk7tEadk
Z87YAHNOko8eVA8ulj4iSk8l5NE7jFEisuWThHVY4bqZu7CXWN6LUznR3l7ycnKvo91S8MpgM84Z
eXY7Gk6f9iWOL8Cg7epr3LZPeyNvDr83ZFmou8zyoMYiMKPKv4xMrPz1Iyv+LlHx1YFRj70mL4nK
cg8x7UHXqaQxyjKfMgvkvExXrXv7RKrMzUaQbAPK6Gt8KiBMZnjrWTxA72jJByTaWmUdwkG271gD
BkN1jg0JKnMPctxKv0voJTgjCtqNNtNEAHNi8Z5JbtrlqAommpxT/l0Oilo7+r+IzYzVkt7HFbo8
yxtz9SmplisEueUGaBcTXHKcfX6OigQcblQhiV4RemQbBcQVdKiRep1kCxsv2BC1t5tUZOz4iVDl
s4U/prwFtabUKK3MAtGeBecUT1ztK0EkIl34vXsTMNKWEHz+RSO2m6AnBYlN3soL8uUAhpKHRR2G
CIXAh6l55S/o8+3MBMfG+BQroRLsVSaYTlQL2qXTAUoI8b5T78Br+NIbQCV84ryllUAuLQ7STwM7
X54MuD3IWWMlIZ6HKqM99ArnSwHrgSgz/6JCK7DWUgunAfEaae+jqahZu5EHGdpJdSMWssgfUVCQ
2iNIJFVKyU5pzhpIXs6XZDd3zMNO1wuEuuoG3QjEoYLyLREeftvCq8k2fCG/SzNohiXw9m9k5jcj
UR4hitEFXCrfMOaXWbhlNFFfSWFnSp5ug9eMtKP2h4RwXMZBpx2VvI4qkbNtqwTIiESHyrD2O6RU
XQPOWjejDOZzR5ZlJeUMVdIznEZXW9qsMSEVjIi1GkQsKNfV+gbDeOYFVP5OI9H/NQU1nNOaxFPH
ILUT5vylywpjfvxaPpKYP664qqLQ2Td0RTWtJBxQYn0IL2+62kzFubvg9UZzsicL6k0ucsJrJ03S
DIteSxkmrej+BN0oY55CSR6QuO61pM698QSoKH+KlJC8h+3K/QailzupG+CNLYU+5w/Db4penlSq
+d19KKIaUH2ubA6c5X0xIU7zMSp30V/b09dsJMBufxrTNVUAA/nryfXKJyaHtAHQBPds7OJar/Dt
ZHd7Pw1JueO4p8CcpK705zvPTA+4v0VT3+MXYgJxfhw2DPQ8Yvc2tH99ZrgoHjERO+0jy9LMo58Z
0rw1dyZ5oV4I358Pmix8tZAnFjHK9WphhRMBgTgs3nq76M5kCKTxAajNg8Gj1oMQUTQrSZjhPWmc
e7Qh1ITRCk+jqV8HhE41gS08dF5ftIGwlGvD+VdQGmlsRoiSZQlWTch/WQP3LDI3ghkQDh3uEpnX
sbu5F+YVWGYtE4fE94m1NYaxSoNFjD2Z61dtCPh/Vgb2H0cE+BPA2E2cCeIRXGgllRglVIl4yNCW
EygQnVPMjnRx4oFMAznOXJDK1XPVDQdjJYhIPDbdIJrKElXlwKMMTpbNbBgOYIcVVFEPbK7oYCeO
K1wT9MbgpFXI9ehi0YavCxCPNNoRt0RXNw2LVsHXEdoHtP2NUOP6POjl8M/81ODr0STptErKKuXf
erwQhUx3hMHUAvwpm2ka+ikWkadLZ6WoxuosafayDVUCUROKa7zlKYN+VIEsFGPo4TcoSSIbFGUu
QoTDQPhZpRBVwO/205YhRR/E/BF/G+XPqx/YuGgsza/h2feOZVF7AfzLWqqwiWJZmTKvZovIyvme
TrFezuvhvTTX66AVCcvmMKPbEqeXZTeH/wbv287dC5762idlaQlVoI5DoT7VqFLY2EUXgMNaXWY4
Fczkj44j3TNXjBl0aIxzFnBa5qt17zcte7xBgxff+ibKLp1JON3jRDyd1ydq+rngRSaFWtl3Teu9
zs6h8q7yYP9y2Cl/jhpT+wJJ0VMAvWcZvqGCfAliETq1/Zs4PkOsb/rFpQ4Kg1i6Me+b/x6zT8ET
wJIBgk0ti00OlwjIbyylq3Q65q0iT2rqO1yZqlxxhYKXj8i+lGsGatD+fCmOrV2GVlG11/53Ca9X
lrU+qElJh7ibejOH2UIxr0t1NikazGHfIO+eF+UAykXvwiCEWxS4eiiWOXLVBIdCxjQf+X6gY0Dl
CRJf4n82VOXsWjAQbNQ3pNtSm29ucJHPBqiP1d/ZEUk5506vTnjTwu2XZGpyV0XyxmfhXD6RDxPQ
GHvtBzl0nmh+1LVyXR6OLWf4vwfTnusRUQQ0YHtnhllm4BUsn5LTv/OW81fwo+QAW7q3duQpFakB
32SaDtPfJL+4pGnWyEPmvQxAmA/3Opk7sfzQ8hZEGuVJ+O1ooXqx5SoMKKtuwPTnFq1GhjVDoAcL
jghAfiqYxDxBZmxz2sRUjENrlpUaFayM5CuNHceDp4Xfsi+fHYf/07aCqENUMyQ5bn2bJOtj33Ot
Z2qoN0WOSPpo6J0UxuCDzmoxaOZRv/ycVU9cpgAHziwsBW161nRHMdLfGnhOyRx4QurFfpUsLtHU
PXXhGgOqBo5Ik0TBEyDoi7FFgVd2Aqol4z/sh3r3MQOpEG49yBYOhNVHW+KIsI1ul60YJFzaIrXK
RDCP5X8m6b7TkP/rlw2vCQIHudruUra8x/L37inGr40BqjbEcmCn/TiF/x4KiapLVOT5Y9pstCKs
+lPgXgxQaOQF2J20+Yv/xx9HAC+E7V0TJVJhXsRPK4noZ/RdKd/5Audd83UEp55PHQMhq75obdk6
tlMZXSCY2EAo+ZLBQmFEG58kCm/s62/izRVN/3BW88JjLZqPwJ7aBiDXv7lyR7fdqf/cQCfSakxW
NUQk4Kgly7tTrqF5ACRK+H4wH376hyNHhemEXS6N85pruu4jHqceCURmL6Sfg9J26FT+xfLiSW3g
kyZZ4sWvDSI2/0o3ZaSTI253XQr7qZ3ftUFiUf2WcQGo11A0wEeov7FOLdODmdAa3IfQIwi8XeOS
TpzsRKVOSamzhbEb3UOmNtffCdEOFRr6hhBjEqjJVMHfaZPaLVqgVN8JaXnuY5RnBeaQK8Xu7m2D
iGmXt7cqBXl0Xg6srXDk+4jDUv8iGS6fZ9Le7JfI+73BYZebc2t5rcyxMo1S7DGKM3Uan+hZfZrq
+39PB6QGlF1PKM10qfFrkZE0v7nQcHqBPLCr4iZHHbUPkXYNh6/91qpAjoHzi0fqDgmiHdC3KZ7g
T8PqZMqKc+3/UC8k7W3LPXGmWJgQDtCnwRdxC1oVCxbxGzRywGLgtt6D2HOJX8viL1cv7kyIZuxm
0jcyk319gAr5sgc5LlmDJA2y0gOI3lesRMHDZHcRRck9KHMEdHYbKFBH7I3wEKL/QWzfqpwdyYQJ
FOeyDuE5F1noIoyYKofSpHaZOQ1M1DKumAH3QggMtP1TFnWnSNU+gPmh0QA8748LbiVW5Fpgijra
shKOy4T1SgBs7M5jDoghrufk+wANd0gfhZ+PTEehg5F+SO4AR9H0FrClxO/7ymhzr+oy/eFGw2Vj
hUOPxRtQGSsNZWiAAVU2vpGXUlP6rkriOYQPr7oFO2A3AOjmlZhdGeOaf4Vo2A7+jniaI3I0dMje
xXXKhqzjWhdmdgaRxRZdoopGrOq8DhbK5ZMG0LRiHxnb7jL4y0RYdgyzk978LFoReGbsBHbP/ZUw
khrmpnsNReZw21yxRQ/hYD4Brl2iWxVCvLLx3PmXr/vZFYn3bms33Cbg9QvPQsuwbUgxzspeL6R2
1sXr4/dJiR+Erc+5WCmyQ3W2olxICapEtrbB2vzA+0zgvlV9P4rjOH+t66UtOfYyd0MSoWv1h+3e
itcIwRVxufcwpwNK4rjeIEaQRjELy4NC/QxUqNKQdo8zeFA0mjc0vG0QL10NBQLlCU4Onu504OaF
5M72/o7d8fu/+X9ggCuXBAxTkghEDLlwy7rW4HaN9R4iAC1Yp8kZbGB/tljCDBmxI0m2aiAHplyL
hsXOhNKTQAXvaLhpcUXWkBryGku2PodCd1+dNJkI5iHBaSRxJO6R/yVx2dwEWy77pe6LxriZLjMJ
dWvMfOmmQGkkK23jcWvX6Y4Rrn9cKaR9UGHz1sAPXXJX7kkyhpRGjHf0iV/cZEM+h8QYN5ddQ4bt
+tuSBVQc1w6ABY8cP06ib0pjmuyA9yA8fMqM4vcDBoYiHtW5L/dusUL1tPncRtzdsLWCJGcSVf70
wQf5elPQLRuJCa1ZpJTUol/C6HxfflFTOHz7bLZJYKTITc0+UUP3fu1OI3Nkco6WD+lmSDRZiHuI
rgLM/x3iR4Hx9KeyFRVxxF8bAbwkQVktPZeNjJelevJBfdHO2IaC4Px85iyOYLe9SGQ467Hvny0B
3K6hJ1pjfrx16a43/CrOCopQ7nVR5n9NtvbYHq00QvMHoO3m05eLPw2nRzevfzgfoQje4IuOUwSK
lblsrtD6hnPUY+ERlM8lIMgvWBu8o3aPhqkBwgubzxZTLBFlDo01jJoB61xlikkFshzp9Pa+plnJ
1pev1ii8KhDTARYim95S0izpMUgary/3RPMr8QK2a+lnmY9i+TCdBfTnBydRs85CAYX0y1cD35gA
I5QcQM97ZZNYd+vvH9R3aQgm5AAxDaMrvqsw5BWsZP0iDhQFrajxFJNMIqb5/hLyzqeocNTc121L
u0SMMW3YlYVhSzR3qQ6tmsXoZSPQObi+yNHaD325m8n1LSvCd8mtF/VyIGoz1Qxm5Jzxl5AK09Og
UTnM1kl4nXbk3QRHUzCPqc/B2OnpS7kUpNuzBeWCbrYRHTP7UTkTe0m/Vu5xeTgTRY2in2c63fXM
C5wrv2+97G64kYmvGbfwvN5iBNdWXVl1rRm4D2jVmw6Qcsg/114YGhKHaZR1ILfMebukXfX8YI6c
+YsErySvlOda3usY71ZDg6Rqpu9McIwEHgcJAzVUwLrxT0TujehZeEvcLRb1IHEy0edCvC11tKt0
kHEO2SY5TGDHqkwK7wqmj4/CA2dKFoxLqU16nXJQyeCm8icapLHdiZlagFpAcgglrMnvhwlax6Nc
vh0OGk4crWq9kUohlkRseYVm2AsWiGph+I/31Q17NGcdiKkE0wEI6FX+cwLHz520nyPDJpghD9hB
M7of63RTAqNnTPHzMK6pZyDHkAath4KmY/aew/0nq5s/InRYrIOnLrF8duh9MUlNFBvVOh/ZikWE
B8hm+K9ufKuMOGOoHsllPsEzaS8KUXTHzTd2kIloalQkAmNHY/H1ldGnG0bIC+unmAZkEhcKaF9F
DjqDubLKX/vebNH/McWp/mt8cShZ9cEELmfIIpxWinF4vJHOuLJMKNhkRtF4CZwcmZaibr/k4u/p
ifY/ppAJUhGBzz/4ZpqNKfuDvUM01u6TgdtUWM/0R6a8/ifY8zTdIMgsyyjqHPfyfiGDM0YDhM/6
Xk9puDgLtEov8+cdFpwqBxLwdHDbI7HDKbyoj0zDpPO3Ta328rzvbvuWngicX7tHJq+dI65g39Lu
m7mVyZ73gMA5bbugzCDZdWpazR53pS3PkzZDk/wjxdsJoUGjT0dhAfya0hsoFhRA48KQNNu0FtPX
WOZIsXVTDue0lJCD7iKdPg0FvNzN063D1hVTSKEFMyBIT9WfzTAMN1g+eEFgJCZ2UVZ6tQDEmyfm
pvNwisi4TR6dr/cgdBPDSkCbRbkterHhn/Kfdmo6PQF27/aGNCFAfhor+Oyj5FMqiRvya4ila1BU
Js7HQzNSW4oDipMvMPoGVNOou7IprsJKHZPvH+2aJh9BzjfB0CwK6OP6kMs1z6V5ZpxS2/sp9D7K
IS+T5JlCPFBhujbVnTisRvAXCySD8QcK+3JQGb3U3SmzsQDAnveDVh9sZKUNo9Hb/Lyz0sMSYz5b
vlXdhdjC0+dkpeONukjJIXa3kVaOVXt3inngz3X/BMW9KsZXLSV3WXVAthPPkUAXSsYJZYPjnrXG
9bw1WpfTSXuOSm65wRT6ILpv0DZpI1Qw9eCWdsgAAX6SW09RNXAPJ6H2RxZrmcozo5FgCVFNtI6q
6yWG85hFm4DU1Kx9DxM6hA/By5UVAvCnM4pweRzbEuBwTiXH9Gq5BnJsI9RIvkkSqlxWxSGYAD93
YTVXp9xif5mBleYC3yomOiDBKz+ewPRbtAl95LV5E2PbKUwySwyjZBNPCu9cogujy0z+awFBrKPE
oU2y1MVqm2xE2VtALQ8MnS6voQits+9v5Ztk6zCifrs5ryEnFrz6FsSbU6RSxi7z1rnBmHoXS8wt
VZFCJH74Prk3xdrddcB80wZ0J2qsIxK1Z5WDUdR5UEVsLqo0uTTKiiKHHnhGWNxyRcda+cqkGs9M
Hh1LJZa+VtBlDL2XLW3ATkM78Mi7j/piK2/Etv8wR3Bmv+Ozlx9HF/GYZvqn73zsByCVTEjdPmdB
l3W3OI7PCanGweaQK2kDriXT4dU2sHT8LnfebRH2BoxOo4jZ/GKIt8Vp6D6oTS0DZ0wu5elbPsUY
D87gweddP3It/4nuj588UqbkLbt0vjKzT1Qg2WjrCr9r9EZrFomlyb46pggiKXcwXrJ6RiA6iue8
Lwm9VwvjlN0Db3ZNx+Z8yQcnn++UFw5lkqvRdWq+IO5h0tIQr3FxOnvwNnc18Y878V3qy1zMTBt4
npUT2ld2oPzha5CqCfLoTC1bVGCEm4gz4e/s/ps0oWhrBURXeFSozWQAK7g0ZRec8ozc6UcQsZJY
t0VSN7n6bB6VPxcn9zJW/60TBLaHAGlsnQ0oyGKMgi3djwh+FBGeuv05XWUbGGY4+DRiN4w4m9WS
LASpdSGP+9+c+F9lKnT3xSnKQCn7T1WnHvKyM2IhBTGQs3dZs+ausJQ3rZkmjP3+dC+6ajAqT847
oPS5M5roju5etgLD8cRL162DsTGFJpfzW3I90Qn7jNkrEBqILbA++zqT8Q8L2T2dbfBigvm4MYcP
zJXnpIIsSVqP9dBi5dQgMoxijHn+rG8Gob4YroY2J+hEXPVQjtwPEdVLwnrW8tK7I4QsJ7IR45to
SolL5jqnEb0L9GrLwR4UXwEnsHa+d8Y+Nk7+76XD/URqUJxKqjCO/hh+QmjP/JY6VKqc/YQJCUzL
f3VL/NoovzNGTSpwUYp2DEI4viTz3YnuopfIfRhJPLB3DZVzdiJq2a+nbI0YuSzuT/cPZR8finT3
/At0QRBsBwjhSy2h7IsIDqdbE9hw+1Gez7qvbimtRwJdU0LQRs9DJrGHRqNf91eLZXYap9fgd6Eb
rzxl8/9+r+9y1pLXn3CI7KsMrjmPVp6TSfn/gKznkRozvAYfz27nhv/vuAUF+joKeihSa/F5scsz
lWPvADi0wjseGfbsn6ntN42YjkwenJkwS3h7+zS4XBReg7+eZZAWjRkNx4Ei4hr+Q0vEnrlQyfOZ
Wa779YOL7Ouzwc2e/GcNZZ4ZVIMtz6I+m3MZ9NqVXOI3AClqjSW0lrVQFwHMudMwcnh8122tBOjV
HZYoNKBihZNxWQkWiPQsK2bfFRq8WMo4ScbWdFHfnJWq00duOB+HBU9XuAhLXpVmhKry+eUWy/qe
63NePjjTp58f97Si8feo/003v7Lybmk4JL3Jw4to1iL0fNQ6HoG61mXEeM9B7Sv12HE4I+4S1x84
3bGAvrX8VuHStFNagVxeLuGoE0nKwAjpyAknz1VBuC+a+N7sjj6nKcWjWQ5gvCqlqHsLfAHwdFs6
GR+caneRAW7DY/akngW+KiNxDm5LLT4QL7HgRxxPwD2KxxV5kmagzxGidxEbiiFwyj0PdIUZ9U9N
MW1HUAEfiOYbuPXpxfW8tXtmcApe3Bbl8WkN6tFoYDy9poNYjZnT8v17Pk6zSptR/fS56EbHbNZm
Fr67otTR52iSWn8KFqbvMEqzrIDy0g/sBSDagRYHBgq11NbtZbVBmXUd27DM6+v6IR55gK3f9oVc
Rk7rh1H/BebHSpo1QnbufTR4Q3PdLTEAKpwZYr68bcPo5Gqqcxqy80DQTTTDdfNI4P7CtB40Jg8L
bZLkHc6FPhIHubY/vs/kuPMiq+RRWKngC59ssqbDT1q3Uu+D7BuAgoqVIwumsepWjOJRxwq37vhO
Zfc06oMEt4siSwRRBXrzGrEmFHfGlkd92sMqsVnU1v2ocn0du07sGHJ2uKvL2YG11VCT0S51WyVg
QBFn4Y6BIP5YDanIspPeVsV3vxfaUsqzGdDr5ikKBq7YrkoNRKTaMWxBinkE+Y3AASkf94QvS+dk
UqWkvUVCLsoBqrpJ/JZsFjAd3nQ+EoB3LyBvA06f7pXc4385zw9nE4WhWD3aUpTNWhovWyOIAYpv
nVuJBqvfX4aoaSghEytnedP59j6mEyivemzz8DzaYNdvggoAeNMt6agfs9mgFPTzvgOZUWvDmaZQ
JH7WrikHAtUV/ar5/oPLwZTZCAh3eY5r1ZDaPmYYOz8Wrw/AR39T3kS4rr074+OwyE1ISpQMCT5X
rYPfclOU/hotkzRzTSfNGGxen6dvt1Rx44aALxSKqgr8QEBybkl7tC4TU01dALka4che2IGb8ozH
DKO9f2Qpj1L+ZOzS7+2gvYjZnljvr/PWWtVMXxuDWIhJIe43dpkk1D8lvMAZWPCecDQpdar0DaOA
yuLtrrrd47NZAw7+fUhCfaTFo5Fsug7chImHEKD/EhRpnodjmMkKteeNzKJ8xPFW9ob82EgjnfRM
qTqWRM0IMQOqOWEglnrBAODCIz1vNtAoBKowq081P8iXCpegf5LAeYAn8uiBHxSv4OXWvIJQaiqH
/BlEKM8rsBj4jgBb3gtfMS3cjUkE33oD3wv/X6Dlrsn8EE7rjB9HQK1vQLkH6fmB7RUkWcV8ilXq
irhc/7f2hnn5DzY6du/Q9hGk9Wh66LuAsXIDntZZBd4HN7bKoYwGxIPn3OlgWmGvSz/OlJiToijG
97FinmNQ2io1qHWBM8/B4DOQL1CGdm8eZNN9jHW7r3fOg7kVA2Qb7w9JI8AUp9QrPHQfogE3esYO
3F+TMyB5jzHqmMdmtcMRXlEXGxTzdkhANxa5vcXAspO4LtdRVZzKmiRH4cihh5C+GdSLbOlUq8LN
c4daeb2bCRe5/Wtn+xz3EOQBNfI4TDF4/ujtytBIEwKXSrV9KqUVV0SnLJ2lk5TOFdMgVWYEZx8J
fhYeUwBnq1fbYRzb8T0/8soKtnEUPvvBSIxcUVQfoTPwnWwPVb0lx4KSbPchZNGJPePOocBR1SKB
J/G5JlgI52OS0WcYz2zSyB1edLArDaPDeJgaM4iDZIKP1NNtAB0f0Ca74KnsRSdlU8mA0twy6kl4
0AnmAWM9U80r3cNSJe1fmajar1FRszhDt3Q7FYqvOETyfcWrK7u25oC+DyeWewIMRiZfjX1QbQjJ
e097xM2ohTJS7CcVzhykDaxeoqdIxx44eZ+TojWRrXdsTK/DWrGDzmxuizk887jCdULW4m2DsbVy
ZCgXFSZj7CX8HZWEayw70r9+Sv352cf5P118wiXzON+dWiwomr+m5xKQsXdYecYp7jUUZuGSCfAG
WF3I3Je41DVOOUE09dbusWPQXWlkB5Da/vFxXdcBIuCRxUM9k1wJWEBwHAp98ak3B5coQ5R0rX5t
fEIZ7uu8C63myAyBNx5KkmXTsxHtUSN7At8wOMPz2gdr2H6w6g3BwkmUvblgTx8fWGzhBU65KZmY
hifLO4Y2G8ZejTvqg8cTky1JUPkRbfk45zNrLGuWe6WeNbrJ1Vj+kZm5xbJogZprZSteT/4hWjZs
r8LTfefLYSPO6tV+5eEwWnW/3S6mHq4+BRx1/+DDDYeuK7kpc0hjTgkOFsQD5e+yxPNkUcr8cLNj
O2K3GjziadX1QIVJ8NbZvCrTC6G1kugKIF15pEm377q8LVWf0MmcNgNQFcelBlOLHHiTg2eKE2Nb
l5dzvYzZ6bjWZx5P17WADzWAvHcDF+ENJW4+H2pj2LaO3YcDTpKaZpzEsr9nmoeX8v5EdGBkq9zq
Y6BXXEkIUS9JMvuKKCaYWiD37G1gJsdIFjFaCQ1XYo+28VaYG8eokqnXW44/lBNcX/zFStEPwcha
Yietwa6ouER2zY/1Vsgq7gtQYqXEErETB6zi26fMZFTZSsbZUUPNtbCrPgYczjvLKfnkz6Mb1rCU
bHJHbz6TLMQnBWeMnLuRCxC9uPciedirXKcPJlnddFYlUhtTkXGWLzpgxi0eZM8/n4lw7tNqbmwE
39W48X7HWXkdIzrAofFQ551dhrptaXBgv2wR9QjX4X+z6zf3bs2d8nKKBsFd3KXJ4LGDs2O7b9Ex
IYO7g0DsQxv1pnvPdVtfIIbTjw4MvE6tdHZIFOjToYSZsmgSY7nTyiANLTvhNpWxiFOB4LrWT6gn
mTYA8uMzONEgJuoEYGmpDR0NAV0SXR9uh2d2uxZNtTGpSft/V+1VIzeJf9aauiTlUfeHZaT2UsSm
t0/M2nZKeyh2aAxy9PkMNN1Vme9/91nBgb3D882/YAKVVib/h2PLBMHTEEHToqSsDs+eEWfoBIiI
7SZ+GEQfe1qdsXzD6mZM8rOqoOClxLYrEt2kJ7MMfQtOD10BIVi4aIEfzqzLRPjdKDUPDe/n6vGr
6T8Q/A+vpVcMprHcBZuRX9ACW4t9MXzdiRkWEBSVMhc/Nv2nAL0dMLtI3+A6VJSioGK83xxSreA8
tynQxOOdRIj8WJLlMJiUHyinY5VYJLx9f6SAvi1vpaLVIOW9kyX5Rt8JpmZi+VHkr23M8cpQ1P4a
5lEL8cs2LJvvQ3c5KXPXP/qfwYfbizC8Dh6qS23oYpbE6w6TbX/M2uCTOYZFH6HPNHtismrNeRzW
IsmC02ZOfmF687TSr7fHlNmSYpyJ13YXXK43iiD3FFS8obTceqqnjJMSvpx3Md3GGjQDXKIxvZkC
AlT97uP6ACE78Tasf3dWNtX9gVKztZIQZbZ4cd0hN5kxZafB3SIrscvldLvRGocaFDmbwEdvmKY9
9zxqq4QeqyDfjRiBNqM2o58sZvtBL5hGu1WHV6+/vHnVACpLJ5w4J3nKRy6qV8KdvqJWZM6PlNTh
q6QtD75lnb45S4Xc47MkXii6XphOsJYaprs4sVKLL7398A5/BCQ9HflgSotXd++t85QipBUdmSy6
GjJYJYNKCI6wKPV6dAtUUy3JsIvGpJXJrwoBatzlx2DRvogwJ0M8MKzftNFnH8vKKBfGkv5JyLyB
T1aw6jMHlHgMBFHkyhCiuaXnG2XQCODUxe1u40cQJcp9DR4w1kKJ8VQPouyB0Y42pCVYIkorkElO
R03oJD9rA6y1tNVVsVOu0U8QB7tm4yrxDjngcFG/IpwvgpW5UE+WFMG1CL4C2HIWYMuldfPJKdvC
+KIIpeJv0yg2FY3jaycGRPzN37h668GgcdK+WUlCxlzB0c29fl4MPSQmbIlhDS1cNUH1oH/MN/Ou
xfjU3FDswj3PhBOf9McKJo3xwRFL9RiKpooDbBKEmYYL3LC2swoOaynIZCSnv4emXu+9BqN8Cg6a
pmhA/ZohbRogOYYzLVoE6yM4qQH9E+5YQ88HkXaIwHXQHUDabLIfV2Ilkjj4U+rjObWKLpX40z6H
Kzlld1UJ8QAaEr2YThVlo023Glkg3GOjfBY0H0y/dySLBS+mHvwUW1D5P7NT7KiqD1imjgaAOobU
umK+nbFDlE9Vvq3rRCnWsBo7jHzFK6RPmm2N/tNxn8SmsVR16gM9JJ/ePb5+7KfCKqmPseoFZ6jQ
y0SnvNSMiCVmziiDe/Scm9K/30ObhjQbWsdKXuodwoQwmyCETE6et8wjAqGJJGwFq8ot5OH12aC4
BNH4XrO67u9vG79/MxNh1ivQFzdNOrEMVRe8u5nTDwi8NB5F6STqVHH/UC9RlXdgU8aHn6ZVElRr
IiQ4fdwda4o+6qMXyFhijFrL3tOW/W2exAnI6SM6U+hQOz6vUVBt49cYhYUI9lXHEJrUkYZMFiBi
tUBqyEnJJ32zc1dgAOYodg1ahreVKxlrRed6bx/hm2+kIM+yUVMwBWZlneYby7VCU6Pq/oN/xHnm
Ac2yyRKGnwOfEb873t+iZFPqwYO2wgi6YOh4o3XVBjYBt1PbWw901eGvabWELpulwYreFMfeFeln
sj0bnGrEQ+gi0HNEnCjZMZqKYb2ALquxK7orQERx7bh1GZA22Y+FHak5DYZyG8NGxRm8MGwWyiJM
6jkwnkno220kLp9AcoCGN8wjTQEsBEbScK8l23z0OIyhRkvvMYiC0M4AZL775Oblga55inwCGHkW
hhbbYxINVwyEfK3o8aI0K7OaDlzmpGrQeulDp++0//JFEJc8pu1uOmzEPZQQHuEnCHWMts4koAQt
J0xeyiwIdsZrr28IEMKt7nsYsV2xKJWCml8IpWhj9v5UoUhwxITv8X7rhIGqwLW1Aj+Tm7a1G8gD
QMNQc7NYXPCPVhPQUqmpndkT2J/Rkhj62J4q4nXRVivLrVLOR9fsQDXQMR3EINNYccacZLQV9TdU
iHUZw6A/LhNNv6LHznCko9o/b2WyR2okBlnBZS1d3Hy5e46IGNQ6CiLbqEOXcoMsUoofwnkpYh+3
VQMaOZeEr9Xt5wCqMcHwk3gGqzMX2YpqXAfBPca4g4Esvij/LexUhnoRWxXtuv71of2L2jw6Hjvu
s0Gd0knLDG9DgIGy8yPBQr15SdPUciFRfoR6+Rmsx/RMqXssfLSEGKbgq8FZ05teaGt5upPf4INP
7MZYMlSpsTwnGrKkctSihQa9kw15ZiloNyCtJmY9V0hJqIH/3r1BhRhNbmyD82Y0iiHuR67yj4Dd
g1tKXM2WJ/lm0ejN0jxr4MTxExg/C+icXgq6VMXdWMDsTB+ZB2j5h3+M3ATr3w+n5hh987GE8vjb
lN/uAzVv4kU4hG2lJIWvTnbuUUF7rLNfYPvMMjmP84kLR5pBwfZcv/W6dD6N3a/YdRQ6q9dqQ95r
RiC5sYwLUYoObwTpGm7s2/eK2nNprVC9qwLufDmHc0V0fQ/M/sThMBAK41Ytekr53A2mVoR1kWH9
tRV9+u4pPnmwv/3vbyZHX28SLZGqw5jLPWM5Ffv2+Z9CSsEQsRnubKQ09hfWC6o+pVgwG2/1RokO
aKhDgGxB3XDPxLL2UoTE26zhw9aH+K6kriBT9svnDziFX7L5oizTDNC7DQUVYBGeexMOz/DqSI96
JaGCOxlLFhUkSBzkf9l2dKIFG4YYUR9cYfPIy0A1evFmXGwK7rOpTk++jaRJmuLdDsSxQsTQKXeL
8eUQvYsSHFXS0Dffc6fjscyA26e4PdCmyJlZVVQLl9mNxPCy/z884XvMbZbwwTVaQePiZpACEX5v
6f2hy5AisthocketrJtJ8+L131JWNBNIdXH3Ie9DpWzr1WUbgpZsDQ6Qa2BxioNvsdEu1oCaPSrF
Q2wHqENLTmNgWmeK/Rm55FHZPQpligCsM55XYx6HEGVUW0jXOQn0xPj2P+iK3hPMwtfzVvn/7Z5P
GAPP69gUDLI4Ycj9TD08h13umgIw+PkkyE3ldMBNk5bFdlZm7RsDEsiX0kNomZsVq22EJzG807vd
ROJ7YUzIQDaH0jAKm+LpAWmZcw7EcCGIABCRbu32nUkhO9HVJEmchenMegXTzJdrSDuwdwCnWY70
M1A2shviE8RmPCQmU8tW/qzYajA8QoB8DiR3BCSxKqfAOb0zShLQHYt0e4gG2ac7PXIo2wXgoGPp
BZl4SbSB5yFJfr9gzXxfstCVNJyIPky7n12k58GtBcUw+aed7WmyRf6t98VQr53zKwpNyEOLbNeA
5Q8ze4MVNM6fOvVVtCVzYSAetjrFo/OkIm7GICDlgDU0yyXPyZKY2L3Mxe5o/LjU3bRZfHjjVE+F
1vozQnTc4WffCeh1bL5XEW+N+mmosyUn/JQPJPQs1o1CRq1fajbga7LggjmJNc7TKb4MHo7TTZzH
ryrb0PnXl0fER3X+1kjmgGoJL/ItEhcxkFzResVYoCG/j3O9FltEDo52js2qhuREPcvU0EqZXr/b
CFn7q+8gOG1X4ZDuelDow8bPAJHF5LGQGVYv3AA/EWhabLP06pjeVNb5VRrj+FjvHKQSy25I+3sY
V8v6+zMSDs383ozwSvIM3TR7f9uHBL9LmZ94r4YXyOihMMuMKc1yisBYUAiJxwl7skh+WSB3of6s
Go8Ik/VaLaXF5uDXe6JROnQHOF7OjXx9plxocerAm8KTcQ0th88Z3hKf15fFms0bhWu6OCfEjXAE
++8T5OJrTS3oU4wlUfY6gd6z7bXB7FD2Y4DpFTLUzyRa4xdraDMBEdmHwhVdojQD0q2pKazlekr9
CUJ/YhzhauSpBxZIQScRh81uqxghUomNMgQzphChrCI+TbSkku8lOVgAvkCs6i5BuCbMP6aBxjV5
ENcRJ44Vosjv2/QOFYytV5shH6sX2vjq2zKT+HUNEVlqmWOYmdJ44EeKFU/xeYLp1oxudTp7hfWH
0C/91QXtGqkbx/WUSYn2+DP2OWHrfqPM1jdJ/QZm3SaEz7AvW0uOoF0juGE7Pum8fs6U3VNNVvWh
IYJEoWcM/PsBlmDvquufBCj5ikPFeAFAyg21oOKEXLnRYO1B2j6kULGlVPgTHayzXBE02XMR594Q
wpBgctJlsrz/TqtwrWL3tv1WXULcc0cxqmzHApcMTtcrBiV+mQUBiZuDOCQf6n83+ePIR4pqNrNl
HVGfBFbFzjv7UX7xfw+dwxJFQSezne49HxFUmddfnq1153whGLbPWPiyJyipjr4ySVQmGaofdGYi
YzTxIDqZvZl4H7r2Ne9kEYhNbE85rHGDIQwYscYDRBuTpCuxWV5yYEo9OoK4nnR96RZ33IoLsX8I
mCuY+pB08epcHZchxIxEn8KB/a9VJCntChJdFJmzjaa60j9xWRwbqz9dJmrNb4hPnniaWQ0FYDfb
uD5r8BwkfC70NtScz8Maaz+5pMis5/eJqOFsjDGwqnJLzi+Hz5s3Glu8Q1oUwI4/2OyLKg9UISVv
VabR9jlLVn8yplaSa05efRsttsWqH4uq0EespLOrai7N1Ii3R1jHmjKWuLjGLCpqfCso9EUbzaDO
K47WWn7mZU74lbdbHoy42nlr37jlM+o/iBw2hTX7/n6Xr4IcZLW/xHQzv5Y2ICfte6PfhLXs/TNV
HtSsuDSshGE82jZYBFzRoamcGaKfLKvS77PJRyV01G+Ll229YScV+GRZdL5RsFKfH6eRHr1s5MgK
ScxYjK1tvH1gTw6ySZJGiBnCo4xVqRG8kQ42qXwqdYjTtmCZMbn7FqtxObTvHJfm0LW2yymLu2Z2
RlhAORG8DTutc6Tg5aIp6Dg8tJ2wmHvdr50Lu2YU3TVwJ7Y01k/uFL9Q6gI8RHTB0F/HwcuOgi+x
GigBt2ZYpX4bsZ/9QIAJcsKy86F7Vx13wfwiQbO1mwcA+dSN31MphwA+IfwhJugOZ7NlfUtF79HK
hPlWh0yl1UUd4QdGy18obA4GELxSq2qqqzIVf0wmJjS/j2LSAm8Z6jsi0o15jg4dLMyCfQQr8rPP
MspCZE17tkkMimrDj8ZFwzglxK2cqUy/8MvPeYpuYgJ+V7NEFHvk/pMXBqFF0hstuvj/RebuAklk
+A+arGu39m8dk4ykjlWL4X6H8mMD2f7Stt4dYJvE9+8HB4EXTE2O6mLoeCc1kcyxA9Xn1ehtET6W
wzn3B14dX8D7YyPBPLRSuoaLGxCBf5gU4FoJbFaNNka0Yz9r23nTIf5Lk45pcHOzI84QUrpz6Qxt
hveZmNnxam3pOzhCR9GQcqzg1aPGl6VfZ8ww9rls0yyxyFxMa4Xbfknf5r8QQufyaPrsR3gmGGvO
6gXFnR+5TEF81Z52su7jQL302g/Fbdy46xgqeIIaqNXdTsnu2e+rlLVQP6LG+RQnV5Bwgf2hEdQ8
Osnjf1t+OHIgrDltaRoYvg7WupS4RWoOj3AKRMG4xXHdR3aMJ7S5CeA/6Dh3wZjCxAS7iP4TUvNM
WXboEsydVJoUiORbVV2l+dpXes5xmcvsKfh702g7AB9cojA3rOA7x4Fx7YVrmyYGO1VyMR7P5PD0
aCGIAzCXTnev/2+DRkyhA2ynhICv8q/2bOkhSjTrG4qmeP6+gQRl91dSVuRzAYFzi6wQN128hGaJ
ePoZC38rNSfrJD6kF05LdMlGhJUroNJ2RB8VEYu4mxuMc//XddfxkftH/yZBSV9vrqEftWVPJm0E
FzYYRfEt8kK1Z6rhkSYMpn5HaTPRtEj/GOCb6FdE5ZQAS/W4b2fNUDUkD02j94Ane5V9zyQiG02g
v4spx5Qc2MfYWYjoev2RnnO5FGBBlVnqlBbw8b59kDX5qVRMF/mTccy/3VfLfJ/bC0Y8kyRG2YJv
Eg8KpZNokflwnntOfD08SSdwu4bXD5OoKnd/YBiGq59zs0yXxqcFiHqPOnqdyNXY6X17nvuIVWh6
Bb+GWHZBGTEs2ow/v/lGBBAXB2kM1FNjBCFb+GriVQ48kj82EY0n+aizY6qTcYgJxGLueABYYafn
W0Hw8GPfwQSS0fXj+eh05y51Vc8H5LFqma4MUXV8yMNqC3KL/h7fp44+8H0SNKrpZMnXWJ7Aq1E7
q3qEUDq3iGel1DG/jD82bOnt4ONRB4QA9px0H3SXJfqfAmERGqJVSVfLMEPTtwmA/+ipSB0EEiEr
9ibJp0SLCJvUIA8U2XlNelmWfLT3ag4Tc9ybKRW6OpKfd0oz06k4y6KAMWYpjUhBCPX9OHVXvBnC
FEMnBdUzS7wxQWeASKhBqWONxxP81BDyyS5U+auRk2eHrVRRGBIeVyzPOFZjkdaJqYFMMf178dp7
Sn5BTaYNZ7EOsIHV/0Md5cUbBv4UquTgkv4ht05e/8UagQhtHsjm/FGrY+zlnT0mSJQ23JDjI1m/
1TZU/f7l+ARghuKUmPVscr8dNnSiCTzZ1hcmj/3uU8V2CxG0dGH597FOYruIZHZSkpagCLCVbVxs
KOpjmmMrDeu7C7tFQMGgqvJ19RalOrxTnZ4vscly3ORTjj83xQ7cbOBiW+Rq5pVIMP6zT0KIRJiy
ngMnhH9PYPhQsUQvpoqOBIC90RtiUT1h2QktFMaaUzTLvJ73UL+nb3IMDDkSfRj2d5MpmwnMj/lk
jbcXaeY+dS9xl3tOic7BoDkDSnqh0k9hgKtDE+qm9Qlgds8JQKlbUFe3Bsk2K0iA1RgOA+cORDJv
3YQCrmehhlYxccDTuUXVlaBObd/59y763Fh0z1J3EyBL5CIpny2Ynl91ISa7bMn9NGlVY0MKNj57
DiRyfO9KXqP/Mh0XMn6HEYZGiiS+H2SCnEdmzHv1YAGxdOWzPle92k8oS5pIdRYFJ/UioM4Xg2on
8l/BQkZjgcFqNM+D7siaAnKWM7W343vPITN1dK77UeXRUwtk3Lp/Z1cymVyv32cQ42NUBZD27Hcx
0EMCNr83Io643UM72r6MuYfsHWs1DrvAwTIhX3wNuDrmIIIk4GYrZFsm8A59idXCWBAkXcC+VBJv
LVIt6mHcKiiCTcy6HqvHNzhuB8H6oa32hPJsvZFXqTJQRcffEpqJE5nellqEKTw5NycvafWESZig
4qAA8PeAfbJXC/c0A9VO2aC1kbXUpZ/cStXuLM42xqYpNY5jkdnWkWu/Vu/nPBf26LrDtWhmLuhT
yPQH3x7DHlfsQE/Anifr3BNK5lY1lUUwZvqIk39nUTEdo70+RlziY82Nx3EIIW8p8SOWKd8t8Si9
8DHKVrIByMOQqcTCsX9Yrd0uts28wWf03wPb66oIwfYcjJsDWoOWn637WhKlXpjfGArg/Gi8QOnC
ZURyz+ihpauR7ZF3GOYfDiHw4fUdpvtUMxahww/34/FnhNXJI9vHz5DyC+t5NrxhH80EKiVAOpgh
bppVqLcaiBmYjoZWNW/o4xl/wCeD9H3FrEnNV/+rEfaMIzKs5NUPIY1J5dS9P1PJdW2JtU3JpMYi
8zW0Yuoj1u2UYWra0fEmaP+oA+SCkD+8E6QIt2vPelImlDAHOSuZaJz6eP6tbUAghx+PywhEmiPb
9Yd7wYWe2bIRaAy8KCegDtZv7FgeEnDYlDExtiD8yy59JpzeYbXW+uRddTZpF4D8NyOMBLGzNOtW
D+24Xit5vkP6jYstyp9UvbsubgBtXSFvqXXmK5lIDo7flh9l+RHEsGkKUkmj8pjn5AbhlII0J84p
aD+LB7kD85LtTCZcaOfSUJfN8oYn6Wj+gDvqQ9ubihvml2irKuF+Qqxa8z/V7eVWZu8AoOH3PaQC
2Cc8Lfdq7cuCV/aFanalKExRrHj89+W3niOXdmFBg2Iw4wq0WvTDqmueWCQ4YE9NLK2/BgPPCGXc
+74tjENffEtqo8eEyX1RHq8gd9AS9a5eFXCdLcHoBgLdzT73Epp5xrVOflQWJPnx4C+hquXIcAZY
sJR7/vUFnu//++2SmaeJPFW40DpRTRh17ROn/0sHFQN47XR1Bd6SMGCiFfPNrmszipuh2Hhg7HYQ
VWe6UF9FZfBmgvR4XV6XetfyDAMO+qOq2qzOZAmKsANUUN1xgT5yhlknwHsJsh2Izeu6aL8M9koW
2bcPLnU7BtPyms9WxE+XUSuu7gwHjLKePArNUco8nYxUzFJFN1sZWxnpnB+FpwkjHTmYp6iQOkcd
UCnmvRWvjdan58Rr0vtfd6llSYuF64l83CXSqmZgVGa/IglmKg2Dpk7QhrRMoqOs4TAYotl0yuii
JgGCyf767EDPY0t9Lc8futZ0qBIBaAEwNwFoXJu1F5JNMfAwlOoJoFYSPkCNhGqrYXtKqmkB6e+D
pXF+t3wfuPiWtNcvh28J3b/3prSHwCvsrp1SXhgFPGHRH4HQrIDj8Qp6jPYj49YEgXHjXz6MSWzv
dJVQqbhR+ZpIP2O9gfdaStO+dv56N87wqKdl7h1oCkUlxwcGTRtgKV4WOAnuE0lk4SCWz2w2KHoZ
mC7b2Bn9xhGUSSx0Pnx/WUgHyBS+x720xjAXRBEXUeLdWMAPTPfukAyhSlMK5gTsIJFrYbI3ZCIw
fgb7HKDfP5YxNloDS/VeredcNQZ5WDu3Pl5Dt3rR/KqU9r6pq/gX1w6hhnu31VneWJkxWU4lezaQ
97KvCSTxQGUWAm30h4nd4SCtX7sdEgx5o6AJmUDKY84Ar3MtLW8GrpWJOuPifGOvekN6HvER1OXh
Pfs7EMDeR0oyigfKikSc4OZm9XYAMiZpWqV6Y7k1uPmIHK9dmk1K7LsxeWa4+um3g+lYF6CbtA6g
sXEoF7hX6B8VT/IuLDUAHNzMcMcj3JFyk98kqN/23in5irKwc+5ZUTIGnRviY041bSKbKM+kl31s
XqmvtwOE9DrreA3/Qe3gSDStlG/ftfc99/LAKNgg9RzqpgayUmjrOJyiaZB7gYAXoBu6O2o4c8jm
+U3zb+7vC20cSVtPRvjollgk9mw7de/loobEsk52qcXnng4qlQec0EQe1gI2IyG5aTTxUnTy5EWT
oHGZLQrqkgbHOvDw0/eJ1Drk+foawCfVuiTRcNhYY0rKufFO8CdwaAY1yCnCp8JKwbhx7axul+yz
oEJzLZ3B0wvfvOa1pNV2KvRvJ+TZo2gKgqwNoGs2vMBKhEy2TNEAZpYYpukwKOfHPPoCYaej0IIz
d9Z4di73AcUTIw9eSkA7viqNddcrD/7WrxbrxlePNHcLioM7NSTDA+y1WQHTu68Zv+Ozr3kOMMe/
VgjtBi+XkLycbho+wBvC+rBbtKGG74ItAUhHovoX9fR+qGtHqS2entRfRkSitTHUKUSl7/kGQrjk
hL+4nj+8W4YVvIo3OmV7ZeE+boUlBDMeUA6nQUlf/KQ+d82XrzamLYhpr4RK5UHlol0n5gRhquGj
aXZ+TNswMOpT6GH3sLd4oxIQiH5pEGcmtmI19q3ul/y29GO9E1g2bjrAvGF8B1uAl6WBoC21exZk
YgSP52znSfmVglVOhzkY51kZ0uLBkWAynfKotHBb897Cuuj+9JHBnhIkvZSVAfpm7Pcb43j05OSA
mCC+qRXccKxc0dLIjROEiGaiK8lJv26LaT62ZRA0IY7zqk8rOuTMGPNyZe/Ayxo/7ful85SQa+4Z
eC2wO6BpBIU64xbSUU69AFIRSVNsqsgY7K+8mRhAot5NBK7LgxEyJRC4SebLnGCjIsXbPXoUf8v0
Rf8L6Wr196oobKng/+JDfnQVhdhDWxgKoFRCMQANFvmUp5ZWUlBvERESaXixE2djnBaeMNeSX3XQ
IOiZ1V2jVCshpmxq3QwlQHQqvljfChD92Ww0PbJ0zgrFCIvI4HnuFJBE9rc2CkZAsbC/Ixrkb1xB
gayucCqvMeeaJ42XTT7gHTW0hSOMPQHuMsfSoGLOJVSzkiVmz42uYbn4Wkg8OtvckNhhZmYOk83k
3g9S8hBMYveDNEIbVp227ALv8fV5tC035hnMNQfS1lVQYuycBbLTupzz1+mPF/lZWZR48TOQJm6k
1/IFlfNmO4WG2nK7xWbGekn5oz9aJcLaub+W/Lbic/KIcJ/YL3E9yb8OA9Sa+FwTdLYtVcegBjY7
amxkXmT4SOtlN88GePO1pxsrboi9pq+CJGaOeLTmkOMtrBk+QSjqVApD9Y3cucssVdP0Yt+6rNwY
RJKZ1O8g6c4Oht4Bi2Wn0/AqV8ov3+0XIqkgB8OXYyBArGBBlA4cpEf4rMFGBpjBKSBsPLxwi8YJ
p0A3BDOmEKf9wla/yFxLdQmWqYz16CtoU2mOWSFtG5HOTsliY6MYjBaBODdHzP/A3mF/DWuocVRd
qohPqItT6DUg8pycdjel6j9zX1IKB+MaWtsknbmnVgRgWy+297qTEjx7jHrJ30NeS0VNDfNTw782
wm7ra8uJpYtjlRt34nsIlDuC6iWC0v7BQ7A5AaZr4RdB0cRRqNU34xUoCZT7s3FQH0v9ZAYNNmBL
hOSBGWzPGhmu8k+3GH6RtRb/Z1opWTTJ5pX74N84JnyjLt4hLwi4T9AG/NmpBqAJGrilr9AdnlLf
Vk6Bq5iChgoExBJ7PdbiXV+5S7VIXFsfQLkgpnOdbgmij4cjfwszSp5VupkH+Mb29WthRVlYs1Mf
QPOeiA5aJXRYzZKJbqW4emVy8ClKsGgzKwqcNO/BFMnwP4FJ/CEe9e6vuh2EpaG7ruWNeWnGSA0t
wPncy8uUwnePWHTQF7h1jeFSnaxxkIit47kmsJubMWzO7nc+u+gHsZ4ltR7n6JpYM60zL+YrAJy3
3HCphxvCsNVL5vyS3QD0QKHd5BJJM0hE2DU7K3hWao1e9JzAgI3Na4mJuLx/s29dgB55v1bwjXaa
bnnbfIbvuLZZNelXk9EMjyoe+YcK+V3HUpKgsRnNu8ShCZ+X4O1da6JmOEv4u+MzO2Gf/skXPdPC
arHSm1VrNaHefqB5k9xlUnIOfieuONIam4IperkECQdrnPRJol5ptOc+WZA3jqcprN613Eq4nOO7
h2XXJbZGobgz+0AAwPxm+eE9dVuQKw0OT3Ssjk1FBVtoAHTvAnyabOVZxJlKWV8aAN+msZmFHo5j
ykV0uR/vckPZ82vp2GvvSEXWPvPEnMnWAQBOiyIqNzj5XOKBBwOqwRyGo7tqzXX30yZUwXpoKdEv
rEIAQfnKOcUigzSXnyFSNBOzUmpPyK7tbnWzxiRf+GkadL3bh3jfFLGxACvofFR+VMAcrcG+XbxL
DtiyJk96Yzhz3rnsL9MEiW9tL+gP/p1f8YA8H5Bf3kp/p8tGHgH5UWEK0HPNeaOEdZBds5p3FwCX
O6IuFvc6rYRzjju5w41hl7P0szAVONpszXX/gYa7fm0z3CrwuXfN7otJkKBhEFuhLsujUQv//vpZ
Za4K1E0HO1n8Zzrt7bMsPpXD0VmST4K84R7fnTTo48pXtjKgX3xDEORDa3nNDhiCcTNgcZrk7ksB
8pPcyRqc6QM7MlEBHwfk+ksN2BU7iegasT55sGu8dh8WtNmVkq30FysQ3mjSMCHsqjI+sF/wdEUq
huRICvMVpR9Oh7Tbo8lDazuRamovAQdtNvdmut0BLDzgH+rdJh4qh5CTVKyItx1Y7QU4EpEWHsEB
DGMs0K2OId45qH0ESQnGMwlnDzMcdDxOer67V6mJXd92nCPCjir1HdVlcbBVqkUmdc7u/6h82Odn
Pb+mKrINpdg74bdU61OqxRQOnMioyWJwmjE0AiYaQp8MyJ1iw4gcF9p8/vuwfHDMTk5+B3eJ79ON
Svx6wXIm/b06L5khw/maGb4YnlKHWSrMyoVlav7QDr7frarCtYF9/Fd6Cn5GboRyRM68WX28VwMl
R8KvTRkTLxbJzQL8c54FH/77ZziX/Jb+RxGBN9TMr7yecra1DLyz1tpwQaMoFPj49qjchOkZQ14d
AdZkNIRkPGqM7lQUJcbNdfSPaJhRWZHFhsIhst60XqhusxKM2KXfL36dm1UqZNyw35ylIJRpXuGO
GVn4mpvRvnStPQmrU7m/iBROOTIzDDqplemQvkjsDV0rx2K3eMViMGkedApA+f6g09HXZOzoPeQT
wX1ShvQBNVJhWf7RgEVP/OgvKz/F6kW3K54ih8ldJ909jIfUSuzPhuPL+DkNINiDGDM8CHReIBrj
KTA1/CsMMGMMxc2UULbOwSrf8LXGW+NYSiGWm084iOJmaf5PuARNziLIQyHrkqpOeS8byAKtXydz
AymMYzGEvFAu/XKxbh9IVDhHOslLyvXtfg8AALvY77S75AJVoeX0OyLhHxrhlA5HyoKKlD7e2zTF
KAkq7Y9C8ILtKoAU/hApfSDGoZaYHo4sCtxk2hMxvHhbOzDRNFE3LMn+69oyo1rGZAXxteTS7lR3
esfOy204NfbV0WrgdDYjf3Tss/qMEesB3Nk+MjCBG38awHaC0/yrgNnqbVHxnFnY4mhW4rFwQg6W
YnlAuh1Xs1/4CV4fZGzb/b/vsk3h3JXSCT4yefMYqrdujFgyNTrO1zQjtoM6n9XDMfJjowJZrb1Y
zJWxHCf1rSuAweYBL3mQrLeIakrusTLhRu5tmBHm4+zEagGswi9W4DG3R3ZwK61GfZvvIOsq+ax4
d6dGNtv8dqJykWMseiroYcXLW7sMe16KjJmYenM0uK8dzddcWmaVUur3VrdYJQlilqc3KiTBJL9e
/tsDEiT1q5aKu8SOj54m9mrydZtAY23wC3VEPScbcmjq7Lc0PdVF0Bm4z9nA32/kqtOh11qK73/C
4gXxLZscH4TccjHb9hyaQucemoDPQI7j6PD+IyAH9ZMzBmxz1VTiwiwYQLULMS4uwYM5SnRqXao5
vk7dq1ZWgFQ4vTrnlpuOy51mb7fbVdvKT4IPA1r6Fc1/GTsyKaIJQuWqxtM08pHhTO0PT5ED+INg
FwN7voLwYN5/q5aBjNEMWVacJv3ehC5yT3jzVj9Gtl0xTgObQjm4Ip94qaUAyZpx8WK48M76k7VD
U0VlwIiOPYb1KVPINP9Bn0lkAYcH1Y1VIGkJWCwgaV4a/2AGmO0BfCKsPpNey4Aigw3Ufqvbiq4+
TECfBsaF/5331XCeqANswuK5cpAgzRMAXIwky0IwBYwdZd+YYsVXGTw2cki+RZQXZ44Se/6Pagt7
snZpR+C5SP28kiAdNv3hxEf0eEQFiEHKeyIOX5XX/rtNck4ljm6ULXbMJpoYsUS1b/H1ijjlzi3s
pXlGQDmv2/7MiRuSLYK7V2J/w6Qh0BhsWBJqWCbm7JQpK098bMg9l0ZVNcnGUOhTDIJAXadhRwEv
MqxY6t4nCXETaxvy8L9oww6AvhEY49CLW+8JAPe7suMinVMyBW8x2kduLZgqlZyI8eCSRRsi1v5Q
XGFF5JBRxpVtq3UcwBbKYzBGkwf6spuzmK9ZhelYzPeZ5eoCeTNgKZ+WDc4I/mR25Ky9QZMNHZ8W
xwfmRZUpX08IT2cH5BjPsujoOdLQ1I23ehRFdnCahq8m0aiuXw2lou7xvM8di1HLE2uGUpYTmKtt
s6DCVfGHjDzNhSW/Y/0oedjcXs3zLvVjJar5xtSsYj9FRyGGMwgzSQsOduok41NktdMyq6NcqW1X
bDGf6zeL+NwOjR+eIwSe0ZZNAVgiI0u+xgwGRYzngTbitT7uPodi4LVLXfPYe4PwsdH7KLEVpuZ6
ONQAuRdiCbuIJVTlD0bvsM7MLZA4gI6hy79G9mzFVhI0fe4HJ6dhKSxu7nvrYSKdp3zJ1nIw8EFd
4VWFHeUeEkmE7LOHwcslJpzVzDyk7F+MhWZUBsABIwMDb96f6q/a3Tt+fiVcqpEdS5vV0XC2mNQJ
e7EYer5erEIz2jeEVisxJblNhMc0Y9R2R6r9rUjdDgyozxMyEjMHqhL8xeM75sb3YaulWZr7coV2
W9IodbRpMcXHlc6eNdiPOhrNA3cimU14xa68Rfg282sFzWMSH/oLjpHdudCiZBoMI/fGDxfeG2nd
z7P4W9Yb1Ute6ViKv5wNdhzPKduf9Kpjv9KOSDfLi7CIXN0H+/rYmXYaXMVVqbuM0gfszSAPewD+
y0KyUY4SUb7KwOgpjROQIkvI/S9n2MT0sOfQAf2GzoAHOEHpkuShigDeKH4nHDe3ZBjOgie8wenB
LefqK3R76fiNql/No6Ec3yxhmYNk+kXQCzqwAmOlmcsMxWDYQi6pZr5bOo0xKxcfBdZ63PQLMcL8
S/mjwX1U52wBjMj4xHahzkOO5VNhbrfhGxyCdMcUFyzhUEQ/hriE+spngQvEKvGfxrCeVKHPBs6H
HhyedRO1a9FXEqKNnaDMMxXd9FzeMEKBuqd+zD4+2r0bSCPvb4dtVL+kB1EP/EeSPOpJolBtkwFU
pG2eUX5lOzeW2la0Nccp6GmJuCKl9tqxJTH7PXr+r3YApZeW9Wb6e0Ty8tXRWB9jM5U0rBqx3g5F
oNsx0sWYmSHm0q2D3gtDlzaMzyHEeVmen36lOU+C+95o8stHwCJor63S0KItuTzC2AUVsN8QtUr3
cLDYts9QH4IlU2eONhuqZsnHxnvrMIjw1OKwyisOtDjdUxDjPWvIFFSdMq3YWYdJGlrVFx252x+i
5yp2S4pr5UbkMTezMz3yP2k6547p+7BQPsEOFBXEEY7GPBofZi9hX9rLBohOknK9Jf8ScsNwL64J
1U0RVNi0eS20Jb7rtMNc7+VPJSixBcAJzt+1XeZ1zwGEh+1rgVKfCRQK39LsWkFQKO8YljzLxNQ4
qe8mVznHyL1ClssehNqt7jfU3AzUAgqsbAV/591s5pMmY5AQKQoQo5YidQ/qCdu2S7yLNGiQMBca
NHCPySxQoXVIisr/A7ceNXaTG67+lBCKt7STf4bZs0VbIlY4oWz8lLSpqWXgnWQ/n4u+MGCkhOv+
Vo2dKsAxjuSBK3phmGmAIxO1/3EhUS7BhRLBnneUIbQsyZsnF+NxB6MIVZWRHSPWu4Xdo48Ech0X
VkVDQ+zov624FVQHAEzms3V8W82Q8udWDRoStGOyTp0ajRhhaaeinDL1XS1lm8+/n3V9VOJTrMkr
2TQzXBX72pUPwUBBKiTnU5nkf0qwVcVFxGsnBEFGTrDr6BkoMTekBM4ONq9gAhWHExBJcqX4dcgd
bA/MrdP9AmDGVx1KypEZe5RLoLnopWgdQE362a9XBmGsGGq2TOgJLApf6CoYsg93bZ9UB8f0pyNd
UEpOu0Ngm0ItG2n90e5HCKXDmBz8otBZaRsIZkSQzwPaNIMjvUiygaD8XSmfZS2n1cyr0bHxt1FT
AnwskQpnT1TXpQgA9XQwO8p63Cv45sxgPKnxT9DyREAjfMbsKeQNSFKiP3DAz6+VzZ+sFzPnMqj5
vKIoZFui6IovtdjenrF972ylMV0izLvCoA+O7b6JrMUzrnTqSNGiTHL6xlXIQW6JEX4xO5Jvk/fY
+CkMstDq3EgS/CEbAdqg7tYDxdw5gZEqrItT1gWE4S/uTItkUfpUh0er38enLdZVe3PMBEgJcbVV
FQmsxeNdrpi/GKdXMXEw4biy31ddxo/LWV4GlioR9fRerwngv1zF6tIosYlIUvmbRiINh8olxyVx
k/6bIfJXrHrOXg2bZ7dN9usEvFC1oSF1PUUPBE70HOO3zv/H2AlNCVoNFh6O0jUyYZWrN9SnBqbZ
tVDksdU2JBLJveEiPXq/EAsSHaCGciMbCCp6/bEJBmybnC0QjHMKdoalxH9+Jdiq/rNifR8xytlR
Fltz1kL2EiY6WAPDM4vtS55X4tmDSzvCMxeUO+EnjqY31a+2pXYE6xLmsz9K5V4TWp00jm47XSTJ
fFkiKSuvRZ2tVKD1aUYNmMUBov97JPDqArE2xo4ETGdbNO+rTme6bsAE2Bg/LXem3i72XpkPIQ7l
WvQPcPxkIy51JZzu+5+8BRINX2J6UD2yw42y0FzApJ4CfG/lR+/BMNimdMymQWTN34NZ6FQJENmD
ME+iiSMkMmWDbD2Qc6dNb/lBrl9qeehFBgCCe5iTkQ9m8Z8RRnFHiyKaEtZc2SRBYrabeS2c9V5U
k2RmWKlLIkSF7aD7hUXcmF6RVpsU+SDTJyO3h5nYGAbgOqJZJ7L1A5beta3mXkuPHoy25UI5iAAl
22Pxoq2bc7R1SA+pSbj6yMXLEX7BSA+Vzrn4utZ4JnL9VE77NS/K2lQUCa0l4U3WZv95NRvUZdIn
+TmJvo36aYKydZIL480Hx35qyh/g4RWkfeJ+siU8HWB+mfZvV6hb/BfTLOosjuIw4z+z7guQBRqr
wlTUDQmu4QkyqmYBMVp+1MsbM71D6S3B3dBwqr2FQRwLNu11jpCFCuDfzfCbbNYfZ7jaVJYcBV4X
u6FI3Wp50oTZE62Rk6GTCBo0OMQGurJmUyOrV2TzM/oFIEGRYCLlg0fE+V2lcSMafFyX+bo/zNjT
vl8wzmednvSaHUQ41682yhp5wcAqgDSgXzTyOSpkjISgcknIQ2luh5KjtWtdLeXElZHFB37UxGph
pAAaa0GfZ9F+6XGYx9QtQqHVp9USDyCpHxdwD2ekHhxxkb1HPgcBfcx/w1sQR7ACJCH4iGRNDLzU
m4s9QGIrtc9fdG7V/wnLB9EHfmW3nAOYDJKzsLS3dvYonQrCajkimj2efUhTrYzWwmveiRoyeCgP
weftiLAfGH8QTQA45+8cjDh6YrISQgDhZXTYaTZCq3FNrN0ZAfcZg6IDx5Xdp4BjId+XTU5Hi/0O
2ERJA0TP/uVxhmVL+2JH2zHuI3LokyUF96w1JO59Ajsi5dZAD5oaPfyPeET0k4Mb60v+avm2YIyp
CWUqr0hoCqCXX/sWt1dFulN1cTUdxj4H5//6g+GupECDDE3M1YUUfzVnHMsYyDVTZIraksbWz3wY
zRm7RDTrv1cdgzyeLOXUsqbBH0gjFToMf1N8/UN/VOWaByyzyr+q72Z25iYyMNsO08MDbif4f84M
+2ClfSVsEjrCx8FOFgcjID1+P6f/rqSLWvPJ2rbHt/5tpQLih2cOTZrSpsa5O4puLxCnTXI94d0v
33dmaj8CFrDllfhCKFrW68Hhb+3Wbz68mUmulaxQpi5+NfN4n/vU8Wmgwnsq7Nclm+pXooINYVgA
KoqqMlzFBaOdVbav5Ktz4+39HeL8Wr8/t2JzjSlGgwJprfPacREFlL16TnkX0uwCA5AgpIJTPiJs
fZMPi65Tr89YbIedUgwJqRCuMgtDnx3+l6Id13j3HfE/eZl3yf7DASViua64e7xuWhRBamQ4N9Gp
wqv/O4PNXTHAcc4VEuHgU/vEvcB0FrmeGHFDKpGUjVWgEmyj9JMy92xY+PvTp6o2CEK3TYtuFXFm
q8YiUOQm7DCZJYWG6soHbs9JLQIRNoBupjeiMIX+ENib/5ydjbcmhMCZQyqoUtwaYh0qapPMwOAk
kAKStb/cCUDPllHE8Mqa0RGUNdjRUZgPe402sgCxPSOEH5gZCDVOWP5VGGFEv5PCsIJ0lkFwtBdx
0utv+FPR7WXmTYWFbpaIUgmWkzIUWX94ztYtNaHqpvQHqCScrO1ElDyYfVIhlw1yXS9xWQiP8dSx
0TLOESbc4N7dPGIyWTXqXYZC93kc7omrzBrzOcdxe7gArNaZnxp6HQXsel+WUZpRhfpppXBKYhJp
aXDXRSX5YigesVwtThRDc6HqeuZsZofX3W20C+4bcDC1pkanWXvcZFzS6BLABqRkfRhtZatlvQQW
fPRlIcAuAEmtvdF3LXuSeKI+zkYr4qQcgdsRKAqQTOFa6hJcRUldApMTwP+R269crYckBcLgFEeo
FB0XYTpZREsCGQHzzQkjiqhbe3m9fQZO9yt9NZVgfe4HyzIkN4M7wvzInkPAGpRITJFkj4fN9jVX
0pwolnPf6SYPJrWwFJb1k2TdUcwW52LEqORjbVYDiHmIFfka5D20Zus6ny9ISaWz3H3x35RZs8RP
GxRy9Dj7u5P7rpiLf3ZpCR+TzxKjMDVeucZdbsm5I+Khcu1LmU6KgCcb7Pbcqee1tMEZhtgaoKaK
6HRBuqm5DBbehdpU83gWvJU9Lxl6x5VqiK41bGgkO/bemZgoF1YqFLN6kY8kRIa9KFyv23utGgJc
/FHfY7rWxCjkq5r3FrqJtFCzqYHWnPolwjSFuwlI7AJ2qFRPJFe0qN8dcr1yh3JBsh59uOueInpU
6yR/Gat/M9eYe9YIngjhHX2/ZVH0QdxAo6aQsqePGkcU4VNcLjKIEWtWwyNt48r/cKh9UPh4LxG9
XQ4UVImRSNlyT0rkZwpQxKDak7MPBcGTnz/nBNVGh54oxh7xUT2HidEYm0qjLOgiAUylBHnPVyz7
ix67yuXgDKYNgCo7P4qtHWYvG3hUh0/llv8tdWtm5TdplXicLKz0j7Gvqpu1ABU4tt27imlSglny
r2sOfDXni+i7lFqTUKGwl29eV6y+CWFvxIwx5kZ6mnU4n8ez05P3/tfc6enDb6KJaTrOiBQLdEib
R3030kOVc1TwQvn+sDZ5Ejo1ayCze4WleEASSYpm8Hz38hVKhGbrJuD2ZU489RlAWrWZiBrbgvL0
E3huD4Rq1ngbB1ptM7qmIWR1ee80ZGPeEtapyl0dQTlGp1Sq5TugHHZNxX9nmFrgLIc47QKjuJEZ
tL4fWq8vLO0PzDOogAkzp21Dt1MwJtXadyrRNVezOdftePOvj5FD0Qh8QBHgUNLbWbmwBVgxW/jx
Uv9AetuL7BKXzGJARWMYPrvMJhgPMHuNsXZKBCZeIypfUv5j1d3LTvrLpCnwe7qK2sSYQaLr+cv1
rPlvFKiYnJcw0Ua74WYmyzrPcilK+vI3yrn9g90KH/g04ANyi7gYAWmOUKYM4ylEsl7tq73aLJCH
S83TQrQSgIGkGR2hsQ3fpGKAqJAVpht8OGFeIxEdEJmlDPrSsQsRqc9SxJJJ/uJZUtczc1Sw5kV2
9zEYkgSdfL2DaWcvDGiFjWR8oyicG3mTv4qW/NxejyvHSYjsnbDGkLBy0jF5v8cpEvxj/LUeW98m
3ckfuB0Xb1SGMexQu8Y7gI6PZCaxS4NWFP0cujOnzvmZ4F8BLSlFEyNdnnPxkc0g1mSvL1ZGq3hT
TBO12PF1iDcbB+tx3mJtJTuqOKol5/kmyw0k7Dg9JhggALAF//VzqecH8fFUphU0Tc3RObP50Eh2
WU8CGwRVBLsh6NyWVmok3LcXoJt55wRxSpxrea2HpPMeOx1skM8F2bOIYRE2VPyp9d8nxqO1i0cU
s8moFNIhFDyGTXQKAubaoyYhMVLjnoZfGZZGiykrUoT0H/2c/cTKjCY58GaYyENS75ohmnwEL0QM
FkY90RdEQYuTRqVsaBwdkz689xfftG9/K8zA3ea/YVYo79VOjoA/0Ky/xfVb5VyK5Df+yRAoOc58
7lJq7Lx809DWNAsi3UP60HUAe5vio/MP6AAostmwfkz9QBpLC98v9vKSTtN3DCqPv1nP5XNz0slt
sPvQNLNHdswlGRG9kpI9B+8RseuGxlMjmmTUKK443jTRqcJovbhsY8Zh/NmXmMlbcLL3yMHrdHJj
/G87pFEk9uAo54zXfd3PiNxkm3FUr5Qfpg8ltq5GewjiXWovVsk2soVfPXGIKWdp9JmVjo4lh2FE
d3MwdRzRbGakz4DjJWMEfULeVcSEfDgvhZiOrWHyrPT30hzlWinD50DyaFzeq2Q6kU4qOW6aBlhn
jvwK5ey1V6rU+9MGxetRCF1GmV3OGdan87/ZapktIStiLwfAPj/0g3nLXEoLnPaMmMdyFdASTLwR
UF/Gv0kVGy9pRtfMfi1RL2wX6AtUKtp6wLErWli6eEGYrpFSFZ9LkMhswq7TqdsiC+8PQ8t+Z5om
kzO1qYVw3mzwBuxC8tTr2lFK86wNFceNzN9GyKiOdXlM0mR0NVEZv4+HcUVVjigvy290PDUFzpVV
P6MUKE/DSjTc4tVWudUbyUdPJ9YHYLuCcDV5UblnxOsoC+RJ4EakRn6EQvzj2Dh/XUlAs44xFkig
4Qf3GnP8Cv+v0OurhjTXdsfUS0TqRKQfLqeUIdl9gpCBbvWIa/EfI/oOpjXZEPZ/dQ4kANvLjdwQ
kCZTQe7psDj8BeXR8fxH8iqaRrh1t8ugwjuBj3/MWG4tGK14y62IQbC8ZRL4NVNmV93lpXHUxtjv
Vaeofo0qeuSm0OL/vZ5YQDKO4eH05bb2QP+fv4moK7ZwsxZPJx9eVV/mGYoULPjy6aIkMvpfw/lh
nXw+5msj8k4sOSsHK4aFOzbHlVkvP08Rmmvn13u9WujFb5nrWiIT0iMb00dZ8uL0Vn8fTezH/xwI
B6Fh/+zvYbhqVKjvQzAnkjEuFUfkYHE7jM+gpPOPlHSJWvTEvi0d5n/E5dZaFhHY9e4ffroBaY/E
Oxay4lLEn86ueo7lV30OqrocML6CpAmDwPq82UcQ8mCzlm5IhD/1k8rlsnA7XeliXiErBgjJ3Vzk
M82cA1im7KObNZb7diQJoeqnjTyHLHvN/EHibo3nvbd6R+337gVjUZkqfm6RdjOiFwPgfmazyDr3
lUn7t9WX4ptaIrghyuNbSErhM3fOnMoZw/XdPL/Uviyx8nlfMvprD+p40+g/xQCOAQRApCVqhP2G
kxtTiXQfu1f3/QZ2BsSw19wgszjbEWeMBbqbpzPre+Zs86uFcgMbVqTUVVY21sGPfydClmfQBw7k
Iyqq4AMfLdntPXlRhglEhvuus9kAfhKnNgWPY/oObcV18xJY1C34jJ39VKgf6RcoKNUwO5evqmzl
SoBY6uFIjO5r5ubSz3IsmiiWCVMOS4iX1PpHmBWPlAalpzO1qY49zozo7apuElRSWscqoq5fC4gw
5MBvioajOHTUk2xFasj6issxq8/NfxSdDvAijObfi1SelptFiakT9xv3hqyAsjzQcCIaKhyA8KjQ
kbfMWE8O7nH2ZhSiCQzGjz8i6qVZfAp+2ZBPyfFE2MDsPRFlskUzugpitED3wqnbwFfXn4g88BdF
TDTmkOuz6SDguxKex2cnS9DxoLfQZ6gMtXDIWcgCES1KPUtiFXjeuRSCiGMQnfSV2FfSP8mIq7P+
2yhXAYAf6l1fO3JQWUC1QRf8XVMIulSiiLj5fStaZT4FEIAj0DMrxn48sm90Pbc08g9VOyjuwHlV
1KyNaIWe/BtiAx2lt1EuiB2gPh5zSOmL4y+jUn/MacxhIui7RRqWbKNBTQtcvf0rEYeCumW+ZneB
mkaprYfMv+bqF2OUaATqvJGX/wvRxJkzK/2l5w25zo4ezB3woRtibN4Zj0iwHaYWqhMyv1+WWmKu
c1A13F7jmNaPRvArZhNNSY6CL5lQdiLpQgez88Y6moDmDZj5uVcY9Jmy7e+hiD0Z/4Drf8n5j0Qj
R57nPIXSwZKUHNRFFVIYM8qXAWdUOFTQfKKJZjy8aEiIUKnq4obHZ91u98aVMYXLdoLL2JTScNv/
AC9w0+A8vuBJ96kexmUIyyjei9sZL+FGxoF8zsqbWcpDc2olUzxYiXs6W7fPMO3PMTmtMqCKhCcx
xPeZ1O0YqZUiw4/Ov0CQfctSE8Dvt+usuyzzB0/COSzIbzryJjge1cxR2ch6fk/zchGJCs7ZcR2E
iWBcd7Vfhq1pugjmkcVFpI4h4Bcfxlqq3qlUt1d/dpbTKdfQEBJpzNWzdAv9fdvHpA+Igfbm3bX9
7yixA8/6Nct5pUv/wXvaGeE0FIgEDON+ICHnmfU/9tt7n4x40SwCl9c++vczC0bV/q3njspzv0MH
0aItSiuWmhHLkYJ+SzNvQ+rgKmchSn6ARFw7gMW4t8WJvfynZcwoi6JqNk935t+O6ZaZQYu5eUJA
LH0YzOWuNc4zOGog30G6T4/XvLVeiSf2mPV7V8yBto2IG+bWALJuBOjcTGdEfpK2CfpjuAC6NDip
ydMNiYiARvMHdc6jBxusxaQRrf9hhq9P7bdza5TBmj58nzd2u2QuiVTRLuA9uBy/Hny4EKuCNITD
q/ZPF02B6QUJzXkH3+fdGagS75HGJVkNtMF8H1R9HqNnbcCUIY1lsT9Xv/cdiiMQCcdNH7yTuvpI
Jm5JlRGcElgmareErEN1GNL0fV4o2nbXKczAkY1WnB9vnIsrW8ZO30SjMLlruq/VHpVLtYkEH36x
4nWhEV0lzjnqGNqy3f4MFWujdzr2GSg2+sKqwkhoM4qTjF+iQAIpKVk3xhX2IYEar6x7qkp2usnE
fglbuIZho0Ry3+EHkMe8lx5jpzDBGzwTKGzarDlSt2t0fUJycO6xs1Pom1lHMFfggTih8NQ0ZzcY
VH4yliUZdj6i+X/WewNpm9gA0Oka5D7uNGsGO2IaTg4Ecl+cvi+88IJuIWW1tpZiDRYMnVrpqn56
GUjyUZpF2FJr/Sayi0WZnwfh+WdZcL2Khw/2xRsln3lJZvWjwtL9CkTJZj8scYxacWBfi4MHmkMo
20CG2qqDg+XosHsqSI4jFLvRBr1TY8C5UIpQoXHDETmrB6AM1FTwfae4Yiw6cKsCp9Rjhkqe0y4f
UQ8zvBTN94aGqyr4rcQnmDF/oN4DG9eQNyRkPLlZO65gKD/0JoOFlTnfsSP89oUq3OkwdW8e4plF
wi053Arv1YlyRSot2GUGdCtA5GmbTVZuxZFuGqg5y1p87SrF8rLlExjElC+ZYtpRH+22umLtDXc7
QAO4OL5n69//0SojIFz2+vb8MUgis46Bia0VO9fBviXHmlf9ryW/FgG+u7TeOBSZ2GGGnC7jwaaa
VDoSAs2cQnduoeSOEUAqFgD5axP6BxjgPUp1KYjMNbYICH+dcL77LYmGizEoVMAS2eIRdLC3ZMlh
mHbXGWFeI8jJZWGosK5xLQaB4FkU7paHrCdHQQkKbX/mFnhYiGC8PiSc/s0Y7xXLtE0TslfuVCGS
uTuagknYJLcHJq6s6MIB7uW5C8AwMry7jg/uXdr04jZ5rXSd3+lelXHkzMa+FMGtZiJCT7/XrQz9
KQlpR9KjIPD/pIEvazRccT5Wvg9zgMi0CCgCPgCOYzu2kEJRhTp34qcgb0W1Ffiw4isf1LUjApMX
p7R6IElGSt4ZxO0ypPaAJ2KLrU+F7uWpJm6/TZbuiSR5qkG3LnukHDxydWna8CAkwArrSs2fNzwK
yGj/KSeLTOp/ZDnh34kFRY4SRF7ZMfYZv7xe52gULLuS3+yASgOOA5kLnQmS0Ii6E6hON1K2XGuE
XuNlpxKSCXafA6o7c042vF3ZYmYl4E28gsvIaVAIHtSb5Z8IcoVXuoTJP0PYcN/eUPxxC8LgkXAD
GLHJuF+HXbwE+pOjad+Z/wjl7nIZqbVolqBbcrW+Bt4eTViLyQ1mXHKGkT7gsV2THbvSApJppeix
eTUBXW+rTAnsegf4F+kUCAek7gEqqigup7WKoYYHUISIfXTsNn2libNCQ9NboQ5vdoUoOVsGO4bl
LndNJ0su07ThPL3qQg5lJDLoKwPkF3xIy8+2sN+WevEFz5pqetVbk6u5ON0rda3KDWHOsHlD2JXD
TBdIsD6yYxmtUSMNWhfB5/tcBZ5xRC9h55faxyV/8wQAeRHX3fWRw8EGBfoHoPL7ztbdQYwPZ+p9
1+msj5H6DJ9AZRUz8OERjla+Nd/ulwNe3m/LwcdquA/9N/iCxW1ukwYufTsqnaM7646NG2TKo5zm
fEVWzLBF5EZK0dg9skIXcEqZMkXKxtkh7rFJ4yP0dQ0xUknsKIyHbPed44Oq16QHHmlToNX4wpux
Wtx+YyHLy0R1QO7MZ8bdi7S2YcGcSI42q168fOaYopRQrhosxhmnHyY08CY6uFOs2cLMKnIiJlBh
R+kN5pwhjDxmmAG+iHr0zWyCCU26XXo1yjSjxJY5GG1OWCDqo/POaStpjxcY1Aae6CLe8Zaw0v4g
ioJb8gwq6pz5fs+vmEg46+ajQIIgRGWirhtXZWEepCYZuCHF0JZ1SyyKNGlWiRKL2fZXihKA1KCe
O0ioix6jF3T5J/cLCFq3Y2FXfGTij4I/JxCe+93TH6gmKaX4zJ3Fn/oUinrNy97uf1mSE4dm2RZJ
nYjNBtQSA/emoumEhXpiXPFwZ5liAJ6XrhkKDTHb+UFI3NvXz6s8FPZL04gPac2z54lokBj52JoM
7OEBw5pV0pWfrT9F3DtVWa83N4EvnA8zfKe3PJimDEgaIflG31d+JZi7Ci3fmBt56+0508U8TNLC
GQ0ndyNkaLYeaW31scEa42S20E+bPRMTT6fK1tKw9GMfsyU3il74RTZRkxKABY9+lWhrhtURHLXs
ootbdO3559kFnymNnfK3F8QDSm4dJsKtfMxx5v1QRIVxVwxNw6gezuCPm6lc/5k6qo8GJPXr04wa
sVIxsXDERSRUZ++z7x+jCqzxaglx1JzGe1KfxUWaph8zU7j0V4qPnim5uLWekj7yriKIGfeOWJrq
HmXV1BQb3nRmhCGVZDkxsOtQP4cyzcORw6XRJ8cDQGtpfMfqXidyh2tIHcjTMllygVc8I/MQxkf9
QatC/9Tim5vkzK+r9B8Q6Oba4Q+ZfwVbQdLww4hb1ZNq5MlFrZg8gFrwM2bHoQLmqNeX7u70Y1lq
OrB/7Ke+IP0+fxnfitxCNhnI+BU0RjnIoA7395cTiT0azZni5Yw4ug0jP/aaPqNM0BLUt/UrCpw3
b2S/sUFURELJSAirXjXH10ePspZuLapLHUWciXPC6U5Or304KnU5AIhX2uTJAxarFDLA6Uly1ld1
2Bf7kDbD9FDXNk88ZB8dyMn8WTswvSlP0mHmS3XNFWQqp+nhdkwcNmVWt8VQzGvNMcjYjLIkgcrV
FR/li2R2jgtJRaCDzlGmy6V/DFBxphT8K9NU3xs5strRTM94SQrsYcuav2WJWVw1Kcz8Jum4ef9F
BAQOuRMCm9ZqDY+TOXR6gedE2D5ONpBQAKCuBDzxNSBlfTDesxXHUFKhZKnePDh2VLl91HVhL3+n
Je0OWGFYOBCKqX++9/tOQ57byZvTWkSlQbMT9ABbHU+TZ4CWph4NZ0bVY9WlKVmupz8cUOn3Wlk1
o+jUXnwwx0iaZ1IEJ4ZgjQDRtXNS+48QGfjB0HnQ6Be+CxCmtv+/jF0HxxIrcwn6MuXxm53EhpR8
FFW+b3g6XVY8wTGUZUn7WOjjfr5WRjtofoYpbcqC5i+gMSeKWklj/MRNbJ2ygkOzL0L1aik1HR/S
Wexf28cbXnBuFrOq4U8hWdSqpzpFD/dC9aKRdHjM/yDgwUcStWbpBZghlU4xXgYQmhi3mBIfxB3a
6grmDkt4cB2o9RTvzLgRou+4K/mtonT/TSLcVtEx9TdK3JrZAejMYdr7KTfqtFb99TmgjBXXff2D
r3BMijWwV56adcas4ZSw5umJLsHAVixNEEDK+CfBfmHV8OiIc+tfZ4R71Uks3T0Nc9wYpx2fHia7
5Za2Mw1Xem5LpDgri7I2LibvkuKKmaGfSSO4OppogdqZ6G2JIXBg13TxqDsua4/NFgLiLygk/QcE
dSGm9mGPL7hsmRfWzCggEUJ2lkMZRS2Y0bfU9rOzYs+OY/KLy4Rt8x1NzDyGVWXWdE2Kud5K/XUg
pihHt2sj+RvR8auRuKFQhYbAxVKKNWh3a2X4VBTKC2wjp/Y8L4GnMevtGUCv9gnQkvCcA4V/RWTt
yh6y4a1SqBSwaIgPH3b8/UR+uKSx8xDpRSDv9K+uEXdoJGzGd1UtuB/jQJzxxQHKa+UzuqNhHf/E
HwRykbWrOHiNsnhlRWC4LsdOHhn0ZzSa4yflVucLpwH3Gd1acjJw8fqIXRXy6OZ15AydXKO4eT5Q
VAtSFJMP9Sxu4ozoZs2oX3PviSGGgKQGRYWk6tpx8KYDwjDyJlsOoV28TWBX3FPylSNpzbs6zSFU
ysSoHoOpAYzrfYXop5xG7z41xJGYSNRyPA0kbAQAg6fuvbAYgDXFrwR/CX0Wp5ykaJ3ggxXIUfDV
6XMiIT+xxLgM/dVEJ1TZDcDkcwqHpQDb1aUXg2Z4zEgyCPX3ipuxtxaXOH8gXTugfXil1SosmQ/6
KjCDafVQouBpRzysNgovKrvbhEQSgqWuz8OfGAtneLDlmI/Xj+eu0zx8gdQepRHSxy1JLcqB/y1K
R9/syXw8+rU/CeMIz/AodpgGogwbPxaRA++t4H0wZlMrCtWosH0RCHU4ShjM+zCZGN/Bhxllktnc
3n2Hd1k2usILNZdhF/2+6XeiMIriJrL/LrFqUItz+3rmQIPvFESz335P/KbW4t1Ipk8ZaWIUpmPB
isd4VDilWdGwDZS7HIelGz5qXDkdTfiNmHA+WETJB2hZtVf92PI/hGYuC1/ueODDdfGVXQZlg8D+
Mxo6azfLbeI8QDGSS9P+k3rhMij7N1AyPti+lRvuqs88dvVD/hRJ7f0N4flest+U53Xk6FIFt9UC
TcUbzWiTdzMDGN0dYl87ayT291ztwFwm6eOJ7GrxaevdSCzNw/ASn6/wjeauaUPzAlJqDhgOHEE2
LD/DJOW9VwSqqxTCTnsLJ4r63TFkzWJ1HXppgAVy8wAwJYOR2t1WzYFvotuscl5ivVPAGnC0F039
F53t9vzrynjKH2lmXA2qk4uVx8pTub/qbU80mM9qnPQxlm+LqCzCFYF8dJL+a79VQp7uYM+9vMf5
FsHaJRhN6EYwdw2UfMD3DNsPzAg0DhTYbOqvjsMHNSWHXIPYcsCzTFxC72LjSvGZ+C4CuckJpeLd
2LVCtS7OuWo0x45E8Wh/7CrVS1pEuE6O58RTDnT+K21ELOtJUL9KadD67a4fgsMMHBoTzN+oSVkX
stJjala6buhKm30Bl0tIKcIoIv8T2P771HvK3KRU4TYN99P3aZdniNbddbGOMNgTmqsqYktILWGo
90vaRuAkB3qWX9VKo6VTxoOPx64L/DBuJTUVt4UmTRupwc7ZdIIx1ilo1/WJMI7G9cfedqUi/KtM
Gx7EPrgVms+xlt+XZedfhKZZDnQXfSExNttivNfluS0j/+oIwCJKc+1GGamXRPKJisq9kQSgncDT
JLHgwhPWdHNvlSRIwkC3eB6CdFjRkUEcQjxsrG/njt2k1nwekpQkedjcAnotUGT2wyxOQdjj9dBb
/UtNKlHu3cRM9EEhBiyMWLMdm+kjoeo8HLb8LNcIsXQiUpA4OPEM0QtPyvgWCyYoszxbE56g/HWD
yOpyNCJaZsXydbmlHmeKxLFg1oA0gsjuflUT3tXJsBhZhAAXV+5B7V2fU09rh16D4yw/7gprQ2nL
ho5lEyh9/j5rh4PLqCTmBvQnslVbSGJ3G1jo7cX+OOTm+VeWNMVRssY6K1LoBzUYrlZZHt3wOcud
OVvok6bgxkFUmr2fPNbd0D6a/Gf2jWo4fDyLyyzAY7A+dnbKekTdD4BHEkkUAwSfgYJkYoewGUDP
ojj3k7dKb75JLB89hGrKQKDFCGmdesETp6gjms1f6wHjdgT96sCPoO3JLSksy6Rp5MNN5EYQ/S6K
46UQz53kIkWuewKotczHZdqXoHu3UDBQblyxxo7NVLjdvJdxener9Tfw6nNujpg6IgLO23zIxGTV
uFcHQMCWCZQiQNUeijdJ6AvnNhm+P3DjfEgc4dlZU4bYlhdisrn/XVHBnuwAqeMFXOxmd3oPhe9L
/eTGrBdKngCZuP0YG4rljDof35fVHbuANJruTKNgsDtbBY4g3HHYlyJS3PQFL32lskvhbZujOD27
LyvddHdJ7WwuaDioH915uinymcc5eKyLTb12h+6JA5nBkfuhEpk2wpaXVsChUo7allfV9gX3e3Yb
xa+HZ2NKX87ALcfs4Y3BwqX9tQLv0HxfLgEZBYAraZFqkQgZDVhZbTVFDFuUvX8PhZni5U6O1qp8
8jE95fHb1BBpPmfGIgU8cAuPNph4Igft+1P5TToPQuB/DSDULbbpW+sr8Q15ytY/IIU5mtkkNbGy
BMuwmzjquZ3BnVCwSH3Dp2SB9b9FFoZtlfZZ7jGAMU97FdvuATrGoMkO8rvuePIokLaIin0OO8kZ
60rvFoCbspmGyPpANEg87btfC/7p1HxE953GRcdwzh0CKxgtDD67qdN/RPaIs0DJzoGlMwgbpDBN
CbCOLaZC7o0RDbj53T0NJVcmr+SS+jf8x7QU8HKv8aOZeL3iVaPKkfFrfDuJHg+vJZbJ7wpAfd5A
3jmnvKwfaLsqGc7i6Duz5L+VgIV/gaVTYn3mxTqc9mVug6Tpi3ML7YgLYr+oBnXcIhTs2IRYd2Dw
WbYTnrn4nsRpWbEbJHIt1ZNyXsRw/c5rV4I7/dPQAfFHrm4i8jEan1AP2HCo0J8lgimcG6UugvU/
uNfO5GKe98o325FxZLwCl0Cq7fxL2TC4NgCmRvH6RQ5UwXGXyLoOt1EwAAWR5wKqxgjuNJ+CyUVn
1cdXnfPki1BP2iAJWum+Rt7S/oHEYkF99txBYM9QPLaP0wNeP2Vg6LoP57TXpVreLvW9kSZWe36H
NV07Ms5Om/1cnxgLhs0uN5wa2R6I0y9WV9q5mxGT7sdthiBQ/PJ//jSuW7J76zspo5FtSBAG8TrV
rAykHE/Ob/VsZKEf1IstiZusqISwRh8jvyBMw0M4cs2HiDLjFp44ypfK6YM3zJJJ1CLAHuRU3Acr
gBNLYTmR4kKgzL+JjiO5GceMBGPvWCuU7bdaK0vlOJ/hgFzcME3XOjKLX+hN+j7h4V/4KwUQyIRS
1XU3k4Zh2WHJDwyoAz8pZ+BfN8Q5BgLrYQ82b+m/3sB1kZVNZC7sy7vsabSM+ejfUudD3MMVyP2f
Uw122FkXLFujfYTNKPVuxxf5fwjwbndGPeuPWd/hulzN8ikdFzrlMGWBI62KixmH2u1zDnVqtZAr
jkPArEzouWSZQJSzUWtuePKAb3bNEYn258Raj3VrZdpEcbnMfp30czbLS+ssa4C1fW5R8Xoujg+S
n5qzh4awYKvlfRjq95lwVoPNoFOxEWo00lSJw5vH2vWIrhfLlDxnGRdafNC0PPl9bjey/5h9h6yZ
eC2YiB8sl/Z/Be8rkZd5URKtb44fe8mQ96Q11jWQ5aTujtFtLMlJAv7ATj4jbRI/aoBGQnkY467F
XKcbhV1mHNcOXjVklCu0wQumsj1Adx2eL/e1qY4r8Jd/tMQ06dq7HRM2XlqXTVzHFBBW0IkK4Iku
b8iDW0kjDTdqRyhvnsQSxZNJUdFTfljvk/RENjvDx52aWwk94mt//58ryy8sHLdQTgaPYhFuvEgE
benR1DNXQkY+bAiBiFHbAMQHx3Eqc9P7mkQs1RT9T9jJLvPX6WCGLW5hYapc6R5VykKPLXsUO8No
wAf0JzAsNphDUGAwiffVUtNPKT1eEvcFplxj0sqTpFh/5R6FcsxchjSbaNMJnEvdHw/iKNqWtFp2
V2qbdypldu7pVCZOrf+Z0klnC76rrLp+z+4ovNr+O17+ItWZDRTrOGQyOY2H2xG7Rw/GAJWTWE3v
VNpatJiwamwZXOY3ts4P0fOze7WuMWHM2E11oYkhr489RpyzZnFSg2jBDH+1F90WGf0qGk/02NcA
7YMgs2hyBf9GTI5NHH87Tq42W5FxBrawoRV3UkMAQgvZ+YGIkNXThXdEiuWiW8XEKTe+7X279770
kBrQbbq1z7GaRwLlKAG9WdtvvngGbdO8r3mw0ap7tEovq9wmbD320389ACqyfBwxKCBdA0GJGSzO
xph5HMux+bkRSzz9I2EpDstkV1+4muxK+zUnq/G6UK0G8zIJoiPucUu0Lk+0SzYkxdBjdH2iZgln
mgjdfWYE+cwEzlNkXNuw0tdtOgAdWCgd7xOo9kmf8kGZrSFN/ffShrEpCrKdsrf35ZQk0IY7W9eo
V7ThtQPTClvKDFSwe3Y5no4lU7Ju9ch9+qJF4ptzT7St6vArqFPh3yu10NjxjUjmELEZET5PAoPN
XgWEebFqtauvmv3ndl4CddEXNaZ8OcF6msqqyxHwNDFn0UZgZ0VetcdlZ0TOGBLA2ebct/YGENy4
wqwgNwQ1qJAhGMa2emJj2r/WsMjr5CagPjDmw9RSM5kIe+e45uEvN/Sq7QA8Grmos5E+N4kUaG3X
UUMZXv5gdDJ1J1Kf0Mh8mIJ0bq8ovhL2E6975lWLWMT8HyIplMzI20IQYnU7T/tRv/1wMGz53EQu
1lHqJu2T+TzAiep05HJ9rUw2vtx3NO+8sKj2VrN0+tn1EJovfqQjVFnrmXQESrSFcbNeX/UeJdhA
SpSr0+Mb0qz3/m5Ais0v9Itf0sQneERrzhW1KnpbVCkZr7BPMzoTWR4epkfnxM6HioPsB0fyA7pR
lwARTC14l9COI1n3BjMl/j8gqRkCuibjcbKmRNT/mvk/CqvozMt1yVR5Gc91Unj1kIgQ7xN7IFo1
rtyAE6QXrR7xxF7pW8SqCB4zYlbG91TwmR+Ah3po4wSIuE9+OwqeOrkdPSzn1dGvB50kCKBP8HTx
LafmXRt+h49CDF89+B1H9iNtmY1l0aiVMEPiZ7deIdNvhuGyeXpIMfPWpslxryC7sPw9vh8n5+DJ
sa6tpy5U3iragsz5xGe3JK9EHxVfnVfaWeUSOMhuJYmZC60uEZAA2Nfm1Kq7Zc0Nbz3deZsaUKN8
lyYNPvaQBR3MWy1PMTrRvJcYa/1mOr4XWN2+af+xeAK2jKE5JtpuzWI09MnkVudWzVJz+G3g02T2
+8fUJOsJPHEglIQBEZHerM8RFZP2GCVslWrk8nSBDnyLit5R3N6bP/e8TwAFrSyDM90zcYE+N19t
MZ1Di+6/ookpn5AGlXX0FssoWP7EeH6rfqjyVwVnH+dXDWA9FwBPpgt8QkZ7O1t6be+glg7+PLQC
xoDc6LTzHF6oT2qhpJS69Od5y3lg9Ze4XBKKUeRXqcmAfZk5F1Juvp8VSCqBJRvciay2vqRaxrCh
aaWJ9A+WZgHWXoFMnHBFI0flRBLwHS6N2by2Dh74J00L5VxBRug5Mqxg+cRRroU1KDtkwmPxvs4W
1d7GcKtGkSwo6PHD0ZjNRxoAlYKQ1c6M8Km6mDBIPStWi0YGu7m7NqZ9HOxKjYfsG51gtwEsYJfT
QQF65OKhojrhUqvq7+KNHxxYHLz3bDyorH+Al3DUZmHCrvuVNH4CUBVBZHLYm+TixLSw4DZePfEz
ZwWeEmlc5pUXThbl1SaGGzpqVpcHuntntQglYa3I/41E08KS68DJTs1B2ztL3Z/FnxU7IKqRuc6o
FK+EMdWEdxKPd/ogWQiEuXhl8wEWkucR+N9ZOg9OUalk8xcB+u4o3YOfa21jRO8FMLmMT1+n+a7X
V/f96bVC1lf+YjyMyoPzWLyYDtm/h5pWMAttegmbI3QC9PTMSdzHMPLOe1kNvlXEEa1uDm4djW4S
EV8Oi/K3lpSnGfuWqWVOzGmKB+C2SgFidejijuyTllv0FaMvnFOpLRh4PD0v5c2NtECk8X58kYHy
TUJTwNhqZ7YciVzoLCe6qBQDE3rhRsyiZir8eKBMhqiQnl+UyZVtupeVuHP4NdDtlRh6/rHZ2dS9
QoJ0m4iBvEdxPjHXr/4YZgYWYr4GjfzYHMGEujoHKcfxaGiR8B8+2tPAKexGfnetOkRJJGanXglb
uajxVPRSNLJnqF0UkqHeBNBIx4z0CalnLJOY+5XigHlxda2Bwc32d9/AfjejHrrz4KdGwH3OmcJg
+9akhlwyYGHPflsB7n1N8IkCXctlrBD0djN7HHvRreS7QOHkuZeM+pXKyxUF3yWZ5fwy7ih9JYix
53lSZOXXXROOmpE/PkKE7Am71rrc31oQNuCXaaDu2KMbsmF+OHEXJwHn664ZZpcBwNYpBYDv08Am
pz5esN4xV+9B5837IN+NSRyRQ6t+YYmsLK154nl8Zb3J5OUHanQnOidx1281Q55w6mJ5ziC9MqQr
MJVO+QP2VsgJX4uIsVjStTqu6LwC1Iz3CsY5qJsnbH9R5KBjUQo23Up/XeYkMyqgDL7X9QbHxwiZ
aMC2+N64UgrQtPkvZ9umi6MTNFtv8jsf8gudiw+mGZmL83xKbj2gJt9FwXxdo+nzHln/eAnTRVC1
gAnIJepRljdhjCaTvBzWPJAk8cWbM2tRSBoiV0UVJxaB6ndx5LtZtSYlSrjiSTHZVxlMCMkzG8HD
6N4rd8/gNKskQHCL29K01Dp48rYDEc/vp8eTShfeQjXFW2YFhePc1cabqJLRGOzWE9xr7xtdifi7
IsSdEPNuGDj5blRGIvuWeo4DatVTlA+c+epIC57V7pmm91vRxnX1BiID3LpbTYrrLZ6lgFqTzRab
zyRKTGEC48Xx6GL+f6+ueKoe6acTSzsP46W7InbTGO+/z2LQPbE+a+lobdvxeAvVkZWeaUIDSr2/
Oyw/yqZajgsSOpQnTfU1lH7OSksLBSu+AlyOrjYVNIHc3HISs8bteXhinWpyX4grzq+FLHPnS1RK
vZxjMXFeDJjPp9wjtQ/FhMbB3uXwlsQDZMEw5jIY4ukBK9J5PcZcx1eIr/vJmA02OF3V5N+/5Cj2
LdrD83LLREWl6OPec9BdG5pVtPqvJpkRjuk/2vpMKXAVR2J5yNjeCJnBbLcikJONOzw67eAjaLcP
z5Y4CafA1ChZh5P2JDgx1JnTzY6ZdjMWucZYumqytaDN8Bx3b+o4ROXjwTaWMrdDNZdq88uNk7b0
wnze8vsVBEtfc0LSQmH50EDMLMG8JXra1yy4X7tC6SZfd8VlP++wMXTTRBZyUoWm06AgY8c8FkiD
CvHJmgkiPLkkuAVSDnALmRoNNaSmSgUdr4WAGvbmn15ZSEbvg4g+lYTBc0AKVqJLmwtU/q3WoCUU
75kqi3UufACMohxsuZ1ae27AdR2UEn+nzIIXWeIRb6w0uzJMM9zo4XE6woIosqnW4kto4ioZ4p1o
IKv9xMbSF5uVtj5D7jsvWHQfU1UdiSl6FxC9EAQsQImluFXQadcr/LYe2UF044C0hImHnIVeCt91
U04uVh9vn9RDkTN33Uk074FU/6gWehx5tSnyCl5gPSyvLJtXQUSfvsSPhjvdLhfwI0xMhM/rZVsg
bwCHII1CzsaL0lI+UlemjrUF41yUoyAOZzAZDAcX0mk/3ucE2ZWXj4wz4vkV2QVOFWbI2DGyDZJS
v7Zd++BHlMRBLtobwHXkuq+gLUxWS54HYPpwyXqWOtFEn08oMqIc2zhdknHaKAi+uFZc1NLh/0Qf
ku4RbPfxrYvMjB1D7ZVyu3khKz10evh0jj77e/Is7dX6SHQ24FVlRij/gdA3SJ7ds0ML3TKOnzqg
EgqRilOIVbT7uuMBBgo4Jdpt7GcAx4JmUP13dnzgW1foyL/CN/AgV97oJ6Nm+/9+xZG6r1AwMWV/
FvAC0u+QlXISKZjxJJasz2ymLPGXkqeELDfF1CbqzjgOUm3PU5jpzqSLQW0PCjqh3XgoMyayixUK
fM3jTcHdrgMY4AWGSMnEmcudNWHF0fh3Soq05Vfezcl2BnmyGwz614CIm3xXQKqvHcOVvLWQ/vxG
cskGawQkVsI5eOaV2FqTUBiB73P8IXzn5Q3xD20xdurhEFZDgS+Qu/tznRoYs7SRBzPmGyfKjDTl
O7DryBG+RPYr4rthfQ24UKuaA3QvzSg5rIsvdzW6O/E6bwMsJtw4+Ngo3VKONo/32XuWUMCYu29/
pWyqt5eHoBI5unbRcxwx1zBoWLw9c17P4c6a5Dsw1iS0H0nZtgkcY3Na2iccHVrAqJ+ZtQyseHog
7SO7S6KJUZHBaioUBZ/zpC0JW1L3ZbR2Si+3RoXM5a6zMoqfya2Lf0UQBHgSTYMHbnZkzBd8m2jI
+miFfI+LNdOuCzp9InhLejPbLlqbN6+HIg5Co4Shi/hLpTcbVL/ER7eXQwYlnbPuPrWxSa0WghQf
dvlNEDjMIJaj2icKTecB1wTfy8wCIjrplZ6EzP3WhhRFW6gw1of75/QYklOtXpEhgJOmBMCnCAOp
jO0WuYF5m16JIZjV+HVWC8vfIkKdiHTusyJH8Pr6jGP1wmGuh5hiUTlQm/jOd7NDEh/mtZRax0N3
Ck/9wpvq3JswHDY4//PrWJ1lbJkBBg1sfg9qbGd0pZ3QzFQFdaITXwYSrePSQZaLy6RhGMlChmNl
FN272xcO4vtKQyBkAvS93ET80P18AoJFhu1py3IdwUZ+syqBOJsicxJRaFUzf/oryo2EZddWZyTV
38GafLV5lyYEAe4Hf3o7Nq8f50WBiWXWjIQNSmoQ7jV7dJVJ8RNeebQJcDUfoaT0Ub9zTSUXi13v
IgK4bBoC34BqAdxbC6ND2ik3QuKhaXoZAT2anxj7urYunoyGT3AjxSRzUWiHL4RNfv21YQPDKLqe
KIsR97yYagQpj3rZgzw0eaEm+5cp+U9Y2WZQ/9dMpo4EaxN1X4yxSZVx1qSU9yFMOdZ1GMTrrAc1
2b/LBgilTPIqJZ9cLpW6+m6A9PzYbhtcfZoe3TGdGDDxo0HiTQOxzPESWVxKOjr/aaBSt3WW8aPZ
igKr04A9F4w6PdO9/6hlFc25crDdy9TBu7YpZ8kpNIq4dQ/S40aluFc82BuMy86prGFQMNiQkEmh
fqExIM7JvA2dprLETeO0d/q28Zig3GUW+qO4H1YNJe2ekuph8pi6/uWfx1R9Ry3KKV1pYdS3pDAe
giG2l/kra414/n1vxBEpPu4KA05XN7wjlg33ecsuw5cRLgVpqOACigrS1Ch3Z8Hd737MoQ39GOyi
e6nQs+sEAnlX2IX8+t36WV4Gfugm60fER4Wq9FWIQ81n81ICd9N8jS8Lg//OwyHQXSkHCq0/JZp7
3JF82pR3BiTT0Nvv8HlPsU+y9y3GDkwrKeqf+YJjRT+nr4P9WtkDu0RmxauiDQaN+Cky14v/2U/F
045KyXJjG3IMk2xnjUvjk4ocFsKXC/l9TYcA0l5GNsliWIQKcVm7Cq5zRSyih1ZfGy40mAZ6pAU/
Cu6cv5N/ATaDMNj/7Y1XmO5L4ugSGWW5BZSIMQGZD2apYJdzDAZZZE+8zZcznTiidEbt0fqKoAFt
y/elUbNhc1YkyFFiWv5odSKmRf3AfI2JqMY5ZHwbbzjNKZMna6q5LYzyQLORVicsnEtqWe4YpTSP
xtrD8BYY5Y26AVm1+2OkVEwPbXUBB4cyeV161YX7x1+A5DoxF0PKeeg3VqHNFkUzAhDfuo7MpjIk
QAV08jmMKsfwoJ4taH2kT4YcsSqJ1hsEB/HwHcAqfd9VWrR7y+gIlSdcS6B1wvcEkojv/i1Kw5jd
wPMLzXJMEtSElC+Lv0k/xpa+9BpcOP+OQ0F/CEiQGPXgFrFwKxVGN0rCCbJhaK3nvcGXupo3e4kr
FigqbENOlHtzFm0UtzS8WhLrWVsnP1MFUee7uM8JYgL/gZvpMUcP2mamhWZLQaneDqQtH/gOlH1m
t0YRTizLFb8DTQYmc0aqMOdvT21Dyyiwd50Md3iC5QM3i0mbGSH3b0Asm0uV0xgR5qrEMQyrDXXU
6oMPuEgtLmi8ypzEz1jpMSP1bxzIqRtOF6pGCHWIUUQUeESJ2k0GJ4VOdSjm87H/prk5rewePMVC
06ol4OOx/WgL/IfzmUWSm6r1zMoEp5BRpvnJvlWmBQSjdqPVVLK7bPx6pFZ8kbudN6X7HEAd6rs+
HWMDRONocBsqAZD+3tp4zStxKbdIiKFjjm2/KPnn+Cx+7PkGJKp/0+fhQvg5/fgr7ZEkPodZ3Umo
sETwkPXjygqVPJye4vvM2v+yqss9kKg6VVP/CZ0kF+eQjuGX5yz8Nj2U1dN9RUHXtFUCMUkufmnt
jal6GOX7tSWvU43rdcGXhD++LeQQVcAf/mQMl1LQ+gq58HMOUOcJEeeUPkJtet75i+m2d2gYig+V
ySvXaedJ9y+32YDWhzYT0P+z9Epa6EVqJroo7lYB60rFNt2B0o2XTw9y7f6ho+Mm3aIkbAnbuWCU
PT4tVsWwd32bGY/ARqIRVYKBUH5SFSedn75C2xu9gDqF0yo0iciDw63ZkLNFLeuLLlkJvDBKmnPL
Yh6BCUEQXzTuJe6yKGKw7BIML+xyK/b/uYvRqUoHSG5x7aXbvkQ86S07jx/xOTOjUgTRE050f+Im
WDV8b+mWOHBukXudTTXsuaJomhzGI5TxoJNCj4V2UOzzIUazMTmKjtNpXsaIXe1HTW63vKqjRhKT
VKTS63ZnkYRaD0stVyObz3PkRXDhC/kHLbFA1VJXBxMdi5vpKYUeGPZUMqp89SZ/IEkqaCrAfXvy
ZZdD4NEHVy/x/H7gpo/Dev+zT3N5d9ItK7+RSTnfV9X1+0MzdYPDId6rCeWb4VLhApJWk0CtK8AU
28KENah+8KDVOi7EGXUAXLGxhqaWVQARAqDVf7CtZyw9sgNzt4Z4KICsRoTG5X2F7g33zzCv3zA+
nr3Ig4fkB1/GrBffii/ieyXscuTmNi9P5wqFhAwmEUHxufOtD4dCHnF4z6acCSQ+mCdI3x8uKbbL
NUtXvsgqTN7benV34b6MA1OCH9r2CZ6lF2d7gKNhZez/pMQrC03NpXs3nvG1vixc6lsU1nhk1Tw0
MqRBArmZIiII3TwdsJ1rhmvMduqGMAVbxygfOiVVfhv5BIKUtEtgyMTQlpjxgZZhVqPJS0DmmjrT
JXvDELSS6Lt9Ec6kKHG9NUV4Znv0nlnApMzgqyetUsHSBpB81f8bqHHz0Xf7q0tFiPsg/ZEpLQ8k
EV4Qs/pXfCR1+fRyfb6uHeJ2m2L+MyOitQBD7TqW+hNxr6BfNF8CgoxzAtVObwRzV4jotKsm1eVz
4CmNdkl+0Ix3RX62yAawAC6yKndHOWstHNV5gzzSK4wO2qIG049E6KyuAQ42Xdn6Edis3JGOUaz1
w2nNZ4o6gF/ZFSy5g37fih120iGahH7NY2E/wM0XdJH/AOqRoON7e6kUp4wYL1JlAmW5G1BcePf7
FaS3GI446ki1cCUU5CzSKTS+lAyqx6YoCwDwsYaO2JOzycgiLQL+oTeV99Nkz/SFR/WohDG20SOe
gaI5RyFVoksaKULWQyReoR/Ay4v4O1FpupEvn+Okzd7IyyFag5w6fCQcFLTnHra3x3ditBUwjq//
5cnwwEnPI1k1GcjO3IvERcH0m561hmIYJWwx3wYGEkS5xMI0B+s15I23Tuig1Ih53xRpsSJWrE1J
BvsVVKG+Ktx+4zwU5EQOY/Y2/pdRnSckP+LqpBUQK19zVL7Qw2oscw0LGEiUMBH9FSZkX8lUbziE
j0gRbHzTkz9zeUlpWMgmW1E8L5aDjxu9ntY1obiPhOr2FB2MfTk/KwC3Pz6LCM1anODqoFM9qFpk
4/lMLv65JYfHOg9WtbBtvMY9LO46EkL8T7RYlZskLwRcDonv4m6QO/0j+o+d7wOfS1TWctDx6Rpr
HvRLKOf85mC+XXmyGhlTovgZlnzje9kUdTb4ibJTrKTgzbL3gNC3resy8NFCKmiAoeLY5voxK69Z
HXfqlgvTbRI+Uo1sI+CWLBttvKJfO1S6c/UgH3W9nY5bPs5vkEkiIFPMQgZt/jX0ON8IpKb8sY4c
B5lJVod16akIItLTfWpjcKGrGZ6udTWzPZ4KtU/5ddAM9jOqVUPzSJlJDrLT0/3uo/Mqu7A7ryin
vS8xKTZOGR6DbpZNfFizg1an+FuK04DK3kPOebg8hLhs3CnYnW//tUWIMwymJmCUSYlBlORAKQfe
YbZx4XhJihPFmzkgPapuj7SfcJZsRGm25tY/GbqdXj2NrS6iEfyhIF3q2q0ut/aGLl2VSfV5IHJs
znfM+elcNFImJSLIrkw8as7JGhxZDHKAPioTyj/YneEPc47Om2PmelM24H0u/yzc9pZ20Czta6fy
PArXKWhmAL4h338wXUeqDY+BEOfLiivsKcgBr56EdXK/2HQfWRMpD+nLWA92yZ4uK3Nu0OLzVAjg
5H9jXLtxX7rI/zUTdUvrPlPpUlh+KZWXdKVdEkTzn+pucabtIRwbbCl0gAlzxfbeV78rKYxS24P1
6k2WdyqfzCUET6jQEx5Ua/wwBPkZV6e98F5FDbfeUiPtZnGMCnt/yGZ6WRoxNAznes/lYg8zek1M
XGLrgY6ZkctoSv1nhqULSIHJBzRgdlhqMvf5vbN5D71N+ig1nFFCxcrbdPlhayYmHQKAManljulS
aCY/jgsMzSl3UUgQ43QowzJS1skBhyvlZHE5Q/BBCSI0syt/NYB14OGxXQmnc2c/aTLAJIt9VMbL
FtV5mEKVSWmZB7I7sTaGdX5Y16DPzBHp3TpabQHVKQ/rsO7SLkgPD4FfL2O8nCgL0tBB6/IdIG5C
fOB5heydFZRqSMvE0CMNWKLXH+4Y62zGJkQjNsPhZxIDM3FdtpHPMcaFe/2L+0TtsWKEaYgIcg/2
7fYIt0S+GV//rKQrzwPtuo0MJoG/oMI3jlk2E0t6LM1cU0HhgE/1ypRhWZl5SmlPtSlJ6tCEx5EL
8n/adsu2hIGV+qTLI/m86n9jaZ/uRQtqPK4ZFUNWnljKqvTVZrZnFJ/LRoWT+zKPJEtiZeVYfL/0
Pr5VtrTJHeQzV/+c9LFHKWc2GQSPSJ+D+WFKrv/GY2mDC9OsK0YHib+HljDGTIl+BdNWloBIvMml
Qvi5O05XH1q990xN4h+4RzXAXuLFHLqV2A8WcnmmHbT3PUeaRuHS9vBpCUAiBXZ1UrZ6KXD+ABqe
bxvWxqnHJzf9z4kcBrkCmmWdSy6WVYyezEzUOkzzVK5bl1Pn+3oteEngg5F+vQ6sYBXaJk/wDKPD
K6Mrvm/Cwe/lWY+A7Wb3JDJlUaTFdahVOgd/8LqjDsgeTjmuPmF5eLdqY1zoe3dSzcJL3hnySCmi
kKpyCKaleNGgYeMlZtbMtBec4sxtuRbnCnRcyfC2TswSoV0iEbNTyeGGVlEEaQ7EZ8JVLvBBDpuj
2vEFOvCfhMmj2G3gMkZNC8km6DafoAGmcF8Fkg5tUH07Rfvkk+6W+3O8kVvzvOgkg8pbDq0gzOp0
2ndowELdt6blzs4Dd8bevzxHifaItWWX8J86Q4IlftPx7H0XRjxIxT9vUWhBCgdbV2vd2XP4HbC8
B6arb5+LkHhp2uBd9idSME+D+rjNHiwK3gQTUidJkpMxXZMEuFp5TjsZCNj3TL4S0TPLkMt/0D20
3xjZY80NEFuAQLbm2kGL33JCwf9OTShn8FYNGY2fsewyFEZagM461H4sMPvc4EcOTjO0tTwzv/2S
W83q7M+/eHe1AcfmXOBnlOz3LN3LVtLCCb4XEYzflMLyZI6aU/0l6EcrlmLOFXwUWcw8o9zkOJQx
pTeKFCpRXXcJeO3Lhbfs16rZ04Z5X+5bHT706UygnlOtnLuD3pbmI+PHHtHFLvw52NG2JdT6QV8K
x6YanPiBkQWiOL2KQjKiOilDg5zI1tBIiTxdzVmQaeAPpSm2YE9wH4jumXfPlt+o9JLu8zqqMcsO
x6wQqW+uMcjQtQSNSSii2bN9iA0aagNslekjvGMnelwUdDZa4vW5FScPTxbV+i5plPYfYmjByLVb
KVGRkC3Wu1zi2XTD/PPXDo8zcKdB16i0il39jawQZnj4A0fLmGfykzCD7c3IfTOgqd20KgRH1h7c
S56xU+k3PJjehQwdDjKG4m4TQSC0giwxY7Nc8KpwUaowU4zrzf12Ilk+J5/QdZJpgB/261OoJrzD
NupEXJUMbi3ddPDGdLhPle5MlkNPdENDqCm5hD77pYjfSeV+jTpW5Lb/WjG0ZjHehcjZ6eWK7oC1
wnu3MHYpl4jnOeMSijn/s7XHa5Lajn72k982gPGmVFhSn0zakk05CQmQEhQqbXI9TlNV8NVK0ISg
0vkZ71e2ZX3+VH1fW4kw1eozbEghtE1Pl3N5lHw3+OHXdUMSvEMlEu3zz94CC8qKHnVIYeqV58bD
MP0GMG9ioxUMKXAsiIuM7AnByx0tn1nNq0BQre0/OdMRzBo2MHnrlosfVcb7tD7qi9KHx2VinJCj
9j7G7W2hvrm5Ssgsv/daTndmX9grtQGnA2NWclAbGSt4/4o7f1XtfrvwjgC8zr6HYKiqt7OP0Jfm
HVLbAy78DFngkixAtFD6pQk/7uQuIH191ybTFqyt06GTchpmuN1HOX25hPSBV8JjSPiLPZDSlUEg
3lNbEEF4F3308tigEkyXCVzbEOJaTWglSq0k0obRnqAIhG6c1kYsuBYEuEVJv0qdTAIwD1BLOShx
+BaxPLDbVD4Ww1/e5GFx7BoGPMfvaJrWPqzYeT25nbk4+urDWPbj4915E4zxQwk2jcqr89G6Zzx2
99ojfY53YW+2dxKjvZ+FAEete1Y5LjnyeqeXG95Iu35tqErZN127zqsjvLTZH8h/0XFycdKSUsXN
Rpqp9iCYYYEh8qjNb1IjGZByBvt51jxummWF2FkEbFF8spVi4O3cV2QgpBmK/d4HgysfDHbc9Sfd
Y8Rn88egQ8tYKJZiRZzTyeyfD7K9s83EPM7rDwaTfmdQlVm9h4Iz7rC8ZYjfDRv+4T2YuTXfsPCp
TxwWGH+9y5vGVLu5Dj+JBzTaFyaOKXOE0VOelLPomfOrxpq3GRvazP6huLXVvCNxQyjsSLuwvDPK
RCeLqXG9Wgzx3MBO4nLHR+/HydPkR/KpFJyDHx/YnQX5d7ApzCGQEB6qau6oNL2REpO/74cZrQAy
cXqKLrxRUYTAnEWY+Uu0bNWJAoc7mTH8VUSR2AcoeKXtPZCrwDb6S8phfjzo2tr8XSxSnVcAbURc
gBQk3EZ0BbvpXxZ55FGURLKs/aN/L+y4KDQ26RvuMr3QV2oHl/Ah4LkPpoMustb55O7gXedlD3fu
lHpuLD3gvqcsHVrLjzKaNJRC8+Ov12y3Ecm7moaE+jd2RBjJxxRZ1X2ErIwpywoHHBAygM5AWP7C
Cz7R5rG6YKS2Ig+zxzGExc+zczAowCMKdBtzG5aw/lLLqOQaeIaP7nlAE2adKjqkiI0diXc0ScxG
bt6Bo1ntfqurltcpBOtZ7qUqcD6oCrK/jGZJAa/fD2ExcXcAS3FuolTzxUhas1aJf7qplvbqJ6B8
6QCqtFp0j4jGz9zxZ0jTzGwyZwdA+jRYi6tFs5jnCIueAI9Yh3lIDGLiRf7ZnUbzSEVp2byKl/xd
TNbKEdmXnHOuXQoZBfF1+2DNyGsxp5yBo3cFcfAC9g8ApK6NVixhWTAjXo3bzKbh1aBxIQgiF/Vk
E0puvqDRNvok+nvOIY/11MxERAjTbk10x44Vi94h49TIRdgWIFnDl4SnwBrDvz/DLrQZ7xyj++tn
o2b42A5gvFxDc3FlC5+7YiQvEEFjPKHxJFuyu9LSOe8zajH5gCh3dAJ7bN+ti0Yqv7ccY5CoHax6
csOBLTsuMSFMCdqmXZ7gtO2vAVlDjn95FpeaaG5TOz2DOp88tdm4zWa5p+xd8Z4m8HmFvQ4EBq3U
tYZbshyy5ETIuvB/9lV2gyIRNaDF4/A6Izg1c+R8sdyfNE4ClHxOavzGsqO4rn1+ovO8D7JNTrjf
XDw6/jOZ1xzH5eK5IsBcV+YhWjkpTzfR8PHLgXylns7qx80147lHBbrwxZ15JQSPeUrTAsajSVhd
uSl7iJIiOu8fdFFuQPqhmC3WR1tUd8jFjrgeV+L4ARgZLQbq6gmFbL7677F1pp1DY2iHc+oWRUZF
LJK3YuJVbzPF2D8a+wTgqZ+782jGYOkxx4S9kn+3w/6CZkfXLgfCHQelRqGADpO7jxuNiQPQxhnZ
9sVaGW5Bxeo1XVY0CxbNn7iH2KKV/SygdseqYCyfrEMwf4yL/Ho7MrbvIlvchKrZ6DnRFwPRbUQG
A+1BmEzqSDL1XhGD5Kbhz3kYM+BlpB+XY2/B0ehUIzVdHa2IxTOLw6CW/PzTY+WwhosMgguItGcz
T8WUdIb4bdV98kmibFBlHfFPyIyA1Yoh713FgsPiDEBQNgnvvee1QXsaJkvqk3qcTM/0BWy/8NAz
Y8QTnRqD4A18IwdObrIZCfSaul/GQqDdKkCJKW8JwiW4wlpJr0SbINJPxo2PdX0NoXcVjdaD8cZP
DzQ1y5gE3iTfbQUszQs+3mezg+N585n0fqudVyH2yhSnImUvroJYDb3nPhTfPRwxgzv7KbtNrFZb
CowEmZecl3GnN/SJB6Y5TZTDmoFGpBFDSPmMvfrwnuTHrL0Ybw15dAkviJCIDnlLn3xSRn6ShEGM
f6ubpXU2fVD0h0FJA1gbcImlpWttfe1uiC5/7pFaAm8nkI8nFlirtONoFoAMM9nYhsnP1qXB3QG9
wuYQ0lCH7pNuAi26IZGNS2SodgumxhZ5+x0ehhUk1s/2ePQV83auhK2mAOJ2vt33xge397c5iUec
u6d2a7s4NzQOpJ65QK0zko/L0B0pxDyjPg+XYGbsGW7lN2u/ubLNEpV1KE/Rh1Fi2Cb4ZFFIqirS
0ZfSHEivAjKz4GZxRgOmVla6QVBuAqUlRLkD6/+l49HcVKiOqrtq8xd3sevmtViz4F4PrTAIXboH
Lb/TcnXt0rwQsHT5cHl1DYSz819bVjjXGHaLmVD8I6Uf1Y7TWT43WnczyNYJ9JMSBhNJ1z/G6vUt
sfZMbJJ7j7e5FgmpE3gVOgHbWmxNc30dR7WtB9ru9fsS6VbN9h4XvD/b1TMwaoN8n2x76oI6nZ/r
mBDPhnk6cNmfKXqEQWnUeKs1z87Gaz2pV5e5H9MPH4JLUVvDvJawT7FJcBXsV+SytjLDEeOS2bLW
ErFinfRki59Usvs9bVaEeGIIvqfX1kV5aZVpoEJ4DEPIvXS5O7KM4ywZ0yS6H2sazz0FzhTMDbiO
wpIIlEGLMXXAkoZa1wZ7WcBVobWeaY+2Rsir8F7lYwxE2ME1En/CAylvUUYY331Kjl8qhIQZuBtY
9qA0qyMw72v1VaH0XQQAbODujtVctcT5r+j6NSm4eOB/lqW+UfFrYUxw+GOeJlVQKbHXFcg/+BUA
D76t/hfssj+JQMvJeNCRaUyQoD3c7LIug0/ShKtsTl4Crjdc9IcAogEIONAz1iKubc7+CZI2JmTE
Mn+9wrIS/HbeYCCe/Y+EwAUhtUPz9RITF27hd71rKNUkNx0JymbmdrQxUDuF2XpnlId4/MlCu6vP
HW+KbBTl7S4uAbnNsxiISGfuk6RMmsNDkZxwMaC/FiUYWnWjMjYmLTemkPhCdB/gz5FjCinIBJUG
EAxBh33652XEwyh2Gn94qRCJMq0KgupNC77iwxAYYc9JYwSSAGI16EnGhlZEGXYD8wkiMG7itPF7
Ap8bOKtekqUt3lba6GuBnPU4GUmD3CEfFsScJZiF586CeFZ5/jFpm3oNm1nka67pK9SfNm545Md5
S49A1Xs/+GkdegmJ3Gv0+F/N6Q0Ii53FI7uXaFrqDlfGW39lf3XZUgXjvM89dsNZJxaGUGravzeX
V7ez4NJ6VStseorc1IudzgFeyBe/hJWrP88O4q/Ix3yZ7nzFj7WmXozsOd1dzd0CV0Fy/6k1HEzP
9KGCtic0SYQJlQjqpGK8h02XyijweBkPvFNIEN4e5/Mzf9W7qJXvbfo0fY67gDQR/zCZMqAumIYC
JIocLa0G4oeqj5O7fHlyva8M/avFqEvpjvUjf4Cudg3bx5PC1xQkB/x7o/3YaFcbGODK77brCnoz
CKCbv3P+C+nRf7LCv1eN/jOZYXiqEVj99m7Z9l+RpWEEN+YZQNZKJzo9dsTVa0lJ+xmfTl443RH1
jbphTX7+MzU88MIDhj3gf6iNKXOUsTak+hn2GzcwVuibWAciM//HTWy4ODv4x/9RkR9ttqiKnzpD
hOXMNWMGXEHsw6gLFYuFWgOapImJsbqjy0R6QJ5jRNnlHzsaD/r0jg246WSzoxXGQV1GghPPd7lP
FWsGtU0eBnvhbeNM7vTtD6BkpOs6B3u3cSFpomKGLAFGC1cJalbGpTzBtkMkruc+G84tsb8YUHXK
V4/yjl25ud0jpTQ0krXj+YK1T0R8o8AA+DLhK3yue7qQbGT9FV/QztVehiZSbJ2eGl4Y2vZmd+cE
rqTW5Os2qyhIRGhV82W1EJ1jljtVIpCoewUFcXVyA5cCvaMbaR6Pi52223MoO8g3NTefrYtbCUFk
PXCyWqj0K+oZ1TaXUGCS54NtWxGA3YdPU9LlR1aVh5kxCI8oi2z+/sEr5M08xze4X9uizhjT4a9g
z7vaJ06gh80wMCJou3aM+1OdR5Q4qwec4m0RBuMweZuf8sK35v9auwn0G/0qRsY8mnGVb9IHouwp
YOGebLjV/B3Pmr2iR0s19TE+IxrntE7KwjtG1OlvWvixRo0xfQsg/EEPeiihbh93oPl7Z4BJKghR
FwzNW4l19r7xByOWR4/3qV84K378BQGeh7bxd4Rz2+1teaSNlg80Y43n3stUof8OeolFc/l9Bg1C
TXeqNJD/1nSOcfG3/59CEA2jcoOT5tVJ0KRKSFCLat0GhAwLPaIe399ikSosPSXDj4SgEdl/y9Pk
HzaZTi910Aw5Vd7qit5LJszYO+DoWS5+cBw90L2qNI+DarKR72658m+vpTmiIvMBXm+3te1hXaar
vDamTeB5iTnVPyiTC89R7ZDI/G3dJKzrawR68gjDOmbt01RvV/WN8HqWS6BXFSKaIInlGp9a6xhp
67SPHcXJbBv6p3Fw9JA1CUWOEVtUGjLiabfwgfHrUT6r/DfgNgFN0mGpdjPgXxESRkPujTpoFtg5
6Je/z1951nBaN4Bbnv6/wQYThOIf9upp5d/yiEBX1QR5P36VxMjfiAFa3jQWS7xBF/f9P260pYLE
hsYY/R+Ikf+42/rO5N70ntOqLK2qLNOTY13GXsSDtnqB22Dg8RAEy9kfu0MzznnlbTe0RFIxSvzM
ljV60M/1GZ7b/0fOJarRYlfrdAsDXk5EQxrK6zYdb8W4BrqRxMzljqL699tN2egGenG4i181cmmq
lfXD9bouOoqhalo+cciMzgoYBcruP/2S+0YZG4Gddy4Kze5rp4npcjpnyQPXiG/tfoUe3k+1jwtp
l4PaON99WAnz91aWhuT6chTmMOw7QAgCeXA1tlSOLjoVw3QFMByapbIadRowluNYdowVVjsqgWaC
6kwsBANTCheHuM1eL4Pl1Z1KK8zV/IFwR2xBvhe1NvoMv2vLcw89nMmQQTMuIp1QqejOmgRbibP9
jpio8Hoc/5CryfZH7NUJN9rlmBtNS93kyGyBbeTOMQhRWJLhcZihnHT/VwEeNuh9PnYQ8DN7EwLt
J5SFTh6Gw42NC7TQc6JgiHpJr4x4nKGIbzNUBFH877tPOLsCFLNlgYP0pJH1q9BfI2M5r+MKTym3
p9K4+xvfb1WcQp+957B0HHlorVpCCVAp2fcEJGFeFWQddxVp/JW7YRxoK51DH7DLtEqTsCboExS0
Hv2za65bhWQ2ctiElFGRONjnbpkeVE86thhCiSxd+6Gz+lw+e04DcSffbfV8dGdIIUsX8Xju3TD1
kNWEjI9K8Q5SAHP+xsgBB5qrVpgGdbnu7Ya2NbB285TKEx9ZB7FoPAfoVlY44lJlbTp8avGdquZ3
GAlhiDeyEb0mrQI0Xd6fOT4iDPSdqp6zi3aKDsIWbnOVRhLpX+tcWmIUt4P2uSutbnLGAojSEmJx
hSAKC8Ymhz9/8ppg0IZFxdNWL1WxF3vGgT5jydoHu+F2a8kkGCrAjNXE0KjAFKcFkwlwLFQLmd/P
NWyMCdqOmEeMvIbapLE3yXBD3nQIKks4f+xNb+CwD7879n3QiAl8z9jCdM6uWMAq8yA6XU2nL0J9
VjuFmbFEXQZYUmUSVbjjK3YobNEuMFuTze5oigNsWMwTjfbRjTYIBdYvIv+j/KgPEScPgsP2a1Jw
gVZJyBJ1hTac4eNq9sp7WeSU6VjHlM9JIPbmykYcYmxAOWxN9X9lrBnW1cduqmhzwcv4vnkJPrxW
vhuq8a9MqblchvlmyYL+833t+NZmUge5KmeYLt1ZP6RsUUuQqaeL30qG/sOfk/5KZUrCip/PnbQW
v4H0pzFrVYnOWVCIBJmT+FabdyKbniZt8w1rg5TGjKCdK3jsUcVa8azJq3dQvBWKP8oMufl9NiJe
g/uZXfaTvThoR281IRBXl0RfGaf3g7NMMdlo5uFsPXPrfwMtywjyIMGzPG8Afn/ibpNgCvk+GDj2
CiBLmtvwZ/TBa5z4Otk0izYaewaRuXOGT3ceOt5uuwJs0i8BndiDnJDDBatpuOw+coiTNt+jG09e
RKIMpGzjl02nwwG61hglzTl4j7x7zbZqRUnQe6QwwOrx1lNsl2PFxg5pGs+/4lVvM7aTL/sXpJ93
nTP9tg5aZP6xhf6AQr4FijN6kYaOPWHImTXI/tAjNBq1FuSf++rasNihsDGW7bizjBc3Doey+ON3
x4X0WjAbYHYfMDgrpN3AMZOFNsGSlp+esBgiTMCSf0j8HeCUnxIgOizV5fh6BbFmymzItAq0Rn3P
Z5qThabQ8dlaOB3CxAVaWTRnITEX8H1655R93kWCKG5cFSHAixJjgTgu2I16SHH75d7miy0bgFhW
wGXgc/LKoZkYUaM6mF/sZQ2PZ9NFu8WU2dOd4sqXWg1FKqMfFct1b9GCLhMeAs+4ShSjgfaGA5sl
k2ZHzR7knGg5lzJCYoXp9pt3sZnOx+dLIyvfbwASO+SlWYeN1kQQJfoDoOGyJwRZ+djZ8KPitKWO
4tswncJYsazlSjuYG37JWKbWR2cDj+9UNMggmoUKSf6JhKhOFIZ9Qi7m6moRn1R4BnzTSle7Rjp/
OUS1OJxtqearVElbovWNF6aQrwNTWEEZgoxntl127whL4qxylPs3nANxD9Vk4v4x4cqEY5zoBsne
MqxtiJCvUBaNiLgjehhkOrYf+8cJfRFduyO5vx2Vf3CWxHSuYKnWipspJb8PChgrAcgv9h+ygWkJ
ztjCLDeRFrR5r8U1x4V0MdpOv0WdZLhpSYTPTs1mCBnoI/cfuXMfv6KAYoMkjU2Y5dAo+AkaNByT
C23zQ8RoP3pK3LvW3ivd57E5D/qb79ackMACi/7mrwKsuq9OTXim63OGY/qdRoaPeX36ZsEINPeN
tedNWKuk3X5RZRhJlV/CBvxE9E8qCFptrB8XjcUV7A9Tfsuez94jQbGgkstRLt1GtxEUOMlg28dD
T6jJI/HrVlLc4pXg0tqMg1r7Z0ZCVYSjIRXQa1jLQhQiPAEdf2t30tU/r+TwVQ5cbWKi50CcnuPG
1pWq9xLPmZ5WIZZzl9JGlMoNnt9pymV1H3oXe2tPGP15R+SDlnWrohZzfWOMotqQ9T2AV3avxh4i
P8sjUH6IhiSxB8EWB/5LiAuq9CRJ1NiJoxYgSMoh+3eAbEYJ40L9gCtg7nndSiK8t1qOhuAn8OGN
OfDI0rBY80M7xyo6a+Gb5rsh7MGJoew8JzyTCbM7rtPlpgC89RoSyzkXr818M9sPb6cLTJnQ8sDn
ZLo66uf/7myhLNxvSX6y01vZUWNRG8lqQOK9FBKuJsSWBFCtg0j2wy7CNk7pYLRiwzkhpdUs1BsV
Q4Lk+uKv3BnkTpubQztzKe872+nemV8BUtp7GfjWo7GJzRUueWLq2l/4zkv6VZrYqRVrsHXwpO7i
nBG3q6YO83s9Ja+7q/gW8y04eRTRIu6CYfESS06nl/IHLWy2RxI2NAEvQWJe7lnQP+3GFusXH/g6
qlVLv9dCT72LaHi/+vak28y7QNc1fDKoE9xhHEazwdr+bAfNqGOra/aW5Vuj7GZl7TkhDlpxDXrY
Mpdc/P22Z38yu+nj37tC7C7e0LYv4/V6eWKJWUg4GMhmIcLasQ8hVu0ab93gIft2KwDCIpomQb1h
HwH962T7V0a0l2IzdSTCcxcM5zWt8i/HjFtsIvse7uLQh5iM8BHdG3BgGF27qaohvtGkuELctqDg
mVv9D86lGpkkUFk+DBfKZRz92mVmLWsfUP7ZdzH+RiZztbI+TKa9K4TGt5etrcijAtPtOG1sOZIm
tMZjvuxad6Xc8kvWoWPEQ9EQ4ry7Xo9HP2NSQOMq1SJInZVzucwEF9PL21VIR/ksK+L4P4ql4qDR
20EdttNOHMqc4EsPteDKfrhHbrIAS6kFyZpw7sG/LJNHTFKHfeMK29l9NqpD77giWzUbpWMHz4ID
tXhhcI39mG2gAajoJq7V2iqlbrWqxgg52xTBUK1Z80VFVFi37Cr3x/cKNuBSohaA79P7Xese2paJ
iGWmNHoY2WI1n+DvB5yZOGteCYizeWw60ypSr1/qUL0a/gFHH7DXgaKwmWEe3uOrbBhsqTHfK9H0
z9Hzn7H7U2Ymx8ANVG0A7QkmyI2hHOV3HvmNXO9G5KMcxUbrQyFxqEUS7edwwdXjPm9VeJFCNjRY
q4Cq+jz9WciW/1IVugewLDdUG872aFooDns3SCWR5Ci+mkCltYxBVDIF81kj2Xx8GeaSG3qwGJHK
NnCn0YPGuxXdTH4voK1G+cXCK2ENNH7zeE4NUYS6apadmOlK/2NpB7otVIC58n+mbWf9gtNlYISW
C08dhD7OK8oAPSfJjE4Caohmm5D4m93JcR+zE+xH6fg0XM0mSSHjIxqV1XqdrUqY0qQESG9da5dK
5PBMeTqetoebh3imEMbWoCjXAjt9TSqBLANUiKZzH4KBP5V7pPVvkaSFE/Porh21Qe4HDAu6p8KU
sjEthd/2v8688fFWu78Pka6vo8ghh3mMFm4yaiDn7QRcDzMqCck3ipNM6ZFcSe6jkb7wWrBOmNLe
6rfEb8XNJuM82cEO6UmL9INLQCoE9AX2oriUZF730mIcjmg2HRUwXqc203PkJnUFbVXvQ792Q5us
X23AQnP11hmBHG8X5J6LFz8SEp/a16Hd6r4BmWs1SSO6cBnallO6oSKV2nui4BUER6yNbgin07Ny
KVCc0MuK89P9Eco/GnfYkr8kI8hb1aPm9rQjJP6UZY8jk6QsO5Y87qC0D45l5ZFCm3hw4C1oQiOC
8l8zBAEqaudNPPBx4B68MH9uJXtoMruLrnicDIkh2nDoSfoSnSemk1WHuHxR6yCodtwaUhGwcfZq
BdZt4aotbRVX0lwzw1/oavHKbtUvfQ/EfhF8cmZ9LZIXniSZggb13ZvdesmDhQBLkuP/ESFQNzWZ
SFMBa5BYlOL51iXHKbKNhjsMx9II7HKtvP6c8ZR2EPT5xMyqiIEZJWWzyTl5DEWJwG8kZG7HIVkH
pbY7IEN4kZP8z8xwSFClSBe4THj+zNBRvq51Unzsk9/PuDy5KCipvR1tCFeNw0g5LP5ue0wQj2eb
kIrbDJa+ayuNikvETu3lYx2767tDvv9B+02m2ols62PXPAhHNWbGDMSMa/KaJMfCtuB3wkQN4ex6
xmQGvNjk+WVRYr+Utv5W1V2TSzp7+4Ko8OPpIm23/KSzIJntOrB7RfuwbvEVOX7hyUDCb66JjO21
swfo5EPwyGlGyb7RRpdYCboCvJ700HVBSL5udf4Y8P9fo1hXAhbQedADra5x8FrhUaGcXl+DUspu
7r7NTWj0xjaI50pCAhobeEMPwZzE9wRjg8AZRxSm/oGVgyWrU9Og9OqJiGBhWGJJSjUjdXlOkp5o
haJR9QLt7WO5/DmlL1HllU2r6mIJO8ZEGitcm7WzqyPXczSieMhPE5+Fc4VPv3qzvxh7ICnxlpaO
BtTfD8rZSiizthewKOFYZqmSd0v8Pl/2wEmI4roI8WrR3pkQU1UrIbKOT3fEvQFfDBcTBi+3D1vK
twtU6UFFcoVH0g15EyOCI38FpBKLXWLfeiQBtCxmMsVvVqw9/GuiR2pkNAl9ULEDlCmwFK/2nZ9e
cNHcM3M8ny2cySw+A4R2YZ4VDxkjDlw2+taGEgOpsdZJOhsewoJ3i8+4sgShZElj6LihHVVMD2V3
K3oNfzZfLZIfYHPjELO68lISRrmS2PpVSATqmXoZ09lBQIg/uYyFuSc5XdACtvpfY1GgRFldBI7t
JLslwgclAbHHS8Fa5coR7OvV95BsPdxQr27z7kmlTx8dqy3J8QImR6ryEGaYnUNIOrZfsapxloJX
NOttWvyfQKolO+fQSoCuGOOy423tG4GuPHjjS1uNlXnZKhXKceazV7LnaJnvpJhnrrvdsi9XGoQZ
WRqr3tl71tHLlxQIRNfXPRU87apCP3Hx19/Q9+vNbTS+IsJHZsnUHLUxNb20EUdEyqSdsoxtr2vX
cld4PEG9TjflloPPdjyJLB0s8BEnCVD+weZDXFSd0u0lQWvRtxKtPXVlPzHmhqwNZGWU0J534e2X
mCLLaa/cxwik9qNG+rQBvGfUZujmTPWq3EnW9zEgw7Lrp/yrulGiYztUmouKFMXfI9aQDiEC3qMw
EwC++HE/bePgm6X+f13OBTG7ra6f1Uy41S9zw+WH8hyE/2rJQhWn13kGAb1ZAADFFy6iUSm1E8Kz
IaBFiWCelXN3KFtiTyOkWRwNKm5TnBjjhzVtzCjZFJrox4Kh6vS9rMaon52UcehWmATNCuD9KgMm
vkIdt/uJY3rWbK0PyyUKK7Aa1uNUMabtOTqSWgpPE3Q0uVwcg113aUF1tvhbz6615Z0FNRPNOGQi
Pag8rn7GW+qiagrziCqdXDtuq6wAK0Z5URC+owm/hLpxqNSUk3LS9peQfgMIxr7qRLoo+WWwvm63
MGKCTjIhtho8UAvxKlUZdrfwQbZ3M0JXfj0Il9yenvsH1d9HlzivJrSqTlaUl/eG9FiMREmfUHTI
aqWf4eq5KJT+T6Xl+Corw11hUzST0vw5Ds8HJ2HxZZsn084gCF94Zj5hPcfaSl+rLTQWC7dXE8SA
/122OsBZDqWknIoUpo4+9CPzJYQ2yyls3l7hkbtaTI0GR8HgjiDwZwkei0pGb+vmjO1UVr3zWRox
PrmrwO/W+O4OOqkd+6AnHchgBnMZSNLcFn/R4ZUEC7dT3A23TPZTGiXTXLtHTO/a4B9kLU/KZg/2
2EzC1eB0TGJ/iwc8DWoGnO9C5E+LWVqSMFCBWxuapFPVOXZL0eaUVDf6ayHF6XwTQ/zXyXalLVOu
DYizGjwck6im5da1bXwmtCg74RySbSUvuMUST5V4Cea3iT1GDNXyfpKHc9yGIYk1QyS4mdYr0N/V
EvsrHmoE5hR0Ta2yeEkITq2Fejmevl2Ebjrr/9DzYSnF6VsKFjAYcA4w65TCPXfiZlC1kP9y/xCi
8APDzhHHEAUJbCZPKsR+5i7/Zc/DJ98u43Z7K/7p3UOgtpguGQqH6y3URWM+89T9zNNM+PbNLAdO
bViGEYcSZZXo/TBvPIlGdFkEcaD3Cc3sVQ31nw0JRyidpGkyKOIyO+NQ6/M+QBGipZ0RUe3z+6hc
1TXjb62rbP466SRNScv3B210pqIYQ0iiXOBZxBdDDuroGlu8KmpkPaeVi9/X4taWnG+3Br/N5wXd
P7MpoLmgG8gY9n3saLNpx3JuYtjRQ+EAaWOJ/l2Nk6PxMDQmLbra8g3pK+Fc2YYryaj1NpH4WMXS
SStq1rqvfu46S8EthETYAK91Y2IxVMtAvvgM3bXOfK/KkuGFAYUmavj9tm8son6e2j4mR3WLr8YK
2pKDv9+rZv1tBhP7lag9Tmy4kbcMDYGoaVQ7n93dSOi33w6D0wExRi6d4l4I/Wp5H2iipD6BSUzs
uci4FwTgrlmOX2GMBcbzopi5QOeb03bowL2nwnO2TabkGrJBiU4R3K3PTmILPvml4nCOqj49+82h
A2AQUMPOB6N83Ir/8bMZqc4gwuBgoAevUwPWzhShZqlzp+Y7gimoPUDeeolWQ1Q/5YAA81myN72h
yOvVyaFbUBGUOIr5AgYbTrpsEKOa9yI9neTNp1HiAgvLbqLpiyKEQZxBXPh/fgZ5NuwRSlHCy7R9
R9Hg5BulDV7HV+ggUm42iwHLtxqyYmX6S41sCA12FMzWJ0I688L+BT+EJEQHK0OVchef+x+iKjRb
qWsexOxSUnS7+Pp381W64U4j31/gttz+RGGCgNKjgraPMkDJTB1XRpERShCGZS4PJe/ZSKyNdDfx
qwirR3y3ajHRsa32lkooSNqWTkTkBcryygK53SJpbNACA0iqFO/STnnCBTXqgiCgOKDfL4Zo3vI9
mcWerM7hHJ9KzmvATpXv36V77fOAa6eNTvCSz9kSUJ10hIhHywIbqTPN0gOWZ42kL4Vq+xf/2OIp
ZFA+XWWDBtQysn8fG4weQbGSylNGU7b4LLOxUF3ZG7OVmr8LsSl/HHgh9/QKKlp4aNhgA8P5HDyN
Ohs3ftiBWmDi2JVLvIZaS8TvB2g2BBUxbH7YVkCiPJuHu61nZdTyHPIBOKf/EDn8reFl89MhyLEp
NDRxwlMOd4leTAXell2E3qv2ecJyq9EAXK8Dm/XrN1LJpRER4FwArR+4FehWw9Xh3wwqRgByy1Ht
X4llfA5BeobeVgDWjnGAgYfrgqDSgM/Vww8EpmVTU3QniagJWw1LrL72DqV9n1s8aDAgYUWym6wk
viae5HcLmqXBmwuYdG/qwVvHaDmY1qvB0WAUgW650HCU6iOouVWl3N4P5PwgNC+LjNIHiCVu6rPD
fEiLIiIny1+dXGcd0vPqpR8Clt6LaOISPfg5RAXHeXpGjRaboNuKHHfSBlepowwO/ZMsY7p1E8d/
/wYg5TFpkOSen4PkbjpsK747gUZfF311okRBBOO2HtNcP+93EQlZRr+gUN45bM5UnT132eeAQnn0
1DHgg0IeVuGlGOE70tThzwoYv03YcU8B0WjycXi2UMVc5qifmx7koxV15kE3ShWjvZ1YJwtvc3Oe
tDUnJ3nchBlxHlS5shLOVEMR1zo3GpJloNQplLi0gFBrlutSIxz7qDXco5+qizT4Jxo3CwK3oEec
Jz1NHhvwz6/dgZEubSpDzC9rdUx+NFUYvyCnXIqdquarPoLodrCDtpMP4p6Hoc4Y3QftDbzvqq37
pz0X0IS4Z1IgQM6agW0Mn9SEAZjoUuyUrYbWJu62MJ9d8mfdrXWIT7eGXmZTNIR3bQZzb2FGwD/S
04UZ2ByK8fsaQTcivfQlAgkPfbKOzgq435wAX0YFkpSw25AKcHKVC1nT8EBQFUXAWpYPIMW11/9b
KLxLkRjbF2Ajze6aCpTwvvaBgVNJt6loQUUwQAAvlMuniEUiX2Ad5C4ww1Xgm1A9qpIsWxQQr0Fs
XhD2vQXVrIKWVsSANNMvhmdqfh94ZRM1QxmBtVl60B8In7PYjfICQUYFLN/HNnULT+r05ILiBDJt
OpCEoNmLgv/iF7UAqZQKt2Pw699Zu7aPlX8kvVj2KVbU+//m8uc6QqG1WRdTYWOw0caf2hiQ0u+I
1tIlukGacI0KhQp93LM0Fly720amr74Bf8HTimVjJ0brfF7z9KaMcKPIFTdPAJ2RD29yXbNr1mm3
sHaFoadWC+LgpN3Nas50TOLRh1RXAOLiSTCU3vtDoIE3983cTrNxhUAOeVoRNL4IWDpqUBWeuIns
VrFuqZis4LsjUBs4ZpvQbE2ycpz+696tYgaNXbySzakwCsktUjiuIUEZ4uAJT+z05uO4r4Kx4ch2
06q+k+B0WxjUxT7iJM00CZ+7aoZYiM5/BxfU2Xeq2OZqiKgY3PW2OSuCPrbDlMSjNKRrj1jgzqsm
tUoeLt254HQMDJ4fYaoQ3VhtCe/Ud9EqWCVKZ5Nrplcj1EW79MW5Bh4ezMLR5WMGrDOe1WFX9miz
92qI4eq2pGVyy+u6Wjb6iacu9RpfQjF3gZh8Z/v4xksdAFPo79obbuoxbmjSEUOSrE4aqMMeQGYZ
uG6fzw0ph7J8+UB8C27RNZbe9l1pqWnnRAb/kNKEKbRreatzzfB8vo6U7p0WX/X8ETeCik6kVO9d
C/yfw3iryhD8J0VUkgPk0ejWmxzttYPXNJsbzLAC7kurH7thzTMnMQoRPhGfOpBd3hMix2aH7BRJ
LQkaJrvQyCL622HAVg1qj8niULq3RTUSTAHRydlclIRWP1JyIgceQdcYDSitTs9qZfCUXwdKR6iw
tJAT4J8Of8N9WCgyxjOO6Gb0qYFEzzM5riVzxMbFV5tSD/NFRVZBPp4gzCtPLAyGGZYybGBQFmHI
rm+9ROdrSG82MJwlF9kqLvxOyQFtrREZNCbO/ipDmuL0DsOAykClPpog9NNJf/KKtMqKwRl769WK
S1yCvwM6Ftzbg9GaPyNjWiAeiNryyvm7MG2l9fSWdoQBO9tzY9Fh+D0SKqk3lUg3wHbsDBaLeur4
KBCe78jP+69nS4mj6ODeWREBVZAUflPn0HPpRJvkTGU2pFPKlo8cl7UCciTK+30kimzivpfAR737
xVwk6up9Fy1rBlW/KbGWPfwxeTD8rRZ/NTRiWf0LFQRv0y0uCyaAwkNTxfdO86h85hl1OSNDz2Ts
lfDCyryTKLxm4XO1AUkDVAP7OX1Un5VdANplmaD7nuJc2zyAWgY00fyK0Ti9vVoPCO/qm4u3cY07
1lUxtJiWfUKJkqSnkN/Vqes8VZIY4kU9m2TNWUHuV2vS7rLkaskcXKA14E8VxSwrnxM54/C8GOC1
XkhYCWyr7GBVJB9vazHr1H/xXag8jrCsK5Scd3sNukL1YIOCrTezzY0WILfQgcKSHL+wqCg2e/E/
xNXh50xEsv4O5eb0pxGdYa++dhayTB15A3hykBfK7sICZochFkB/B4h4ultWVvgL+MmtrLj5sH07
o1pmYjVrlXqeIFFeYqmV/DtqueQ8R8OswFKXazkfXsC7Fr67+TMqNSonz6Hqbcg01fEdi+h4cCht
zV8rzd6lEF6jsXCUzMUddoXidC6p4TyRBmXeyoYyXpZqOJuMqsrbPkJrOuiF9g7ja0maEAJz0ejz
bXN8Zzai0sqzx25p6EOXDPKVc6SeL3CTp9DdUYKDpDFndb3jzmbPWj559INtDwqyFuZVn3YaJQLZ
mQ5UY18QJHwvG3E4eGbV0PjS3vZD8+mxQToa8p2UtnPPOI7tYMvB+f3UHWXXqkzNTb9C/ldLZey/
p2/UrPz8yq0xqu2ga+Ptqe7GUgyeOjyHxJqgxN/BTNvdBxLDSMHpAFe5OZ7VaxhlonphuQy3ipML
hul09up1UxkrPBFSe25xL+iLCLpVMYOLSu05vB3vlPgzA3zP+UJtU+Ik/xskQi7F6o3XeVjJvlyY
C/5s+tlbBgGufyWSq7uQWF6wlTWVonGzRa9hy4gjKPZstEMiroDhOH1qlM/8WVlDFH8fMBF6K9ka
nM3ep0CfJ5Srvdm4UZqch5NxT4o4oZ2oUgCwHrIMQ0xba5Lc1707/dANHihaaGWGmuY/InVIn93g
cF4UaYryGHiiO0baecgiPXlwPzKzmBQRbgjB9GyHVJ1I0KmApumdzAShagI31FdNC841NpTxkqO3
yHY/DQCsm2zPbnWkRGo72CRdg6sMjEvIkBCqh5yDbBqfbxxUIKDl9er84SVrjE9HGmkNaYkEdhT3
o/Ao3cGr/2e0sJ0Y9rnjEis8MfaaElNXxjggdWOip3ZESfe+kwj8uSvlWnJKkkvXts+iqSSC3OfE
7qDK1mR8xiirz9hweStbLjDFf4ERtphUIL0Hc7OJe2Vp3W5ncwRQAKOn68hI5C5ac9Z5lAetD8+J
2ksGD2k8YszrkmCVJdkjsXgOWkus6o/Ldu5JQSZvV1+g9IuWkhssXSg2gNEgPRDYxW9PqkJPc1D/
5TF61Yhkau4Au4902fM0+uhSgzabD8o2znz1E4bK68Huma6r+Lruh+CvHIlaXh7T0d+MEqrRKE3/
iop9VNOc6Vt78e8YOD2pI1gvYPaX3lF6DfiqOrgf3M/pz2losf+Es0PidKXOOCN6l2vLcEtDMVKV
Bwi5ncsQTTQ0Q4ffSsrzoU8DBtQ7He+CI/EXBtrSIGCQX5jzlXbOR5xOyqLNYwuGGn2+/tP22yxw
NEpYxko902q6k6tOQbvLsHZHnw1EVv+UmVq75OCbQy3aXSGevrMhgAL4q1pIrF8622mcbJn/+aYv
Nl5cs8AfeDNLTMJ+mLZ5a+u7LuJ2WNPHnTW9jZ7wmLs+ptGRMHlsMXSmCO/upTLGl+qf5ACB73ME
aPLgcXbd5nztKurGKWf95osPF/Qarow0YG5ThtlvKPSqjsFt7J8gWnMUiQ7p59vTV9BMAb38OpDi
KU4Ci/d7mHad6qLQgx0nTW81d7anaLvcPZgMPhR2ZrldlaX+eGVNQQ5Onzwf7SmUhdAzln/ogrtf
QfByzwiapXzTE9jzGETe6/YvGfqFEdUxaum2rA0C58+vifP8Ctikd4d5+6xnGLDq5ZQpWJHHhlOQ
2GulCuq2SoxgZlsA1lGJxVD/yRpuJL7SHRgQoRkJB40aoXc1+rXIJdkMDRDAmvhagorbDlxXQb10
4lYypjxRQzWi2CnGGWvQ6NAMTJv/O136L0R4h/9WK/i7aKVtnjoi4PZ/toemYtgbnyrm7mbL9rcx
k36CaaltfRAVUfhbZqLm11c1OC4KgKw76u9qsRyVriEV4QUtUinbAtuQGhSV+gTOWWlCTeEJmnu3
YdZWSoESAlh8Q6LuFOCE3+X+N7EvAeyy8tDu2bUFvElCboJnZoAsmpoD7BRxTXC+D4JeWX7smRtS
/XFaCFHysEHlSw5NpcvtfMJjzAO1aMKe5h+6nA57rMBq7wGoDBArfXo4/3szvH2FJV/GUZj/hV9w
7gMduquvNyOGixBmeAEBmh4zgBsCMi4tt0voPHwn+pYb0GQQBpJ5T42lPyRMhu1sCn0dWqCZHn7H
8O0O9yexue9fMrc4gipsVkI4zWxl9SviOi6K5dna3FSlLubTDVkXSyzmhD3+UpN05FFoLy41ND9i
pQqPjrHOIygjRKMOXuNWAm7cnK1uDoM4PUrra0Nj/o4131JqvG5RoLg1G4BdoT+qCLfYMFXUJL0Y
7b2GaXQA0+wG8rE4pXUb7k1JnczduStcDYnA+XiPFLd3bBWfGBTPUZh7plhHkO71+S0pOqOVs8O8
/Dg7CiUw56Yewt3GU1yTFCkKUyq5c6aNtPu/5qvuuMC9SWOrbtP/cgPfsGhPA1IdEAKTM3FXmM8f
PJydrMuTDFVb3MPCeF0Z45tIKoPs5kcMQv05UJHDGCjkgYYuEp33C4Fsz9JNOAkjNbWrnbZf8fcW
3EdB4P40p+YqS++mrNuD7PzZ8RDiFMJ1ezD+54mEMr7BCcQMeyiXgNGmwfs64fNNqfobA+z2cWr3
4c93q5gO6TBWChEDYdiuxYQ+yO/Bk2oAX1npTKdGK3sAE/C9CQjHKkQKSY2a4qrz38I14KFNCDKm
eAnZ7Q40k/0R3ytklwnS3JETqxw+TifHAvf2UUlXUTabjX/B3FFPX0prfwxb3Xmej6hL5OE5SVXX
LJQMvecZXN3z/eLoN6mQUJZFJOIb9p1UfDOEFKlJmqbppLZt/RUZW+Yd+FEmpexnlX0h7AWqMira
OpQVtLSjTZ+f3ZxNbSyaiUM2jOn4vGIPtR5tOkrFm/aBBfM4e03rDE24XG1DffVZBE5wt9wM+gbd
PtE9N448Q2PqJZ2O6yK/6MtjUXr8u+ENhnEYVXAhm96A91A0/QE5QdU1fTObqNsF00ub/5GEDn0M
7uODsJweuWjscMFhWV+LnKCe4NlzE+zJbZkHM6aqbJ+BJ/ReJ1pr+5OHMwIR2lzfw1T+PgUI+iJs
9lGhXiW74NRgWPVjNhk/Ua3wHZRRPNb9zUmDC1e0F0Xvrpuec+wQWR2Tl3dt5SJlmxMeWejAN4+s
1+2qLJ2nWUzTSTNFo4HgpZ1ObTPcMXFPwhfJHOILGHHH09FgyspxZ0NQW1aCN00IKD7IlfIZxIdH
4oexX6gdsall/nZRR6zRuoijNBG00NsrusHKdUAcDDpnt568cA3ySl3sZKs+KILquwT4O2zFM0ql
y9G3d3bCbj7pVHEeeuEeoFs+enPAaBiKPafZdQBKdfuJ4WvNCKgKdHhdIUMKlZDDjC+Yc8VjL2V7
KAwOaot+UcSPyNF6TsQop23xfAKmTKQfpbAQHGFn+3rCw0yZR/b+SH6cLISRHhtXVSzngLGJgaoU
NysfLnwoBJX6ZtWaUyBS8fsqrqEWO+KCT6Z+zeX8tpI8NziETFxbpxr3SLbsF/BBHwXs9IyNo4xO
NRYJwlhAAj+zN52YnblvF1Y2LeQeh8CfFP7l2X0e7ZyJcYvkxO+rxs/Cetpy0kn+c4Ipk+PBuERi
US1dFitFbPMkje0f9rRitlfUVN/F8AriS7vCM64UZigPKOV8OZYIgLb1kv1b4v1XYcSx7zxTc7Om
ibd3GUjyZq0Y7pYfVbtO45i+kNM14h1UVokeoPDPgRliwlTb2SgR4gUZky/DcaGyGFn124ZskmwH
gHmsrNBEu/lKxUJ3cCohWekuZ8y9PeZckchCu6Sf0uZnvTXgrVhEP5Dg63GwpBblHJYjaCoxNxSg
qroYyarVTRWyoA9THjXRPmqCY3dXl3nBJgDXR8/evEJEWU/nF7nKZREW+irdhuH+lGz/I6ppGZ40
w4EFcsIzSsBD+6jJa3cToLEo08lZnxRkts5G/DSHpHGV6Wc+VaMeEFkSK/JQcOmfkEvL93pcQ5Dx
fEnIeFPYunvIOEbhRobnkJp39pifTaiGBgBMhDmAX77Ddr/gBkh8ki9YFUDHG5cDEeCiXKYb0G3I
Ym5ExnYcAd35OAwcVMHEbiPaxjIJGsFPHGuu2vhFUzTfTcuZwU8/87XqWTBtvPoP4pg15tR7St71
lf/o6hcVd6N1JHGLxXP56htZnvAHyfPWLdcZ4Mopm99TmBZbS05nbEbXJHOqbkxBsdFNnjk4j44+
bdahNf7n7aezTNISC4pux22RriC5HcDiISDtno2IsNuQrt41FCZiHCwszUfi5J9wdUVB1V50QrYG
EwI9WBlSPaZRB0yK4JG5JY7+gONFZbBnk4QCtrAV5ma4N6Ae6+vboSc7beLSvmzkRZnW6OH+/sE3
rSqBTGwOYBpcpGQsqtFLEtYCKzhvqdXxySDHfe8LmMa/doQ820zHRLFisLPvDuncY8McuKzNWsmd
HEW/ncZgnyN5d7p5dGfOTUu3V/s7h5I+cRXZYoXCm6VTg0em+l+2aQq7MbEUDyNbbxsXpH0qyub9
nYihJSbKOHDrUX5/DkGZR7UcOVXqXXSHAC1qGGUfMCtc5WxQiGckL8IQLmbtRxnymUzA8bRp6tLc
kvsQWltZEpLWehJ5236bsf8hKPBx9LPOMF6rAWTxH1G3yjYnTQPS1IvaWSOxhNvLdUyZMEr6DHUp
MQkdJv/qvqQgrj7EBQn7ZZiFm3RCAST1oql3Q/NHN9BMv1LocoZp/U3qTWtldPdaEr3iYXXi81zY
DbVN7zRjXgtl+ovtxP2irUsqUuejf0VsjBNOWgAN6iufNNKM0+uSuohg2LFuIL6y0gZi3b8UcRY+
UPHtLOvAh8/IjkeM5keEudvr3HSEv2TwueoBn1/lXkOBKyGvrNissyjfC3zkgdPNM+Oe7ZN8lp73
I9K9nJO29XQmhSnh3KnkA9fmV4CGcEodWFGIbaTOVGY0HB6DXLIPNCluNQEpe+ZQFnk4/sUzJ1RR
wycskQsNoW+g+BeXJYSZ1t2jBxp7i5lNwKu64DCbqIGYuCv3jqPtnETvXw7QPYOPkJ86a4130yay
HW5m/1O5cDXtkxSS9szB4m+ypfeKu5xeexO+3Z/Ed/NuUMGw24dJiB1e1Y3UmYuEHgKs5Cv72GJ5
6vdgOdQD2imXM1+O6+Hz3bNV26F9ocAl7B9B6tra3Px8EtjPQiQDGTdmcx3/CccgFbafaVaCkb5k
I41U1WcUtFwxyhpQhJpzqjEEo45AAN669q5aYcIuP5NNXakUb8Kv+CuqMHUgdIhVLbSLrVYtbRlk
lJ22NNAn5j211eI+Bc0I0eNB29km8RGizjfg64syzMoFiv208vsLI7hBWACp363SFpPVS2pu5PYO
qXmdBubgXIRS7vwo0MV1+gcKOJfV7CgLeKMBo9xN7d9lQDDvKaAc3wnCQOIhO7CU/HQE/YPtUx3F
uhkVbrGtKP5Rj90/ZPaVvW7DdDi6rGzKekiZhIvyKRC/JTUmkFGRdCQVObbrUd67QmoUDXrVE6P2
3pmTyUIVakgFV0MOiDuXCszvr2rfjklHL6j/Akx7s6vymL6m0Tk9UEM4maXAjQEHNKJG5cd9VuiA
tyt0AnVbIBPJWmJI2gTorEpQJjAHC1GzsEGSvWqUPrVzfcVxz68sgRQLQMWZD+zxHpK8iVOz7iUz
PaqE0Lz3FFW/3EPq1xxNurNd62rCCFcolwVWPKk9ipV/cpYgc6PONsHj43Kn5CnJWw5L3srbl1KR
1pKVHqE5xi47oDhIyuUE5ZDelFh+eecaCu11iYVpiQWADxqKCPO/cJ/cQss2hzi+M66Zxi1fIOS3
qqtQbNxg0KrQpC7te0y5MaMN4SLAS25x9VR9qMoDayplW2tsH+KfoLH6CVs3yHzx2HLxu16MK4BX
RjwKt9wInF+uQ55GRlCCI4/lmys6GlgskXINtItgWd0pb+Joh32aG6zbqlnBZhwQhs2QKXBZSpG7
yEKd+PrjN+Q3pKKTG/H64fJxLO4Rq+cWYEgVONp75YW5Qmje+ZnWUk/iy6OZlAehFUFjSLw6e4YG
wnmeFy5vpS/oxm5mkzr67NKkAgUHQgtj4+OIsVRv3gKCNkZ4ZEczdAB4puLpgjCMHVd6dQrJxotf
SIxIsHyxIK8ZXw45PWN62dDEX4ON9zOVUaXPm7AuURO3OVFGfiQ3AEJPXWtw030cwkq5vdLf+svt
NAhOT/l7qzc3ubBBepqCnAip5/XzCUV2RIiHE8Ux1ZS8GWZH5j6HJqzci+YzrODHu7sbV8nVF57t
5rod+gcFbV+EFzMEF33Tf6w4JxVnwagYVS3KvRcxOtMXKEnDjXzbyj4uofVDoza2rt6zvx5RjcZd
38H8LgcETi4+Bl0jhx9QsLpuyyD8YraGtpRM9GSuWF1gi8Yl4AyPlfxy90uH9fxnfmkPVGg4KHbI
Y+RuBlLGXd3u6putald5TFR6e3JixUVo0UYU5zIpcEJdYuetS6QUxP1tNjX86vmilf+nIFzi+dq8
/+Yh2xR8VogBgOHouqkWZrvlooGwAhLWvJWQeUeI53XTAFmiR3ZIvXr3Ij2V7bt/CefmwJDlikbQ
yj+gMPOmpcO/jymqc7sF3W1lQI+ClxDli7HbRXDmenqc4NuAd1ZzmmyrvT5ulvvF/LjuBVykfniL
mpxCsWLw1wWoabdobYN/WeqzTP/ajqvO6MdqUQyMYxyK526mJICs2UgQW8JCiEqkGy+lffieKdHT
8GgGULJmZbtlEhNiZhImX/dEIinlKlFBNSTtbNndiMg/fFXOIKHvTCnWagTs2LtR6OmNu3DHMRGJ
owH4DWsZsU5Ndp2KrBvmNT6v6Srvp63+v8Rz+lI51hCgj6gMEYN06YlrovunrpeKFlp+6isDd3bG
cmf90e7fdERdMhmzlsvH2oCVsHlQu9km2uh48DSHVAPhekbDEtGmX87a3hsHI6tUPSTgSCEmWQSs
osq1pPZQAu7DAYa3HsnQBPh9dGcEGSU0N+BybJ59g1fus1dggLhY2IxkRMkLf1tjYOp0/sjQvMep
y4xoa6kJQSz0OaMTek8b3ySDL44F8Y1q2Ez6pCGKMNBYCGfdEjfi3KJHOgaV4sfE3VoySqCUW6Q9
1n7dJbNh4ayMAqkDoDqF3Rhyz/y54Y+n0hPUL9ONsEgfsS0Kk3bUfvlFXMEo8xi+BZioeYmnVyxt
WLoHf8duhZJ0ZPHTMhIeOwYg4XGSRauzUCo/Y8lHi71zSz5GTpaJgbh8LwM18S70BAXH3T/zgfrT
NbhmRcuFvdsaOZcz9CHeVRqHKri8xHu0QK65rFykjWBSdVSmn0kpAicAXkFyc+E3sD5T/2gQ0IvM
AcJZMvBWWiYKhPQJZY/7KDQWcIcyegANDL0lOSmP6BqqJR1x8CFnMcz3hkengcV1urM9sKF7ACHP
ASH0Y0rE+Z7DLqFaBQ+RdFY8HJathCgXeYBdScparGoGajYzfB01KwXEFg/dIgGlGcmI1YprILDS
UCrubDwd754M2rzojnHClT/XD+iP67Qcq9qPqAd/OqoxwK/QvqNb3eCypszv/8BfkUYeSFqjfPUf
7l4X7McUC0wnMQz/zK1HsDNvVjEcvnlIr4TQPPH1PaP8ix/73Z+7WUayMNWm+4fe+LIbvx3WYJ5f
tV0ymD8MSrjtKRY35Uv4rO/P4OYcHPfPYCmKRSVBZV955oDiQhi3U0BF0chZw6wSL025rxbLnbZt
m7FtOwNa98ZGmT+UBUZKldPe7jU+VW61pqoIZFllpxkhczBP5gUtuCY0UZCBU6+TH9y10GA1NRWW
Xzvs0cJ1wOTi+qfjKzmEwzHUQ0VN23HagRWomIxBnaRhv90dx3EdlEEJYb7KIC1a3N/8IYkNWV5K
8vU1kBjWgyCBNYQLmEoX4smVEuPKeg4ubw1Wsg+F25BHQ7GnfCSFEUrP5bgujFekf32p6L7OgGTD
5v9okWyG3MH1NlVkfC07nqSedOeEI4fMLlchiXh55hWb3KA7QAaGkf0wWT0wwcLFWy4mqPN8g+OK
mG+JVCMBS79e4PrZXSDP4Wsy3n7gsZcbYQgF7Np3zIXq9YPhoyGx4YC3dJ9T2eIuVIqFO7DC3rDO
W6I2H9F1JukhGjCeNhCCUiikXLNB51CviZDWEo89EY8064+DrC8w+Hq1I86fBQSYWC0LBb2Vu56B
DQU2yNw69FryyAyd43p8bGifo9r0Fg3fMS5wkg/wPglkXoO1geLDHsld5jDpEzVPYhRffESxqoHZ
RbVnamFmMVDlGv9dbysftX8McafPnKjOzq+SMWvP3V+IpG+yTSmmgIVfQ51qQjnIbgD3db8VVskT
ApJLKvVzRuhfwD3FrRCFgOQCqNhRtawktFNv9YlcGZzWqWksujr4tIG1VVp1QUeSQ8vxW/HMI3Hu
YDIlRu2+Ou1ssX/j2+oHN9dZ/rMfE5o7WmJQ6St7tiWRnizi56G9BH9DAFdIsoKkxJyykbM1bSfH
RMShcjndt3CtS9QJ1UmN9gKh3p1EbdeBtmfFpN/576P7R7PG466Ma2ihSnHF9MSsOpKumvs0RxGF
hpPMcE0lAzIEjOdZjRkvbML9/IxCjlJDR2aB590NCxw87STVfMxpYqCzsecwpiGa+4Oj4Z+wUI9U
xUlCE/8Ys8lVubM57iRU9yJ5tZDXmimW4WbKkQy3sZSIjfSpOH7v1oDAwJ/Qz1meDJzHRAVg1NGN
BAZF9lxaBA+fgVdl2Zuq/X0K4z4jAO2TK1Kf8PMXF+NwDGtzrKHwa93zo82QTIapTmrDcmKSpMTJ
pKJpDGZczS2rGT4iXbMGyiAGHYqqz0A0tr2pn6UZUB5EhV/M1znqwNWdvPJMDmK3L/gxWeWsviMU
l/kcpu4yKLg/ruKvXgzDZ7oAsBYUseAQgNPBv3PUIVNDSQIEk4TRDyHt73dc1ATKKCJNmnjVBgfu
pQEWEYUBV2Kehq8cRVJSobVyaabCwAR38aTE7xs9MVPaFX16Ah6HX5Z0mp2hw06vCQbd+ty/4QAG
59V1behDfdq8iX4vhYgXRWYlA1SD+FOH4T0y3B1fwCB8wMXkHY73o9WjYxY67Z6+7kwgTD6Vmn9+
DaN2Y2A37C5IJJSg9b30X5kThTmzp8PXK/N3sFDSdiZ05BnBBwAWu+ZVSphnmTZWUy8IeZ1a7e0J
mGo+cStXAKqqfcAYLDzs4OJz1yJjBGjgElSe0fxH5VH17nzFySvHb5R3RuSB7CgIF9//EbPmWEED
/34h0zu4zWUNpdBAZgPLbRPJmsNlJ6qrrDVDz4V9Uw20Lnqmx9DvvfgiGiuMkZG9qQcVWKYn08Kt
Idw2Ols3qB7ONV5L5gMkR+h4reZjTz62Fmwnat+OWCbvCEVvRwen77zUwfjQ7iocybHkM5x4xs7R
5DoCpK8AN+xQKBKeMSyDbl0LgBG5WMO8Ln+9ONy6ocF8QUjyAwocgdkLVxY+FDUduncgPLy6w0f/
ho92OC4KG8mrBAeyerUeyW4JuyXIBEU6rThSBCGOZVQNFsW4HuXNgwlaJkflJ4gWaX3F6SLJdXVm
i/dV9sEI1grH/mLseKaCJ9XAKTOK2Jezq9RmOrR0L/bn+uSHdW9aSkztjF+KrIzGkCUKl4D+b37N
ECjj0DOAwCoDTK3WXY6V0dJNNgan/rlqGqsGX85qn1VeUre533wrh1Fnd92Ka899DOF31rivTLm/
yExTrMvfMyaADqo7BwRSkxM2Qwk+TjvNb30fyu7JTLe5EJ3MxBgJgna42h+MP9WIwAeh3Ah58tB1
N+Di9ZELul+qduKQ4/ebOCRphHe5z6F8nuIPbb8Pk5bV4XJNuxPSDGmRILe4qttXnZ/oxI2SnigM
ah8R/JZQGi/oJLZMUvmjvZbPSJyr90oG5tKX0tn2dzuRm0v6ChzBVCiFIMD9YuocoR/c2zTQTzib
0F/SJWNclaICv3JrYMeEIShU6MPInYSu5kHe9OEv2GymbOs3GV7M4RIu8GMB5bkMf7akAnFcuXGE
diQt4KS6TMIU0pUdvzOcdlhCHBM9EtYTEgrikEORqglvcbtwCDWc8XydSLyTAlsyapyotg2cy/ca
MvvrtkSEDqG9RGJlliD3vL8Sz4W3EyciH8tse6oTkCtW/CJYyTsUwcPs2ZRbxK08IChof0LRS1+n
lt1Mc/yZWG3W24ZkVkgkCaXFB39OSRGxo9kbrj2CPEXMaKvp8FU+OKvkpAXOryKLq3t+WQtKPKG5
kkYTcgw5DpXjyC4Wd61vr20oETTwy617gb5+AGR4hS71KLw814XxpLeDjC7TKHP8lp2Coh/G5MQ9
f/YpqMG7yGuHT3FwDHt0RW+TL2A8DIpE+/HRs4Ec/liO4mW2Ce7nhqFzqcHU7e23TtFlr/mUdXf/
mINiAEdjiOZ+o9Vi0o3qWB51tQ+kTZn1Uh5EiJ1ddY93TQ6yDFtXMCJrC3aiDfU8JuWWcuSzUHPa
TVV2kqzKBTN33ATrsE7nS1Aqm8C+773T50IPfL4XpXs5sR+SSCaa+R2NrrZZzdIrx33YlhjJW15x
vdEugcbUL76Y5b/s05O45uxLGgTXrruG6qOd9w4KnjN3DTGLptlGjXwLEwxJwt0Q7SpX1DUrhKe3
HMiwYxJf6CThtTKw25Rr0yvEA5MnJewRy5//ttMJpuYvIIsXH2O7xVURfPSpybZ88yF2lhXiunFa
ZAUFTj1nx9KiCcV0vw0J8eZd9hwTFjYuykJUobJER3/8mgXNanoArsmN08aB87DAuKG5UeD/Qz1T
ClQLK8S42UOQrynZovJhYHGc/mDwllxx0kbFKRZ1uhYT8YUHapAImmY6Mr5JYlRdbckgC7ikud/4
cxBpfyr+iF03jtpdQ7i/XT0cNa5NmtQbWdpbDwpId6bcvq1oV7GZ0+nPtDBtwVuCoc90bhajq/jy
FQ2V/MkJhonH5/DLutmDHtMyGrQXm1aaF577/uOp5CKxO2c577C6NHqNoc5zYwRqnGrFLwq8/79L
UKqC4FS0P0DYBIb1KXZi8zWsmoXNyTScIpBAcWvJrtKwLBWaTvLJyYzG7vuW33DFCQQMnmVavWrB
YKpjZ220h/e5FUHnNzfGvaqdR5bMNz1X2JT/3kY2rpAw8gxHCk54vsnjN1drvw+yLJcWcNvrdi0F
kpoCkRupsvML7GejEbyvXiRYJGgSSc5FzpPIhVddatqO0GXISvf7Alo7qbVgp3VoJxEtrvOwd8ym
0A7WtZ58XISvHZxaBTMeaow/L/CVugZXC9qJrqBF5ZS/08TtLxUO/Ws3QT7Bf6oCWNMRVRnyzZiq
bS28yylr+pbQV6hGJXbN43wSngW9kODJsXeZoV8HYURn+j+n0VKF75TkbXFISUJcW/nHF05VeK/Q
RP3+yF3S6kjqA+vkmwDZC0Lk8JaRA5x+6QGUFLgH/9IJ5kZK6H8TiWu+aWKDbsBx4a0wYYsqgZ6R
Rs/mhECMFDB5XSEO12jSyu/J9WjE+6rACoTpA6Mwfs92I2eyN9Fva5GapMuktqB+tXBnJbogFigw
zO3IqlVYfuglO5LDROWd5jexUC7Qenmwdd3rqqSzK/Ry0f3+l5LUzsKkkxCIh+FlSC185j1LX76i
YY495SoGUOIiXrFxPjI+zpOAlclhzrEcsEJS8eYBVqhUFMrPwFmDY3wMrEyLNnUgaYu0JQn0Pcla
i48JYKidnejsNB3JCBg2XCkvMaPQN64vEvkw7fSF94LAhiX8usgf4+bmgw1aqAHoq5/iHr9dfRCa
XWms1OLRJSfS9SWkEGj3JUMjEAsSr1oJkWivIIVjd6TspBxiUKQ1oTyWCeB7ZOlUA6jI4IJuttu9
Q8R/ijjokyI48KejGpOFuMc14JZmOAwy4cgq6fiW5sKLPAbomAlILuAHVkpkrcr4tZ/VcqBTOI4F
9Uz8Vydj0saYxmjABuCrFs5B7/Hop8zLIYbE5kU64YkdUDMU9WVT5P741T4ryDPiAGbr2+bdpwqZ
UOC4n1YrlsxDAGUgFz4WVRAYUtwQ/RfAzmKwvxl7g1W0YyY28NwJTcbP0qle9TFrbVSrkSgX1K0s
47Rh1SPWBJ5aAXDBlE/Akl7KXg4OjEQZv4isCQLym3tk075xBEF3W2LUcnDBXlryx+WwXkMuxR1f
QyXzitTMF7RY68lwT3w7xbXSKoKCOoRTkejMPrDp9vx6wN80RfTAg1WID678FsMeW/ytj22cQue8
sC8aHNODtYVNny8y0UC8knSkJ7h3LViqu/1PSSPaNfw6u56KptDGqFg7gQpWfpwRz+HmLqLWVfOs
g44WoJPz1UhwuhXFEOSLfzZgBuMxX4B/xJfgegacHm3oNwn/KKykPzJ5pY8WrhI/fXIPOEOztmto
pIPbhMVdA4Z4HjUGTtJpy9bCl01pkf35reFXp1iIIlIRlr2846FjRWNGh2+4bGCRFdJgf5aggw3H
8sPMTJwkPEuXofSay2iT9RgdMePIRv4X+Tl8b0vKShz8+5XTLurRJwYOO+Hc2uZ4nAYfwKSX7Pbw
+PHv+RfWGTgdSL28m2akaRKTvNPmKoKuXWn8WZDgmNjlmOYY2C2f8MSBecWvmDJWRExwqcONetw3
oedtX5jPL+L/ex4od1IlrF0EYsj+ZGKuYbNUzNbKcWdGz9Uey3l2EcUrAiZcOTnAinPzAzO36q7w
ljV6YKwyh1ijIkPrZ/cBU6SmiF8juA/DlCsndmosuh/clgqpbhY4O7DivmRpi68uLolMSAKGxokn
QOcsqrECK/WgPgQdYRAaBOjAuM2YWJM6ntpEC2TBdrByFAcdbqX9p7054HtJ182vAdIlRMvzOluq
CmyUgal8e7yvwl1LeqRqS8LaTZ3dfC7A1qCB+80dxvHUAccbNDtKCPFTF+d9HXGpTS0TbxoUbPjT
eoMFvAvb+l43xCTkGiW2z4o7nrLbSuYN/ac3zuEDN6mS+mW6pWlQ61HsfELktKXsoKKX2wtuC++L
Sh2qpJ+yvX9n653ItX16urrzD93DtSoLG/pqLP5c1jCYjm0hcOz1IZouHewCHeArofh6fZtRTLyM
ZrRYw0BuDpUqQqQlcl67xnHr8jR8HamY7XM9iRMmZvF1KOUvEMnRmuzNc34yKT/FRUNk4FbGS5/a
pTmnhLhc3gGHDWkavafxm7Chpi5nefEt+RGqpHLNZalJI5xjJwPraaItpEznwWl0T19ARtGDwlJw
NNt4eOMWswDEwIix2kb4GQXquHS3a+xvmgo2E2vk/knl9Eu4bWs0sRzbeM7wo09K5psrbtFEKr7J
VDM4g6wQ10Zhx4mm3hAuxBt3Wr4yePQXWscDZjO5+9z1EUzWhZeVjZwB8z0LxyCnXeEhgS5EFFwv
+1yNeRwCUtch/ZgfY9cpm27+I3eeUiFbZxBWUgtvWv2RhkrdwukwVn3VeY4uqnOITaiFt4QwDs0S
BnEdPM6d7bd9mDy4DUDCxbEOP3GFlGD32u5ObnV4BeRSPnveUjFNnZD3GydbtYUpQliWc1eq8xCC
WLKxny3dv8k598Esft39n8rjFS8VnXUVgGLGkw5yDhNn7WS3PdLa4nkJch6jpWwdM5gFfqZiEcS5
XS9/wY4RaVhNuqKVwXQHMOZsbRhb1HABhEscmYgs0m8rnlGQmEnUGduJGstVwJ4y+4b6nVbrrpl5
CWqIG+1VW8/etoXHL/DQoGCxq43yt1BV8CwPGGrPX/+RvM7prC02w/jyfqszrpicndOUjtogo/23
6jebO3xzyGoRL5xp4e0GkxcEFBSptzRywobbzOvFmrpl2DyJAykqT09Bhv/X642F44OUEaZDtcyV
p9D+3NgIoAXhrmNLPIoCxX5JkTKW1ru7y3pjW9uAKWFW6aXl2OSfJTZmRqk0u2lN7jZDyfjzvcbt
xWYKMqg0mIfsqbNLNpIMpuAtDWbBqCIkphkfXKEndJXYnYi9+80bB8VqGpMwQD4PxOM7gegqhuBQ
5Z/7WWHXoVa1cZPiPkY3BtmA4wdwO0GAX4neok7gVBtGzk9rerTsTZrVvYKMMFCX0nKbbVJJQSIm
swjX9DdO1gih2pfbbX+kKLehGrUjqtCVat5FconcZCOrjl5yadNp5Gq3mtk7CVZklZOXLQcnJf+9
JoFUP0qZICbHlUex8FMXWtnHy2VB1ykNpw4WXSOmfMdHqt+69n2jWiQ+HhxVQdXDRfnuYLme7K+7
U2nRy3pEVbkcFmyCqE2wKrILuKNXXRaHNjxP52c4TAVjRZyLIXtvJvC70pP7BuU328pID7hTmrNL
zQVB10EVsIVJrQptfXRkMtjDIPUBx2OIAN0j/sl8TV+KzrWYMiqamWstmAS06IcnzrMM3yuaSyK2
UpGMH4MdOmjB4FQEol623SAQicl3L+9BSXJLSZTl6EMYNDvKEeHizIcCgbNtS9rinID6XFmJyjhP
r2VK8IfWK7C8dVZXup99h1y/xJX0Xv5qqqW9CfrgdOPiW0Xlx1Ayl75umzJdxsUsSagB8zdvd1Xa
G/zdwnBpEjzBBGmCtqsh57dbDdDw6B/91KN+GZLeC2cbm4eC54dxyzvm/ze1VRo+zEZ8gy3R0iBQ
GHNjXJrfxvf40IDic5pf3KmiE1trl/XAyTTJDE8cYDxvbzprJWex3jQQHODD4tYfDrtSQ+F/Z0Mo
4TjpwlcsWN39V7VafrCvQISDypLIwR8ywLtJUl8yjOF5wWXkyPxfx1oNSmAG87DrGZaKDQQYNeCW
b3i4QImU5V8v6cDVqk5eA8Yr5HjhK0Smtoryf1wPmqXHnhE9o8i67Os1FPIOmtxvzvm1n5BrbkU3
U4UiZMQsmskv3okrjV/yK4fqh7zo6UU5Jj/F5/JyFtX1zmBHWQ3AwngH16xeNpoj6aBDAyrrdEn/
6R4A8NmQmlxzT9QFrzBRi5p/OcpYgrp9qI2CYuU/oxJ56hyiHwW1hTfGIM39cFMlVZvjNaX32UQR
+BEgAn4ii1JbK42cCxyR6s7+JSsK1qWDPNdeqWHnJ8LdpvKmYaA4aFQyCnJKfZNosO1ilNqcalUx
HcCtNzTFdfi287YrIFDjdmmm0MoRiP6J7y0RcK2XKlPMU/WsruJV+jZBNeLbDQXUMICpD/sfxTYm
t46Cgd1XVrUgJ9VlzdmYAV1RBufCiPGsgQUm943j7mApfulbWC5BSNEDT7G5aAECHzjbpt/u6GUD
ACE9AZCvTNM26Y1GR3pbxyHNDMmKTNjDwba5Epjjzxac3nhcJQunkSFZsWkQt5vZFdWSRP5tPrge
6MOFyYhdxypxPQWmSiK9L2S101v8XkgROjAFutYt0hnnmROFcDGDAWDr9pMA4isOf7pDl1a0ec2a
s0lfUbaeo2F5vf93u9vjhn6rvJRLdHsTqotUKNqESKpdPkLpYK5khV+O7pcSlzoxvh84wSz6t1kh
+VULN6oq2BtUZ90HEJR9IZ22CQgMxF28Uswrf7VcjcricP1vav/mOE7F4PccNA7R/1LZjNY7b95W
tP4IBUdH7wsPxsKY+HFlQWgT+Qiu5kkTi8s+uuNuyDf/TywPrQiq/NX/F5BwWnrHm7BZefrZZnYq
3CU2YWOXqN4LpSzmtfUXWp7MquOhpZyxFHX56tswY2wAUZrew5b9LbeyFexJmxSQxI/rRsgByG/W
+Mr6fwYfLHrN8VKKhcFWtP6nPGiGFGnAl+MpQVsnkSAXCMBVgu4pym3nwec/CZu+RLJohvOgMmx0
WRL746znKezVhIhkJDVaG4Zgh6ghbvxMnf2cMUpWEwTrHZn9C3OIyUh2W6e5R/XMqzWH+62HUL9v
D8qTfR6q3WIG9NuKq03PTG+hfSFR6ILn+E3AJ1DGw2pAcrfL9OvFTWUeLuDK/18yIvo+1FPnsexw
8HuWxI8+6DADO8etoQVWJy28MfImnQdLEaXNrS/S9S+LGuE8Ln+UQkIntkGL+dHD0rRra/5MxHfg
fGtZ7EKVIFdYAEWir/goHKpYjBJLZvWHiXgB4TI6/yS6DtBukXYsJE4w0bi01ropXEvZ+FvGIoNR
fQNRG8IK6S9FL6I4MCsuNXnm50yrad4QOZ9iNGp2z3q8wdquFCm2xkeGuqSoWJmxZmoZdcni1WaR
XeJnlylPxBG73oarXTXyo+BrD08LKGQUI6i9HOynjKAYJfhbcrXqqnoiEfc5iuo4i5dj9wnke0gy
mK5CaUlYgokejSAsZHwz9D0seIGI7ezw02p1YM1Bact+s6r1LUi8DUcKFwnf2hVQt+RiWmp0Nfhp
coB8OjIzMpP7Bo8rkePW85uv3nmx+yaXkaUtgQ9R5a6Uxki3eyxWDsydzYzs3Md1DIRanV9GH2Fy
P1qhEVKsewKq3NKLl80SZMkDpKeIEHA1YwROKy/vp65E3NM/9P47lA04YmK4VqMCuUWfp8WD688K
wJJ9qw64+i5dmOHbP/DOe1DNDr1s57L0ZYTx1rJQNTdSHsZYEJm4QFYdg1CPysbwstJiqBOl+uTb
krndnE+nRXlwCTJal/29oPDf9avjtuHnqCINlvt8ovQVDWbVv5ri2RwXLAJG6g+FxEsT+5e6gAlK
gT7/Uzr54u0qTnH/TT0Qtx9CYgc8BEqOR/xABmKNiNMix7CtFQ494OLEcy4fShGrZ203B5bqLp/R
EF944wm0grAKXWsz6igVvoXV00NglA+FQBF8VnjihiruL3Q5lir9eDZN+iznOK+aUaIAAKm47WCb
P3/lZgRDbBx5+MYM4BQ8bQG/Ery2LpF6TlLz/24uXJaNEW7PyVbenjF5ewN2OBk9SVU4CMTXshP4
6LqOLqUIkVBHELiDBAFEP2wnW8L4FvXEa3I1Gr8sxdSWy7AzmYAOH7LV1N7wh/nagia0sU9Ub6K2
BpEbR1dO+q6RdM0bdaG/RzrgDfozC3CEEi+muzZzNNVuXr+DpmfxkYpNVxzdIMGVkEmOF2eN3cqW
Q5iMpbTCWrJpHQ628QKpefzrMo8ILGryRTTqU20aFt0X7Lu1cLcqyzo6PvwR74ylFcPq3VqQ1zDJ
AwLuJfbihVRaVZYLyj4Q4TFeEuGMfQPLNMoOl/Lp9K350GLBinzQUuOwaGnY0qfv+Wcj5GWYr1mB
mn5NB3ywIKRvzNAcUy7DsMSpK4fvliMK+YluCjq+kbdwb3pVcfsFiyCFrAbIC+v0KlkspTBxaHNQ
17121UluKLMFTRHwRTDFyvTTKJUqcax7eZ6YXxetsXiUezUgm6mI/iYzp2VO5DMh16dNKVVSGUDA
T2t/V8mTA3BcJMFRQ+twWGcALLKMo8w/yiA8+EnOtJYG/zJ0LaMsd7aev2yLawosGHW4zgt+z3+2
dutGAiCFjemFXM1u1Ns9n7drZy5D4Uy0x8dmKehfTupH8nh8GooWvyZgHnczEPqM9Gp3DN8oMtB8
ov8kt3N2J/KLgqKX0NzCIEItnqUF9HZvUVkqJ298vkXPMpoj3H8EehsMnd/Ptb12A5QKzkjN00nu
VFWXMWVylUC5P/WS/ZhynfN2QRxRd/nnSYf7cJ+B2/Pf7r+FRTVJfcPMFFI33Q308IZ3IZijz+jp
bn5/QoJo6cEeIzKbhv1FESF44K1Mwyi9yjWBIpgRUOObpZmYrdovcy2PpgYxMjE26s7cffT/HKWe
e08uZbEzD2fH5T/wcF6xkdEFeMcBOXBoMjPSRVKTfhIey+KnrZ34iFDObthHsX4a8dA+p7jNsKGM
mVDG4z5GoPz+CAtAhYiuvizsHvv5QCQrpBR1R0SXwDcotGA0pREUPJ06mhTgEOpEP6ESuQNFhS5E
2wWqOYY+MA/U0CZAOhRa/dz1AdbjOFj3j0eWbgTEEed5AtekI1eK6kBHLHdawvxRhexgHVBlQj4r
HQ0EN3Z+E7u4NGF6grmZK/iTiVtWdBU6Qk4eX0O/XmNoQ+aDGXnY48k2oSDFzhbSOgO1MYpXO/Jl
nPMAfXAtj9lsxVczNNZuuZWOL9UWKXGc7SRiVoUylnRAe9/+tcEiGhWYtQD0vvdIVI6UE0AWPWKF
1rRmY5mCDrr96lbBZqnzXqL6XKzHrGrZVM84sYJu6qMvehbJ1k3dj4fn7mKFsRNPnHJ9yZfw3P9B
CBEJweBwmg0kgYz5UrR2WFgr5PI2xFv3IdC7O8zTSzRTJ1QRvpGdKauRjjTfSF1SFlgR67UH6Qru
ucFDEHzYOLmyYurYCJKD2C6r2+SIYSC1zwBlC9RYOyyOiTRwfAlksuCBQpfxtJRPOEmYjh1o/vmQ
HHBszxjnrG/qkafysJD06MLaodTI5ds924TgiBUabK5pcxEJjYG58nqqYEvJY3Qxltwahx12u1Kw
0Bx2jmVQWVDYS4zwohWmFOULgz8pAhdUdnGZZcExFlNRMf9VhDwp8xmiFqHJsN45fVdq1TMc9+31
hKDiOg48PWREsmJjMwfut2t4uSUpLjLIwpGhFH9njR5ZYOvcYMRVe9bOT45wRaH1fTkvN3FY8byV
oy7VDLsSj1czVqJdVjcLRrs7JA5bqi83DMV/VjVeFg1+Zm8R9XUAbJigI9wk9Sd5S8iWhxw8p/Tz
XMS5G7AqPGwnHFoL2lNkL2ocKu+/CAwVAaB0y2paqaW6XzdTd8ToNB8uvLQzT/46KmZqbCm/Evp/
32G+C1ggZ52Zo1kRSzUFfWQ0sdCgyOpQ6XDQa/3SQ9tritdlyaRDMZE+n2R3DuEE8RPZQlpmnGax
GguoEdyGA3aZN1gdjcgf/7Q1zR31GGa/wJ1cd3PAR8XuZvSHkIAxgE3H31ku7t1IbYrzIBfkxnfg
VgQWL8jCJDyTUrXdIlNr/HiLwpiKV3IkxCHc2/c2cR5Pkhr95zldyC7OeoE5y8KPCugmJmxHckME
IJWpW2XCA26Xp2K3T3b5AZlNrYvWxIjHTHsbma3G2lDdPdlugWAj68J3em3RqfwYrW5E33ARkx2F
aAbr3DOk7X6gq6SuPUwFvn7EjQH0/QS+n2YbLZ84xn46K7YwnkxzIiCvtX81ep08Itlir7z0c01n
nIF22kRbm7MgBK2jO8+cG4TLM0N8Ner2IqZx0O/Jb8dHusk9CXRECTL2YDdVhFJ4e7ySOtQMg3uv
+bbk94du5MKyhVniIME/ClZmWMCwk/CeuUhRsCjr+boa0We6XKPNyjEFZwXlIeNpJhLFdkwUtq0E
c8MbLLkgyCanNfuqWoApfjbqvw5jO0MKk2ZZX/weXeW1OhR3oGcTDLVHiseHRbpp7J/Vj+px4uyV
OvNVpaUy7rD1dwGgBSkXpdRKx3w/m3nWYrbcL0nfPdVNLAJlTI4zDowOVcxDHUVCoUx0h6TZmU+s
O6IFCoreXMM8SZaeNfdbKFGso86Rz1nfZNx2cFjXHUCp728M9uR8XoAPwu6Qtj/HHe8qFjf6QNO4
ouV2dfLrB2H6jflcVIRwa69sdci0X5cXGloWYYsa9mOp0Pnnx4VkesD9+YJeJ+gSoIwG/QvLmZxO
pllcHIFFTfRyHIXWaoGl99VDxRxenwJ9W0kFqzv8tHIlzLNWafPU6xg+MdIWOgtePaqxnDSbkzH+
vUkqU5dCWZJZWRJTDKWHlBzh6F7Y6VS7hnh3W6ZRv7Fvq3XvZ/n82BthaKAsGiGk0FRBrtRPRdSp
2wPPcbUf9sdIDWK6KNCaLHfpCL+NQ7o8e1wiFce+tC9ezKE0N7gWDrrd0RwnE3Q2uc6l6h4ofQg3
E0NCYkxqGy3ZiMULFhktQksFg4WXC65tZ2yrfdMpANsJQ9qjlbC8WOtx37dZKB/pZbRPN2aPiOey
hojaupIlCAv1dsgcSfnfQt/sJb9X3r3KTljcM8Jq8yb1/qnvUeCUT8Vs18X6oi+UHTgb1QpVmpdm
AyjWTYnm3e4A7f425qEkOwoJujI2GX7H72pUO/kvy8bW9yqRZKxyf+w0fgPeNM7UU8FbEWVmmBW5
8ZIfPwh5oCXf/mLnJjTaiT92GrHbNoQjCDVdCcic1i8vBd5xTErlwFR9NUer84kdSshx+MaT1+PX
b1P9FTdTyV9YEoNoNNLLBmfhbSrlDHxlEHoiXym+ZvcrfC+xgaNYO7+6kiDUk1sbUJ+7x9W744gY
716bIgOHWklHtQlBPHG9wQEEZx9jaBTclARIsqQjXr4OHrn8NJtN9VRLGgXKTbxRG13r4NgT4QUH
FtwCV9W/iMFgrYw/eE8VTJXJa+5raLTdHDMLe6UlONBE7m5LvaEodl+emakJ6Y8rqyTvI5KpsdZ7
rRTYOqv+3oXQSnEGKs4ZioN2w6wsv71HKQA7VGvy3CYjJ80zDyj6Y++5LsklaQPvNJeGsFuopIqI
GGR89TPvucXzTycJtGGRyIaDYJis7RApbuO2k/KKvjqTiRD72BMDdhUKBVTbr2jp47xXxROWOp6x
Vw6OsRx30sBHUOzgHgBfHiPYFClkbZIOwWhmCLvDZiMC2aShOIin2KZm1mDl0GpQjWuFjx6oB8Cr
1PQAhhNbUHyiLwgdRG5JEjffZkJVA/rbs2ZY48IrptMAustpOAg0wPNAP5AKm6k0Ik27Q1yiw8n4
cV7AzkNbvcO3Q8PEsU1La6xPAGRm5CpYEJWpHlOs4UgvDPKxRz4AoekOc8m+fLNVE23c2X1AnlJ4
VqraxuKwUZnoQNkav23VT3zzEdczYkqzzQ9tXjug1dyd/XtbUVHjV++Dn6pn2xFaZPqRKYXS0Z0a
Fw4v92NoIjX6KkwVcaomUd7DQ/Zm5SuwIn2EGcnAK/pJ6LMhsyAqtasR6tXCnFnbr4SjPvXIsgvb
JaXm7YCicGT822CizWiYxFqTUMkzlHlO6hfpqQU1Ls0VrnWBKQIV9TGvcoJUimjJ4Hyqyc+U/j7j
q+dzsSCYHEWR30eZ8lc6WDHwnqO/jESgX7w7EYTTZXPqrc4klsoWcaAww3E5tQSPuaHtfuSN7dOi
uJdLu9iP2EhwcLq62aQAgqtvXopdK0PBuThiy1QnBBlsYiRxGgXAnkaw2zl+41/NI1kAQbRSGTXm
q4r3V69U0dAulgB901pAzJ9/cIQWfkgwZ3bcWgOV+8JcT7X99L8yFc+J4Kl6vYzyeVKW61zMSHNj
QRm9L/Q36IMBCPg4SokU1QwMJpvLiJGQfiFyMECo6qxW3WflAHh3dYNXAerHYsdS4ijiatqXimYP
j8gUzT/qdq+Vp2MzhQ26723HccqYhJsNjBFMM1CRYZYLjQeK2NEXX40mXuQRX2z4nWuQ8hrlQL+0
zB85aV5IRWzdHzLOm8E4DwY3YsSBtc5K+wyItAPQRMH/wGmNE4nc2t8QXL4jgodTyL2DfHwWj+Vu
voeiS+oO1rAi7DvGdVbGEdHyAWb6VkhiIV8WDFsfxHco1Mo9e5OlMcjJ4oGtyHU9he3n8OpJHd3A
1HSEpSQ54hLKxTKzJYEqo9QzGWpzNgRUpMBhf7nWm6JZHNrlc9oCnaoIwmEcFCabJKQcvX1MCnaD
ky/oI3/l1nTzoLRT8buPqQQKLPbfJCAjzZn9zK7PzMQ9pIXw6x/gqGhbvLVc6oHw0lTwaBmfkPqL
CicbpWGZ9TlDsxBLgTWXmLmmqzqzEk1jqWpwnNJYiueUeTEuZ0lAiyJzP9PpgZBPntC3SNg4IgS8
RKwS0nRM0dastCM2nJ7lAKRgKecLxa2BUjLp3S/bp5MffD+W2+11JnVhfFFL+SO544/cxWH+jfZ9
HyZakFekO/8T0P6Iv5vh4UK1zZda2ZrKj3hsq0mPFuOOtGfwwKrek81XNiDt39VxZacymRiII42S
VKz8fqfkXjSne+4ZdD5kV+Oey+DG1eYnxTDne8Sc35VJQ4aVM4agxlLXc1JKt6yFaatS2MMW0OFj
3xaie2N0hNieanH0QT6pfxRFi+XnZ8lYlWXe7K/Qa23nCwj/6Q5NXgeE5WfdIdmvE/tBnirjmeOb
ozQ66LOS951cJ8A91KIjKgjX3DXijIrelZVYbmNoJqktowTVfSMVlZ2TtpZdZvbM84dB2gv8gsAs
JIMNqyoifCUsId7C+0NTdopEwOozKcOuipT9aI9tqmOwh6oIyNQ1QqVHq0tN645lqJYm9m26qsJ9
CTWU0GhP9VkB6dUAH6BgO3C87Bf1evAUu59kqAYCjT8er55djzieuzDL6DYStl/pIEgo4W0epzfv
mHsoo4cL/JRK/L8GwQJCulYH4HIP8Hyhtt58AwDaVuXtcgv7CUhlsuzrTUCRwoJ7VJcqZyuvgr1n
5fj9JfUZvYQ6DO1AIYqHsseV2LTHD8RXFAydJ3skCss7LjVYC8cpPPqHx8enqmQeQ9KiV4hHFex5
eF4QxPTLUKV0sIIR2l4ob8CKKaBh1j60Ph+Z6x+JI6HsQJlXH2X9fXLosyyJzZHI8u0JSGlViH51
kzaa3e0KoGBl030Usu83pfsT6j72lE+uCXvFyRSodfYanW+mTsFPjxVd28Mq5RmNYf+NSvbfQlZG
jvIxZfbfftptqmEP1OIuZxJN0r4GoY4ZrJ4V0GSGXojzBVzMkUFNaYG/HBiVPBOeqyMpSYoCrTii
5eGodleUiW6uEw521rUg7juisMHDi+JgCHHrKpNcvYJF7a5vQGo6TRuYRrHie0ZOQBtfUmeG5hFK
XAIt0iWg4SR/8YP5vahlrePR+z9bJ0KSjt2/9AZ3jrYEWKb+tIM3knDnuQhJmo2hJMZtommBriZJ
WFh26QnxKYkGw/2pa+yyvzCiSwHCdrrYrrNijFQXlpfiN9znTO2UTb6xEoEgmx6zlIchuq6oQ6cD
hg9XJp3l5f+7Od9myZ9tVZnRcpstzoKyCr6vSFrKFxKkrDqBgebcIdOrQMwfFUpNtNsdhyeCfEGU
68j+Nsu2AWeP01RyyaPUM1PHOpAtkvpwponEtmKuhQA8wxWSKAr8AUKhtjt524c5N1nx4NKht/6h
F0TCX388wJQVQH4ivZkjNlj/PpxyLK3moTlE7FfUP7rjF1zGmMph53B7UEmBjrw3AXPf+EWvZsld
vPC8pfoLvz/wM/jx1UBjH5bJV2PNlm5QfLd1Exnt6E1v6QCxjt76Ose8qEVuhszrS+jU2K0hXLS8
FSUBHFLIRxpB1vkPKztPLzSlbVUXlynIfZ4mfcMl5b9xQZaQrzOTiLKuZ9DETjGpIIHxYtjVDIMG
uESYXcq4F+4F7fbboRaJyXPP4svLfrbr0xeSCjt6mDsNipOfASFHvRlxakyDtv+tmfucQ1URKlW7
s8R7vuUBujbel3kroZBMzpuUluOL0bEsOM35DI10UxITAt6B1z9MaW0oJB0mdSOJaBQcHuoNFLgq
F+Ovz28php2drVMJ+XgjkTR8NnkNDmxPnAXxBl+vKCF7N8+I36G6oUDFZ+VPLfaxvKa5fa6YglhI
oblJW/xdd7mlhi+VmK79xhL5miwlnrmdYKvK5GttAfxiNBg3P+L/60k90OtkA5qDrRTOqWL7Nm6E
TzkJHEOYTaMHUxYQHhnL3Czc+KPbOCTBUme1gVVUU8q3Clayuo9/ZL88bc95wnmJqvI2C0Uzf54u
SrZSnx3NAkGMPzQ8wEIDylKojMZDBz1+jpQ2udSE2o39Sh/OM/l0UvQ5EuVYQam0fLwcUQq88+bq
e9RXDAtQI7STDkUUd9K3t7DXqX4cz2lK4ka0BGtSuUbd3Z8sB3zpWtACBnNgefdOodh+B0bmJB5R
7j8UpPrIs6rXie7ayJFngAWTiLsMGpEBMzf3EhgH6tDBsaWRDGlIyLy06MexX7naJ20BRUIL8+mu
AQgaO9rmmT+awaNuhpfJWKJjH6BkK/RILsZYtx2nfi68ZMb+F3BDEa6d0YLzkX7uuaigNXPSGwCb
w3z7PU/qEszgNu5taHDSiOoc7mhM1zeb+73L7N13s/h/C8cCdoN44f+rj9CKmUgXlSfNUXWJrLlT
ERVRBoenMK4IO24gd7uyNXs9U4teVYXCG+8fIvF6/NMm+tgSBA5ZgolipH/OZhXRkY06iC+D7Zq7
7UD67U3TF/17g1cDTbB44gS1Fg1xGP+R3eN8fhQz4snSoQ4XJL9ZJmURLHA7f+r7/pFTqiA3SZ/l
n8NxGj9TDq8u+gZ8xuBGBxp4621D+zuUEBd3ZqWGtFnUYh0A4KBnfEhCfBW0WHhS0KXw0ZtMghCW
8Lk4Vmh+WbXKPR5xNsmsiIOW2oTOviDv5nKR9OhlKj9jpJ0idSg5lhfrY2+1+bLgdxFISppjSxpH
i70IYp0IbGJRXSypw0Vbo0QiHT7Oi0MyLfwGJFzBGeGKWyYehZ5OGGCkYX2iWrsrgTD5BKylz2/u
4ic7YPw8/FTGskze1QlcClfW+rtOW5iLb1UTkyyQCJDI/CL6QorYrN9BZHb88dF08m9U4VGyJzzI
xWoey6FNTqroV3v781gxGmEU9EbQdqfSVpkC4lWvFtyT4KqVGPVEvshK2zFK4DBPFP6r3l0x5l0q
ka6gEeGLchsW5BDTkF/EAdFHVYZ92B358//j/0p+GNHHV6rQp7l184bttaKSJM8T1BQVVTtPc5nQ
iVgqZMcfLXUUo64RZpO1olKdR1jzLB54iRYFw7uAZopZEhyBOKoF2bnc1bMBORAXRUw0mq43sKUG
dk3stNlZD6YNt/hZAVH+AraQZuQYWNrrq+5rXIPb0x7h80di6XLouFA7xcJSkkimTyX7fK1rLg0V
8UVQB4CL0H6mp+RDMnOXC8lfo5dO3kigL8hSBdOv/h2wesF9kTKa1kQr9lu6AbGStiY/ZRafd+Vk
nx7yx5CzRC0Ib1XwUsRdKhIkIoNxzAS2U7YFi37Rh1Qkiz5AMN65ZssfLq9ksUVnO70PFKNu7+VC
yEz9lNRRBcE5yOp4jpSNFryMOYbayNn7bReXvijzmIsMFFQffxZy/m9cCCHK8AV4wldsZNFF6T53
zsgBJesmuK4aeEUb3R+SuLA9/QrNySx1QA05zf9QStI309LLzWyZKkRXnYgpme9JcgXuP+bGgmos
ymaHTv/QUX36J0HLBbktNa2vMs0dR+Xs2wC+B+XXrHVdTpbh0fw2glUKcu1f0hS9uRxakq+NyMbe
tBQ4dR/KWU1mTe9FLA3lMX1YYGmQ9c8vBkyc11YI1tM2dM5P0iA9VWAQvT0pfG1abTvEqDpWAAg2
Sfafx9nQG0CK04MyZOJZYX9r6vBK9wNPBHE21N0S7SDh7SDUSU/kpNpyBCN6vBFh5Uu3KbskObKJ
vdeM23195oP73BLtRcvsdJd0IXoDXTbd0I+TOiZ61eJGG2ItATAfzh3aT0qYPgswuh8c8SDb2A4E
rAs9H3cDaSLEPX5BwvVsKCPQu4hpRsz7JJx+LtIGFgy8AbG5Z7GLRcLe6Pc69mV9lIzuS10Jpe0e
d80HHu7YOjwroXO2OVI3VXWR1KFg3AowZGnYPYpSQJkpFhdyPCI9oyeuZqsBRv2WgLvHSxUA/XW3
shvVW/KuTsIxq3LWFYO0knrrwYz68rpJzM2OxRufLySftG2H5rrPgarIUzbPw9PYlqshPOYx5Yxv
pRyvllJLNZkqJtuFWWtkRdzdu4asAs9lE0rv7xCgV0OmmwuwZMs4WY8RtMw4KSt4CuAKVev23txj
p/C6XB7QADaX4Z0uPAXj+Jps923Z8Mb1f1TQnAOqlUn3j0xj3bAvi/b5854bqigo4vuI27yFlyhg
f5lZCOrr82NQTJBzizN2OwraP4EOPgpjXTCcxwr8jSFKjAUxNVuiWYRQofz3gNwHxo6IsjyhNfvN
uhpz79FBxjNP0rt4JM5acPV3I3sfB+yyvnxvHZppF01lGApK9ossRd5nCTggeMToYzlsqMm0pQ5T
IAFN17nm5tp1loue5qqPk03fdQf6B9Mv4O8pdeXKjX3GhiNZmJCA4iDQauQiI3jYnIuSuV0TDNXD
gxNMh6NTvyboWzDTa7rzVqtd02q22ew+7GHVqQBt/RK+AA614ENTbmOQi9tmlHfsUQ8JFV9MhjGN
zedFibgOmOJkL/WjDZVtGXMeD8oDNm6zqOudfoa0X624HMEI2qb/ho+xXWO0m1cw++MqFWwq1Upn
tRbJ8kNqEljhptOB5TBcXj6xGeI4fkflgumBSumozcLEZNeMmtxtwK0RuNg3+ikNnbbjQamNIf/c
xu40bZlOwb2shIgMYxy6tscka1vG4IZolgVR9hZryM5KpNQkYUgL09xoi+IBryH5ilDfxjHC6k6o
CTfYiER57PDBI9R/aWKM9zfzauErouv3+xvd9WEoFwVIe2IsRnfvBTOZtZ/Iqm8mlgUxhh+PYtxn
0TVSDUQHTcWKtcTElirILzgHbHr6FDnrz5q0T9Xz+VnA7j0sLpYldJZs5/Cd1OBZc5nAxYFULoQa
Tjia57fMfLBCy7T5dHC/xFRcJXYkbHfuqfp9L/nTbz9kC1oyAuRE6Ye95b3AQ0fEzC1q/o/mIkJG
1/u0WRLKM3V56wwSTU62iaGdmYBdsM/6Yxx4LmGuYOM6IrWCPatxlk5FCt9x+D0O6aek5V5c5MFm
KIRgdSXl1OCtAZ0QaX6DahrDKDWVe/OPCET57SxPub0PDuCZgG5+RmPvou3X6KhsAoZbqrqIDpyq
EtjukfDEjP+QTq8YI5pZS+0N/YIQ6CtGMAmgGa95fjvq4djiKXBH6eN9tfep7wwMe/ZJ9J2tion7
D9HFCFRSlUFT29V8/u6eQg0KnpABeaW506HsqZ09jR9zcYfWBFS7ty5yaMD/ddt08Y+0biaCtg96
gXFm5bZcRVkb9b0IAnQQ3ZVZb7xfiI4hyTZQcSxd1VTjiXENZtgD/GOQc9xjN1oS14Ei+kpCXG8f
XwMfkPuLI17LCi5q6F9PJD5S2FozIN/CCqDlgoB6e4TXbiI/tQ61mVjlA+mUNa65JEy6Rluv7/4I
/Omkpw8+XzxOUBxZlGIIfGDU5tb4NsJHUj4qfn1C+jOwNU7oSQHZM748hU0VDIlSg1mqNK17MbMB
UQf5pZaYPZ7fonkqDHbbMw5sZtYv+qJICGdlBu8mT6AjTwvEBhtyUDc+F9CUP+6Cg9oeA+wiy9d/
3+fXO2Rd5z431L2BYtskh1D0CdnVKBxKqknJOpa5II1d06rruGxTsDQQfwgaca/Uy/gRHi3NbIz6
wYPnyQJ2GzrlirjOTEO5yNwX7zdFCidfIvNG3mTUHXjWqryDvc2j5o75jD4R7YPBGIR2T7wpSK66
nvkVrdGOQMmhbTXxagklpEV0t9oG65B2vcJCGf+njU5yMEsbmAAoSzQuFclBGMz0pDZdOxeTNMi4
ZuQzG5Ai/nTcK8V7/bJ7CjGg4EzggvwHwIC55vXm/B9t8BIN2Obh/XVA4xs28SteeAlNZVqq4eMM
lzojo31U3Tc/whBvDmR9JyAmpKVbmhLiQIl4PMRCfu8ApFd8oQkmNQfaUa69F3JAaZLBq/yMm6Gu
8D78IHb1uBF/kqviZYwhD3gJjICCleVJYkQMPNh9qMoM9rHzbqnXRYN1yEx88PbTfjevKBcylBAe
fkSTwPeUlkOSraZZR215oln1natx3v/dwLoRvlUx9i3d8PobIlqAKvusNTF34eHsLnyXKU6cshcI
416K7J2nNUiXeE+J9AgYW45aGoPB9I1H7v5bC8RFirsoyq0PbX+caEuyxhcHHwLNqs+o1ILLsEVN
O4a9bKYhI5ujF5KBkNN5uBB+sgE+W7+UsDTBYP0J+QR/e9vYWsl8C+D+04FIzil+lgh48ZTcEWvE
HBOdeIQJsX4V+qUh4e+zSBfmaalzpPVQVhhoLQ7vGtGZqR6nDYWPy8055qpHULcjazqTGT9xPDLs
tHzr/AXmnmyvAQod3txgUei2OX301YjdJng5j3MR5Nc2FA+Pghvy084WTI2j1EqjhKZ6WdlxKoqf
L3mUiUvwQq7CCesihqWPGvej8jdSn+4O8IzpcZzw57v+5dzQU4iVkN1IWAkTxsWib/gum9ydEmgh
1UDcRa/s+hGT6DgLv6UcsuYeuErrhbkIXLGfd8eTldhA2skxh0S/8XcMOvsE70rP22hlXXaCKXVb
YNmmiLt7LjfCR4i3vU0YzfgMxF1CgSy1f4rvQr4BoKEqGVdVZIZkTkpDtAy/09rU9kwWEjgpPoXj
Zjb1/+mUVRhvf7P+ph2L/fcAFNnxS0hZKXWvEka6iadQe7yUN05Rd1VURawf1MSAyQMg6Pt8+ECz
cRzCwM8xjKlmzjHAItxAOBlpJEaIcCBFVjWo7CBgmgIdec/csMSPGOl7nhFm66nGh+RasoblEILt
7iNnvT2Y6THP93nYgXosaEfaZnUysP/HsYEo8tzrUFuSs8PeBeHKJ2k+uhbZk4YZMm7Est/8549u
bmP4zEmCyeI+biXvBgDWAA9CNQAUgXAD5Lc7d3upxcWmyjihuTi1jKxaDC/35yRA93FQ9QWARtz8
FKW3FOfnP9FzTp5SgdCrzZBC/JNhZHsIC1rV/I2frwOkKHMhbUssiF65NZh364xgZTEgM1X1oNXY
GrFKyV2NubWyh7AnV2S45bVV2cXo5Gum5++TctiguWa9q2UOKhZriRWbTsrQ4z8mCo+dm+taVXMI
QQyD6VCx3AbzXDgNVT4QVaGj0vnpkzuHzY5WvnFdImDZldUrGI0/181+QtT9vHAbFR9sC7RLDkgz
3T8zfEz4V6eWk0z+JzU2vLmBecap03SO8WCnYZhTdODJWaSE/5lry+ksylavLylr1OHYRnfafF07
r2oMy9+Xoy1ArVVA6sKRKNCvEpXc+Kv15hqylJ/UaGIpeM7c/fQGqVV3BGtPClHNuM6T02taIGfX
e528AmKwHzEOHcfQdEnLvD3CrSYDEZhXec+rys919mRbV9kw/oU6/K1yVxKHdoWEcU77MssclczX
4H4PGxPW228b8vnTAWGWlqi3bGHIlqI5Rnld52B5I/vpGdX9PG9Q8mc3MN4EA1xykMTtjwNh/XRy
EEk9SOfnZgKq7sbsmydW5sOu6Depwhx5pNxqDJ82Vcw2Y/vKg0nCLIhtf2UDJmAtsuRWt+Kwp1Qb
3ZpVb5e8pnwIHEdoNzW+18m/vrb6wn+blitBUPlHfGVqfTObG17OB72a3KZSt/kkSEIxtPq8umCr
48IalbeG91PoI0fBkVGpst0pMeMFS1YBMh0V2lj6RMZ8owat45i3bkwszNlCnhri2t4TDyfPftpd
9+THWiAZhLIj00exVRgargvzUA25rQqsMc42P13O9lfXUxid56IHsLbpdMFmqbbjgVCBBMgCnENX
N/eKqjCfBeR0XBx/WA6KRZRH4SPSiBv3oOUW/WrSAaRiVEqoh6564MilvAMgWJnMSHr/sEohpvVU
AlQGKxCfv8zwWhE14Hprn0pbg/SIk40PHHBljDUwOW4GOmu8/gmJfN3v/5/9TpyVRf5qBLPZ1fcB
IEY6+tczGu7zMX2ScZy2SJvvzgdm/DuEDcBvxLEu0XdcUJ8gtfhnXfGSbHPjGf8mkPiGo/oCnkjP
+85HW40aW2uspqg4y2mVeFuXZfZy06juENBlWGLoc20TlMT7LTqBgeuOxPuOzXph3klqn8onUKGJ
fYjsop7lMvfCcTTHsyPYEQIOw+G8SNb0KB+W90hFQ3qnd94FPyQnxdlTE6AkK12DwDrhQZobr5ro
9mIQrVqSucPKCB5GZ931FppbSDKsB4+6yV9X0cJkwNkVTlbs0AEl+O24WXDy8+nNaEhJF2AXVI46
OEmxnicCpY48aahy8FCa5kbfJu4pxuqL8mPdEalct00EhPNDuuAfGgpBNwFapfTLIPGA3H9Z1FEE
UH7xaTvX0rT6f1erTSHs8LRRddtDJk5LCd65yRD3QLMCphbMZO0wIX2pFLXtpQuPl9puDO/UiL5d
Kk2rTJ5yI+UDTNgDdB6a6VlHnc5hXAGIxFZjZ0UYZYG6Vmv53egEqAJvXBXtGK3RtT7ioLrf4dW5
lfMbkGxqbY8dKcXnlTM/MsxBcOFEap/QhKy0GrOxuup4uHqdnUGsV9fG16Gb9b0sYd/06if3FI88
Klc6S2vJyg0rD5fDU53doUnis7FHy8gqeectaGpYiXpDDXOf8pAba/uzUk2ent2BUFYFD1XwgUu/
P3HgRHrcYrUEzsMZcEXjmQl/R7ioqdXx1vHznKXPVC4LNMbA6M7o3WPRkBt/OdDuSIBRXFmdG6S8
7bpV9lSvywub0AxCVQRReDXM8TuRa32/DBwDsmiueF5WTJT3ITZ5Pd+HEN1ABW2ZlXPfRcZOXMns
KvigThep+oNZzmxPKVLt1zIJ5BHPRbUXiAx8zTxjcC4Vv7wMDh3u8tpJhtJIsoKQK0/v0cJQc2vK
oDjIu8ZR7ezXqyhhUtuP/CDwa9vTVXGMBy2VpUorqgKS9uhy59XLPLhAROqNGLYR0OqdFPF9alvZ
pjMBZmStpXxzDHqdwK+bMUts0crE6aUyW0SOqk/lh8j7fKoRpgMZ2e+mzrEv8iySpJSKtRWR0X7Q
3/KGieB0/ujyakeDHdZaPqtm40d88kphM9QlMMHm/PlZBrriduzcNMJ3sv77ls5X1ktZBt4CdvTe
Ly7fpZuFzAUzWptgTgIc2vdwQ6SAM4tY6wMZw9iekAfrakfC17mDvGsoDC8zru/SwkYHqk2jbyHC
9z/f0Ph3vVBX1FTuRZPdUwf95J7VhxStdXCjYyo6d+Fa0dC6k/n7x3l7AGhQCodSy5d8nQjiRuQq
+j3WavaQLiEPkYqzLMgCj51X8yafTvSZGKh9qhFsrcLDHbVIHb9zWh452YTtrLHH3aktspzwX9+k
pyETt8WH+39aLXVIKZ1w21wavqOP/pk9PCK9KP9CyPIHc7pC+alY80pXZDEwrVeLLTz+43Wq+Fz3
KptUoNeQemCz17c7r1XD7dwGktyb1fQbjqKCcp4BzV4CbAEODtLq0QxsF007adpg0GVH+eG23s56
XzALw+tVVNdu6IP3qn83BIetZVFb/UofFPd+Wm/NwcoxsZsZTC70T2j9wCOBiK7Wf9Z9loE3H4wu
ARJ9YTI+rS7Q3ad3vjoFKCQOurfO/tyYylk8mwHnYsX1vmpx7nU83TUBnhoxlr1U+B82VVhYdZFO
Yw3QCNJDTX6+FzKRgIg/LoUwcrDoFYCBAOK4Al32j1RW1W9gn5owvUsTJS6A12OLlFFLacIeEOGj
2vSeiuZUEmkG2oPIG/yCLd4lmhGtaW65KFq2RYFZV5x1SH1oqHhMkVC4uspy5ZwN7d1pOVGDy7gd
oZ5CgAW11mnM+F5ZSEVQiGaW7CAwbJonlmeZpUrg6s3goztpCsEm9q/dvvXLi3jYJqRYxCmEeGv6
r8+heeqWCC6xrIxsHpS1ukTii5Ttsf8YmuUwBCn1L73ccLaJrR9AaL0Eik7l5sM5oeqVm9QWSVkd
S9igPR2GWBninY15Vq5TIk5TDTPku9q8fIyO8lX2m4DSywsB1UhI+wZeynMyiDNzlJeQH8QrbSMB
q0C+pkghI1WBKFdMLLhibqcMjWrcka1M/6QTcx5MiuxnJsFqho5SdGIZhT18Q6KPUQOwPGZVtGdH
QM8pNfAlEJF/NitWXmhwAxUajj7ae2AT3hGZwWU63Pi6ckdDa4/wu0pEr2fARUIZ8+mx0xHEQgA7
merXJSC9qzioi9f4hrOJ08HKUzGzHIyJIe4Z9/7XujM9jv4vSlAAuqFcii6CW/Ao3pUg0iGHFJwI
YdPVJ13LQPRAE1ECfk8l7/QorjhqrCP0xVhTpotauVmBA55RXh+9cmgKKJaREkDE8rNAsAJSxWkx
HXZGLZjvZf5fw2iDZaOXWDdb8mZnNs2A4xm5Mm0oF35YL65izLo2F2y4zzmwzFkf6BLffwIYB52C
FTFmahR1QNL80gCE8o9YnYTqX9RVz/HCDKhpktFintQMGKS2Gj5AGo5Fo+MZ+dOyMivYausGdXpz
URL9Na9KMbD1XrFLdII6awKHoY4DyfK1Pp5fRWyFTHoOqLZqzUb1GsoeS2s6QWXGul+kIKRh8omQ
zFk5ZXgSylZFbByjpTH8Ic+fBqJfcQADm+t+IpnBIOalhobh5waDY5Ky29X6WIZbapKjnbYRXs2B
EMTrTO9uhxa0RQxzd37ZstTMWWt/Mn7Aw/UD8VjtDWU349EwJvW6JrpdxUTSyyWVH+Nqy1Ob+6E0
C8lyh2XHBpNpmOoZcPFeu3NI7557StYln8vXVcbRluVwx7uXItTzqzaKki4BEza4Wa52XuhpckT1
hPQ3fDsCUHHGiWuKBAR+hY5yZoinfOqRlrAS4Qb8E8rVEk2qrtJeBK8ltjPYmaGUSCYO9oLoGVQK
gnYMFuE2KhU0BYptilprzyTX6Z1c2gtw9OJ7Ew/wBlhtCUt5eJX7sKbIWimqQgRyBb+GzmE7ndal
aTzZXr/LRIKM5z5fNDf9qAlO975HxI74Yu1DJoP5I0nJ463lQD0M+PkIzlZ0AGT/qiZB5uRg0VF0
xwEtFJ+IXBE2qKL/Yq6ZZB6L8k4g83BYQ8LNFEJUajUy2U2WZLw0KGb4t9au9lD7Lz7SB7ocUhvU
B/KPqcolAQ85sGKR+ghNzE5UgBtjH4BxeLYw5FZe8hiztunlBd+zWHF/8g0pENzDPmLPOeGa1GPQ
Fiwmh1XgHrUXWoyYUKkBffsQbrHioNpyrJ00H5+gAz9uZtHH4cYrky5kPDM9cZGuaYfBbFjV7uCS
CSFnpYIrFej7yuXYs8oP4qd/pD0agIppRHWmfbkEQ6NOgxifX/+FfZB0op0JjfEoX+xfd3Exd5PZ
XoqItm2BPc7CkMlxtj452gwNtizi11ePmKWrIh6lVmPZykmzUuQZOPgP6/hyc6PlPbYuswY7MO5Y
m0Jvt3KgisTw1R2XcFAK5YLN6h5Pdgt8wwfnT2SxOoQm8VcXuHzFz0HdZ4ap/Tp0pds/dcyxLhAr
W+8rxivUVTo+eXPK5G0b7objTZIYBqDgzkgIvWUhDwcuAtLaacBdeFYblEb8YPuBNh6A15oSwcFB
7Y3M5axii3a+h7sSC4dShXwHYOwgnSrhEkQez7IGZaucoWy2/0eAx1t+xi4xd4YR8wCMc+L5kY2R
0NJNl+XR0lXYBlnwYfgYDUZeryek8/XZIpkb+DobccvYhyPtRYFWS5kH2rUPOyowqgE2SQDmym03
DbSQ2NzpkMwh6NtdXsG5X6kL1mO7wb4YPGHcTIoTnRAMocziX7ruLnQp6VS6geWXZXWZZUSE4Niz
qzuVoC4WIKTZe8hqZNAn8ABsJdlmQjwezkM2vp+vCOaTbf8MLzw3hz6uPSbZTTIiDft9nXxLlohB
J6RuLS3Owwj9GqpPLzqUB3H0h0JVE6JXMOKwyeaiqXLQg0CslLRzNx1lqpa3VQughXHKRUNollfO
NcdhIhp8US8hNWuFjN8coOumIZZs21/1xt3G9AUPrYAVAARJZ8K3z+wYR5u8v1mFcylhJkLHf5+I
8nWytjJF9JX8Dd6RTY+7LdRN1ZlvWCXlKeTh6qcGYdvA/VFt1OkcsUYst9Iv44QxC1Bc/ZfB6JNG
ymS68foi9NWo0IdYaUNkD2x+iKQTYGMDfrLeFblgJM+gC+1DSqbNQYsGspqmso/WBjv2h4/LvKux
XbHApBdqoRWWCwl5lsa82MdOfz8HPNxUA5YJk7AmG+1HwRXPVg0wyd8V0AQpbSJ0kWutyNi+ipN3
R0hPwibzPAK6XcK68/BhauY57vOdyzD3jXZTtUDOiLP7XPfahEnoRSgM+0BcPrB9qXVyMVi8ree6
Cqz/vAkwTlEBzAsWBdD4BrLBWBb9EvTQEpuZegzqSM6P/6JqrLI/UJl0hdMCwg3aeyMMlAMeE0sd
4luPN4QJXUiM+hN2EUGunT4kFPsPTjMwMuXIwpxEhPkHV01sE8RNi4OmbUVybaf9k4ecHJECNMkG
LBSgehrnlFVWW1V1/6PZjKqADD0J0FRx9HsRTC2YrPSuk+T7CWM8MFZefNo2JvcHFLLXjvHwfqju
rnfUhSo8KHC7wM4raXSR3gNV3gCzom8F0nCQqjeShvzD95gflHfaHt2Hi550hmwOppdR0NTTgPmv
qCpfILiBLYqHdNdP+AchEbZwDqUUBeHyw4mfBVK2VpYI7LxiI3aX1tevk27q4yLuLVei+eQvkJPg
1Gx6n4LrUU+7K4CLP+gJYi2Mh9dZRZyMapNMw/l6zVnnNsonvZeySaJDGvjE3ptpehFDimLkdlgt
XhPMEEBFeQob/rI1+kjCnlTkC1jWMaaGK0jYLoWdm+VokmZNdA1zOn5gM8Sl5h1NHJAGfOiolqrf
rBo394DDAcL9E2+WG1CdJgP1FSGhjg/KjKAAVyekGv1JCv/C8lhP1CucUea4eLETLED0eN2oKyGs
tNPPc6No+sOq2at+8uUaZihZtnpDKsr1jb2Vg6oxCjW+6vjFuYc7hIlkooGkPOGnX/3fRzHYN3JT
h/D2THfXNLtmOcy9hzjuaMbOmp3ZhbaMl+PIc9iKMUtDtCK72czZrlEC//30DXs3gbwzsBBwBfAm
4VP6h7wycsHKEELqAP/dizGgb0A6EhT29Amy4G2dCoA3iWzu6nZ0fKyr7vMH7EQRqQSBtaUXjKV+
47uIeZOAc/NP6L0HgWUFn7p2yU+6q5DvJeZhdHaPlAk2Wt6l8OkyD4qSHI5ZI0KnTzBbyUaY8GoD
2Nn2bV5jLGL0d+pdfx9pGmuV3LhK6ZGW04WREQqbEtPbL5KLCEFVn89IxeEerKAI2xgxLyHHffl0
vNQwD5VLJshKQJTbX3Mol+e24f4N/OnfKCgGT9LXmQUv1i4x42jKcYBlenMJWIO9D1+lK7f390w/
W4+DM1y1JFzNfHJgvc0b0CkzbuxSRdaG95ADHU5+caS4tP/V2ry7hXmcjAYcekoeccMf7Mpak79s
ECwjKOYLCmFZ5Ig4+gXrR5m2BYcnd2OGEfYYLbFTY/I8xLTkA82boVYzHajKATwSExR/Vb04q9fN
gUOgz+IJPC1I1Q8AlZ1QN2GyE3sWQG5XcpOCH+5ugCx/oHRCEmhlPCStVMgMSk02xDwnMv28lEM7
fo0cz6cvBEc/mBvmtgMq2ajL8StSNVGpa5kWWkRxKKo3lMcGFJfxSHdn87ufS+CpsY2AyTMqaj7d
ZxT9CVuRhC9hUHRgyebNBr3URiYQ0zPK4G9DdSEO47EGUu3UxUSW9nrZhvTocm4N+3uvQE4aV1O9
ZFgYuaSgxbZ5s7tbhJXZi+FvIVPQ8R0rWtw+UTSuPXLv/8qq7ep2ETVpriANQForysPIQ4MzMZgl
LpaUfrPe/48Hut92Pi0eKb0OITQE7yhDu25INp4jZnCFn586zvVDnxB9TtseBaqeRWdlhJBv4Evf
YFtsfCVGEKAT2w15jLJZ7q40oxYN3NnFVGpEuhfl+cN3HSe1qdVDszbpaQiY5FWcEyOGc8c3yK0x
SPrL29EWRVisVGlyxRNSmCiG1Fezffcg+cOACYP9BSX6ge+i9/h8TjWthbCcSJntssl0AGToMmqN
OWUc6hEVcb1wEdEZ1aIf/G6m3EWELJxsSzU8x8+/jETg9FfVZ8wMtOBi1ZujO38qfDvu0XleWilL
AkANx1NP5usfq+QQHiIRKX9noCQu6YryiP4DJWfgstyQ5cLrlEDuqwssJemcxeF0VOPdMHDFwfj4
3x2gOAd1XMZD0wlFyLBL6S8HgZDfxtdnJ6dNq35Xx43DK+gP2GtREOn2PlPKz/BZqoeQPVLYvmZz
BxAy68dfArkLUw3nBMIeYjvSjbkUwIobGHcTDMYadzmqObCaJUxFsT0dy4o2cqlG3QLfJ/FqGiPW
URLoQH5J0798X/+4z5BnHf/F/1EgQs5M9eBxde1Fu+Yk64sdwJjjXFyHw1omnaV2PTdbHBNqg7rb
kCjtTL/5OGxQaISzzv+gmx2kFTpBpxhiqgWtKquJBqkRqwA12asQJArJHy6BXp0WYbFdUCCEOGAw
KGFlhvJTjWnVqipyFeqKpDX8oJc/3uxvHa96OaQ/kESV/4bRjLHQ0vl+sP+uXPaLGVm5pDl+h6Th
G6kDpzt1dEvWBO1v+s/dhEzOdcGD1byAnwLppgchvZabW6p378kuEamtv9zQmCI4xte+qc0LiS5Y
6iUGkY0SK7fiMR5/grIhYGxXA5B5QLpb2/xzbAEedmhJl4G5HDGQpFxN/Xlp3dda+tZaKxwN7TYu
cyIWEwLKkuE6UyNXkphdy/K0hFCijB0XG/94ra+PiyagR5x7yhrZD94tpDedIZhDWIGoLh3shzM4
z1CVjZ2Qw5HFy0mjeZnilXef/ZDGCwDOzvNrgDOZOthTBng/+0KomgIsfwBq5aiGvaAdJbzmc/0a
nyUYd1y8GXk+5OZQ95GT977yNiDlYLj1IbiC9Z1NWmwLAIn21H33gGMHZcul4VdenxXPt4ZGhtai
/L85fyDkNY6iQ1i1cMUgPRW+FOlpcovqMqIP4vxf3SeHRvU3uJfnBQeVs43QEqPt9h7Wh11vCsIw
aKYWS6o+LlX7GHiWhSPcVX/2VtJrWyTT0VrzCqd8TCcbmjmg2cTURhz0oRIwZYqg5lfQI4zzXYW3
sSz6bp2ommM0BPE1Rw+5anIafVzs1JTGwRxxw3cbKBdr/UDmAbITxED4vILDuC88+p/gGqRrFnLu
qS6jyap/BSwRnByNnIjVT7ZPMmxJBMYuCHitGH+a4qhiEL/Fd6S6Iu0E3QEhIq/eCEj4yEg090pf
EEWm/VJucWJmgp09rkrzKso4xalbTcKHH5mq+zFTWaAaPqPwpFJTKLT3BvTl0Dy8/6sf/w5YMyLN
8zzO0Xry+R+ZO+jl67VOPogh4X0Tb9bstGUxxA0Aoe3/XgveveZM08Jv+XafB3BflTgWHHPVMSIG
dD7ylFFQ4pcowTyWD3g6y2Tc1rMwi63Of99urCPlXuAzSLVv+tsA0gDD/ObFqZDt0tryR2YT78EQ
z9rPAbCSEzIlv2kpLqlGMMBB2sDfUuBL3eqSi2WIR99TsMzsv4ZjZ4qWaMGSz1B4qz7mY5nlPyQJ
A1MsjU0Fp91gORDv1yfHx9cyVpWFkUoCO5JH3SV+Y2ah49mWP370gvTOAWgcIbF9LKG8xWpkTCNQ
AJZeRojgcBv4eT1Y2x5cEnDzQt+QLQ0G50DIKSxtbxmWzSLkxmfhMqfXVJH/iRludDvavInq0CZp
HWhXDFDQ9zYlOIp2m6b9IAdKFAAMG3fpvqpdOkgRnujYxF2j8ofPNsJLFsEYO3MAsXEy9Qyli5iz
RWzs06T31IFOoOZKbbbNp3NwhcwSbKDPSAv1f3W5I8lOZQik5BNLUScF4SAMnkKjV/TzG1KSm487
biARdCtTxtKEMBZ4XhF+HTkgmBerWwOkpvOCniBNGpj338H1UUvcFv5QHJgzH6YOV9R0VrZ09UFI
W37/zyLxHs/hsYuo/pmK7KBFSlL+1bTnMUJFD/sH0OxvOVRT/6OhDikawAyPwwnVe9yd9MWxgOIP
/FySIp6vU816PwBgGDQvyQgiX2J/GmKICBTg1ALuT81FMxL3AeQHgsei3BdT+5L9lexxgNI5KER4
tyvT3tO52zEXhgLf64ihUjbb2ObE7D6MkWFI0wNL8JdGs2Hqxl0hOlKuvlgeWJRceokNoBd3yzXm
a5jDRhXZd5BUMLaUq4fUX+nUNZZ4HPI7prLyHbxnAHkn6ys0ocWgniS3ZfScM1zv2JuBuDIbIUyn
GepUkY62G/WIhZwN7I0e+9YUYRU0cac8tJK/j/ClfMbfp9FgRiF5UhlTxp7ab8TGyuVFR1C7I/Oo
b03qh6QfsCAqhGrc2ZlWoy72ZbCt++395Zrcuk/eR8Cn67bZXosXZO//gT5221AX/LRMVl1Mn2PU
F/AwU1LS8AemCFDx/ldrVBy9nxzbQtA+MshkZtJUk4nGt0JDnqXwDrQLpnZrP0qsDa/56IJGWLfM
qK6OtFG3Gk56amccwqohK57UAMPQQht9NYcuYWP19XVg8q9VyqT2pM29wec4ZFnTp5KGC3MuJfib
J/c4lRjmcRuP+0xJM4J1KLBczRHSj6MGHq4ZJIW6hzne0Wk5VU4auL+6KXLH2r7ymCgDtkvmWvug
AlDHWE6RAcxx0DvnWM5StAa6RwDpfhAFIhPnKTfxeVry2FfQh+5ShxDm/Z4PJNqkEbKDkg54/saU
hbNLfOk0rqD/ZbLyV4RKSLj2iSQ2Z8y0m3Z7brP6FGx5HtUm+OPZYlHnKKN04i3YbQx88KEnuMnB
T+b78u03js5qh/9FZkzW0LR0IiRn6uPADHpWwmFiGp76qBzAUyOnM5Pk5EFjEzsQdiKxhg2xtPtJ
l+VNMLykmKNd+AelOMuF60EfjutIBUVgYTb7yXAHOpNNnrERCB2FNTJjrg5xc27qYvHYvhnIyVGg
x0Hj5SUhavCnMkUhjGyZSLlw0AH+1vwTRfFAV6V5MInzlo6N+V+E1eojOnionjngUlVKjyImS6Ys
o8p6allL0t2GXthLhXD8w4ZsroAGvkG35sMhmefzg4tqAeLLaPlJmEfI2jE2czziG8u4hoc7pViO
eL2hYNLw3IrNA37bnK2EJCmoUp/boc3lG8oJwUx4UnzLarhaVcuH+GeRk1a4LNY+qAam6oODH+IF
IX8QUMH7Tf2HVw+DdFcftN6rQ3u5Eu4mVAeEADWGy1Hkin6b9LBB5u5sr/x8UkFD+eGa5gCo3csi
CizeluC4FOyyWRvktBkqvcr5DOu7y/M7+pF1DoO/nur5A8gGGecwakE3KeBiR48/VO/1+m/ePzY8
qDH7uPr0Ghwx8er6L9T104rYY2RJ2RL2fkQf1FTIgozU1LxJYYGDyXWQS2gTJbokg0IUp38KgSEJ
79WhloulzpwR7PO9bEdCzlERUmRJFDP7TLwDMBfu6+k6+nz4Oagi7KA2nfzwW0E90lV/6MmCHlYY
5XWHFUv5FJeltT408k9wITiJ8AUsoCwfFtIFe9VuG/zpbRmAHAcXdijMP3QL8kTfecSpGy3uoxvJ
Ta5/vL0oT4WguuewGhT4KLwL5gCN6lF8bkLw5IL/wkNQWhjkn+Bce/wadHvpT4neUb2hxDO8f/+1
0mOtnBQSNcf6o3bVfLA2TXTbNQWMKNZi8Wv8Klame4fzUZn1E8adGRhK2PAnlEVUCjmtGiLWh3jl
+Nry0rNAblF9ootCUdHLEa+C4nkCNQePpaZDSpJSI7YRdc+B80r+BRSOARa5cZY+ZQn4wiVUTqEo
XCcq64wpKBzHhsTPaws8dHQGxxzOavgZ60P/MQPZZyrpS6ZWwJsHiHtblenNEfF6NlIlDCv6VGQf
v95P9/t3uj50H1RvtzijIGjLMTHd+THFSj0p2qbgH/rizxVUW0+k2NugaX3Yy/uI4B/wAvCLCCCo
AvP6Q9itu1opcp/bUeeks6/KzEDCxrhjdRPUZpaa+O9ziWWbyE3rtnYuMzN19PZVvX7wjZF9I4Tf
FF/qRYGZZdv7bOohaY/Ml9tr2scXrFThiBqyc6UzAbRyY3E7C5eZ7/0pb9urazjuNwJtHc+yc2F2
V0C8jfw0Li9hor0CrMmqdIWh6zLCknTs1ytK9Uz131kN2xGKnZsPUs+cbFtXl3eCJYIo5i6qc1iM
AI4HqX6NYfWHciECRAFmiHYLJJzwQPKabHanfwvjqFcPkJ1J6iXq720Fj3S/KN7P4RYi/GIIz8wb
B5cFv1vwzC/aIUlqxPiXYxbkmqbOb2FCvAwV8rP4jhR3stNKU9nit2IHOmqOWv+OoyBZMZosU7kH
0fVFNOkrJB/pUnyOCje9DxFLyRK2d4c86PV0YYdv4dKORrjzCZem24MCBM6V6McNaAAzLkMd8gdn
Y2uVThMe4vCJvyf/0rf1YvcRsLV8EFJlVpgijFt/ufDEEZgVvodkPQzcNfBHs7ebvnrCczDBit80
2vM+im6oO3TVEoVlZXFfTkZJ0b6Ujj2+TaX/g6L7S+h7lgViQ6ty1WYi124E8be78t3RY5la1x2E
H4f5TaqI7mne5VGdnv12nlCeRJzzOjmeOMnbvjVEiXMot6csra0gbJvOe+1PkWW7wxrsS966/T/B
GbmT+zKCgemLHwa15POkbSqw2SsZG8j14yfsbwxSgB6nlNyWrKb2rlEDSmFlI9NlBkFzHBn456aB
c8kBGb5KQVjBGoQbebkuiKuN7pBIkD4wPl6K/OfyBhiUt/qdGfvy08QWGtE0QQAbr+PJbFY/McUD
AEQABgfmOiR+ZocYj6eYkpYs5B12df5c5vD5YqW8sMoxMg/KBshEXwezsKq8WJMUukjcAPmIEoQL
mHaSWTxWH4hlzMmXuoC4sww7+ctaZLiH+/TizJh0g9WvO6uiv7YmANo6cGUhlb+GGy4jSaqcnMKc
cx/87GmjVK4c9Q433p7Fa76GJ+ARwesXTBqcrH+ODYipC68y/RaE8fxX0eWFGdc6WgtDy2ODeOui
XMpk5OdrrZh7WKNN1fMP4z3hq1x0PCeZDGRpa4NPRBgQW7ToBEaPnlmeoklrEG9XOtJfWZ6LKPiC
2sWnvtlqVLUfpgFdKQcn6K1DEFv+Ynru0Q98cmEXkYBOLBnrMFQMlni3oLWiTU1Zvt0ooTdWuJvO
WYlwsiW4akoc5TeCPYG3ew1pkdlgGK+giof0eSELD+LQpxph7kY8/r7JeeUzH0Sf0kONwlas3ZU7
/clQ+q91063zEqZ6iT03ljkNaTN1wxf42uea1KDGBzKB/FcS+bIkmx7nf6xmARMVmH7rL0tJcrQc
XKi6rUIKdTHO3JOSLSlf6X3M6aEWFrp5GQKYZDDefi23TBcMXcowR0Uyog2y90OJGgFu+lpRZ/E4
aGj8s2pNYfvTDR1thmitSUNt3FtDX/5iGMBsa2JQ4O7/yjcBOviR/wOC6SHBNxo6C00o5cl+EjsA
1ErKcsnEMl55QqCYXS14PgG88whPiEka8rOls5WhCjrCzF2PcV8XwRyP/0VPE4RxoQrX2sIJjwz+
5Og/aN8c9rnLvykVAc0vpGK2XwBSKB7qO2gQ6Za19wgvWShuAv/VWu4iUVc8737ty2YZFFpW1j4l
sDN6sgsrjsdIXXVK/ckyq67hf3oZAMc+dMRK5/8X9aF2EH4FcH/Jf09YUmiF8wZOcCM2BWWsTCyL
5nfiQd+GwiUHv27Xufw3N+jgvAhg4Q+WUQMhbKDpANKcQF/2BFQyJeguCOUHcp+lURoghwCpnOUH
N9d7+00BDQuQpY2vNdy1QshD7bwjBhjhov2/dhBakynCsdbudhrLdwyhkgzJxOXmGMEYn2OulfQJ
Xf8rnSyA1v2MOj5S7V1I1ZfUj7FKWq6sy/c16/a4IaN9ZGfot4gIvHWPXkEMqF0OeLUpad7WvWk4
G3HLYFEO1cA/wJeaK8syaZ2A0WczGU8SYdLbKqmpIXgWbNB6/pPAAYaN5W1NxQHQHVk9+xvMJBO3
4mmskoJABf13Vg8PNBaliBHA/w9yVB2bUefVK65k0dumrqaCJC1+QWfWjOFg0SfMIjGykWjqAYBt
nnCArBkns6dyZpHs54x6z5qJAbik/PN9XkcikSbDJ4WHtRyR9krtqiQhLyBK0kwxm2w/6FaWSA02
VSbxbV6lqZexl27UtzekC/qwjnf7/hWx/RGDF7BmrwVowPPHTMJqzHyyvvHDdk0F3llhfCgniPFM
qcU7IxSORN66Mc3gZmTl6nVVHJJ8APPzTBmBMKQJgxntgw+GA89cCUR2CKgV13mwatkp8ZaUawc5
myPdKxqF08R9i/6Wbtugp+A6kTaOjR7ta5W5A7lHvurVPMy+kdFbwYZ5NxUQoXJ8qiGo9VXRhza5
K8nglCS46rvB3e+PxmPeu56b2hfZYbOn7ESNaeR4ahBe3Eh69sUJ7PAj80OljvGaAYu1W8pcuKNi
Cpm9UnMhNiYPPuCu+DCyTZXkifVRrnktGUvsvVNUVs9Ai0GoZdEXfuiRfI2waxpvD4zLdqJs8OtM
WcaX+VtkS55qqqRngBCF7PXJvZcdAokA5PXdypctvuaNya+5KTFOMwkxh/aMCY9MkagF5WxkYZ6M
HKxIPjlHyDTi+Iub3pJxotLeqop8/rOWkqkoT00P1Q5pH2LNkBagUHNI0CiofmLu2z6Fjo8xVbe9
nEdZrJSD+RHo77D4sZOjZepnKAEjSFt/nL/IyitbSXlNLMtoNCK5laneKabmIOOu+v5WVZNB06vs
hIxxYV5Pk3CA3T8y7THYLSijeCJbW+8QDknZvVyssi/Z6IdTwyCOdM4fm82yoyahShv9pADTDDMZ
jDqr+FcxNsWnUjg2t2SyZ6nTPJAgXsPdHkQOtJ2Uv9mi56gNORiKgmkC2qoGjf6S8eHvEVuDPrWN
DoZKIu+nFhYVtmvbvFZpyjN3Bh246sAsST6C3NonL1YzYc1FtWvannwWF19h+JAunXThdcfYpV7N
TEAQrw/VAxZvQTsG9iqlFUnP6VlkGDu6YKetChDMzk06AkHKcuwh7f4FH1F+tboratghnhZU8crp
nCKx7XRk+geAXpJCgy2Yg/Q41g8GPT9Cil5SLj0bO0mShPvJLtyghknf584PkqXHXwVOtzSE92Xc
/mTgU/yEG9botwWXa9gUEe5LQaNCHnwhX6VEqzRtSxEjw4GWjx5ev3q2VKJyMe3fc6WB/BnUWl+y
z2pjrs9f0/SGhw9rw0lVAUyZYDAtiLAdS0HLk5Esz1+mv+8ecY6ur7+D2UlIh4o2URPRTk+PAvqF
J9S/N3KXHq5HgqU3o1I40CmnqpMi6Yj7AL2uTUj9Yqml11UmBfapxRaqb6NQYrG1fznaMz3ayX4W
AB6V8jli2SClQ27yldNwcwXAE7kgHtpfAAspg9o2eBULP12fPayzaPPtAq87mnhqO0PnqO+w88+Z
ptsD9E0vrz3B8dZMQaYROgK5fPe8ID0W3LYEl7ewzUiHh+n3qG+y2FZshrg0hylv3c82TNDdr4d9
GD1mRJZ4+/ir/4s9sIPcsOqAPEC4iEPUheqXYiMap1V2rpYd+YqoYCTOxLdxlQ8zDrY1r/QE/TXm
ryZvKKAGLXL46i0j94rpN5oWHgCGPj7MGreACqoxBcDgD3cFFCqNXcYwoDk1gAlELSNyxD2gFzgD
kyC6xOWbFI8S8TqLp6UvUgvWFiguUxM8tSxDjpEIxucRZ+N7L8ix5+zAVE97qFhcETEaV33OzrUS
A3lcxBe9PFdqa/2EWk42jiMeo1or1+4mxWcXf00jIxawMOvDL1RgvWB/aI2D5IvZG3mnU9RqDZr3
EvN1nLigXpimnzLEuv2qFCn3OCWZK9Ymg3mekvemOMOMt7aD9HT8hMu+vC63vp61CtDssp7IXlYe
pMfkbmf8k+biu6YlRf0E5JpPc1DZ8YDZ1AtdiHNING49TJGFXBJ+F7tU0CVbYbTFSi68RHjZul/P
n67uJg7yPPOc/mvDSHqY/Gr/oFgcuxsRJ4tfH8Eun9EvUWroOzub1KxvWbjjm8BkVtEnR4MLTuwN
AETa5j8oKPRN8s4rSiRQPHgdYKhNt+uQPi4wQd6hfL4Xy/s6d0TIWIBIL0dpiFZQ2T2CRVb0a+nM
B6SXDtUUz5yMkl6WOw41LTa70GW0bpHC9JRI3+1WvcHuo7bVTBxOQpqNTc3ooUeMJ0z8HgrBberE
4DyHO086QRKT5x6jZYpJBv7W7qAzOvouMIXqD1trlG7zE70Jh2CNn2STo9XPXamCSdJmloZLWzLF
eyQSdsUUCmF82leMD8lDBpk+eCxDWHuXurTsE0zUxsqJp/K3Fhxl5MVFBWoEI3veJHpN1eFgAGiE
xUPQ6+OAN52Cb7zJMB7V49NLireUs0NfUxH1cNOMNoSeHVJSHdRr1tjBWl7BHy0BED2KWuaODcSD
MOWEENBYh5fWPGMAzttcV4Em1QzSDt3mXZbvNeOkhkPjKyK3z4+dkCBtbgnuQdRRtOXz1NTMLegg
On7BN6xnrnxUyhTrJDKHsK6rMvM81tmOmPG1W+hsIYgnxEOIWk61KqaVuAeJdjy3vm8lW4WXZaCL
vZPFkjbtSarXGqWhiovoDsNa4lZCHQC/9Kw8C/7Q+296Shv1O4sX/7UztQO/DlopwWlL3Uaq0aiU
XQUygo++RR51cazKI+1v8N00fMBSTMgyR4khzbHO2yHGoH9pv+M1svoozPTyMnfmdtlDKmPT2Uzu
NseQbcQ0s1Ut4Ksza29IowrwfSHFRrdAKj50jGU7HVU3pWRxhyPszhKaKsQr9rb/BXw9AqXeVjyb
Vk0xynOBHwEh3WmyTZc+eB2gW0hzP5hzJDAipu8jSQd6qdizsPTmaJoG3GCPKuAVS6BaZYNPB3Jz
hT0DjCYO4Gv+KabhMYxKWiLtg8/4nsILVZq0Rn2+38gGvFOe11Z+FjzFuQXICUAbTymUZ1BMdIbS
Wxg7sLVQyHVqwSBrmv41+zRB8laiPjv3jwKWVCTPTDk93aSqsbDOfcPNJRCj7rman2S590e1BpRb
RlyIKb6V5TwgzML0DgZOKkEqGpDOv96fE8jJfsPtBTf/VF5/yqWQwwumiySxWXwnzev7tdqfxjsz
eKoV2bPMkiLqD51JDMoC40z5LFXaYFuM+FRH7OOh7kDvwit+RKTkklWSQsp3Vol5jZOhjcbGISWr
1dZzxsTZwKhBnvED/I3xhab53cL56DhLC+iIe4bROahM+Lilh/72WUWhVOz24NuzMITfbfuoXDDQ
ZMLHteYzxcRRdx0CiDekj+u0DqZjvkzrmiKQsLqo//v0gBfvSc4eFgvw0DRn6HjpNb6L6I6EXFOC
9SyFd49a9a49ZnEPvaAg78XFVw5fhCp4s/JiMUcjcRZqjHuoxnhJZ6Pe08I9Kz5m91TUtmQHnSWk
hLtnrLSv6tAi3qRJsmDbsIsf3WCi8dkG9qFFsdfkDVTQQVeD80Gj38QG6Dcl6BVqK67Cb4maF6ml
NuxjYBWutSEicm6RERE0chqzW0t4DbjO1Dl/LJMx63mmLvg8khcVGckWG0URhk65bDFMuReOo+VD
bKYpu7rTfEpXmRcsoHHleKXA7wi+NQ9ZvdLGY4gaX1ynrZSHQODl7tDLrdoIJ0Ggls6NPwnthJAS
U0fkKGIX/kuDX9+mUVquctf/Rvm8Tw+ZruxjMa8nS8A2lEbaqQl+DDlZxfa68Hmjcq1WhjRQNpNr
OAJ6eRnil9c0tnMsRjCIAV772paUcbAGR+ubBxdgMLohc/0HLPywkvGOB9ZmnmriwrPxy//1ZOx4
ZmjnvuQHA1pKEgUT2yFILTfPymSJvlOl53Q2EHn+/PbsJZ8a0BD7tbJgXOBGc/uEVs4yyVtKfuJ+
imDzx/GxI5wi5o7TgwqSIDC4wDSM/44wqdIS2Eocs+hAkTby+XUWoa51AB9/sB3IGi4/Wk13FZKS
38RHyo4QGGnRtYRmWe2NEgyxDdYGRjK+hkZHRdpTHA/1FIjSd5oLCaVBmECeLNOTjii1RwBCoCKU
5tZZlDDsYWTjpcPpTTisEQ4iGurFIg80fiqubB9d9TbMXSHQOxCI493IVqTS+hhY8bsov+3qj6Lu
NG6eu0kxYRWRqwWVmL9mhaIk/tjxVXNinktkcmC2duh1t98eY7Bu0pUCsm2Z15wX3rB5cTftBWxw
03R5FrKSy4/j3aw8yq9CX7JLvVYUGAQyQkzjO+Wv2E0iVodqteH4ZlnKds2NyktFiZBProV2UP7+
E6El7cz3nyf+N1Jzp1CNOxQeW53/W6BGqa/Sk/vwtfeihDlXQhQ3xykeIc0hkcujNWXzknE1l3TE
rpRSjqW84upZPBncp+1D4oh113occYUnz90Y02m5HRi9JVwpsGRapB8UkBEfRHt3hVKtpaDsR0fY
arHCWN6YJUpwDSHjd88ncrCnCBf1iJWZ0Pg3rFCylCXpe0LpWx/jOE+/aBe4stjADPy91QDqkmkI
j0J+XlFu5IbU70uPd1HMwb3x5j+r7WMROMlySdQCrsr/n2nCKuRrNAeXc1nfAM6MT5yJkRjclCms
bPvy7FKVCuPRkE9N6B4l71n8DE+nCo5AnSvP5Wtv+4BWK2OvridwE9ZGLs/WkbGMoSdlURkDdqCj
sjfbz8iMY6fnz26MUSDrqX99fkGbfOWZJxnUbYzX7fGA3ETwOMLbJIFfRiTyOInos3Exg1mfQvwq
5gDFITKjOdO83flAc+tyPaxFYYutsiL3s3OorGLsQVW1uaJzBXkBr3sDrcVmdIDx0EA7uR6LKd4O
sUbNff5i93mnHSRt1V/0S1ePPfHHC7NcVTdX5Nr5yaNaQX1946ocvGupdtD7CTucdG3RoomtkzIN
g2Uc9+/egbbmoDNX55pEPf7HogXwIzSaufRkNf/3dNmLyWnVlDFjV8OqhlvOIZujnlLwNIRhI44e
PHKYxVEBVLGA519hZ/C3tyYvIbIQKqWRHdorCwyH9/fpiTwOgbNdDCI90HtROWR11rVx95g1TEsR
O78PjrD/iWF79C5zxDG7ebk0o7YCm2bbXtYuL9IdJDZARMLjDWoZol9jcUKJQrIsImcxhVbElhRD
hQT3un49/GrhCnBPEAH9zVddzB1c8JW/fMPW4FzZHo5HEjTu3I4AbK+AUvmiBbnQIMyNReF3Klab
Tc62aW1Qijj10hdooFGtaoJH9NurSGl15R6922n8kMjkk50z051XbdDAbq8w+H3VQjheaQXm4WgT
dhvA0i8SPFG5mZwsBphV9qnwe+1JkFDH0cgmFR6Zu8YF8mhrzgW7wQraL5MfaVkPsftqcB30Okh4
+8tNc4oMSKUXWvu4HOMcauV0tJzLUCqAATEsUi1gNJFVCDAbiM9SNNHIG7/3eqxpkJEqEBPtbRpY
/b0jY4m7W+vY/MR+vRCWLN4rQZNYwY+rP4wiP7/g7dKbQBGONBT1qMXTI/qO0dBU4z3VAWBWZosg
U6D7++QDSwL2VfVmTXVQmpbqWY0iKngzlZLzF1+gA+qkEvwpo+6t8MoP98i+eao3CJC10Dr/vdY9
PAqo41JPFnG8n8EoZ64y4g+xDqeCZNJtUonXmu5QPAHex6mlIi/VKHzlyMfPGem/SJn9F6y9KrM+
+TTxeK8h4xezGL7mfPcUiQ5ajwO5AdWDNhBzbdWzPfUBedfHpd3l2tH4fSOzpEGEA9RUxWW27wO8
zUxN9C6j9V/SSiaZJJtgpnQnTb0MAw6YUPq3+7IPkQpJqRv22nfYoTWMynyC/CqNOutWgwNdDMT2
68b3AUPWCKpwslWKs3YgtM0o/lwiSqJcWNZKrbXJ06zzsyEQrpxtqeGf7zZGzWX+nejsXO9T0x1J
ZJutJ4s7PgJFIRSkIlgBp/FEdop9Hnmzls3KHcjirERa8nzQTAZSE88a3+ic2/jFmk427S4h1tut
ERaTMel088g0kebSUThVJ3CXVr2UuwXRymBOjBvsBmCvjTqJ89/Dvu8qVpansoIiqO9VVR97zpPb
OItBkxoUi06LZNxnoh0iAnGIerNykzXjPVABAKKJ0aYA5jOT2QctvRAfeIIzbRhyFoNC80zqoQ8U
dvjHZXxSOEBmmwYxlvDo9reUS0HKmQslZbAJwK8pKHZ3GpmhOSdGzLV4fjZ+sVz/bipFPKPx0Abq
qLYJo3j2K0sgt12ZCep4O9ueP/5aRxay+nc8wjmOFpfyV27lLsVbhWq1mqcUApmL1E9qbvm+KmfM
gteyuDTaARHL6MAxfZa5r2nN2/49QznUNeWrGrk7/wHbsFACOgcQE87KQNlawFsCCnE8MkJQ6E9e
0ECQ7FPhy/RxxcwO4EuFDDILJojhpMT/2B4aJ8fBausTJZxS+RgiWzUbnAe0xeEuCVKk6b2p4uqt
j7VgdNCNAGp3CgKrS/EsGVn7B99zdMcxkFoRQiRBFJJ4K56luq2JWrBfR6kLSy/T5glJVJxs2hD+
oHWfaZTTzkhZVvPOnK+uOBCfrEvNNj5A8ourKUXqW67JAs96poCTrGEQ7uGFTfwIh+B4wf+RiASI
9/L/BrTLkMkSAOf5gugn+Q1CwiCdWfNrhTsCSxN5GtHfg6oxHCfNSP5Wfb/E3LY0lIHSdRNdEOYf
WFz+Yq/fD+bKm3eCnZEn0gsGQzl17gzACBDYxaxLfYJ/otbZzBleRj/4E9TAAlVpizUMIKlp9Yzg
yh6w2qLj5sZEPTLYqTJ56cGAUYCLMVbOZrMJZFsxYU5P0rJ77x4oh5v7GNurG0I/Rx0ixUsGDDQH
wwJQyO5tC+HeFJ+FknEUvbSRKl9CKD5wNLAuSLwkdNRDjKpYG/KzEi825jrDlQXzdumBYzjrDVQo
/H9J0Qp9m2OVkx+YAkVfVWXJVuVSpPfQ41KF9Eg+fPbTPgV/RjaZnwcpUIXpbXnbWj0YtmSnQ9LD
7CE9loDOsBHAfrQC4oOzoo98yKSGPJxar39jq48TIOb6XSM4mOtNLQGr3rjxkjwko9WQyhKu098C
xQlP2hGd6ZGKS0cSZmVZaAZ15YQfsCH7t2R04KLEE6LpBpu/6Vs/ima6DyRPdqRtNUHEd0GqZenn
CsUip+6nJP9jGBGwHi4GRRwpGTtBOIxHYBgcVk0IP2Bhuzm35SF4QRN4zX1XiuPwBe+6s5dI5MGA
FIjniVZYPuOY/QTi7F9R8yz4ZEYvZVt4WvVJKU09TRIlAxoaGdLo9t9+2iu6jXqqW8eLvp1JjAE1
UwNq/043PKzsCs6gU14z5IUNaRDUtJUZ32nOxvE8azYPdzrpVPrCm4/RANm2glMP4Rh3dyXLZeG4
0kStd9B/kxvumean452G1zsUmWyEgks+QMvCQp6JUr/t9La1pz/FxDpcg5gXM0WeygWgAzVdLhFU
VrpV+VigoqWQec05MHMwxY1NdtoUhUAS3TNxqrvJXPmI65P1XWRYiIKKd+XkTwbYY+usZ5ZDcg3u
Ue5csI7IyrkkFsrBBYRhg7Uzpb/Ksev9yakrj1YRCJz4kzW51ZcS2KDTb6aRuIQ98z8lyQRKWsh+
o7aWl6tcNB8Flq1tQWCRsXPerKMlKAjg46TFSq5fXEgsSP5eXg015IexMlLCfCmZ7WC0mjK0avjV
GnZRWkHK+mbP+0QtKiiXcGPJy/Or+nG24vnsRZOuclB1v2fQTTd4t/HWL5zY3B23+fuc3ztqbk2M
BhOKmVFzbbV/AzvhErPNwn4HScq0wsOhnXrPsOc8axRjCc1f/Ek7XNEVpLvp7dFx2akBCKgdyxS8
fGDowi7i4PFmsxP98j9MhxJxg7HGNmKQq7R/PDb2vZwFQFggRlGLknfY9d5tvuoZ5aPf2lZZBDXq
U/p6p0ApXyHlNjYwXpru6MmQjObyTwS2NRGIENaiQCBowf8tO+4B/wgkToZTirBgr+GAyIHhrXOU
HxqYihF8paQt/SJnIk7j5bvOPCrcMeT7Y03nTMKmAlOM1RPZ1Jb89PrFoOoVt0zoIxZmLSVnD90h
TXuanFQy7sBvX/WsR1S7zPba6Sr+i3EmRu0U+tfBwn/hH8IEbRLdIUYwNIvazELRgk3OkpFqwSCm
3k0FyvrSIzGtGorOiyTcMAxVtL/BHXK7DYqYK6so7KWQeERPBS66FxFIrPRbXUYvBSRHM8LeCAvP
naGcUIWNydiasJNXgisdPKC68j4Ro/jsmdvQK5uIdtmz75RnnZSOVczaZnAqdRBL+d+102uTxFab
sUdkI/2Db+voW4D/SW+v2RHZqhCG10whjXkfGf2t/5NS9gC5gdlpTxxxtTLMtfCCY/7SrSPyJr6n
yS7klBBgK/ucVBtcZaDWaGMj4FCx9Tw5BDn0B3lY9kUiK4AaA+83OdYSGvF/nbjhDzroA3oPz9J9
N1fQuOxzpM3vNmp92xZ5w5nedOvy8wOj2qzE5cBo1pWL7lBHXUwfSwb8p/7QXnclysUsBGW5x8Fi
LMzJFPo6ZeXTu5F3zp222+jowPhm0w9Z/ZexgU2o9A/Gp7vnjWimmVdYl+uYzSeIvPJFbL2jA9Eq
Vmiwq1I0H7CS3Psc3F8yub8xiI02jnQ3FOBmeMPNPQtySNOZdo0MHi5J4eh6oDVx/BmlzpidB3UN
RIdkXSE4a7c2t/j5opFdpnQEX7Rp5lhHMwCsNLSwaXLjhmf4czor1EeozwDWNDC83Iu5iOUPsB9K
LtsvTYl2Yk97a0t5Vj4E1rfbQYbsjBH3StB6AlholHUV36+pPmcoSODPwZ1XDinjexk9V6kOXEBC
FZX7j8z6S8rkrK80HJL2ou4QfJul7tHNbHUcbGr7wOkxHQ2k410rqYtKh1EyXGJ68VPZ4224RQo+
kJ8s2qozOhRrCv8MTcO3fEC1s8umBjfSlWno9d+BsJNu7j3yslqrfecvnPzXWyV8XuIACC2+1TS6
hudtWDy6eR749Be5TSZkwKZVigjrZ98gTaiE+jnorvn26hjJns4vp+UMfQPj8pi6P50nxWH/+31p
xMwBUJPLUy/DYe9x4ZcAdtLatrGa/tDW7Y0mVKkc2CQQwxDSzWLmrjYBqEujeIKU+TyzUDBhrwHW
RNVkP6JyExcY1H0D9hQ02jkB1Z6M7tJeM1qBOrz+CxGmEbdGNko2EQzBVTRf/deJs9GBXfcnEW3H
GvN20UgFRn4kDdTexbnR98Fd95AbvAwv7BbZwtxmyx0cvDbRP1nh9FcqbwHtvqwo1X7PnYphFODL
4kEdO1Sg4T5Ug+wh2JU7NFyKcxclz4UWo29gLxbqpplfUrL/wmcH+bIn3s9M5oty/X3jEukGoB+P
X38PNQVkHb1EhDkWHPxHuuYRxdL0zgf3D1FyTN+DbmwVWmO35H9ttJ825DcAGTIX3rgMClQxMBLf
tAYtvmjpVsvYJnST1eyN7LPHqQSimp1RSJRngi+6qGRgAJ86QVICc8fZlZHJJkbH0o4A9XVARGLo
TvwCHo2pUwsJKm0V6Oe4kUoMTx3D9vRTGHDJz2WDpFclLuQfYmgpELTuizZ+LBrxihW0MQwSU/wX
RKzc49fGS3U39lHEdd1lUh/0/o7/QgZ0/ZwcaG9qK0A9I1NIdaYgBcF49FAwqDSaBHEZc8n1IZXo
Qfbn19wtygfbE5cwawPZnHyhZUdM3lhotTuFwwEMiob/JiiJHy5jFg+d8L4P2fqUCI9LaKAKF7HF
QltRnBGMyDhcU55fwKbFZAvnFZSH63N5GhDtRNyLmeytCtZNQTyW2TvfsUNDHmIrLstmWERbJ/Va
e0gLs2OWiB1yNAVJRGIqtHlW01ZkA9DOsVCLrX1Peu6TITuJIdoppbW0cCIclK6HoctgQ2wFXnEd
pKCFUeFJHZaUdx4iEqEjPM1e0e90yHnK6I/udNMqoXd1AeWRQhL5NNn9C/0cuLsXYkBAO5HeT1IE
AX+7qC+hAr0cE4l7ahj1gDmRg1MD+MW8YAPBajSaS8Y3ndd0zXIzaPi3yuWltZ3FhhLwO/BJxzw8
VWfn2uulPJhgDzUtc5UyMbpMy3q+5I8Y01+ZSbxyqc+fgnkBZqMLJvV8xliYR4sEnD3xPwvVvoHY
mCtEzA1lXgmpUxnrJ3SqVcWhqEzcw8icZ4Vfjor7XXahwurhHSAj9W/P6XoNG/i2BEZJmB4Sie6K
YkTvAhIRm/vMPXqRKnEq12HBmYq8KLdfCkRAM8F68SZj+fapXF9pojY5qajx340akLe3ScCQCpdk
HFatQHGRgmdDRYnvi678czF+M1RSMiJcnh+JeJowhDEqqYYo0578KLtadTdPdHUINipeQgW5Y4aM
EBMaaY2xuJm/97a0V41PiEQop9t37asV/HdBECB7fJxY6gFB7Gr/qzK4JuJY4RLD6hJzBimeYBSb
ripaJxoSkkyAxHJepzY09beGxhLKvCZoSVSJkSh3CHrmRuJxqPF8QOOxVWBbAwy4eUZaWnF0r8vj
ijoSz8uem1ahVR1N0o2YGQHnz7pieQnKrj3NmIXiP5XiZpVXc50WlLuT6eCrFAjJoB7wp3kNBSKN
d1ksDU401UWCGJfM872x6hSv1qjohFygtuFTcM0rAdMGqOSLL2koyuv0Son/vXz8UW25Eej4/r2Y
0220d0PFKgeCmoQJ7fusoysqU17vPQ2eBVbgmqRJQeBU8pFSVa3Gd/VKkQ3I12CrlMA/35xbdkJV
y0hC5R9h6daGr/bGh9MfrLABDoX7Mif+BEwkVjMdsoPGzKuKSIiBBn8fy8xmKBrjCYJnBJ8a0L0J
sAdR+1mkZtPypoHnI0cgewQjdGCzGVaGaBXKsO9CqxirZW+D6/R1d8mUMkJ0lKj79WlXYW9wmEbV
DtVpF9wk2jXWDRFig/ijamudcGqFFNFwjdoWe+3EtlvriNZbSSPLFRDvHN8B5Y5HwlIVLe8SM6aW
2EXgOhA86NNUGygOQPyWq1pwk3dsCU/h4hOgZFe/OtKZYU5275kCzHa5oH5Xkr46J3yaZgwTj5E5
sCUaoXzwLxtD863DT0JhxxLn0XYlRuOEP4YBSuRhVAsbmzmUeF/VxXUTIA1B/fIWe8Y1YfsLXO/T
cuiOnXurKbZOUjP8wV5/Jdld93p1rd/hn6UHLkvtL+TvYQv74Sn+7f0OobYcJ7tagni7+V1zglVh
5jF6BNvQz3J0flf55tr/GUdHoKaW5wqETnD/CvAt+2T0ETRQVKoDFiGcuXelSthjztlhora4ifOU
uwToFEty0vkJKVV2LrfqfVyF3NLcKQgx/Gc9A9/KbyHjXUN9S5yxRtWoYv7CG5ODtKdSP/PA7jX3
y3PNdxZPjJD/5XbF0EaLnGi8GdHLCXQ82h2dqEtiRdlpcp4RGJBGiEYjhAUR+4LyhpvBIKuQhj+b
YN9hx/7UcLQnk9uO8mxu+a+DXz2bazx+pw2G7xzerH4NA1uPNCb0CXqSeFJzLYkb1FTz7R3fuxFn
ooCJ5XG5ZfgH8gdm28X1A07q7LO4wVHnRVcxLXwqnS5DICCmiWduR1dY2HqCB55ZuIQmy1tbs+Tw
YgbIDNrnJF3WdNHoOlgpc+Z2d5bAGLBGf7Nd6jPgYqx6hGG3iOM9rs/dOjWzZInHFfry6+teHmEY
JAVzXdIE1R0KsFSS+7IYBStFguwAaC+vYcE1JNmpAREknCiv5P7Z/CmgYGeBRtBTdpTNRl34su2W
BR5/VGr6Y9PGbNHIovCgcy/5c9+a9qTKqPrLXIw72IV6au5Ms2hiSpPt8RnHJEb7wMMfRjXbVBZg
BKPjB9ElMjjfFY8RgqrwAVp9c0xMjerhtGx4+AvXXCQ+ZHDybEic5royP7ulXR6bEud1ja6m6DGN
+9KPEBpsrpUCQ1vNTbNiQGB/EfNo1vQkYUHzmjEziI9YgGbDFRsUn/e93OI09nFlKMe7N17llhAa
gKGh6XjlDPRO4CsANfn+OWHE8DcdwKJGuk7HYoik09D0o9IyMUNJoY+keRy6SI4djF9685VTnrJO
Hjf11yXN5nde3mHp4zn8xG76yGIX0d8fcayofrw82ST3LEnyzMlmdupO1c4AZqVHXecjAHiAS8mV
o+KTZUgQJv3JivBgZV1jtWs3lJIaUBoXS7sO9P4QSN9nzBfQRwu6OnLEl7QdZYFsmehknBZzFb/o
CIIUh90NS+iARQmYHxOrUtZuvbrA8+XHItPctJevx2SZG3IhJ3rthVrFzgFKxrvAIzfrSu71ToDd
W9+nKSeEmZ7QKUFLVjZvSUvoEGSoy/of8MOTUOtYb8KfS/P/fdEZywsCyzesouaj6I2qrchYee1s
74fB3ErqXHlf2BfZE2ObpIlAqI/IlF9h0KVp1mk5xW2ilXolYc6YtPUf0sJLK1hW1GamjeSyeHM4
8cQTyH0EZQB61l9uT5pgWBsr1VTzGZrBuagQikTbZyjOLFjub5USwvTd0bsN7gBOfmcmmMHth2lZ
XEtbQlaw0CXnwleOB88kK54RnW5G1iS8J8COiv4BIzcYvJ3yS2zhvDiHoVVG9QlU5pqDgugo9Udq
xfJjFXPWsv/wc2Yfe3RMK/S+51ZlQ4svMA8s+l4GoIya0uEG5mPRWxBJLkdMFWO01+r1Ie9UDQwJ
ImpdFzn8zhe53I6uebNqz6JO5yYcLDeu+HZiIkckpd28YGgt2jVdbzB2eOB12CNuhI24iNkSJhr9
xooj9AnVV4ogSCZZZQQ3+2jULGgbA190YX2mSrs4Tv4MQUEUtTNX9NUSWTRfqdjz90W4gWRa1kjs
wums/IuSAuNswAon5cUsdyVllVGFG3Ii0Ysok80hvBXzcv2o9Pyx1x+R0qsqht2uNwaO0sNu4Kig
8L3qK2rKs/OAaeTGRaMtQkMg+vUIJUT06MAEwu7MsLAXfuwC4qixKW2XllSiJsghbaf8KyW1uqPr
cJpXgHsTeJ4zPFLvfu6TxOLGS50VisJePLznONyra3UpKL9uC22aXSksbjJSPyZe/0aT/ray+KFI
gym7blR2Ijo0YJnhrTPWY11EhjjwvuPJTTR+3aHGEzqWidhAkGyeEinuHh0xtlGt8Ohzt4KxUXpJ
SBvawloT/YuPLowzSftGWw0veKWhA36JJujgaSI87nnyxalHN0uu4+FriFDHBtpUuZ8lC/sSUTFX
VvW0TNTuogIEM5yyYzHXC5SZtLKlnreFkhdGc3mT6Cn8N4pHpA7bWJOKpY+oMmoqEQdWKsCFBdZ2
aOc6/igMkIIqlkpjLBPrujbmeTfuonIsldfrsYZmvKWsMh+MeL1VkhFhzQ6kjdp9DKshJugH0zdN
ZySoHMssRcfZW4o4+FS6GZjfBfSELUaXn6nJN1fL/fAxZ6+1ndlR1i+gSjj+7YdrcSY62vuY7r/Y
xK59L+a8RtEgPheOrZctnLqmuzH1LLX1wbJvejR/YlpVkFVAoXaDPz/Em/0hfY0GB93gIna9cUkG
NgGflgYidNbpPZmQI5g+UHgmnqe2oLU644dHe8GZvR7cNIcNC2brFsDYN8Yuqtu3zueQ0f+usbBw
bpc5911P2yAHMKE8asdZY5CX1Xz97+mqXGzuuowf17dzQGJWgXc4dkeXYnPKiUb7SEGizd9+FreQ
Z2I3B8GDU6eHQi4HIbqn+vF8+5QvgZyQGW2NuJAcSNUswcZUobBdw1uuGvfeadMP4vLgn8gVNTRc
wbcOyCKS9tbjMIqdIZi7MghkjTveT9rbXYUBgUTqWBFljm8wUEfHkdKFZacRPRr0upSAWCHCybJA
bE8TvyUXYsib/hpO7cvTDKno1yLlRzAn96n42cTkgr508/7LnuwIBYAawm78A1IGTxPB9KYewKho
U4cfi0YP7l4VxQ9O+icgRl89OoP0VTDKPOb85i0H2TzxH72R+EQkk47/qNBOiL8UWtwgCzLg3R8A
OLZYiMDlnopndoJF1AEyC/XINasfaNtQI9yFP+vY+twc8SImGns5QaBJVPBe8zbg8k9IU+NDChS8
IUzNftRD7nD4k2ZYz2dhLm5tdTfZuvnJITZiSNBeyORhHJJzAW7BKVAxSNBoCaNjXlnPdelAmABT
9COgjRW6IR2RR50bOdauRFa6l/wStRBrGV73PI+a4anQmjiNFvDJi5p5DTwO2LNqFLeosMGGQSpV
2C4ydWK9Kh4BDgHghrwqCWpn3dOchJosrnP51I4sYeRBsC63/eHX0OwsT2BL4FF6jsWWtqXypy+o
JuHF4RYUR7Lak+V2eLhInEhAa3Tr5ZKe5urIVAxw+5lo+oG4dOGrlaLxXyxnd8LmVC54eZler3wA
zSooSaZIf8b1q2DV1O/jNgnhs0nPXgpVBauLwWIJ9Z5jnN9zvDtt928PaK1nDwbmRXPczMVBmBXs
ZnXsUMnskVEoe/eZOYcNJeiZYpbrAE3I/5BqFRX3N5LGJgiLyAgpEzFfZD5NLpeO2zfPbjVSibun
4KiU0iljN0fZ4fQpIdZwW90XblTOBM2zNBHk2+3LdmDhjt8wYq57JbuxBN/5+NHPL/BIUEYA3HK5
c7nAwwzGeiroAHehgGIYnJpv49YwQirg3ORxg3wW0e/GFkKQ+o4gZMcn4wSFylFzSxZVZF+wIDkH
BXl4IltL7P55IaHarZie3kkinsi2XAslIJqlg3DvdnVOIAxsC44mPMwwi+Mg+Lc6cYPTYSh7Giu8
YgBeHoopXQ3jCZRTgRgbOOVavwhhSeZAYmeYJDb/iVn0BLhMhuJ974m7JVieYFo3Ss/2LpW0+Ucd
U2AmpBa8hP+IWMHk3SIX6GtKtwJ3SDeFOS3jfSfwH6NM2mZ+9K/Gum3SlGLzKxy6M4H+sXFAfhc1
yTVv6M2YpKVMVe2yTp69caiMvZYnHY084jlwhe/3GWG1PXRgGR1EnKSpkLGBfM/QyTHoZDhFTO+z
QR0DuMNY28GVhLeYHRgvwtbjtp2QDmC/PYLMEyHy92XGyvTLX9pCjA+o6NZin5RLZG8NiEQqXcQ9
VTVv8ARLdkSbk5eCfB15WolnocLa7pvcD1Cl+GbLGUxGeOGXfiTk8xo7N51oVLMQeeK/hBNcvnyr
s6rZGObW252SSoCalU7k5Sx9KAKE9MtvHUUTM3y+CI6tZsrNcM65xdR7snNN3neGU9M4vJWfanr/
/C61O/okJGhIVcMRvoYzpjXKozKHF04Jlt+YxdG4XdDKDEm6cMH31ly8Q8kQx5Dko19ucqi8lYGf
tlVj3mUUeBYsDaS0D5KLnUW3cy9WYkcNXqWlY+MB2CPQIdpofKo5Fn52ktoHkcPbyHdFKy0e7QjJ
nw069LEhIHqO4Hp3mN6GdTShY4j8fmMXNwabVmAEKJLgOKj7RWnsnCb/isiQgJevaNZ7qE8KajNW
HfxXGpFHV9j5Ze4kQvK+y5w6NQxBAFbC7OunT5cc4wHhduurTqmLqkyzgKzgRjBYr8wvIxrXCi4P
cQAweCQdaqJ6lJi/3Q8hRo/NrEoIC6H8Wn6JcCS8mAl8j+msFy0UqFy4uzZU3Y+VUC49EO+5JH/Y
EdihwjBwg2rreZZG6RDomEPfkVEBg9q8g0CFpG3qDUxjAOtS/w56aS3WG4CKJWVFnxUvnuNvid9h
a4XDMjIQO6yc9v6iu3UiEOsxoiWGjqTKGscSQHktyl1qP5MIw2tFBsoNbMqVlyddQ2+2iaZ6w7ny
j1wdt9hbLYFS09t6ECAg469yL7Gx1zReTbAgQBCD7GP4OZOETbYEs5uQcKHqZhmDN1FCPwIyoth1
K22JE51HQhGs2Fm+xZCdzNeA+o4y9GzWkGQyClABbfYCrIji4+Vt9kbIB/oQX9Uu+/8nBBoLqVac
3ikDj4cVaVLkqRIFezIwTEBbzZsm1Q+IlqQRuuO1Ch2g43ikVWEe9H/U0UCv/Wm6cE1d6dxAeCfN
w4V+rOqSeRV680ZgwAQ/uUEQn8tea35p47Qz7dCCtjeDrnzP7h260fSSjJu3WD4em9BClAB6wDzC
O+1MKQjo3s5BUPy9NVqZaobzBFqOW8yUFAyJmiKvsQ2cNTYREKgcZZ8JubdHbvuGukZM0Tk2j/bz
jqrZ0BOgt7rVXrguuKFtJDUMIbOBYxtjdhzBpqR1GRRJdrxeu5LQXUIh1OmjaElOkS0HtA7aaMmO
dSl9QbldX3Mzs/sejzzZ4uyNgdPx+yZ9h4G/XtGWf5UQrQCGDzyNnWKbA/DC74ZWzGQAtcECGRsP
vP/6TC6x02GCo5IQbWmRdGDGR3+sOyQb1UljZRWbcfHioxuGJQAJ4TxVVHycpPTl2gw4uK7Q4NaK
WvWbLtK1cCl5UbZlRGs5UCUpwsiYL+4KA9xVwlIxDfvbqKZfdbDSo73lMwxYok0EoZIL5xu69x3m
FkgqSOVRBfAzSZPA9wHx+Ka31qHTNC4jlbPY0UpObkyXJsn0K017oPaeIoyzpWb3HyaDnQnJqcfy
RE+LwODdzWjHj7xmCaqHFKQPUlzcJgEFfDlQPem2gOoc6q2NwIiwTEa+f0S4Qh8U0xMX/p6cW2sy
mS3j8n9EtH1CWXhNweISB26ax6M3rmvPhQYV9Scp1fMZ+S3OAIzWoaAO0CipaQTeoYJe6l8Agg9e
j6i80wgddH5xJDgEM5KCZ5v/NRbL8LgtVAWwF77pnesN4S+spiP/RY0xDrO6xgmCKGWeH4/LXesb
LcExNi8ZPTXaenWjzJMj6GbaAxwiZ642bs+0LnxSkhnK9Lcj1upDndtjgmxlMpoWpmI604cCLF4f
2fXml15hVLVMSr4wC/t2+425X0E22ei8iIR/HYciQSuoHZ71/4JDX1Y4tISkwht8ig3K6RjpgVOS
HofJ/Bqdp9H9aMM3pb9ydLw1Yay6sw5yHpkK7j0xHGeMVo95HKciC2yH4I/hpW7VYk7ITAXUE4zE
UA5F2s73j18rf6wSV/ZglfUrFdExHsKChaUyXeUWxbbOfO31rjwUa0ZbQoznf3U9/GBuiGcsFowM
doh8bK3Qu4U1WNNqi27S+isfV9ZTCO749LJK3VqfarZwZiajZ99rJAVtNUqILzL5ZLyvS+BydjM1
CGeqS0BKyGs7nZOmwIrrCichAryu+xzAOVj7eC6rxwanSkKSdvmMydzGthkFQcV+/0BL8tA0zAip
wp5fUAlN6OlDL9yGnQImTbXdX4I4aFxAL/yffHdFPABIXMI7n3G1qfW8IpLZ7YDZtR9cIzpPdXag
fguEN6006V5nFvWk50qq92WpN4cHA6kNC5Tv3uwShXULONk67iYWMoHEP/tNA4zZ/Rz9QA3JxLfA
Wr+argoXvPoSHg2lNOZDySHVRp7lnQavxhRgOf8jl7MdBUFoAAjqo4azZI8H7PYcsGm/pFtNIg/n
EPCgm+uo4Ip+xCZvG6q7lHKl8AE2318kNeTMQVAyCQ8UJ2m6OcUce/TAZgl8q5tgkvU9l9VEqHhp
GNDXXWMF7JMXpJuqL0ZixZo45/3w5HD8prqQCzqYBei9ythOTcN/M38vJq/SPWhvXV5xqJeH1JPS
g0mGMMJhetSVrefZeD4J7z61bSAd7RA+kW8YwuYE5KL/GBNCcWmQe+tk6g6XU2ajex1Qy643dMBQ
AW/U0gA3/0COAL6OJfB9gl+I96gLnaxN5ILLuw9G7mGuoO2WBIYGRfTgLQnn4IeMrfy/ifEQz5ww
X/R6xafMljbDcdxavo6UK2vQtUP+Om/J4tA2bKxW/pIZ8X+qUsHyVRBYDYX9pDNn5Osn9KV5/5sS
ciua1Fo9zT+GWW1Yfo7NXOOuLnqv6u0GKaZz4Z8uwwufhIYWLiT1KwCwvMF06J4UOOra2wn/UbkW
fsUioLmT/CUlmMHT5OULXYY6qtH0zDNMQylaDvXyeIFwLs54IOSo/Cut/QM+WStYGncU7t3bF/tt
nkovrqE5Tm05m6zPbEkeRZq1bx1T0BMtQsfLJialZPH7HJhRnDVf3hlmjLqWFGnKnb33g+DfePwG
CCz9+4MW/S7z0l/zYJVW6qC5wl/Gk037an+nRWBl9v+tJcS53iiocdeSyleqYy+p+R3h3l2KPghF
At8YohhrMatmtsWiRox0tDY/XKbclMQFM9qQ1Z5Q/5ltaSInk7H0zfpQ3zBVvM/7CbvvmtuLFh7X
2gbhuocc8xN+2fAPFylB2H6seLxkgWTdH/ugjLa8s8RQl9Krm0J7PBhtcM2QIc6CmoKU4jCtVQ2P
xTOfQ8uwrAzAriky/EsTidrDpRHqNcj6/BUtT7ae3pW0TfgLbwqPJn9tU4tBgFtPimfQJHISsABA
NGhGssrPnST5If1EHIyXMg80BcqHAgNRRdoOjMWCLUq671CzLoKVwxPfOtV4cMRSc3RdIVYqVuwo
YUdc9A/oF1qgC3vra24u5WSVBXC1yjHr4TmZ/ibf1gxr/924WxuzSrpk3eygA6/ckYIwoG6tVFzr
4EASi+Bkt0iYTm/DLVfOyvpc/5MBHjibHslxPZILk14o5R1oRKaL7cHegV/mpO71xuEGaxHjuV9v
XnkigWXPWB/w4YScSt6oa8F2i+3UsPhcUHZHbnXFB3tenBM5jQ1QTxE2X54Y4NiUqqxGWnXjpCsk
osUvyEyPT8fpRMw2zwxO6Yedr04V8g8W84xVW2/ZvUj+bLN2o1NRLS0IqoKDCD/NAsn0ccL9zqZ0
eRVMruGczOME7OtCrpr09GPXKKqyEdzLg9HjakY95tbkUhQkdcGpetk3ZubsT67CMuPt/MOGwHyP
p9ZFhFKXWUfNkuqGVjVpDewL9t4TK1DnfsSXwvDnjDaztBL0X+D7w3idAW7PhI3G56cWwWVf6CM0
MrlOnQFKriTI5x2Dfm1oVqXcGeVvXrsLDQTXAUtAGDxBDWAJr4ys6me0HtHlnSiD9rohA1a4aE4b
5E2PYQ5bNrU6lKn3s5GZWHDhDOpd9SES2Jh+6EGVZqsck/w37SiIivxQi0E4RLYBYz3sB/4PoOdE
YM+FoX8Amuuz3eIX3tKxYLUlF69k5XFpHqMoSDKLs6K3P8dlyv+fELJRJ2q1QSDHmyeQeO3qQZ36
qR5tifxiVoqrMgJs4Uo8wNrAQsrvYbqkN8pbjBkymspOZR3W2wL8VSBCqqlJ7ENGhM47HXmvKNW+
uAaxbzyhp+8Objyun6bvmvvb9lID71DtQv193XeBM0TADhj47t/MG7eNOUWqfos4WyvdAr43WpN3
EmWumy0Iqzu1ZvGrJhyeFZTWHh5GrW/W2Hq7jC+9jdPQyEkcJsXoNm/JSykH4xirIZbow1z0oa1h
/YkR2r0KdkwXd4ghzFC9vq/mYBwItFa4qDYr+7ELMhMQ1j4UxnpEEZ2gL0FK3MjBW3E2D8/xJvnN
kD0CzYzVDGijJN+EjcYYcVjj+A9BWeJBmnuo529BY9yj7YlVwgE3lHrX9CS0SFRlMyQNfgrY1jNy
YqJFO40hJOu8YsJayGj/7ju0j8/gmdiimZU8qG3hB4AWsMavcUqNq2dQzZtvXOftdPrqyT1GmuAv
0F3Cya/2DOM/2SScw7CXw62BJ/p+q5zFzxETYcdj60UjisAI8oIjUjnUnF6fiNTHOUWqIGAf+5FD
ZHPd4Cynuryw/Npe2rMcdyGmOr/E2xFLfI+ZQaVt+zqCVXewY1BoO1HhoDfDHqN2em2FWk+7llaC
4PyvMPYpTqbV+lfh3lgmoQmsa2fMJ9xH4He+iM/B7tYBfNVmYSF/wsaEvueoEbpjWDbC3kYeGFiU
8++48L/qhe2FCYkWY+8P4/w3onqAY9WL6v2XW3e7ag+5sEVlp867cQeKjqQmwwlj0wq9xPW65VeK
dKWqYuUEH7CEcA9z/poOua3v513QRJN90rwHug76ptmSB1l3zGubx9/4PbiVtB7B7/gaKE8VYvGv
2P8gxyc8EoYVu5jaH3429tJXYyzq7rVJnXtN5tp7LJ/fMMvIRybOKN9NUnn8v1vX5C+TCXnC9YAd
Wk8dZIptUk2x09Mf/43sKzCnd8tzYLSBs6wHshjfis08BlOmKSkhhXVKE9TE0ExcxKRuYiJY5vdR
EpUbDQfjOEpUobD3e8qxR8Yh8kb1bMz03/G7rG4iAhnt7nPr+/yx93/aCfEKx2V3pYYxyes7+OcE
58JWcZnkjFe5XnvMt9IRWlZXvCYzmZp5+GWrzBF6L7cLFZmBNZLe7aTRO2v/G6klisF+7ZcDEy7y
RRZMikLEIuueGzysbkHyw868HoswUQk8ln6Nkgoz6K+kTsRk+qWOqvTjK+3ti3kA7u6D1/JWi7bi
r4Yi40Ha608ughgMSOxx6EXF05NT9E9+bvPUGZdb/GZvks9u/qIM4ZeYlUlrXAtOelwjyxd18Ovc
+UaB5Fgp5hAoTuH3V//NcX/CY+xn4cNycwfQygbTC3QtgIKs6FowfDUmnmAJAFne6jY/jc1SrMfi
Ktqj9120KvdH5R//0HmGzXUg/CNbCNh/pVhiAvgemkzgvy6jhPCyXwYCDDE8j5clP0PATYYCtcjr
VdmJTpZx5LFfpwNZAOcK2R8g2aCJPy9gIVVvYKdgEkBh7ibHgy1iOuNiOiIJTliOOvKdmrYlV1w0
Y6dS+qhfqhb1UL9rdqDumsgKcGp0JCCLMuR7HSyTWRJcHMq92cC+C47KXrFp4w25eFP7gm9DjcTq
KFApsyp+B09qP9iT+3iAKnbbS2ci6wRtZkzPnskQhkTRry4KsKjpGiRO1RClmDi2llkCusGDOH3l
Qv3CgdnO3dAqnYZ0buQqTJgfXHLWY3VNNY6xTydr4Cy8az/8BLRdgTTOOqUajM+1MOwx1ooWqG8C
VOKjGTl40k641re662w0B7RFFhlN4a3R1k0EaZD2+O+4PuRBMrUIDl6k2yZzmBThyDhgut/E0O3Z
aYM028ZSibanUaew8kus91d0LSW3mim8jAITv1LX5wAwUcqspIxtdOiw9MEK4tMJOXiAom7n2fPS
qvzkJITX7aUJ8ESq7KnqosP07TTcmi53ayd038Q8oY/qPTsh9a2HLXj6lWPh4ilOaNY4l+BXtnWP
IA0gP9/B+cVYkshMJu4/s9eGEz/9vcJ7UPFQ1oVESKbTLrqu8pp2iTios2ACm2qUNhX7UQ/GhOUV
1JzuYbIMIWOTDGmHyusNeHI+loB84CXDemsw/1yHto69gxU/JJ+TvYDgP/HBZTzp4/0DxsrTVpqi
ASd9FHt2E4+D+AjHodf+8xR0jw/uFAw3Udsbm1DA7RMuVc6dUaGks7h9EDCDf2Ju7uhAVfXdlWZP
IXqm10mypTCShK9sKBfPmWU6xosDhHaBX6cB7WHnvicUG9FwpeWbY6o+tFcIbcBRvfG86E3nixWX
2hqIcnGrH02Uz24Ija4ijVi97q+fS8vEeDJ+m+C1SFK5XX0MFlfKkmZW/ihNSrSTHWM4DZ+xx43I
WY3Qb8JVTtbXbwW2HHw6PAQ7v1r77L78fKPSm4CQ/hMAp6XZCZV67WD2nkAWOiRKJclHLZQl0Cn0
dSvsNjl/zHKvwkhAXDHo4inwrhdBloCgRxzRzX5t/Re7CGAhpUklT9Yn2PFHWMVZOym2pd9nTU4U
4FEeiP/cGm5XF/20qdTCMHu7r7Y5Z/qZbxmRBGpLSqdg7EWysDBRXClbmn3cIRotAgS4+w7FWhWM
ks+zG6stHpC9RCTEtiDt/Gad/ysg+655GfKh+AS3gAxaJ0VENR3Jvupxz5umZ5auhEyMD6r/pbVE
dz2OFY6ZniC0h3SsMEpdmKaEB3KgHSWbOei0ye6/3rmWcvjkSd91pugzzMIIbWXOiE8sogGyI3N1
2ufbMBJBw6R2k97LOTg3ujxUS6sojWhUCjjIXN0FJLF+vOznh3Hhs58hkj5LO8X5t3+vrOGw5vYh
MidaNSLh0ETJkzbY+Rcz9YPbHQLsErYZ93vv2zlG2alzFC40v7fFKXdFpbPrWkfzicQYlRtUMWvh
MLyENVlpYIM3LJu53iQPbsr76tss1qmvF/2UyXiPbqv0RAYsw4dIw57L9JY3XbX2bLM1qiNFxhvs
FnASGPQ1wg0R8KPjazceOYP/m2GLFt0xd+p/8wcoWKEO7WeenKLFwUd+1FFjBLvL/ZjZfR0WP4/g
mu6QSkezX+wiLiY1iMAWFXp7RzAUWFw5E/9vkYOUXzDiBZeUgvCTqZUIh5YmaUXmHaN+sNSl5Czx
0Gb/8j07Quhq77xFCA1DhTxkg7eiVL/D8R5i8ZXYpZElq/3O6tm8J3s8ppO9EAmAquustwOnI2CV
848r4RzzP1cI317a07/57CltVMKvS9HpnhYKjPB5CcZALyOWqIVP6Tgg4EoqKoCVSUZNMJR1LjrT
Sv5EVsLUHtbxoQa0e0+u3R5qFiLPHAG+MZbPqz4In3i+LsJnDycY042gkalxkOuPS9XvI6qXeaH+
ftUoNFi5TsuTpvS9ogK5DitjUtn3l76vQmNhgZIKhzmsiqteUE497A5dtEbFJYDMfUS6XZl5sjJW
NmA24KUcpHAE/oGkN3AQpdmzqCbUgFWAX4DQpd4613OVy8YpV6BdrCGHiEp90ZjF9MxPY5FiMC7h
qJv8b40N7sWe/GZfvg5/CUWIVG8E5OQNt5gJnKJBhfeLiJAm2gc6ap19ibONq9HoOm2h3kzlf6IB
cEBmuLSKOwsHs8ebCmi7P4y9tyun2OI+a96aA6z/YkQBXplKuIn+rpUS5KT3Pl6nRJRGX1OhWvNE
48ZhsRO9t7pmjcHAJzVqqyaE3II3+lTmreX9ejamhB/0Qn1J/MmdNoxoaJSSj4Fsxg1cS15pV1bV
Zd1WzUetKLNG72MY6k5R+Re01f7yx5himV4p2oPE5m0A/SnJCtNUq24j+CT+uRKUpHP7SVZitI+g
j3TAy2R+EztYN4QLWr+OtpVf2LJT41B06YT67rkK0l25TOBOWhhLOWHn+HoRSQVv9ETVwqBHgkGM
2TWf+tVjYSH55OLwAXQBqONCuJTz0AFExzo2zDD13q64a8ynNwoOPQlWjXPR4SQnM1zM/wSXMcV1
dw3JrmK1E27Li7zFng45PowpCV4RtD0nZOapWpae5G7LTjXFutIwOtKEt1sN3zwF135yqY1yHbSz
vRyyRCcV1VVPAdywY/LXdfKCTEVOeAmXoUgEcNjhbyi6M2qbtbYx19DqiASvsrsharD0ALKDV+OT
Mh9VbGV8VnZvN0ey/VCHa1EGc46wMp3ZaNUMcdsjdB+7f/fLUvhSXsHsh1TODC79rawEUdxHxPjk
NjsdAtlf4THF0n47r9BG2AF0UV2HTpNU0YHdnL/LheD64VKDOmPaY+SCtI+k3G7IZHxu1S21a6Om
TSF+dNhMY5i8I6hBizdtGoHSrjmCeEG7RJHvfWBr8/+AKwu/x4a3m23jUPjbAjhCwGxJPRoANULr
Cc2c/46Ee8TUZWb4TQJQ8eA+QaezscpGjNRaaBelGR3LHH3e1nvhAVKg4SbPmgAcMTUGyUXN8n5x
ug3j38gzboZjRkGiyOjltpY77Mp858vZuhCCfcouNNHq6R+ETRx/axnogXOfpjrEeqY9BfSYf2U6
gIqmQKJLnN4GbliHVE824Bsk3asz+raNMMkxJIXB8Fw0PQ58OedonwlRQk+5FhsFunTK8Uv/pQOZ
GLj6+f4usaVPFjrd/qfUZwq4DBV4xXcSSkXFyVNe7RU3tzodNNhNCAtwVrkTE15RD0fgKwVSpnoI
U9vvcj2gfNSE/Pn11k9Brs/akQQgCmb7d/wuuOfXTEcubEIsNSGNGBMBr2DGQwe2JlTCXAIW5n58
OwGLBcAjGRrH6m69Iw5H/QgmEwnHJuRleN23uCyPiNWKIYO0wudFjAlLtAknntamlvnVci1Mj9Zv
wxNxZDwxEsfWe2KkPJh4Va392UIJY3rq+Gh6ZiiIcrBeqYZcr54o70DSLZ2SsmNG01CnmfH16Bas
vqGhZq4CYAnk9t5g3ZX6He8RKsMny+L0MHL4fkLNSwYoFnOKZAeYbK/3oINMyCtvBR09iMgKS4C2
vQ53TfV19Svb2yJq8+RCHxvUDfADARg77qhpXNf6l5aPI+zdrW7FA/G2YTQlQpZ1B2CXPdD6R/Zi
Gxx0vAJM8pyJZ2K+NBuYvqeZAqNzOwZXKfULCMfNkyBCvEWb3ZH5t3rz3GIuIdGY3JztO9bLSKeq
KHq6iv0hJd46/zLpgST1s8Ne0fFnAHLqJRkMVvZDnrv1c6XPJgDwJ0TQZTOdaA9UKYLbNQGE/4+s
jlOGWxuay25aFmIx4c0qS6sG64MdeSkqVsX/V/rmh790RytpGEFaDnFck6r3uj8cu+6HDQNsH8Bx
lL3kPLYPqiXqNg7c3qWiZt6Ai/r7KXXQ3Rl7g66SI7gQVAy6nfCB3j1GVDwxI5IUJLw2UCGVmPDN
6ktzdDqk0CpaX7Oe55t0eWhI/k8dY+6F6w//mLmO9ggo8Z8UHZJEKv4GwKSX3g3Ykg5rm9qaqBPG
ysjjzHFBfvtxspEsRiSEADb0MAC/I1ncL2N73BHRT44E4NQVe6BMw78A72+n5L4Azv7sgrkqnyqE
3jkxY1c9WaQwS5fRmznNSDtAHXtnlvO72G8owiAvTuX99z2nz2OuaNdn8Nr2kJPdvS967ZLGB0gX
XgOi/KkkiCYw4xkDgbtjObXsn050a6Ms1yG9R4oUw1fmyx6RglEDMiUR5tJBWw7LprgxYQ7Qe3Od
IWA9/x7peKCNiFhhHnsnXJj9UxsRhc7cjzfXRmZMb5vKR/bCjGortwBNClPJYxLIpEFjiwR98Ahv
0hP3rsP+4P8uQ/+g48+hZurXn8UQO1rj4urmn22sBMatieEVb5XuX6ZYRYrl5+gujZ+rUHJyIoHC
XX93jSNAWWI5CjzMNs1aQePve89xvC1cmMwAatJwvk2rKpCIXyGRvkLjqZaDy4ydyMaeFY6YeZ4i
tDpSi24pygy0F2w7v6PoLylmGYLS++T/3KWn1XemKR8fUAztq0HUwWHCpUSKNtaXlDec+KNPXeG2
lE+49d8Z/ugpT4HHY9n+0u+uVkJ2VAFdaywAVzLGwl+5r0mv7oP6fVCcUeFepQ8lW3Pq7yuOU270
8065SkJlbFH2zrzH1dDVRay+hUTIpofUGtZ1s/2FddFlF5KG/2bNNvNbMwLUtzAFrudOyD8ZeUfN
QTkZQmLyKrE0FMx3moLw7Va8suQSeC0wQuLy4uxYI6zwNuv/60Y4zIvMDUhOZpJD/VvivQA1Epqc
zE38VoWDKOjQ3jaJAbqx6D9cUvapibRut59HODNwKVY30DRt3qHDP710qTCe3f5nsFT/c0FyoHxg
2EHT9nPqDLXVTM4dB8F9J/9ZPQ4g6VsU5+CX7EyU8eDn/19V+qTQTd7KUwgUXzQEZt/yvpkWNCq3
ElygHEy1FhAaBklDVnfmL7WlzKyMghw4WpReFocTyG9HeTMNI/kIl6E5jKUyHd11kZqoztVOc4rO
tNPL5G8O7Sp9MVMmrIEXPHHQgt9Y8Y6rjZ251L889fPIKhfi2pA2SPCtCCySZQI2hSr1bwHeyogK
igLK6rH1GhvjWZ+rooOeSXWeZfzIBJJS0Y6rCoFbimVtfTSZVpcJhSDiSydnWR0X65e88cLcGkxw
DDXphLUUdPZwNhD9E3WMV0ATk7rxxX4/AH8AnT4ZjoG/5wSFXP4cC33JGvBKK5Cztp0YF6ncQJX/
mPfGnfLWW1G/2U3r5LD3LBOWRuLcxvuucWjoPVXTtqH0egQJbCFbPUZXFihqpo2pQ6PePTd5moeF
pSOkVstmlrx8W9bPVy0v/h6ozOuI4uw9d6+1kecgixjL6aGhIrfMDRbGKMYiQRICf6HWmM0hB7/X
DK/uvSKETG2V7pQ6wO9wybp7rzp56u+m2XSaewdUOuXB5UwXIs6ii3ig8NVKftVJqgjRpcalDF4c
8pM05vJpD+EkiXInb8rXXmRZLk4Uj70gO+H3nFRlRCb3Iq4vRtFxpE7PUoUZ9cL4NB+1Wyz0n4eJ
qTVnpr1+FPvBSchYYwybnAYE/ZIr/SIY7OFW1kWB3IG2MGyyPZDs6FG0RZ92bW25mYPrxCLYd7P5
gEwScVcuULs8bxJD3Rik5cWMtaD1oUzxUO7bGiRC3i8sR/eXlAPNvPCVOAzVLTJi3pF+SfX2vWhP
J94qi0Ab5HXG7gVn6aKuvEMZmJiC2ivi7kXZYU7vI7k7FxzDJSbfEVWHZDjGk/bh3gE0sDwExKqv
XE0hX6NOdfecVgCiG6cow6hnPrwtdYtqnOkuDdoauXJIOLc4A1kNpSWQjnyCQVDBp6LvJoNf21aH
6iE/YpEaCLRzSXS2VIX/wN7B/878HcIgGvvi7LrdEt8NluyIzT4cLQg4Im/rtAE36mRkI1cS3b5f
dE6TumiqHs4Y3sdygGbngf4RP4ZshUskmVvSJaTCyndoyHEASQF3QwlutzsBzfpAOkbNb/CB3x+p
QMfjRHuYGVSj0J2mnQfRxIy7e6M8m51qyr6jM2YHnJrm9UMDXfhJkmvoJINSDODnXNNx4m4j3Oqh
gfl8iNrq5inPjiWCM+MN+EPQXEv8v63rUDg9KQf4OGNnE1IkAmjdcRcaEL8d30mViJnSPS+gHeo0
FvgXopeZ1yCGRF9JsxZtK6KC/5WuOuUclt1CZnx8sKvaJvpVazoPvSyFh5+T+NHeeVfNIgqRx0rw
fpDaI6dZTsUW+5j+UNuzzScEozYNtm9cBGGg/QLcVHCTIxj3djeQ6m9URrM39GY8K3//uGJuDGgR
iy3jZcQmcufrLfINh6cPsefMqaTdY0/DYovwMz62aewn203RCGupChj+feaCjO8sYNFBsJavsII4
HfjbvvtM/K4n/AoqFBglTAAMq5hhKEG6SHJsqwExSSX8hw3aL7+RjwbsC33sJ9/6M4L4vyIShIKO
Bsjj9vGzFF9nQRRY2da3b7gdtcQII+h6mdXq3ftQ/tVmjMv1T6+o0qs+U/GKnLhfQI2HM30tovcl
KM8VyDG/WgVC+x7/wq3VCoGzsJrQUfRh7sVboXRA7zpEBS0BUhN8+VTMPIk2hYBKyI4teN3KSDIh
12XpaB66dKfk8RXVggLUnIYV4fHBMo8x7s7KccAqisGmcD7Z7sEX7Mhl4F/atRQdKQUi5ewCVeZw
FwxSgk9eXIO40BkbSS9SGfEUxHifvIvPQ/GMPuLF4P9BzOEZmbvQsS19+TTuWr5QnTSr2/F42m2O
+PiX1VF+IWJlLW+9NGhuE9xt9rkkKmMF/0UG4mDx1442FWJibmcYYX2brJrX9HTnjfwuH888IQY+
sIV5TCzbqqMink2TNDaZR2qHklEjbAy74m6Bk7eIPzoYC9K4uc4DLuMI2RClpnhe7n0ugCongXJG
miKXf8ZJQ7+WX0w3tq7ROHrLIErqfpFWODAjY0cQqRhr8YQaNGEvcwSwLm+efyRzXg57v7Ni637i
HAGdP0WxJFUX5qHAGNUSjDXEsLMbwgEsIdLtAupbN6d0W+ElK9lOUDB+tDqFDMhVc5GaTAHqz7h8
IQHhMWqE4icPhfhc28/GRN9SEf2yFdbwV4IRmDeG1CyQl+BxobybhtDN/Cx2gxfAkAh2pnKCYgpt
YF66fH8+wdEVECiP3O5+fm+oe/O2HpZHi/+EvKVO7E6d/MoWvFlDbnqduiGHaGT9Kb1TPEqTjnTt
RcxqKNsk9xkqymnPMsd4dU4QIQTtvNamAM9ouXSUeFWWQKCJ4zGCnV007hMSAZUEVrlqP6tlICV7
V/4YKBnbZvWgbMuU2hOJdGdugy7c2o1pBZdnXkt4hYm7KykZqiv90xLsayoP2cU0gptqPrAU8l/j
hl7OcnG5rcXtpFYT6WHN+JUucKIX6B1LPSX+2CXILE0+e4ia/U1RCNxbUmmOQP68mz+GVIH91p+B
Uwq99LZsyWYUZc/HIplWMlYWxYAU9Rl8DOH/16yEfdzcsMzNZ2CpVC3WkuqmuDjbVQS5HZJYtjNL
WSrfUq3cHPTVB4xE9BrnbIiYHRpt84cuEZ9ZiPU1OCRpAFbOw/MSQe359qneMRPNsazrFkfXzkaR
AAEwjHJUFko/KY1tUlGdeTBNi6aROAXfCdPRFvRNdb5ae7WKr5yU/cOe6PW79pNgDLZsU0AxUijJ
mnKlQ2pja2VpFTUl40kx8u8F6p3kafhQe5iFkERR1oeBoro80nMP5YOi05CM/6a9PztpkGiuGj0Q
jqMeD2yVjHw6wxRrLuKj/o17hRfxkT1WbdbNEz3548JazbRsFmOmT8BSHlPDeqdERmD3uuXBeUkA
gaRxj5yBuvvLcjFzOcrzFSz9+ccUqfVH+CslUSytDcvAgvYXB2aGkvpVu5GEbjaW9gcz/naSm7qB
D5xaRUKwrCDRUuDj8jf4j4wQuevjkXJa3jp+9HpZNOnnQD/tQeFSCJDLhbgU3q6P+PFB5ibHmLr3
qmfMHMapXR8LT+Htqx2Q2AeYB6ExFkdk//F8XmLvjKWiakYagUElUEXOjp89FGCom9bThURKIsHA
rt6cGaw2u2NuNZyekFh36gpkVZBFjntvCdrUuRTUtNgq8g7rIaudOCtSIJLY2HIgXh9hs3ajpwkL
Pd/VDl/I4V13xrs9nQpobuwlr5elBAXeqJADEV7EIdBfqDOEK48p1D4yOQOZYCi3/D8+g42kk4Oo
ENTMevhUeSg0VzWTtkm7mU00KBvbxP1FUdBqkOaBjW5GmFR2DbUuYh3p70H0DNaRMILbb6QnXxLv
kZ1SiSVv9Ym1kXeIdIP1ZvWssEPny+hwBkBn8GXxEqmQ967oX+GH1Z6kKGQzFG8uR5+bpbiol92Q
pgjG8Y5+oQdNGl9/uL4UeIg2r2nS6tXD0NPq4fYT0Dd2SqvfriK5xoBBeudB1Vg/EtDOnYfOSTfn
anCklZevhvt8lt7I6+n1uObSBXMMeEjzriunpb64oIV/vs7qkTEjkfEf6REs5ItMRw/gfc430kWa
ydUZ3fL1QZDUImB9uFL0T8DsYczueh8S/Z17LPD6rpuDrFnAcx7UQKtjKDOW+gXpc8kIrt1bQll7
hpeXQmfl6STxIxER5yFp7jkwVTfgBrisoXAN2v8bjg/xyEyHEnJdIsnwLaxI4mH2xZHWYHLLWysZ
RM410rRQ/Yxu6HbsRm2KCa4dkA4kYikJhTYao3TgyF0fmb44hPTseVkjXEHq8o0a50JAQdrdshZX
YAW51PjbcpS4VQhNa8kRWY9iY6WL/r97Tjp+Vd5yrPFtKTom53MaFruJiMrOEkdHqRkKjTy4KbAm
BxE8tXeFyE2v0GBtSuQHD1Gb4s7kdOgK2idCvLw92j5l43bkPgxY5QvQ/5GnNQWYq4nSG04OC5Xt
MQGJoed+B+OR0uOeQEfbJUDXLodigO2aRkMNMYCGW4QCWg7nn/RQeMBHpQZZYiPifhaYop5N4PGZ
+q2LhyuMAJX12R0sOHljfMhWsKSt8Br9PO6WVx+bojn04PbMLs5REC0qQfCDL944Uiuq9rr6FRoO
3HCqdJprXhgEw6mjVzZlelYlKUs3DPYFk1Vp1O95m9RGvsuTL5ePJnGrAcNzSpAAHtJqK6XKzuwk
ZVvIQYElHBLY6DpqsL4BSafAmEtYNvNtOq3slwQj/e3I9iDWUeJ6pOWhPlOnZ6ckbpcsiAGVvWBN
bHtJNNfEz9HRzHVHTJlc0rAQUoGcFfrgDyaS26R3l8KkqzYPdpciyRPj5A44w4LYfqhsGV5xCzQa
wG5wylgAE278O78wcCLHtrqeu7ph0FiO4En4i6AKifGQ0bbIc/ShjKXASvUqHBETaRWaqFpTf7Ju
MBfZSfcHKAhlye3WCqT1AgMORfWrxd2/Do7efdGKQIk5QfG9IRwAvfAbVEwUdzOsBF3UQnmnM03B
L2wtiRsPg9Hy0sAAodnv+fa7Y68HagkxOjyKylx5eZSZG6AyxfK7gRwb4CKDMS4//Ai5HoqB6s4i
HPJZ4oWxyiebi/iDX5GwqAhJm2CLnr+a7dUAXyFsCMKjDJUJq5Jd3+o9e8vl7aHRU50PSq6ELj1s
2s2FeL/sxDSo0YFbVGWrXWmrlZwn9LRZ2P8FYEZWdtJwzWomlnCGfYXexJOJXPv9hmqJ87RXbVGc
ba4ipvsOxKWbyY0mSk/AAXoCzT+x/ugKHfSArUiSxCARI68c61cRB7WjtT1Bs4hDlhag4D5aJXzW
X/vT8yVKTQJDnzJYntoyHJGDCDlOmz6ZyQNH687XDerytv2s6I1/zQsAG+qziDbfxCCDgDda65BV
iG63/8CIp4O9YUmti4wc/SBC+m6bWKXBStHx3v3yOghgzQqvrik8xjkpablIEVHuq0XY9Y/pOT5P
nNWTDJe6b6+vCD82aEWvOxBzSFbMy5F2BUAB8ad+DVHk99KDI0JTVK24TtbkSD0WmdKpDHAnKKPV
khhYzFFfwrZ5dtFXIYz9nQRZ29jVx41G4Z7l7Sdl8JBBnk4keqSFqRrnIeaNUvQ77OEto0pSHQBD
KfqGROdtBt9LQoEyAbWgLhpqyu9CHEkyCzkmggI/BMFG00CUfzG0vBa7prJ/OmBvzIdPvaveOrl2
qlE1SFzZu1JyJxZTisTpeAhlNKaad0mc61k2f9h99ZrGycNYO3x5HsfXaQAC39MnGVNtLxks7dI/
JSpnBagmBxbmPbCIC47S6Fcc2oWK41VLz++u+p4REfLV6Scfk4SQ8FCl/iGPwbKxWTinbycR8rbR
O/U5z9a7LqJfHN8W4ixY17APmmumkNmxth1FHca1HvmFxX8HTr7SbHm+I9r9it/eX1doz0egKkU3
qkWZ8/53iyPXIhlVFfPxzOGK8SBp7bhMPFCcxaQURIJhnzg9ADpCxprEvvhTiEyJacukxzbQEB9j
zsF/F8vEgaBkyYrjPd8qg3rIvUeMq/1mTfM6D2WsZwk877i3NdfETW4pxNz60diSPkLuvt3xJhIc
squMM4OSSPpdpuGwxXhcFGBuvXMaRDvoYmx9lAu5LQ6Wef4v3XyMw3BRh/8OBo5pLGfKmC6xOeSV
y5WsaS/co54uDIMvQDDVFhcvZxAgEt2owIWJzN4uAbToOzw07ViIk6g1nEyyA6oZ8EAj2VDx8OYc
/Hc5KwCLsPT+NhOS6Oo7VyNdDiaDVYhArv915SZu7YtPYij3jGlgHuuiMw7pgldObNoqIh8Iu6wI
F9NIW/AYleqMQTQ16+3wRj15Z01xWNKQabhvPE5VuubVpnFMoa2lq9lO9YoczaGxnLglZisFhMll
jQO8dOsaz06GjLXPhEmGSHr90cf1+9ZWq7z0eTFUs3NCXe0JACQHihbLl7+4zQAK6i1CGbDEGZoq
T2vfEzGmBhHPeFmLKlzQtKjafNZe35KAxeydQz0AZyknUH0ygPSeJ94ConE71hh9e2Xnwc6hkjWJ
hfye9RBu/3zvVVZ/dfG6uOGkypzzElmALhq0OWGoBXrAPlDoWgIrr0Q7nAifQbmMl5QI2TodIUOM
X4uxpb0K+9j4JmyLTCWgNhRZo73QNAX8SHh8MqpOXUYee8cGSA+SaKppDwv3iBjsPnotGkAa+S6L
D7sqp8F2K/g532sA168Q26Sj6VM/TATs/PBeAtjh97+1iNYBJeBfLTC+e0KDaguwKpL9J/vjqSVn
TH9c+VQ8n5KIM9YHWIlfAkUgWcAd5jpfFsJd6a0+dDLIp4W36ghQmRn+lRFIOq4iTSyqm6fRZFeU
2Sizq/zDXHYZu6Rvks6mEqI18bXBurulBl8MJRlTP7DXqHKIAybHP4hnsM9R/LbRQuQbXgOqblno
idK0rNARczWI3d2bZ+8fbnaSiFG03554KkHEhYUVNP536S1RRpHaunDIrOazW6oXGlrQqIlLMkVV
LBU6bu6AqMYXmyAM6RPBiGhPqoStTKDeKTujvOSpnjN5GN3Y++fEu1fwzI3cwCdOxljRAIqVpEbG
15rhtAFOX3AgFsfgCCJShxQpZ+u+9GmAYlpO632Q6/t6f/sXCJG0oajQY/glu3mTKK+dU/j/Ojlv
I2IBL6YYdvKwebUqGCCreAWjQWwUnS/XqkBaZ/V1yQr0u8pger1rk7sFuRg5xncyL507iVifnArT
49byCVvx1TUKHkYyoEOOJGk/7DMJpLwfKAzKofpsIjMJgawZmvUxvitn2NQPaMPqzC31kgQe/nCh
L2IPLB2fig3+DK/1LFmf08MnUXgKxbEqpGoLNrELW8TozOeRFMyqZYuPRXStySffiyWov639I4O9
QBkR5NcF+EBKexHwn6WR+EGEsI7WMKqzbLHNdJv7rlJqRJ+VoSpWa6mGf8Iwji8nyG8XTzam5I5w
hLa/OX0YYy9MDpEeaIX3fehlYVG8Ujiw5iltrDrztdRML2A25JhkgJ720jltIq1sInOigwWe5rnA
BEQS5xOnb/tCpKnQwRmOQeqiul1iCd4qyYtNv2p35huY5hoTXvx9P7F22K70A+GATmMArg6TuvJX
L1cj5qMhXRmC8rruiarWFZBGWuMabizb2RaqhfG5KG4wTLqRvmZM+qSQr4V+kWDcfe1H6ovxyG3G
fabKZ58LRTbK8lEvndB/5n2KXUx0GmImq1Ef5ra84/PXjV+BZnvmgaiYs7X9ZW/RePYuOZCQj1r7
wcmcdIv8m6NpngKiJISo1R6yRaqO5ooGbGvU1MPfdWFVCssYdlk59fz89GjPLtL80lhQkjW8or/w
p9/9qxppvwViySq+dhisU9ST8WdG87UZ0G3UPuSmkyVUfvvnEQu9LdTQCdYGe+DaIi56xNLmEwtm
zYAXDrTtckNtbUYncwFa2jgCdpCjX6W5K266PAc/ESMNaGL5wQF/L2Rv/euqX1F7WivsURPmEhOt
djdsv95Z6DGzQhYbeBiAGfBa8pBFF6o6vuhlscFt7NCcK+E9dOMcpVXYdXcx5/oDTI4nQWGJtHou
RLgDsFg3M32u9U9AoGC6wI7ml1TW5mi2y5dHY18BIElsrsf6Qp9bdn7lR6yg0E4NzcnpA7wpgWjd
p/qaWZ8XCNUpPNLc/y+TldzLHu5R3bBp31ribYgfpzpEwkGmsgnOvXScBMPpNd3ERCkLzVRAySsd
pNe0Oo7V94glHkFiQpQbbW9knLbB/yMAetL3PgKJf4EeDu5hWTwft7UrnvMmsBdMusAHP9ny77WJ
ql9AHKqxh748lIk9BybFf7XQJLZEuriiXY0QLyXlS9EgriZU7KL3L4I2lkp/xlYlJT3ckcNM/byw
owH9w9CZYGObR5LgT9oIRo2Qb7ithNWvJMTyRbwFgeY8eVSRDc/6Wpd1/punbawxvYl2nFboGl6H
HY8vgWotDJdjyo53+r/T3PW7/NA+0wG/0B+sd1qhfPys+3JTbpcyrShobK5/mNha5M18AqMtckvC
5vTzGxzCA7eYtfsDmD/XAWCDoa3t5JetmpiIGkMcWbAvGg+3IyjW6/SeOveYtWLMKXWCZSmOcaLa
vby2FZeiSsE9ucL/jNgBw5tEty0Sa1LIPTpinARnn9DYmNd5gRAmmJEH+0ooScdFzTtmFYImCFX5
1i4RKrTvl7A7m97dNncpucM1h2FrkHBd/AN8YQncTtJBU9ZCtWxkThpH1yzbIhNqzgXwCZUdpS+j
c+IIDUHpx3PKaR4CqWL85S+Rh+E4HpQH7HkTTMjtF5KLh21Tr9V5D4Ru55DQnMskLNE+DIeB8yiq
iCMT0FqEnl65Ma4UwWzLkqguRypk9Z3yG6/HdViyaCeh5resDZW27Ip8a4ofUkc0LFYLg6teMiFH
P8gSUZu9qkEtdFlinZva2ncRwc6leWZKCxgOxAMGYQUFCw+xCKK78FnbQpaD1LdLwbpSo0dQ1wgE
WOo8F7dq6xW6YY3qdRyjDGZulSYOx/OhVsQQ2K2qf7408sfeMZ5rjApTQ86rjMtCSVFE6fx9uJh4
ByPWpdmw+twFOPbrY3IXcPIml3dVlDqbMtxEzgJaH4RIhfYktL9wDep2lrTrURcCN5KHsLttWewo
BH/kfEb0MdCp6++0mJQ4QaVl+V1VzHzyeQ/yidTOuA17af6WAEQaeGFdKG6112rCci73IaDH6aBh
AVWvGzWihUphl/1LCX7BUs/R/XlZr5N5BnXmv70KnrUxhZcRyAaD4LTqCRIKXv3meIKB6orhoVY+
IqFsKdCirtU29h4li3TLMgEENOEKvNG9x5VCrLlk3JHqwKT2RL64Korddn3iZ9AreVEQlDIWbvLW
/YR9R67jGbIWQfs8E53AwGS27IQr06uz6wn9XjY9h9vYJRKU7I7KUSZbuB6fGxjwIiSgmvU2TLnu
37cflwCmTV7Uu1MVq/hl6sHobI8LQUwf49I0bXcQqNCxoe2shtrYPuTgu59Fr7Iu40PxQXHm09P5
l34YH1yb9lbhur/ce1izscfZNYA1c6w3f7yFvzfH0CQPIWqIN6w96gCt+NvXrVNEHg+vvTFpeYos
Gha8Lv6tcqmOeQUEpbWV4E3ytLU9Zhrfvuw2g2AtYEalIvUpWq3oDO1kvPk85i9SJuewNnANB97B
Skvz1zEhFvxXvO1igBWBICGrZHU9EvKfDLKoXWaqjt01leKB08uObW/NSZoVlhk5F2/Uv+SIZSnQ
SoW0osEBcf5VIYAxadoI6fxqa8P+5ANNbPJcjhxV+II/R0eKLm10+lGK1w3l67cF4wCR3rAhuWK+
/ZpNZ/3J3kIs9jEREhEX4yAIJTdeg+ZZsgKGLhs5CGqPQuLZYgZFp6tJyOL29QSfIBZ1kcgO81l0
V8REbq8E5drNyE9GleENGIAxbPNwuVYHV4+dMVkJy4+l1nmWbnRK0kB/IGJSP4XRHgOmHeACuBdo
RLNjmekEkoA3vkR4mwwd1oNyX23jbjtJhTixbDocukwXV4XAtplEk3Kfi6ukx0MtRQ+789EO/yhT
OnKUIYEM1cLix59cUcB5zqCK3dkivnndhF0Jei8TxO9wy5HEGl1OcBtNcYVDKFUMXaNMz2Pz3okV
0xIf4EFuR73ay7n7MePEkb5cbj5nyEUBtkf/1FaXOZ69JETN7b0jlbWHpNoUBUy7Yy4P3EbAFaC/
lld6KYISUrB0LOpVSOZyEtxfn6UAODwk+yYQL3dqtGR/bVUDi+OjTMGqIk7yT1L/e91WHopBVthi
dS4EWCjWu5AxL8AwV3HERUr3fGl1WBvKpGi+dqCOSkutKpCOhLlwB719Al609u95DqJFN4xFQAAb
Vu6V1mnODfP0kFX47CePBCyZOaShrYF+No6t4JRdv80n583UM0ogNWKHshXAsfyk0UxlRw4Pv8A7
KJM1IM/QOgBSQw9FW1L3R5SHFPZCmcxNEv28/n807v4VAcY8Y4l4HG6ejgaepfEsXQ/McOVVmTaC
QTIug6aNBZZWHh9RJ3yMiB45SUeTyk43gVj1VpJUgXmzPqh9OhD+OazOa1QAc51Rt+5w4/UvNleS
7kpkM4JsI+Y5LP+/Z7l5h975LCXsfBXdIiGRj9p/SFjZOKwCeCWP4Wpzs1Ez+A+y2y7MFxu6i3oo
TmytqV7fW2hAhkuze6zeCtL0S0qXdo0WGmydW+PmxZAcv2RdeJCmYhnGB/oaKGKxpKHflFGlseyq
NuEVNDK+FYEWtFaujC6JwIcM2S2DP5oxMswj2o0hBRTJV90tjGeCijahr4tcEm70TPlVdPaJND1p
Ii7MHeZ8J5OP/P4a0HL5vTAgDHwRLrX6A0v8QuCaUu5DpGij15usWeM9DE0cNyzqe24xAuSsg/GC
nBMfr+kcW3fiHXyZ5LcdckMpD+Zn4BVWx0sZ5oYoNLwDuT+5FkJb5dsGTNele+65bYAz8EutM924
wpnbEWKtLFEITvUIB8AZ2RFynNjpyMR6fmPg7KJlIG1l4+YIXu1GyBKEjU7Igb6Lh+2Zgr1Kq0Qh
R5UFvM9DJQff054BJe1TyMBVQrM8t/jwmObVYmnfN4wxL2MoPSWq4F8Ij5f3g5I2ooJbr72azeh7
+hNcBTyz5PIaW+UVE2IBqPntSb5CMHO4eIxOvw+HMRvLmnAXllhFt2rbc73f41KcA7CRSqbHWnil
5na5TNa+xcl116NJEh78HAUMkMSaVZ+JUi8A7vdYo4pOZpgtLow6kfvh5ozE9eBksxwiUJokDhp0
pcacgJvwP0quioRXY32plUUDLMLW6PFd+fZCJdfeOYUDYXL9K/GmBVWRtpaU8CbSpn7hVy9Okt93
dwB0gjfDokom85D0lAZzcEUFrnBvlTc5Uou+/yVTlg03+fAkcnHEezWbEF+0/q0EQeNGyE7DsMX/
QQySkpwKA0lJe6DJiqQCcAdttUL+dZ4GC1I2cyEVWpSLcUeZqazkmV68vplAZqMjLFzdljMBNH+w
uta5bKKgJiJAVn0c6IB1gXrcD9jE9nww3aiba8FfzTJhKXPwTnoX88leqo+yQ9KQKtiix87JePqL
IEjituoOoX/WzTQ5bFzC1lduGwjjEEiFILiXtcOkJpvtIEuPrZlxLATIs9m1H5WctPVIdNzxVD/n
4el8mUpUefgZHRdZ0hrmikBDWU8ZArrbPxhmumtFyinrXl8p/bNaKNtX7PbyBF1BUhiz8D5lb884
/+B+aKp6lE6O1I8WWBA+S0E7+Ovy3ivkLvsyfQdInqKz0QS++ogEzwfF8eQF7eVyw4jEmwawhGps
K7n8+OsZ8WA0vR1W1A7mkjO+/r24qbLX+scFMgk1UdfF+uVPn0riUb4QfRanDKkYn87nAxyk9t+C
aX/C3n8LxoSRBQNVchi6IPQTEjhnxD//cF3V3bX3Hz32Z2d0vzK4VDxiomQjtTAhJF2RVdpbwR6G
jOrvYtN9VW14yMAjUOPLbwaKHH1nVgZMGdgs53SVE0hWlLjsEWrktN7/4ueRtcjmCrYTU85srSMK
aCVBydJhjwvMLsdUJXJdfF2UOXH8ZFvuJz8uBaoW0DtSwrzOF0h4qU6BcPK08cfA3/zKz+wQa/0y
QkTtpRIdURwifcXHSQeD9Vvk7EPgV4u5TxCbrPApiyMSgh3yb692A5ODnAwqcUa4LNLw0lTZsV9q
5EUf+609YrYamOVGBwVyG/5kefmHOkLg7opsq6H5gvqnoYqtqETAwBotjMjecKKsPSCf6VSyopTF
AgrXJISXd2Q94g1YJ1bYo/YrQ9jWdcFqRfaXaCOZ0icbWXX0NOc/pPdCZb1Hi6d9QUuIBFV7IyXY
sBqSI1Y8ZGAQpKX41sk2GpWoQtOvdJnXqrYhXPjWQX+XAOC1byseifUfIt3rU4MboFHqWvV4SGC6
Lfgxt6dKQBl0tyelF6bCsWfhx9jljP4exbAVW0+BdhVLGi17MRf9OsXEQbjN34aCePcYa17H8RJY
PjHR3/NMK5AftBBP5P0vq9WAgXuAoBs1oSuurCmyIr57VD9QPJsynKc143EXkbfzZFxJyd4/pXb2
WR1Tbx+WR9rB8omXhBppYlh8EuYzEyEPkqaibTQqgS+bR9oxCFXAEq7tA5Bn0et2xMXKwEl+/BDG
rLY76cOYBZsJ0BuUJC6hJPrPkrtJyATPKxAWoY1itCJDpLpej/DmKHD4L4zPBrpqVAZnF1mWZfKr
T8Uv3MVzFLQCuan4P64n9O8QBOPbJudshqVbiXc9EBYomZm9wINkfaRgcBdi/gD6CAhFlYq1q//c
M4gVb2p8LQcjBESbMQUafNQGexrHxs5WuBA9D6DJVApQeFzvE19Hpna0fVU76fNiEentxEBk7FdV
/d77rYHXMp1hdpAxwGvqE5o+Czx59qnviQbPbyCtc3iKGbheMPNtcsKxLZmALXRGoAORi61VDk+j
A8PJds33hwbJ8zBHHPhfS5CE/NfJ/t+fHrzc8lHuTRycyCpfgE/B+celWydG/3Asyt/F1aJex4Gk
IfzXOfnMV1wHsp8iAXpGDrwT4hlDhMMAmMFJHY4RhZw2UKbfunmYKhhVMI6g7kEwg6q5Z1Wm2568
n1At0ftgEgHylJBOEAtl0uabpMDJYwdxEsx5Uxrf//CeqzV4EsWqlzu6g5zlmbyY1xzHMs6LHROX
fqrs06WTDr3eUN8XEaPCyg6TRJJjy13SMmcDyuZr/d65XWbjh+q2iZb4qdqIJPHvQJ0LEcxSAzoG
MSRRQNtp7SDITNbBXr3J4JpXay0Q/V5vGjGN98yQOSGmlw2Ma0E8fyfYhiOgVjLbkTtE4o3Rry+h
8ZG+RjUh24L9bDYnaexYWDAgTtxiJaXzfAKRAVKTwicp7u6kLhNVdakFXPU4sGALL8WuUmbutylx
2/qDtSr4p5/xBPWVJDXUQrW2gtDa9b6JJAYD5byCyWrSC32hPhZzBNrPwlGVfVqb/5nbuIFur5zh
ERavsy6XlOhAS/uOm7ZRXMJuAw+7fp9mcp1g2hkINt/OcxFRvNvjAWRBIAG/AbSRItm9LwcYFOCX
58Fb/XT0CDVHAXP0zNvq37uYvpVJcLU5nmlaMgoqae4VJQQUbz+6ws33vjBwD1MnBl+MzT1RaSmv
xij4Ew7osPMabi6Yc1A94qiUC7uVW7onxiXX4eCGo6C4pmmVoZJDlfR3OIF5YQ+HZ53261oBvBeQ
wQJahFgBTXGv2siSE5x62UVheei0hsD1gkeu/nZhoOyrAG3a1wxQzb2z1IbQpJ4hIt7+S+KH42CY
8UZI7XW/f1tmkhlZlzg2xEq5jTCQAKBoenxKHYk//42cXYBVt48P2AIaVq6eTOh01WoQXIJ5u8Bp
qhIjCeQvmLzLe1wkuqb3ZaHiF6Ch1L9Nq3HpbMsmi+FUxS4sr+bJSe0RCYT0JkjbZkt61yWXS2bA
PzFcVM0HInHAiAmblTF7M3ieB69GZiq88ddXaqOeqmYJo0w36L0qP05lxB3Ky1RV/pUx/OAzWjWZ
iJFPrwZFGKIG1gLWuy/Uv2gMhmuFhNuvaG/YVpn+dLrU0NSSERQG+gU+BiA6Xg8sSLxYsLDsA+Sw
JWzta8CJAcB1pkeP7QjVu0TNIxeuUNnGf867kOCpRHuUosuLYHZZC7ZsvTipW4c+9vwXzu0NrOLS
rrVFwvVxXG5y2CIQB5pFhsvKR79eRwnH8zTLc9ZeD2kginb3uH8ygRaNhKh6qNbDC/brAuB5JUBq
Wdcw+eOOuiyZFD3Uu0aPCdIZmTGqoUR5roPh6HqdqvI/qlosjUqThr6tSkyhbDWkQJajx/wtRYbk
SjA58r/ALW2COvqyBB7RHvAv1mS0RsvdgSkgudKJXd1TcL7Ghg8zyJ1Fy/oGshz4S4WtVDOtGsGU
ozNUiA6KrUwU6Cs+0XF8Dtu/8I8wscdL9ZlvMgfuZDw4vQ/P2nk2jGqpRGG8PjbKQ7gQB/PK/cmv
IcUZEvEx4d83oGlIXWYJ9tp6Fj8G1sXpvVNsYsBXnUCtKfrz/qnwhZxgKpYkPJFEJHwlWPgQPnF5
XSXunKvO9TcrZ9NIT7v/+EgZllSeWn0Wq25ltYxzzPK9/ooDYpOL20Ts00Lgmft8qRNJXmbpa/ti
JhreJ5+itSQ6cEGEY0ciZmWh8ty7E69GOKu+qC5pzcmExHw8iFTw44EWFIpJ42BbU9mPKuzUnTJR
TVwEVxkHvZr3mOAsMx5YBVgxAkLOFQIHNH3n6gDxjzCB0F7sH3M8MISVZaKtx3kB1vG9HuBunHq7
IR/D7s4ODd1poz045wCT9yBCgC9tajNsSBgeNjBkhUH2kQjIGB0atIl/tb451Wq0j39ngaFDhlB9
Y8xbEJQyP3LJyZDPneFbFGNbmO7cSb2M3Uya7fvkLXW0rebdqERus5Di4+TG9FsGmN+G4JKn+CmF
VD+L7VWtNQ0UcICQklDbaqNs0cgBC3XO21/jYlD7Kd9CFZmdXhLUqdQlbNRFTTYDFEXlMAAJgCEB
yw7aKlWH3ZEpkmcgZpuuPMBUTm+DEkJMST3ALszlw9Gp4WdCTqU2DaijmxIb1Utc0RBYIay74mLM
IB3JQL2+f0SAIzQXyHwWmG8HKRevLDzxcV84PVUDB0NIYFceDf6rzFAotPI+ZJ0YLP4IwjxXFw6T
lmPjNDZ5dpGSWRNrUfV11Qn15LKbpQu3RMTTI/s57fDDXVgu1OpVe1fSlesq43QArL1QZbTYLMk9
pTByh9jNlP6FpopKIUO3rnLRF4W/QRax3im+7XI7lQ3zSw2/H8d//68xRyEV/e3/zv9PNFKkvFHk
/znTf2jxHnt3YkXmZLX43t3ao28Ifet/DXmYLU6F1/wmZyWyIdU4kjCP43zSOl1fvKDCKnoazICq
GTXwqidcM8kYhJEAkZ7GnGhuVA0hnnaZA9hvzzpB8KNcSnxV/Ajbq5Z8dq1AkjUHBBwXc0dHy8eS
yJ/sBgWiBkfHhhgWPKRThO9a2Voq8SyN3c8GLcsAofngHlQC+JepHiLwi1FvqdWaE+LEMS3X9o03
iJguU24bjo8YOWqBDPtC/5RRwm9fUl+k0GP6aqFEyx3zFY6Ykwz4H7mnjFy3SyZWfjrEpDmxgFz9
y/gzlN3dn8pOhRpW0V1a5ehHQEeWcoUGepVdTtBXu3mCs7T7K7MiyQ6supRwh8wVthHaKiG69S5p
13R3N9lltP9PWNcrbwHH7vxozqWBjqA/iki2ZcLp92eV/dSJ6c5aCmbpEz3xaWZGsTSTGprr6JIP
vGyeSxuFym7T+4HY7K2LHmVu3rnI4IkJvi/I1J8swwqWSeuKQUvUWXRmuUl5b9UFYDCST+pUeGlN
WmSQbHIHymgIwO9E1fQRUTuJzTjSYUkxWaU/peLv4Lyh6hF8b0Si7aUhc6CkdPP/BKdWFvRyAUC3
yyn2ss8HDWjikxvX4sMu6v9PxWqegZafnbvqUsCKoB0euLEbrAk3cg5ERj64isWbJYk12lzx2YSB
0RzHqOVUTcUi93ZP1eFPwSgxQX+pxXxQRe5AD9g21C5NrxVDhJNEN45uWE4rY016j8g5HsudNYt5
75bqzHH7kGhaqL6w++Psi4H7XFxpAid39Sow43LQ/oGtplTa9sBsJlQk0pDKBNKZpWKkkpfvI1Dv
AThg3KwBfuI71QtwumAaHorT6vZR1f3PhYp3hmJh6/40ki/6nAYlwDVN95ntlFwIfbRW7/BPCshq
vbGHoNVv15uyM2+G5fQCcXNNRGubPtJ8BlqBKiGHRLRQKstkEEl5v4mNKEWboqFerI3vOpiYb/wN
FLfavr3Td4+PFtGBYoHn7TajKN8TkOBZWLwYqjPc2hZg+RX5pSBW/CC3b+6Hv+CDf064l253zQcx
8xXTZwE6HJsfeBTwp2amHPCK5QNu6E4GiAkZlBcSP7ygBpRet3vJnCmbLr9x49zXY9g7WHhlMwZH
vAp+HuKRxi1E0KW9qdVnUsEpNtZ1uK0ViWrt9h9Sai/nxnVBnYHZEG6YadQrWc2vU/iSihaMFbdS
1qBObXzJJ9f3qxeCrRtOBL3ASs24iN8BRYhU72sZs6rCb6S/mzjljtuQQmwd5Q4jWHeZoyMnD0KQ
IHXdCZ1wr+tmcs3ukKgTjgGY8SRFvKF/7QXBHynxBjJJM3UXP6I5o46qxhzf4e48i14T4Wo3nmLt
dHJ3HwvjvyiSYd8Hclr+VIAaXiCgdGFQ/OdNtGcm43Zg2G6KWO+XKW5E0hx7CnPiAVygTPh0MtsO
UNL+7uTkJ5/DeYCxTkCov2NEyuSTc4+Q2/7azQ4OX8JeQfNmdjEhMRms0aiHyGYwY4K5AW36s9wP
SHMwO/1dqcixt75AoQvrl6Ds2fXgiUXEg2EOQcSMGKJ54uf2F47zDFdglYUZPjAFPYjS8TKbIuj4
fTcgxaIlyZU4sgoVYlB2jTlNrFEy+U9eTz2wLphpL7QcAk/dxZ1CR8lRM5SMIeADc3Kqnwru6sNk
zVHjYeKKpAIBr/tQ4hbeyhyCQBYcin4/RGySrm89Xn7T0c2ccK23YUZKAZNmjrqqHjvg6DQ68qtJ
tPW7LvKBvEUhiRlKQYQdpZVekFd1ujNDCXBhEsdSIfmhFtPP9AkdK8ZmK6VAeMLf+jqwiobMQvH5
RCH/zdAuCJUpXpI1aLM/szb9qg1tBTTBPp9CFmXiTehFjEE+BvuNjNuaNBKF7ejWohUEsmo9pcFf
S2v6Bt5Jatil6m9NFHVz88LjLfA+xqYbdzPZp0MzonV4BeJk2XBdPtM9CS79Y0e/J1eE8r6+E0tT
pe01CxRu4EIy4YJv9Mx3Y7EK7C08jsIjpASRipaVfdJW9pr0iwSQ6q0/C3zV2l2KqxereI/3CQo8
BCOMulUMOgB5/4qjsXcM6yHgN6eCHsUGTyRtfRIU1wOwkDlDU/vwmrflJZaxZ+vMYFz0i2D9VNLI
bm+klFPWULU3AmbLUxaqcCy2O1wMJiT7NtNjdiI0epYhwloFig30x6cxCEZjATqaLQC9oRFtbAu1
8c6/GJ724O20DNI1Wy2AXm2h4PDCXxWlHCKpnM3T99bgLcRMxKLZH++1EhSqwTvLZRasbQP5BN5L
dPFPxVaugnc5xETq+j7GXnqMBHrVnbMFkgfja1IWaZ/g469IZjOfMFwx6EtxueZ3JaPf9SOMZ5lf
8Oun3+vDJ2tAiqvif9fETnZNMROw6ZlA5z5ufbx6djl9bz4kKiD4ZSRAWK9uufVqTrlpLtFD2lkx
KVEAVzJal7OksC1/zzVlWizZqRynLPDTbcB1PxLEGvLbdHjnT5CW48z1vPatGkvVkzXytaADwxcM
56RCmkO5rm6zrx4l+HnDQpr81fQA54Kji6CR/7QP/Lr3VNGo68y4Q582sieNoHFM28xdIfKP4o28
FExxd5v7saXQUNr7LMvBSwTBf7EAWqLOAVfX1+de6yhMkDWOBnyQrBzglvApbocxw5FO9SNyIMTY
XceS8Vtig7GtQtQyZ1qBtEIqkjZS1lrdRTjS/i7sHD5lnKEDwJk/xcC1U9hNdMMSNFq4oIt1iOKK
UMlsCCBMzf8GXACs+OCW0LaT+RLxqspDbNx9W7fSpRbniD8mfJ+REjPCxTu942HDznjFw0kg+m01
pEVpiloQ6C36d5IbG4/41aeBltHtWdLxojSTKIK12r5w48UwQyd3ew8sLLybB0aV36pAzCutUzC0
y8qR/7h2H8RlrrPERfnrRh6FB4kaeLILtO8H+5kCk7pxoZEBEZ2FwOOQLHyDE9LF3sqtEvWiuBIn
JgvcX7bf6xN9YbHz+FhRzdLMUBuOMh11s9YQpBURJYhU4WjuQ2Jro9XS23o3NHlE9yBJMLd4CdNV
4jye3W9rULKNB3g50GFYyi2fMjdoGgQgtR21bU0BHrq7YoYnvaqKtoxvKoOcHyIO+uKgJQxyeSA5
2b6M2wvhKqcNdO9/wDeRFbNyf+a1G7nj8Wt3TVF0BLlciBn9/yiAQw3AtHIsG/zYhtgPJciCd9PN
9UTepgIlwabglSzg9Q4dPAil1D5jD0Oppj+F+VLEmR7p5986cDjILhhKbPtcpGpPoJhfzNrS8hJW
T5G8L6TJPc185QXlLv+BSZYbEWzQIpFRpSd76K0qKgyRmYFfeXYazYDHfdZkWYcGIMb+g9oNfvRN
xSDHdjee7B+i/U0jBFnNTyK84LatqnWi1Vt5n4w9m3ggCosu7i3q665GRHGP6z7hC6fL0ztSz/b0
3QpL9hfUIsI8iPjSriPmf3b1cUj9Z/wiVg3g8Q4QHS8He6YxhWFGAlY9mnMisPphpSt2RqGrigXh
3+9U3ORsn221vFJBx/yv4kYGo4+ocRMljM/XLnKcd/nSLsnsezVPloWEV6izmCjFd54kfHbxleQj
IqpAxdSBSrp43JPrMoJoqLol/pBusLkh5hZFpy5/aBusjR2daJ/jrkEe6c6unYQS27smjWp+I/uX
YTD3jBY9R95/+vB8BZIiQw2cUn/UBlh2XkBKU/oMqWXmT+mxQBiwI//J4giRmR9aJZo5M/mOna/J
cG0gPsbhJW8S2wkl0NyIdfnPm5vt6fge0lbLuioJce+k9Pr5nkOwmVDc59DzP+dEIsRB1oREs1HW
Z3YJN6LK4pY0z3GKe4x062/euL9aDO2A5cHzmCr+mC/2tMO8AUa0vXVq/r1wnoXhVes86RJ50KaI
hXvUUHBU9FKfE0CCziKTYFOmb+xh7iA2zoVAPG9w8pDCO3Ti9mVUXZzPmtcY12luFP0pibtM/8ZQ
O8CatDYxtOk22k79tUZmxbbgSc6NJksuTUoWt9hipxdHfAhZfcGUe9keohu2Brherus9wbUfrrCU
J++Atd+PkfD8x3SlJOTvH5WsHJh93OMlBBt/IRXAD/4FwlBd8JY67rhZhvLghs/E1Dz4OHzKg6YY
gXatp1MwZxLoewD1ptGgpIEx76uFPdkAJykxQQ/rKz7jwD3K8qbtfjqBFQiCBTnOeNIcyJSL9Ok0
hmg/oUndcAM/OySmrnYPgek3ja0NCIcZqMuGEvUey2eb8f57eFtV+tJDO8GNd7Lo1tvB6GhGoHsu
ffMvy9KoCyWFNu4csTj5s2m7in/GhIGOI6VI3inQWPYuP3X74az6LjL+bIbwuMbMu+Bdr3Tjmv1V
V2W3F7YMMDj4e8bfQmiXI3PLCjFIuulLHaIOntIJ5Zh1pKEl5S877dFKSiCj2eeSjXbecfK6Bvn/
UCnckIbpLUmnV/8dhwXOnJUrbwTih2ZTBz0KJYPTBrqukiO1qDRDb9OC927lMkOxSUp1ACB8fody
HZ3rk4LmuFovDp7SAmAW8X7ZkvjPIFzCdkBWhV4KyserM8AAgqJcqI2h8cV9OtpHKXKU3q5+gweF
yJiCaiDiNBcxLlR+8gzYQ6KZdoBFx5b+fI1dAij3EXy18GhEH9do8rWQdm7iJiTgDtOIentCayTB
RRYRVV1IulixfzPyf/2wcSEh1PoP18GtwuxSHPG+ziXKR50tIcZJeh+K+VMnfAD6jQvAWYVS7Czc
7YbIG807T3X7iBZhNtg/Uat5jVnmwqWmWcCCY0IoMFp1nOJHBEPlWItm5eYhpFJ0g9MQ1ouic+qB
uwbSVPtXlPHaCBTXaDl5r0ANF7MusYg5zaQ6ndgKcvQrC5AGWgovHwaUplaeNNy8BlYV8QpiaF/R
dXawksLeXNxWIsc4mmJleldaOS/RWxDka3AdXzdC5WsFW6Wym5VipitrSFhNIKmsFnIjOxCfb4Od
uOqtgeUO5N2C1e2H1dcsNtq2monxvLV6nmpMafh83AkP6nZzws+FucagZZDuYRjzO+wF6lW27SLm
2Sf+jOEhfOoutd4u+bMomoPnh53MhRzf00tPhfzzG5NiERq89GQvXZLJh06hXCde2uIEP20aggT+
lliC3Sr9H+TJTYhPWL+3qex/GUVB8KmC4kuy2IaiBB4jrb+ryGTOBZsbfWtMYqbFFiM3FebHuEMq
kcZUKnPqx7/4gCEnObpec+vt9H734fD+6RsP7BmMEiT6DYTjTS+hChHF96agJ+E4iJet3Jxgc7/U
TVw8h33Fz4Sif+eRQdPRKU2H3rF8o3NfbZ9MRTNWPnjnfRwjmNYD2UEASyCD5uP2svmp87TjaOhB
Uyv6PdonDnvxofnNdd+AHbdH0HMkiwQGbgLmFaEQ+C4n4/T06GTpy8psSPM0mLoyOK9M2Ru8Pbwq
+IgIPSSOuKyB5gx8+TsmDbqyD8trj5D8eIvmqoefiyqX2btVs2u6kyAB0rRhAfARF5z6P8b5qLOY
hTq6Pp3dgThWGUPjWHyw1J3vDmXjvtpyHsfgYmpc6g5IAJZfsnAY/FTnNKd/2ydf2HEXi+XOmTlI
4ybcP1Qj0M4J8CRPJK3iGo5jAdqiP0BTC+lLiGFK9Xw6poWWBpuvBEsjGGPd3B4V/o0IDyKuErWU
ZFCi7m79niWqX00oWBhG9ZwrSGKp8sKyG+Q624IA1mdNmkrgvPObp9/W74b4jILqVp2IbCzNRfrZ
zHOiLb1KJZfQ/b5CuwQGfomVtUoWiJwG0pVMI3lo7Pzwq2oADVQg2f7QDejye3WOWyvRpmPS18Gc
B5KRd1j2WBBFzW8qOqAtT7GiwgvBV2kdh/MANOUEZ/phINSImTJiQ7/klZIEechu1KYZAQKyGKy+
VuZebVdQhf36tLMqL8FmwUwAWLFrhWzFzhgQS2CEtMw1x5ztsrITZAgXcpK8420HjR89w9BUJ+HZ
WLOiH8CKSOHqTbEu0Jh6UzreaeFjposFSFCIsY0sLAL9nRFnt38iEOsNq2wmTmQyKWIKHRLnKRPH
UZKBb1i/0pyiuZI6Xb9pmdXOhL4e+i9m1vzSfRQjzrB5unzv0kvYtysOt4+AgNngb7e9oBj4erGj
d2i3Ro4x2cJFl+wZWNDLisobbkIyDHWMfDS1tT2S5oFRlMhvs7fh4rVmIYdEX2sXzC1rZrEhrXtn
IdkiH+A674e6Q/MA4wQkkqe2bvnq8Dzdh0MEoz5L5RBIRPGsvEvYdW/aQT3Vs0x/Lst2R0/+JoiE
f2OWCNVDajXbSdytgTbisa40FPji8DUsLnsbbZbb7xCa45VE3BXJSbut5Wynl1r3oZt+o35RMaDe
aS9aOtPml77/RvG72oogwXfhDL66r8vxLl1AXT7xd7Vw5F1f8ph5q9OmGoblJig9oXl8mn+52qqQ
E6KnEOAoXKkrsqxt0Lv6aANwltDyfl1OT2SvdN3Vy1+4Mldorf+yx72/kqjSEbsDPJKaVJiANXBN
++DHLKORI/qOsLyF2zbJ/jBX9Li1GmAyTC3P/+PUe5BiMDoz3l/EWF7qnhD5RqX0QroqZZPtXtH+
5CW6nDt0C8Eywa69tMKTGX6trnlmCKscrMorcdwbwOSyEObfoe0kLIUwtjojzHJzM0fE/R0/s1m2
UIC9VwcjPIlR5IdaU1znz6/qsSVIj997HAiKlSC6Ns5ef+t1pM9vug2TtfgWb5CZ9dT5HU4EIEOD
ygdTWBCH5KS3cdfMvzepn8MfyDuvDw90AbM37zbYRftB3CPJQ6IfBTxWERYxSb0g+gkRi81q01Jc
vBWVVGCmZoxAJBLLYpzxMB7lRBVUAmBdktj+4saMKnXWOeI7uEkJcrAaMinHqiX+4FVrrJZEW9TZ
i/3DCuLdLKVbf00di2Omsd+2RF4Bqu7HTqywcXXamg1fzYgdLNNteOhXcfspKt8iPnZ4h+xhx/8b
lUGuIVXNxjPvR4GGv1FhOU4eg0SXDe0BvRj0WXNqWJ5iWsgDzEz2KunzbtfLlpMHYP7s64nwOfQf
hSAB3nntBLiW+LR7xO6n3fpjedtErKlal0F+Eex/IakMKVy7SXHDOry8R6mWNlP/Ym1idIE42bxD
Vt6fsNtTRV2T105uYeNZnmAHKaNV2SJxeuQKJfinRfMYrXCKSeDxjcXUKFzH/AT4190LtvnX3B4v
xlLdB2jPOUPj/rXI/0Lhy16tReshF6rG/PWYZzMFkwIeKrbAm+25lPlYy3dIRyQAwZHZkU9e5THX
Pg6SlD+ltnCOF+STTIPSzV5lQa14nAP8deohE9fpsaJjTSl8Bv8+nB/VrPDZyZ6xdY7+qABdNu6Q
Owmu37/PuOHGiouYlSAt0eCps9RmONk96Boq6uJmk2Kb1ZmrYQVVdK/WglL2mAKxmhWma7gQKVur
i1S5llBVAqVThXZuVJysaWYFQ1aTvo8tRogbS3Ul7GxZMgLN3Ow76by3QdrlXk+1c4k5fMrGOR3i
FOOPSFEzEhHRHkd5se7wxYUQX8hwW4jOQL/lSj3B/iu0hUXoSawx58JUSgrra145/pAviymv2gBQ
hT0x7VdpYR4EEW8oAPu8j7waJM3cs7dGnpPaJszzjc5pJlXbQOJR2sPLP2hwQkZGzxLjtsxS0FWu
w+bvJF5tQ420wOuVzyMAdBSGhFrKuDgLNvobf1or21cAgwI/mRpJ94F73hCPyPNBKKfS4I9mbbuT
s7RWySVaI/lC26DINBZd80jj/9FlP7pKmMRcp+F2mooiLNtDXV5oUM7TjJWzKbJHv5sYn8uyYmmF
EqFZ6XzOVyJ1Jqg3uJA+i5e32ufR22Brjj1JDm+2Y1IQeKkaOvgWX+XSs9eMUkQaIBufTniJejwF
HuyI38lE3vBTh+lXuDsyHtcGrfPedL1NG66fK85sq4jRHJ1uRXep8HqRk3/GOlLZsGV6/An0xD4w
tc/Wt6PIllTSmeJeRFk/1Yw0Rv1Gyrw4uyqx1FP2/VRuv/NQm3lyHFztcpiTf+AGkwT9b8GbaSer
8Ql54dlG6D5g9lgNMf+wruxS8a2iNs2wZVzR9E47Z++AlAje1o3uOGWaVoUQHM3YAdIhPfUst5Ul
uqB9zVeD6WU4ngWcw2xFAD+g0do07WYcZ0SX0q+QX7fugp0s4Wa1SHqRkiATIuQZl3es6ZRoc6uT
o3f/3lI5kPs09YNnfinnZmFTNEbMU6zZniSwJnXPdlD/N6cePdTGHZ3wH1ts+DI1cAOFJaxQXohn
agNnfhiHdr08anEzmUp9mKBrizsJvYs0ci+X3Dz3sz/4Le4CpTDDuu9JEbsDvz+Sjm4wHsuhZVnO
hgFaQuN7bXUvT2PvKM+174bNv6MZpbA/PbVEIi/adM4nEjB/enrGiyC/qhtvfHa1PT4XsTcvIAvY
M+wB9KAxMiauqUb6TLabGT47OlmbX8evXfnYGTsmkHcCyFoOK7FrrxlqLrDg6j3uzE3s5Nd5hV+h
uQGwU0PHy4deRo+h5r+UDYG8wp9w7Wkxxh2GDRmVdskvuAIl11duWJ/JC3fqCGWXVfX2APKxQ0my
uyCn+tVDXc32MlLV+434UG1L7zK3uJ2K7rZZh0N7cyyEYd9uEpeAHDsHc3QKXuoXbo+28Wx6IjFa
9q8wv1XORIEJ5anD5xoAdr5e4nN3MSBnuvm+HinnPEZC34mujywt//fIWf0CFEPaeJTp1JNo+Ptf
3NyyxwGOoHnE1VFpcaRUw2GnzOFUoPqYM4Va4gU54C2Is8JjwPaG+RsygnLLIArIoF4EywB9o6/m
r6/c4XTB/IunJdRBD0+dGx38qKaszGpcfjKveERBuqEmQsGkH6OT7ALx7lF+m/+tnpL9m6n0XYGN
xBzuGpQHtezIp6kJTHYxcMkYu8ndIUW6jiAJtDpDYjKZjxo0aSoH9YuamtG9HdJU63nrIvOLWTC6
hE69cycemKHi6J1YgHB36qLgFZOpS0pAp9kcR2boa30caQoJsorlWx2d76R/BnIV/M5j7JQVVhEi
IMNpHMqB6zQH/QNPfvK1+6Z9m+wbJ4SSpqkCRV0pbvGYlmqHc/EzL2omZrGQGWV3voBJanygFj2J
hyhQo0IFdUEusb8rGWU8kKgRy+scrQ/o0atKPVDBxADaKjkglh+WqQK2piUQuqg+F6/4goVMKfgZ
F4zMRmGDduQRlIWai1jo1FGRaUp5IXn2xVJ43/HQfOgF0FuhHTLjdb2+EqMM49igdyWCr5nQU7z6
bqoxp5QJtjFnkvnhynMKH0TJawz9aOQ7K+TBCYRfhxG+fnGTLnvlDpNpy21c+570g/eUB+e0Hfc5
pOhMSgtg2ikv+cfLPawsX5ZojdKq1DT2kZoY/hCzbUsjdAufom4o4NOdG+N4qvJ74IZZ77yJVCzv
ZY3XhXvgLmJ0f8sb87GkoqX8sAXfyypSJPNuKnhQc28KbMeMOvhw1ttgQIFMAZlgrUky+mYVA+dL
mlc63nIqSo/SkfxRILveUiAyDk42B0pukHLkM3Uw2DIMiwKDYhqrRTZKvwN3pmofD1Bidx/CiG9O
icY5IgcLI/Ja3GXf2HT8w9+AndPr+Zbq6SKIQ4agWEXGBnGEfeg2b9dntd+h2aByheXfVsNgg2JB
PrJ0rOXZ7qNzfuhln5aplneFjbg3pCtk6n18L28lWGBKgEWvSdwzdhO3Pqxv7phIFxa8LrTeD22a
UhHgc8fuLCfHrZvF1cZtTIBnS0PrtwP4mZZ4ncuGQuzrdhCyibnZznCSJtUO5i+N3N09chKsNLni
afZKmgj6rotQnGxQs3OLhCmGt2bFw/MTBgLdPTPi2QvX1iSsnruxMoknXhNdoOkbsns93kXca/kt
SXfk6TUcd4Ji1Npa+bQcvbzVh7cangxqtmZtz+soHytJ6EyxcjPiOKwvqzZLWquhV5I0ZRYlgdH+
auj0KRCJYGSAdbVxObLxX2JLtjCKlPOGAA2pjlmILkAfyfjth6unIPlxIoec0d2dic32wh+0ODbZ
Ctsujf84JHBVdC82cqpQhtnUabzKlWTaFXKfeggqpNinj36MucEpH1HAg77JPyiVTNoLQg6kYH7t
OdRCWt/gT2nsf4fW7TK0HqiJx1HyR0w/jx1dtHKTIhSC468QyBVpa+xUF037OsCH9GJMzMGej9/2
kuQt+eQYqMs4zmigkEkct3qmGiuO/qn/41VODmUGo11oB+xFZ2M++8Fw4zPO1fQVAuR1HJ97dK1s
7RpAxKwCOI8ykKA/7vtSnrx4rtXXMD5/mFzudYV8O5CWtcx0rAhPzSDy3+ZY1jlsxITo1+1us8/z
g4fqthodq+y3K6almkraMy9xdRBZjLEoJlZGqUDQ3tD3fkNZpIZaVF0+pKB0WbkLeGQZUNUwGJAz
myDQh9u6nnH1pT1/PTei+dV83QxMzrNWCiZ3+1fyeHyuRt28sZy/DHP+JI3hLs+KR6sjE2VHCzSf
1g6rcCkDP8ZyuJ8aVtjxnaSl1kEyTHVDZqfMdyptGj5BtyB2883dpy21yWtXTqfmKIl/8DsZb2lK
MO8TS+POWwd+Melg3TvzkGnapuIYMvs+LydjXpqehsRZq1SPPm4YMXthcs8xB2KjeY0Io1nagagc
Biii0rRHzdB1YKlK+y9QhZZUKpQF9elMqh4eiltKrke02GN7Y3bNLp76Mcp1YqMaKSOBV8rfA+Dc
5YYIjdU4hmS2NcR22LUCyM9s1u5FWiadRSO+61v7dEsMwTZrBcnEcsajy2oZAl4KngNxHLYdZPxl
xD0t9YcNJAu2DF8/38SyivHNpPg3ilzmY9OaJ4rgh5Ju1n3icOJqk2WHyNVdWalnJkfxuMmdDcTo
z1IGoNgoR6BdpMLnKtEnhb0VGB3h4PELVmeNFxvlV+auQF089Otvk+oUp2qXznv7N5ezyMHnOkxh
E2I72PSoarj3PWoJug4zab82cdAdt52OiVkCZUvzabkaKh+3CGzOLmoFLW0gkVusTgysnad928Ey
UqdaFdxjAoo6A7Tkxpy0Ad1c5L2AuMQBMMuLupk4/DA73TTGt4YD+523fOmE1ETuuinWqkoCum05
zysvr8oykJHnqamMbcuZplND8W6UMjfnBk7P7h7nSGA9JVo/G8GPnnr54/QhPGtsLQsopwaHiVhH
eil/c9TiH4+cMhkIO1KdLFJdQnZbflFQn9B87x3RArKmo4MStvbUVFa71kqDlcQYaL7Opin9iFrY
IA0qIXKTbeptR+IjDdfvzHbfBSIhkAyRrmGETqZxnlEqFpfLg/jx4wT9XKajGS+5nHKvPlhTHDIh
9qg2M9hsa4fEa3lVwnh7u0c0SRIlOJXtmDd7Pd/M4DtlQKG1XwCExEpBjg1YhA0s+lAZ9YGaYgB9
sYaEf73WQFJwAdh64u8D2XgjLccKFlBBYeWrBqOjSJQalz12GaDbPKoRllDYfDiRQaSnT49KllUi
jdrlChwz1MVh33dKFdfiAw5bG1Bj7p5wuO0sjOZBuWjw7i4iTH7CpEtHimmyYwPj3lT3uONk/VVU
xCdVRpZtUBJy7UYzZCIQY64LGrzO5Mkni4wzqytCo33FXOS3hoKL+RxQ/tvQOFFLakBIGe6m2GIk
7ZVCsXuTga/FUrqLy9WYssKYn/Qghi+2jDpeiM3MpAM8WLRwczLbC8icSGbCuUr2ksFcnjbJVnho
mPdBOZEDfQ3lcCBpMVBCIBPlKAENEqwWILtpsCfeEz2vc7zcjwbLy1TFzMxP3SvmbxDh9nZMg/Qs
erNCYIWBSFpdfMy0Z3Q1SIdJYWMxeU8E1Rh041MG76DlBAEz96fxV4IuDKhhAMAjVnGTmGCydDUt
oteEZXU7vQYoCCyOixJluXbeCl4S1mAJbKDxJfmba6q+EuCsrisw5A9RgVymof5jCvFsC20TBa2I
CmEQrmRDRZYFjxMZaBBaV8BPBRl/ovDab8Os9K7+XlBwfGboSasDaBMQ6c2NC7NtoXIHqTiEH0YW
o+nNO4B1NcaapcTxtsQHIw+6ridNVfh0+8fEobr2gR5yZbi+ft+TxiLtB4AvpRKSIyjQLK10DNX0
rbejqccz+Y0ZzL2iWcOWifBcswGGf4aHqBx6+605lCopbJvMTdj+wu8U3Iws4KEIbARj3NIFtpop
ENGaHjM8x/f35YNARpObnnj1LJ8U5TUIpqCuFxnDb1Bsg7AwKr3ogXe3c0D7rCgQwG3dfo5ZEo8e
edYAUwedrHAgROLuqNTZOF5+jbjAM+4OHg5IALi3xTjKYpIzVHeMTeHcZHele5a0NfvXjFWeW1bW
PH7uKqbze77fxN9UNPEBe/JyyPuVUj7bCSeyiT48VvyQAQMamMAX7R1Z8wppF8+Ki0tW5jbwSzEO
jDPoB72BjlaJTbtfDPWg3EN9U9OAgZdwU7fTyOFUtRnEhLQmUMPrBdppuY0E9QWZlaD0yWaaxpvq
NQ0lRF72ftbfnH8CHtON4JEZhPkAgZHhDJxlXcOpKaBGl/0WXyfPKsCF5dtwwXXz71CHakVBeVZJ
RfHdKDlAdbIjACUm/mUGTp0sFQ4jR/ckZg8ysa+c9d+QNRj5WxdXwNab9F0/OETrJTbfc2SJzO1S
W/0e3ygCzeueodnwsSZE/Y1BSnTnXd0oI/IddcSX7TTeUPB9MaHPLmwZqqDeuFVtkG9BDzoZYvOR
hBA6ArpiDirFJXppdHFQWzvVwHRtoTE6X3TFk2gickFqVSD2Edk5oRGBdH9ee4EFvgmh4EErLLF5
g/dNMJogLoylTlK+FCQZ562ycP3jebpkehn7L2jpF6YswYf2NttiTtyaTPlmlDKZi1v5OqIR78xP
6lk4E78vOeYhEoNgxnlv3hAIbXY/dhONIlLPx5AGs+P4Jqh4/l88v8ACmsqxip7aZ9+vhPnFH7uS
pbOWCkyPQ0CXrQziQDM5pklL3cyyyZJFvbTP+0u+veaFBC4AO0wOM0vARvmyAurdLJcbK9tZvy7M
1z4tDrZHjacBPTocmhL4cJ0GoUfPjlmgw7M8uukcyrAA0P7zSsRV4a5+0OGhce2h7V7dGPaZc7M1
LZ6BWZIqM8lZPDf+sIo3k5YX7TW8t7fpLRNfabqagEjvHGL7LMx/PqAsdw0K93plCsnyblJmA0kL
uAhsvPonUdCQD29hBiW5RHuKArNQod9sH+Zf23qL3JeiX+X3ncfjq08cswRXKmTVTOEiwjrIIoC2
eRTlKzL92Afi9+Y670YiJh+3da9r4a7z0Km3RunnWckUSEsaWqqgq/KEdZ7ZejNmmu9lPCkd/gH5
jkMLNJY6jWfp7UyTWfuI2Lm6pf5HKxCEEEWlwtxJeogp6S4N0JOgaoMwct3zqjXHIwpmqpdpY82E
rGBsdZaJOv2PYKQhTA80mUbqG7QIQMmRgV2OEVq3l9GVk5V3vBeanLMbTzKdR7Kr/oX3aG0ZhWGE
+Ov2NedG8FzSuT58XPCWL3DmkfDkEXV7telzBi7s4gmIIVOio0+qRq/x4k0K4sJTFl8QidwK8Ib6
5m4QCmPR+ED0vt3PXIQohW9IsQ2KFVWzm/B3ySJgVGeP1/3dpTbWoHV9ZTx1HwjzMs2F97j6kxiy
QuURbu6H+Sxiv+Xa3cmPEsA3bLMS4JS1fdtPEXvnqv1gfrJy8rGfcJEgtxlM6k7PF9DXr4ljRnmc
Vi6ys7uVsKmgAwgxzUjO1SkHFUVfjUkyPXOJckjhfAlnfd2oV5HF8TwCZKXjLttn4ZZoJ8OYMRP7
r4olemugCZe9Woj71PY3m7FF/iHHvbvWao0A+EA0mdEOneQr8zlOfSHn3m5vRf6EeAe/3i1w8l0j
riEoVbb/bynw/D0+Lup7dQuC2WdwNdeQ5/RQkk5BWF+bf0MBZt9Y7TC+l9v9823k4GQ244QI05Sh
Hbuv/LiEUtM99UjPx9SXa5Dh4515HeUa7SaekgfGfiBrexN308L0tucpStt2KkCYFeTQylBe8RK7
P1PRdUuRXy2BfCEFn7WhjXCbAHOia1akxbsgW3WkA1PA6cWUG/aV5SUSsQuGmYTBKdyVd0v6Zdsq
LWyufTwXCp5BrGbhdoMkcHDTZQp6/dTkCEa12QkZKCdHv0zYhjVaBVNk2K4qYbkHfvpBIrAnNQ83
M7p5mF0MbWhF8h4if/LMsEz7DYC+T2QAgd2O3uijINJt8yvfG5FG8+Ps/kinOhtFypbKAcqBRM9D
JXuhiFgnG40mKAzBYHwclU/iTde5AdvNnVxYHyVEEj+WFgHLppMPaDTtEWvXerx3YhjzrcCba7hU
qH+0E6+mfXVtRoC/7paJIv8s+kvhmggO0Qszz7ckAddFMchYrGvZMVX7sIo/uJnq7Sr3FLfpRSOM
1xVLpILKCAl7W3ZO9R8IHji7O7TY9kWLPFFvR3flibFmhrom7txGIFD9xqb393ra7J9UD5Meckpc
bUbOvyn39CxdH5pNet8O6bZ4AE6cUwB+rzvwE2OfyfRQxZDIH4+dgCPZXJDsBElDDhykQHPpzLJl
EChxjhrO9Xb49x9k/qAOhQ42JCipegjJ5L5huUnR7Paj5leEigxVN27Bq0oyG4sGNt6edRMVu32L
4b4hRr3gR+Avr4ecJelZ/3w55bCDjntljn6rQFNu2ZOsaP0OtjxXHA7GNgTkqxAJ6XEw6HfjyVBk
GA8MVDfhW9lWYnX6kCaF9gYh9yVq7FPqCxXOVegODc3v+yTWwJqMLemq38hIpJstAJQiQFKrSMj1
9gru2sw/NzQtSjzQQn/m0/488gQvZTpcKAaiS06dBnRrRj7CpJuwLzN1cDKcIHIEdkkUMD/CIeyo
vRNEzT1/QVOD8MQyX+tQRCdvvoe+MsOSYRx/XlqKesIzuMjIhaTn6IHNJ4KOKZ9Hhsaa0WZ5lzBm
/1oUMzZKFtCMFw33BhkwsbiCI9mj71gwsTgK4NNdGvg13wK7ya3HWhRkagJknNX/34W9sJnHlryj
c8NiWJy1xNdiCgdwnx6p9TdZKHMkl3/zcYkG9xKuwZTgHx+qzjyIH04OP8D9niwNWNishQmexHDh
CxBqlVVUt7cIUOG1qx2GKC6Lrb0WGz1A4Db9z/UesvVlGVsW09zwNKe98UIg82HhYSapqPHMaAHm
3l5vNXzEvdQrJL/OGWo85NTswYeUbxR7Mgdm2dZwfwH+T4RjwDetzwRiN448XkXohahKK+jdCpYc
r3hb/USHMSZaI7r67xpm0yyf/u3OpI+PP/LTKFG9IXHQsMthH3eBSmvRgttyCwnFPmfyCnbyToOP
at5YRWWV9lqlraMRMDve27fHL5y7yRRiHiogSM5u9t6wITTHg2Z7Ptsj4yLu+8MTlB5RSsfLI714
5KWdqaUBhiAT/gepe4aIv0/gdgkR6OjL0cnrI+OziqmFwme5cC3VxTDf0KAX+d2QvkXkhB9NrR9W
xcTEjtINRL3joDOxm0SJcnXhvPjXHq0dLpvOygpHz59QEkOro6OcWFP8wlytcqXZeFHJ26qI5FTb
MhIFCW53Rd+MLIt//dq9I2/XHxYKlxNfe9MDkdSDfBdNK/4NTfQyOha5rVy2Eup0EIl8MVin0TGf
zj96w4RaiKVBNL228J1s22s9R0w7CSCfkqzuH0leZGPCMP5NpQbR5JPmnSIvw+16NKGDG5TW+i6F
Lu4UiIyUetaQAaw1J/n7cNEcOIfu4mJhq660CxxoJz8L7/UHSyzJCwtKH15kPOP0gOG4Egyi9xKY
cF/ZzLaXuVpZ3l0GsjmTBEjV8z0Lu6k77Y77EWJMRIH/8dc0qj1HtaRq+eyKKOM6GPAxAhWfrm7T
urS8ANCxKMxtILM7zyPnKjeD0BF7DGUCQgQzuIunzQdbo+QTJchnxI2cCX7aRsULSY1iikw8K9ms
kooRvKLfAinNljEaSSzdArA9Yn+ozM5D0nGWa7uvWG7S79Tydi4MFZHG4uaHYcMq+qbQVpbQ9cA6
Tz4RAzVr/MbPL3/uKH7XKU+skU5I08Bxp+ufQ3SIlQrUjq7ru700N5JhIACJqMvu1RleD7LNyhI8
Bag6PQHuQOeb1Kap1/gMLLjY4oWG1ZZfLW/MXqSKCQSnAi+YB0VvY+P+4zHiG4tbTMHOy8FDiyOs
WviVRTsF/qQLLH3+zJcKw3UDzLHP7eCmkINNbjghtWJ52NuqmYlQb3v8ero3I80F4QMTIHIgip82
qyrnqpgjCWjOgX/S+Lb5DVcx5CXhlklqeUEsKDWJAUGI86MEu92eyCEmt6FMBsvkQGNu38bkL69k
sB/Wo/ghvjF+dO3KCMCCTe0FLoig+Az5iWauPnUgVSofwOQQH6s3uFNdmdimHYGwBbD8ZuviLzFj
0/rdOkUl38kfudc0xrK+7TCH6y04VswXSWLdlIPhftxAAF3FGEQ+G3K/W8EnSkcb0Rk5P9wxJFvf
vkm6t9WKrpT3/YOidfR+nLyj9YeuiAGi0zGg0wKMwBWxFQVHCygm4XXZDLH2nLcZqJfv9/G6GRwt
Lmh+aDBS/fW2PfwWsvBZ198kZarrzirl4MJvEEP97vgwXfhcD1BwtNa1/01472EpjVdadB/YPhqd
QmOIUBQcxigjueZOnJ3RuXRVUVKw99jgPvjWLqytmH99my+AxqUSbw7jje3ucPxWqe19+nYFVqDO
ORsoh3G3ybqmQcIrCX/4zM/Go+k/tcHLF+ZEvjQvM4RW842HWYZixQqJbuq6+rCKne1kkRglEMqg
jxawAM6G17vXu2ZHUSlq7AYdSuZOwlEdEgQbGK3rAthZLj1lPH2EjdEUOo/7nkta7KYgg+trpGCB
laNuWJGbovECG0swQOv68vHiadk50vw1FwSQDsroH9GfRxhVpbQdmGXXFqHCdRi8xEpoCuSC9WL/
OJs0FDHo7ej7Q3+ofMD1rAWjWCVFAqsx5DMhcBKIGhsXt7FXKu77heiCJgf2KOflCQDCqScM5CwX
jPyaGqlG+9kgHErxW75L0w4k6kkUwlvUXI0Mfy/gfcGmCDuwyqiyMBd6Ia+HT96Fs0uVUn9YzEz2
pDSoC1l4q9B2ouRG9x/nlpKIojUVi6OzbAb1uIAlnUXsSSq9zy63boALrFWBItCwPEnKnSMod9hk
OshHDoBhMUxUkfpDsrS9oufrfSbmChL5j4LKgTlK9T0h/iANwVa8drETofydnxeiM+rFEAYMXEUO
TneguaT/KNiNIoDuDyEunzUjdR843/rpWh0y4+fLlmu+4YbgPRXkc4moPb4YLLjtJSFGfIB28Soo
gHAp5zcY/fsiRmyEx0gNCjIAqnytPeX3zZdkTPoATElETZRoFsY0+Ru6SHGsOwjfWQER+Oui+Foq
cYKuThvVppcSJQnwJvGWWdp9MeHSN5lBSW6mXiWcdaDfmyt0sd9RwZ+MAbdxgmYoLxKDh3Y/7Nx4
pt6pCc0ElFMuNj75jEolmFSSDFmTOskkit+oVYYXafUJiJOWLaI3MOrNDfd7Ed3vaSDZOwpYGxrK
nZ/bwhYJhcdM0mwf2aEVawguaMpiAjqqh8irmRTeLhK/rgZGnt/klQZzjZz/AJM77k95k6H+gv4+
mED8G7IzoL8ta36kzDVq1132WLX7vbyYnmVvbF5X/B2R9nOQidsaWqTsxfGyVmpe7SAyYIDhQTJb
AyxPu/oX1Bn0prgdo7JOH6Mlhb+g6gywE1eh4exiVOVMtwdDeRAXkKyJbArzVNMaz03/CBPnCSBw
kqPaxxmhx1rsnvFRr6gR+Ux13wKYcME5mmmF6bQHJ88r9dVdlHZE/oPTULTAMFNPjAxYhvnCglG0
SiQGRxD/WGh3pIqxC2pb/Lr+JtYGvF3QK1ev6IDLhdjMhI2rH/tp0NMaWlOCQmWQMCGoB3sFQzZM
FKOlXkYldMJz1ug4JHYF32SsQdY8nATXGhMVnUHfn8ba4av4gI+cskfwad7nkPl9SBZlfJhy4koa
mSM68yaxXVLOtmkTV4v2P0m+bUnasQKnNPa+wTbRwT8HDMQZLv2oek2XnFo8sRpZdgUlSlEbXgMX
0O+HdagGzja3QrFwBFL6JBuV8P3Fcosh9tYwSaHEki8mHoUO00z3NbGLffxzDrK55Zk3A43Z07q0
0DghJnPNvwH9NiK5rPsHoHELIrahxOwT0PfkWcVEcU0iSA/4zWZIx8aL2x2l+mNAYhAyiA2RskTk
GccCRwwAzihqe3rq5BB/Unn07S7mozO2ApAYV8lefztNwnYk+D0oZo1PQVTG3oWekYiFUC4n0RwP
BPoEdekovxq20IZ7yLC6suwe91itlWt3Bkz/vz63VbH7PqCqRU4E5aiA7Txta65szBcleNq4s7FO
aMB//R7TJlHv0hfacdsJAFOxW6Nk4Xs+d/D3REpsM0s8TaxMu4U/CYabAhFfop6pKwJst4VO2/Zz
AXowzGPnxdKOeaL3Dtg/6OkescMDSFqYkTdwJ6oYRfT8jpJXA+GVpazgJpNQImq9mEhPyi3Crm0d
M8UDOUGKsDGS3bEKPfYVLWrEKUZMH4+eQkL6bS24PGjfuLUoV0k5fd4QMMahnFjmVI+NlGB+ecOP
Iu5a9UrU17rm3vGq8SRY5uCSWMTm188455GiOSQRBR5xpPfk0S5SDKZ5EetkrLksKX0tX+trdEVn
liUQf3BIrK4bWIRqBH+K/g62HXv2mkeO+P7ugv8QNqzxHkJsvOcmrJ5JEb6Q3z4+AfIahLUEV4sA
5aIDho88qJLqd7Bc89o5D1+pnlJHtEEbAFC9cPnWm76A20AOxAPnrN7SrMLu3yZTsxsi1WnBBdjH
ymrwMqxXoSz6gJuJekpqmFQ8VXuG0pvq+7Dqq+lc/HwtgZVy1RDYGgrxxDxpqUFR0lavM1GqXRKH
sbsSLHxXTXVqprj/gpZl5RWyUiNkvnUF3hQ7kOkpwmPMDort+mYo/ZUf5yoZvWKRerHYQbHcpzCO
l1+mWc3wCr8FtPIji5bYxylPs6NoDeGiIl5FJz6+ifmhRawyfe4JdZQnitLb+BVKWNW5Wd1bJArt
oPbaYwOkVib98+ZdkD1ltyi73cYHgeEA+ql7tCPCpSqjOtAKSrY8lYKaQPmE5r+OjRvqViK6syQq
tcUvnFwu9Z/lfez+WXDylzdLv/zyfY2stL54xu/xSBbGPtGTUwr/cGNtmK7gYOTTFrl/I8A0vRF3
g3bweBxkmQEVbl9tOflN6tt0k3TTO8KigRre9XDGZjF7KZQvxvGy+rR1AuVMit2N7+6E7JbvDZUf
j6ZavN4jkDuWWQzVcxSzT4Fs5Skd9bQuLwK8Cp81WnXK3Nfa3U/yXcBApMtSzY6RQq610LmJ5caY
LkRibRsMW3NqmrfgTpdUtRNfEh7A/04nGmwuj1UE0kBAhuh2TQSTALjhlDudE6cm+0rPaPwQy9AI
4j+eZiMRj8wUTU7zwhwJ+Lvz0GyQWwI06/Y173bXAg5GNQH0RMVHYlxP1W6yGorVFi8m3wnfPQFd
pfHlWgVRHTkDOqnDmzFtFR3pN8sHMgZi7Wi0bGh+j7+YFVTRmGgU23RbudCE2SVAYN+azbxBiDof
RM4wni0136NAJqfrkeHd7DY4EVO3H+llTejQG+vS1pJerDGL1OePu9r+vj6yd/IVklz6W86DxcGG
9p69nM8NxLe/UgC59QkWOk7mERYHxYfnK8xdVUZwlzBviPO/51s1aHyraP8VLrLiLUlHudKxZiAw
OURGCpyTiLe/yat5W/dV4zGSigVB/BdDmVK7TybT0BT1myGvkDCLrWaeW7phiuq2Q7WX8yrdWjiS
spxPDgZV0o5UAuw65FY8vilCmyI3nZZYhUYQseq+hAVB2lEAgRC/jwAf2iibLfbNaldYIJLiMVU0
mwBUtjFlGXrcDF8u2BaXPVGiero/2V1Oc+7J0X83wQQSwDJVCfe7lz0/tFHmKXM0X9uv/cJuX04Q
jseysPMA3cRMj+V4JNPSGe0ws0ub8V12cc+oi9Fu2PrPSywUjk4sGPdBuEyCo4Sr7xuqzvhkUDzn
uzxsk+nBAsBYZIC+P38aeF/U2H6Nzui4HDhj3NwH54tg74C1ym724kFFIvZtclNHl/ZZtA5RNzUb
V2A42yGB9dcLvxpwpEKxvSgHfYgREmW7jT8e3K0SleJK3hu4QkHo9zIAOZ3TDJ/xHcqvl6O15RJl
gns0Tu/RGVIAJHJMmBwcgj/MMM1lPPo23CNOAk90VVz16cBuzjpiP7Grbhqn648hXWS757M0XBxw
1yCtR0YOERCoVdU4xhcfjViK5qep2WBx2U04Nz5zThDMvHPU8UngnQbBJkzrHmva3KdoBcWgD+Wq
KMH1JMcRCuj3UtYpW+gQMf6gnRStrfCfstP7yc9Rym9dvABuFDIgklljEWOuHE4p4yLYsJ1ext5o
mW5x72+yijz+B5E/FnlNyG85gkXYMb3un4Ihw1tu6zNUKOT9rUVE73UnuNIHWkrnSfQQiRyki3XA
oSIWSgnZ7RAnpepqZYvbqmBR+5JXKZXZwVss463eKdZ0+6i92TNd/M8fLREagOwxFAzzz7FfAW6O
2tod2aVbJYixEhxlDuhALqgF/rLuow6lIqI6QhqJJMHz+SdXsReOB9Xj+7NP0vJ7MijYZK9c0hNq
jUk9kytGto4Uq3CL4/tQ12yo9vHChQ31yAMvPojvMbrKvr249EAc0HtYyHYhGy9CCCtngCgCQkVl
FZaZVkwMeanheRtUyNTs0JBP4uqL4eialzcbOt+xigwkj+h1DyACr6ujc3Kc7wR3hZGI6m83L7Ea
+D2wHc8bq7q32wadBOFZODGhF58IpJXf3+BlCWIp3uzn6FiJtDOo24Hf5YJFo29xOK2AoB5LqDFc
wKVrzE52uWy8yUmGudBCgR3YPXtEo77gNKUAXDq/wLtDGFTUln1qdxEo8Klp/4JPUenuH9sqr20w
fNUmxniNQ14RtHySoE25RQFYYFUVDKhhh4FSOlmiOEqR55OH2ZyXuaS2C1018dWdoMEgbdBwBDQQ
q4krpB5N8jbK4hJEiecsg+qrELPH9s05O86N+j+HVQryNNPHORxb6jD2B6NGJS9nh64h7GwDm60w
6QCPeM5uXwr7d6eajOVUJmBks+e4dn2CcX9IzJgQzx8DKj/9oyHeYobU4lLszMSOjr1xopMHdC8D
6JzXHH/KzjVROybdgFHjjtspTadB77UUPAz0aPcnVApJadMmklT2ArOYULdB1SsYaHELA34CoZus
8BKb/Oami7Q/0KrUzkmOjI0jDXgsAtN3OBNwPYv+ibhVk6sHV9Z15KRNpQqG3EddOCsoU9YeZpSA
iHJKdZP54Z+6ynhKALEefRRwVAWXx//OETZ5hvQGWW1tlMIVkN7mTKN/gFYocM00X4UvxXIogZZt
IMjZd5EEDD269pFBQl2aSJGS8EwoFlyQJ+ssZfzkH5yDZwvHQyvv59bAPhFijTMrpf5SgUwcSvRC
G91WmkiOIntFtdbZtv3m0MFc0+QjnuL3XBvkwJh8JaraMguJf9QfPKTnp/YRQMgJOb2o9j04pz3l
Pg58oWoM5YC02ZSCt/K51q4Po9rQV/ya32goh009qnxHL22DqhIo9TpPwnC9EKsHUI/13CIQ/jX2
Jb8OgdbkiqtKHvE8qDZm9t7U5OzNC0eIcStayEuEICyar4hcBeVgFpGluoTWxb5yrxmkPBo1g3sz
yFWhmgxltpq6PSRf39+4OcUQhSKuYtcMevkf4s1qbaWUjqu6nKVsaseNzsyXzJHvMqJd2tzF4p3l
IxOCf0EUZdXW0gWydCJ0AbBT99sKcMcJjso043sAeNXOGnktj4BCkMrdYvdvfww4S32pO8GQCgqI
PZTWCpI6Vb4tR/AptB2XpcsYrEAClXFX+zWcna5NrkSxpkre4GAp0HMG/PEksPZziezEyKoVS7Vf
UU8iix9glNvtsC73PSekZL+Vc8vfB+yre88+Rg6uiCTDFsFEPuEPP/mNbsrSCbvVI/0b5HHhyLWz
Csg51VO6bhII4dFa7V6dp76mdfLqvsvs3OfmrKR+6aCvtFJe4AzZrdWbXlQvQFw4eLXRUm76xph7
87Raz5uXz54ykaDYtE4q3YnsZ8euAn0mxQAONm8e+/ubwmrL8KEwSAwjoU/tLNT4gUVe2aJ7UpKs
+JivVq5U2eaosJQyPStwufLsATz8K06s37p6DO12TBZVzXrob5TqH5e6tlC9bxEsW+J4g/vuKR1d
7V00uMnpDYbebR3QJeAAyaYQDxtm58OTZKWJBVl7BMuDjMHy7O+2UWzrL6+cBTufUVTka8Ibgliq
Jz1wVJIp1o/LCFzxP9gCf9d6z1skgNq8+syM9j4u0SQBEqeGI3lMpQfTBg9rI+4FvS8lNriiCr+O
5xJSf1gEymWrAWa5WlSzOlr5P1L+nxc1sJpeqJDpN24smWcPMGSEOLbzA8wC427Hzc6QIqnB5+Zs
5ckzZ4se8kUBrMrO9E12HBlOouAnspPbzyEp1hJyS2QXV/bKOmoOBlaYs58JcrW8fa7+D2FvueDs
PfjMfJBnQkIyc8Rz3dbm//TbkFv845E4rTkSDhddoJE7S5w+vlNpm3xmHn1Tp1OeX/wxEfMsoLuA
ziyGiTn5WYfL98S78faVLeciISdGwF3sJ/7xsWcc3s92gR+zCMVhdtx1dGbGkB2Bj5lsqXei0gp4
IVs7ssebSNXZg+vK+FfDBTXzsCBOn0T2DArYgxrgMImGjfW95z2xoAAGRJ54mJfdPvA1FBwfJvBW
OBl7pKBwOHAvkr+lkCnNyg4N0yHtkq6WLOdEuj+KarmhMZCEWGtIa4htv+vFcr16X76nd64eTDxs
j47Hh1kBobkCDjVSvg/G7WkjRWx9k5m93r8PlPevxnZ9DfCTE/7avuvCFJPxCKu5xcgbhjvyGbk7
PPnGcNZNnQXygt+s9GF9T6SgS6e/MD1fXbu8nsPG29dBK936yTnuUVB1Fz5zYc13R0ePqvHzZc7A
ebQgosFXmVaIK29ZvgQbiyqN9zRsuNbQN7pzLw9WfjKhNfKyg+98mrT1AoDdVAXO54e8MedWW89t
zrh4v+cc1DQqFZhyUELChTWEPI+USZjlw1R5x5basMftpQ0xsgdY9TH31wrGyL9AuJIBiMiVUYeL
K5Nnzc1oD9uWl/oPSaKGW17LTaOaz2L7yAYg70GlOmmFEi/nOiAjxBJ0EzNOuC2wD/1+h8C8RAsG
6+nd+63jSGRVJPp3weg7OkaOQCedK37HGRmEnfhgK5+CHjbmVwcBEF+Fvf9++XbWvijHp3fJIQPT
bKHpZpAg25djiZD/iROW3DuKBe0fdUbyrAkaseZDOnbWxdQT59o40Il0B8DiEDLKITlyD8MhwxOv
3QbkwUHl6bjWAm8BN5/Bsv837TRu1+ZrYhYyMRKs346LraF4wYFt8hlcJXjLCmB9PpdxKBqaMJCH
XF2zTdVnc45vYq4rthd1RdfrGA6AQHZr4eeV0RxLJbzSQ2iyqJasfSt/n8O67rQl3RBevzOCtpGv
1zRZrMDtrosF+wGjdQyz0MPLeAS67/NCLqXkJYecpid+axTZEgd6pV+fORqSS2CxfyQp0DqTn45i
0VD/kcQFpKDehQSPzyLWeQrKvsf1JoilsECRByumRKOSgdYM9s+hPIohcZHd5BiDMJJsWOq2dnju
tKrSuepZfKBDCm/4/w3Ik+bMqkbQv5Dw+oYNHaAYVUeiZ82TiNnad+Buw3Uip54Rh34U/jHMU674
A2EyRMVEVx3A//grhvGicl4OL4Sl/sOA1AH45n9XwOX2BT/MCmj7PTAvsXUtHTnqzuUAX4MHpCCT
zbcCpfyRrd8XaXBfXURYRY80qHf/n5U5xhUBAbm9BrSvE6Br+z9RJj/cVaD6Od/8R769fkiurVMZ
2AbP6Fp2aBILMrDCGLlNDnblyA86EEotwgm2MjG7pjA7gGdLElQhy5GlHOWiZXhHh7sjNQoCDudT
93KaNYtq9ATA7vl95YyXyBULkI6mrwnGTfULg9xa0/TGtF5k1SQdVIB0ElQGijgQE/sqtbm6KPjg
kJYigrRb8JsdlMaSL9vt0Ikj+4E/RRqgOk1HMI7DGGBE0ORZQonXqVzBNBczMiT9kAKxZCKdj6za
o3ShqJw6JPMEHXncbWV+d3oH5LuF+gNybCFRpm4m645SlpDzr7qYuhcv4sQSTTPnKnMopD3gBMlz
uV63L8or4ohNWSg3KDhWWFv8EP32nxA7XAyR8OjK91/H6ZCgRCXnhyXo6hF17uJ+hiR96GVw/qg8
MbcjB0iBmuKFziPEyRHBnGQCLVGE2g6XmE6gBqBHzpr6MEWnvkwa3mfk5BQ6NwdsPK/vyE05M/E3
LjxfPVHWKTA8heUYBlhEBJ+cUzTjqvdvi6K/Nz0ISTCdEbxlWHnWbXA6X5Mj/vuClz417epavdxU
fMm5v11sROg6aRJQUlM6kmP1JZr6+Ag1+9odLv9uTa8o/Za6WBDGraExQg48tdQpczw3Ehappk6G
hbN+KA/V8w6nIu3ZTtBqcRZHEzE0IZBoRNhd9btwE81tO3bdOki/PybATZeoKVXeL77ZoW9vp5te
z0n+S6bG2vud6dEtuXSb8OoUn0aKTg+wDTsbvC23mV1PqdB3hKyvgTz16aJoHhA50obQ9W9Gzi5z
Gye01VY1GfcpDQ7dM2okdLUElVahl6LvEB6UHGayUoi7yLVWo56pD62cJ6uz2EvgJ8o0+rMK02zA
+Dav2rwmqCAskTIkBzOyUe0UEFjWzAVVab+LOGcKQV3geRxe9fLBhGk0Ad7Zr6Yorpg6b8bsS7AD
O3l+8WWnvVKA917u9/p5Y4QbJldKglTqLiOGRLmmXpTrKkQjzGplpeRT2aWR4hLr2FGapwstKSCK
c5kvSsfSUIwVO6Kvdcj25Ge5ErsRGJ4L7AzJ8wFVoSVhbDaXc7tHe0VaxNsBUgamWBlafU8YrzIN
PZzEv4BtyiEtMiCCWU1L67ZbJ441MuzMXOdyqJwlEjNrFVk/BU/siEYkMPsOdjz+DKcnTlxxEyw2
KWNQolfdPhtCQz3YfTFJUhgs3S2NyONfCeV7bCBi3fed1rSuy1d+dLqjiY7cHDMrs1Xcb8Ujy+YD
WIpnnSO0Jh9OUIcXaq2/fpM3ZWOAMPRlWhQCOqTzvO5qOXtvvVFQpMp8oM4tlOdanKxcWVfeNju/
OTCBfdZzyWTYyi5H1mzGe8ENIQ2d+/FHUyEBue69sfitiCH0pnXDmCoe9IoHMvMlimtPqetR7sjz
vi93Zqvq0zBupw5ScVdKKgWtrjEgU3+JVBcMOl43QGt4eIZMkKES+gee69P0yLDOHOjG5hanbcWn
hGDDjK4gy+LNtiO4R0eE84qIQzbB6xf5m+Kor7aJpXGK72BGer48BRA5NhA16DwTrElG+6aTV4W0
OaNDBMzl9ynPJxGZiKVXQUAHPmIJQ1rcZ7E4BMZapyMfyFNcZ1zVFzByrVjCgR0GXQyKIs/BVMgi
SVS/yd9CHmpi6VvKfK9umq1clIcQY3oh844w5rvpEoP0tkCt49G8e98KIQ0kaTnTXMLy4FW/aUhJ
48s/TLuLQNxzuSSBw+gnmS8zzt/SHkEH4o8/ooKwsX/gV0YMStXrxsIwVXptRC9J4Gits3fkjg8A
/ft9UKBaaQDIttifqdoiMxVqQyANJAa0m5GzAdcuB7pt9jsj+ZHec5iaIbecFt5HuznFxnKjmTln
3PFQbO+65uPzQK8yFanW5UVZoO2BlQZyT8Rut+yuLQTblEmN6074L7KfSTzlIobIlBCAmIuJlBQ3
6/gKYkcyAg4ImhH591yf3hmT2JyMcQjbyaIe36hAcB9+b7HXhllQYiYZdQGXxuQWefM1Y8cN1eEj
Yln9nAgalxNaQSCnmr6Ga+T3tpMvxJKeHk6cMqnEDHngnhhaDZ1ioSBqivW02uFE9PjdrASs5NYr
miUuwKGKsgBVF1aCuELiq8JljPYCTfdB5TyQ5erXIqWD00oSEy5Akjk8/DH+f7OMLrLa3KuvTotJ
/No/Oi8X12gBlCkfOgmQP1OTgA9YiCTnc4DSH8N48H4pS1OrOhRuxwk6CpXg36vN3e3RE5StYYrY
2UunQM8dtSVG+PgbfGWx5WyO4JoIPRrVCRsxHr9r09BjjRBTnxazl1J9vdfxj2MW9LkQbIW1JKYU
5gpc+2vD+t4TV5wOl1xp7acy7JICJgn5nHDHIqlGPf/V53IwUHB+Q6zMm9NZqR11hE+rPCmB0iH0
dUB0FbTT3bIy+xqOcI/FiAg3/u5+Mztm/w4h3CLFRLRDVYVyMSHu8heHPtXbuVqBlavgBuLaAIKt
A8lqwIwojKlF9cdEDFnBOyeX34vG0Ru1eqjebvgmYyiQy34fXqOTkHVsktYLQbAlAm270bsjDgEu
nzlPjJsQz9RhCCadxu7wmE5PJANgYAm48CVchHAgxDMP1xZSeMj7YEuB6fp1fDBD8LzxvBH0jH6E
FatxpBYDJEeTdUw+mnurTflWw0/oDl/yMJ4qE17/m6oMuEz6qk+NftixaZoSLMoX+95zQ1YrMm4y
G5qKos0ZlnDCEYpS2jFbqmd48wYhqpAzwBvbeJsLT1gu/NThLnCGSm2FRdOBPYi4GWVp99zYYcwg
PmwKquxJZE3OExlDBYJtZPYCMonQlrAhDU5uh8wPkAlxJGv9/LVdGqnOr5ONwbcTf0Rn2tdWCQzx
TG/4G282GnO7pEmrccH8qa2kNWhakpRGKDNmQkxdchqOh0m52/B4zF8d6+tpr8wU7Bprw9rvOOxA
XFm2TI7pxRnIFFlfZ3dBu/NimTarbvTGwWaENTKXJUJTPSaob180q67cVyxN6lGk/sQm7wdVpFoQ
UhZ3MiKBbNMUMgQq1U4Uz1CMHdD6X9gkOyM1Q3sIaV1/BQYLqhbI9eoJW9CQisRBF3HuYEZMAc8N
wQ0AnMBTTPVsaO84T3JI7+DBInRPChOoUZR1t7B3O327NKbPi/ZOrLBcz/2BVHpo432//WCxcizp
9U9+uGWaqXHKm4ZNhcZQZtxGuof3hk2MTUHN1uqeFnnpjAFPdaqyyHYu++dlhOG2UFPqA5Ug0AaP
cPfH6Tyd2kDwsUPvSOpOsryErgrG678HVsRZNKTk6pxpVgI91FOp/89E9ofawrLezs/fh3pfg1yb
eTdbTcWJmVvujcjZaPAtkOdagj+WmKMIXlUmRaP4hhtT4a8y0Er8HtcUw0FMNEQDvTY1aBNen/xr
3os7XYoeqs9zRU+9xHByO14f3mzJ18i3mIWibXCUEglgQxP3c66iq/v+uzthSuDMk1S6PYIx1/f+
VlCQlJazTmALb/wn81kEcciIPnQwcq26uaHg7MzHB1cl7DsjnqVQoa6MasH2eXZzxAHKgJwGc0YH
UgOzM6uRZ5v8KHU+HD4Z08iIm9T3432UeJ8ueqX8+imy5XseqZFFfOaRE+wOw2EL8StcyyFfs6dJ
J5HxmttEsIXd57Us2D4o4q3KqGJp8yDHQM31L8atS+atg4JXoYEZvhkRJFSLd+dII63c1yWZzdJM
HUYTi5sOjkvCHo1p73h93BZjKRPN431scV7gkQ6fPC/eRa/zzHKh/N1yyarzHthHpPOaCFEZ8fAj
u0odlmcRfj2E0cRDQVxZURaoETRVDpsiIishhmo7/ir2XyFo7JmqGSm/k/mk7gtQmeL5ttA7Dr+E
MLnLXK81goKp3b3B/qKHIkBHN7TnnWJDw2BZMx9MrN/XLhkF5MzMd6F5L9cKxBC3YiHLFyEZhUbG
LsBu4GjjeXILMEz+hZObV+kEDmlia91PpnyKnBnFm5jO9cVlJjMMRF9KheQTS/fOipyFrg97HU+p
iLnfPkfRUqSGgHB/J277J6H3uv3JEZk6qdgeY14iwfNi+LwXHm0l2wDvHb/RoBvCwboUS9R+xxQ5
Osdbu9eqEq333wHqPMyRXpitl6+fM/J6VBvBQW5D53qL82+KwgC97oKIwsgGc6Ac9SCMGIdYvik9
06d3H1LLfrtfpi3Wah+S3a9aYf6q/bxISBSJZTNCNOv46Plle/rB1igbLVTl2HrZ2qfiMylPTcbd
P6DufRWKU5Ygu4lrx+lWqr2KC/gTtYUoPHrLeOmPay61ty56s8NPVJWp2lDdolc2z+CbqTjy2rGY
6w9BiE83hXW7qNX//dF7iQ/DiHx/uJG/umrKbm85dLb19ohh/S2cdP9L5fmLAcmzxWtt7YvGQBMA
yuub2DP2MLmfR/ROBxE0TFYlSz/l//Wjw67oV8sTZeddrmhEC2eVC7yWr/zoDphBXEJSY6ojTncq
ylKS5kZAyTTInC6oSlfiXEilV5ql04f2+DGO/TBpon2218UgcP3/Gvu44TEnDGNs20Mtg5E3pumX
NfKy0W+h0v7azOLsvBiDky2KmSUZxcE2DJxUyNGiP31PslvSpbY8gGbt1VcO30zR7fxG7PuIeRxR
wqS9+VqRTGjHMLEroCdETr46ERzCECWh3rqHhrrWqw04AgaGa9D/4D+tFkbnlrsD9BwCehxB+k2c
hIijqR+yTEd7ADvlfitP5KvXMl3GNOHAp16+xdogW6gI2ZNivyXqFc7Flr6jM+X02C/CKfBGAwS+
fkA1s09tyHuDiG71r16tMPl3NOp7LhqUFcHJqHp2ZcLjtJYnyr1Kx48nOdriDciyOqwfC2I0XAhP
ObAzCEf/c2WHDt3EiZhAaCNWDo+ulaa/keToRuWmqwlPAV1/75osFUrBK9uw3+W4TgGa0YfawooP
4EDCBhU7/NmXa74IjQSl5yORdNDBvEhmuwen5X/zN4vlOaVnA4rMm75fkPKpscmoNO+K1nqVMGXF
MVtPx1rrJrMgUIyi35VmGQLVIwpZQAAEBK99+pT9kZ8M6cYz5Jyf6wHZMnytkomdpEEWXpMmHuaE
jTFE4GBC53C2iDlFP+AQL/48dlKAD0qd68heia6UP83eusvxOFNME7pyDfPqEhJa0AWHKfk4Gj4v
NeEef8ENiCzqG6QwvfAyKt9rvhYtve96svqXKA7n37VipceYMZjEAHR3uLA2yvSnB5aT9dpzVto3
HDVsS8WaTKUqAb4X7W7fYkxrhcGlNGDDYZk183ANEOB1yWH1HuSVD7mgEcjWrmwcePlCkbbZ6hFk
FpSOlOqk0DFSEPZ7e3i+wGY5Hr7cJtpuKMllpHbGzuK2ltaKDUV7h327OWLe2z73vFxiJJ1Tm0mR
7VPTxAyGZxbGhFsCmOXNhDLn2HrsOs+5O5SzNjLkjAZAUtQe3bOgSO4VUISsG3igWbFW0adAVo+z
JV1sHQ7qMhFJvL64T0I57bLprdYlir3hdV/8qtg9O7/vMSBgQmtg8H2yuRLSm1XqDejeQMewkcuX
XOnz/w+pcgI2HtNcKRrcMl4pIIFhnitH9x37TTqPeG674pHqHuahE7a/ize8s5PpeI9IGlLRuPKE
P5JTtzPZJptfpw2RG07O+sIMAhA6PSIWQ9eju/TChoaU8ojwfbDDmp2wj7Wk3JCepvsHkdd8k9Uq
EDg2qCLkY+zMYmm8xJ1q5yTPRV3V49xwBwuPy5NfponIIYnZLIji8Ff43qbZ282zYWACQdwD+sU4
H3boxKiQ7Bzlx/GfVuyIKNNrtPqDKlf8dZe/u7mFwtMNlcjdl6klL644mxso1FPze9+7TPW2HfVI
B/I+6BqWcmbv80WONVrArRQGRzngDclIuj4mtxauzcaKnewc6C6EhTENcKGoxTkJUQaAjeNAiwL+
RcW21D6yg3sZKtNCQf1Tvr7rWK+AHAaP6XSKMhRX1WrHeAVg42EqPOFHd7XFoTrXODoLbee3UrLK
uUKmoIDrOEY4deULl3/y7z4Om8TvFtF9L8yhhjiTpnbOTNG2hrvX7ZKR/PFQZlhDFboXVlBkmf57
+tY8zXldyUEpVvDCD4qxAPfyeP3sB3g2PfjnMeBCbyj915zkWxhh36aFeWOX1lf/JTdw6M/1YfeQ
vOdd84Sr7b3c23xF/THS6ThjKCOErmJZ5oElWRiFhDriOHZ4SvKpIayLZeO408V2vIwwH2fLBxV+
W45/jhKKvp1j+CggDjUS2u97hV2PwVq6Jsa1rBewb4Cdik1a6Xeo6yBPTiq1YlYwaj7d53RUX4l6
pGFn5BxwjWgD9YmAUuTv1xDErATGz5lI8+y6hvpK4zJK2UwPWfampf8A1j6xYgJ265OYoiH/uTUF
IK8Qz6jnY6EbJw8YmCGDONXjY30WIK/NAsOGovak978Pl7ASLZ1CMLuLd4hm6UghT4s61y78wIPT
NdBuwGnW79JkeGtRXWW6P8kqVOUvBRyO1i/K3eNyehjS297PkQQVnd8HMG33BqkoMUgQhEljNcRK
MG5lTfxzO91LUOW/479VOLwnSfXrEXARGh+u0u1uE1ewt8/lujYpEQGnzAtOqxIdSFXkeEGEmZys
TEqzDqTh+kwHNYRj6flM+KhQlfERcs86HqvGF1/2rGSAuHiD41Vtr1dc48Dyp8EVpYI0GxeBfR0k
lv4HlriSmG8zT7exx0gNbx1cXM7RFyxQO7P6VB18mzpGsDcV+k8zTTxejbu3ahOMoJWtQXzmpo5y
0hUMe/BktGssAXRruNarROUphqS49D7+IwypuupiVZxDeDPsT4NGBHxiIfz/XW3HKzbU81PUMN42
j/MBul5opu5sVhG7KivnMP/5Ix640+uPXEasUQEw9TmMdfW/OOrBakQpn/elP2BU+PYKia86qoo/
68GSXwuwaQK77+XipwSA0ZgNHrw7/ZAs4BLFKMn1r2nrtU+BpUvI92K/o6zRrl5HoqbujYnSg3dM
8kfg+PGEezjGjyeGaGnK+GVBMUgdxdkgbMwk4lmuOAzRBsXcUL631fhaOzyREyJgeVDgEmiiRcMz
UTHwi+PwdAyQkJksQ+XeTCFM7/p9jNOdDa5mtcLjKljKLMCijruA/phdAXmKWenHYGgYSf1iNlGA
OEQlBz6eQBfDkmGIqzbUW8pZO49w2ITjUmrjJcXpSqjQnDKEEaBHVa7hZBVQoQEF2Pzpqf/XzVRG
s0Vd/taEbVSy/JsevQTgr4q2ZRniBpjOtz7qelWD+hEGq/SO+w0ZvyRinuT3ak4isqY/OMsO45eJ
YsPOVBZ0Sk7l2EGuI6y4go9DiOaG+ukrE9fIqxjrkiTLZcjt1CyHmNYwIdGxPYcDOkd3Lim615wU
gjs19hXuERRo2P7uh+FPtN6BBo9bKi7fV9HOdbhW93ibz9zkS6MrDp0nrlrK5JncmyS99KVOefmg
b+tPFX58aQ98KSC/wx9DlVSZ7mWCDJSQae0Z8pxZiAYdiJZR2anj88ypDG0vnSpWs/rCmHQ7wT3S
lT//W5CSk59me4RO4wHpQ+UQtAgDY4U8y4jAWBnU/LFCrC84i2n9rGr7E+xzu55tZuKGir3zEKap
DSK9wVJq5Cdiq61GL+8PHZtNQQgAKKgh8MDNyjtjCmKyBpz9+/uhBXVqG0/ALSzelmQcsiAE1bhQ
BLMcgtMINzW/yBEac0c6DvWnKgFxrPG2hIe3a5bcm/036vGAnMdkYrSfYX4o5w41g6Q0+anvjWJQ
TKvYFJYXheXgbUQnrt4zvaA+8cWit88N+Y/ZUPL0Q47MpLAjEMbJCb2OzCiU9KQ5VJO8Xq1xWPr9
cM/sohSGCzGwNP012STtJQJ7VZzIppq2DWLwTVxN0VnFcZ9z3iWve+lukrMANd++Qj/YHj9PWwrF
uYpzV54XXtVPuLGCNkwBrIPEThNOEutTb4TrL4JBaqV+jRGcQG4UumR+NBVn8AaQ/bzesogXKH9s
8UFr+38lbZPCafQ+zo/JxMO3tV0zIt6Dg9yTwrJOk77qJIiTy2j+GO7+7cjjMNGJZv+OR+Wje2Cp
9ox/Orp0moSyJI84Qtbzhqi3C7qdIh866KLZDF8b6angXDZ2mTXrXioALXrJO+Et02PM+FirzvFI
LopyFNYvhP62+zNU9LrGyN9+5SH6aAbIIRJY3CK3UXJCfJhvSDzIiuCFHU2DLStJ/QAigrwmkG+l
GywZgJrD1PDy1/SK/d27zXaJYdOCm9SwrwNekQMSiG+8O6PT9iwe/vrb3s4e9OCJ5FM4pi0InoEk
TA77hTI+zdbJ2sEC2TKqVsn5quMemXcNQirLBVmDexs0/eQSGEkdxXR2IvCUiaTsyWthyKRTDwZp
lKPk3Wf1l1AihwpMWSHx+9apWtkDviwXUMp58GBsNCnMW7aek96ArnPb9dTqNBjCLqp6sEFrWhnY
resT9VXPTCFcyR2CcixxlIeVLBj4zK1G079hOlN1EGJdxYQe+CtbjlYrO7I1cdOSvURN61HtUVvk
CyLzga1of4p9kN223AvKF5iVIcw2sq/n+/gzoUbx9rGAsGdkCau58Kv1aNbH4AYItAGozaeXkLMd
QSdf2ecNbx3kiHD9px0wOBiSD+Tp1nvzHGTZOrb8TYGdpacKPww2v3X9/5zLNcIxjWcr1q7vu/Ec
XU0Y8KT7tS9pKgtMYZfcLzRc5nbg3qxSqjC/IiHrds1FCrDl/dWHWRnPSKX8i8GcLNpO1DvAvfFm
xsHowiig3JvcqZ8InDgUS2/moFYN4GkL0jp3pIfyCtoECEjzhvuSWcQzcIqLxfPvozyNLRdhWGMu
lifEQFirvSH6Ltsq/AN9OQaAON/gNfFkpPBoaPCCMmlLXhjWBSVxeKaY9zfcBp/zNqCLLHjC4QJk
3WT/No9cklYgMD2TMZWhTRbSTAJyiim99USwQzrnpIYR/AIdNfYcArSX3PqGRYg/KI5HNqTd+LWj
TjxtEz1ER+P5WepK4poB677U+E1xD5RUjtDNwlmXjL8FzF9VrqO37zDWl679dMTgbAEQhkAE/Zqa
aWQmW4Gqa62lNZ1eLOHWrs3SZk6mRn8N++qem58YyGJLNI/BQYRh65lV1JnxU4dzHw4KTQKK86gq
FO45H+2hSXArWthxg7J1vdoWqzib14nLrBXy6KSDKi8TtQAEXbX6yta9oiOy+YWhInReNhFRYKTC
aPr4iwdNKwNihpjUgqwqc5otUoqIhd9lUn3zezwNSa+0cweGM9s/pA3+qqJejgHGBKfbyx5odi0T
yA6wMjRXyH2n7A5Vb3WTpKZuNNKwUJYM0t52qDq/44WaFZB4L7B4U94aXwGrReJrATNYrrSOFgDf
jfIWtl7cDYQkg5R6cKxgtEhZFbJ2lZGBCyj3QBz48CfJP/t8K8qvjv7zh37wqVB/8CshembzZw5j
hlKbhDxrzLPTvuw1Zmxb4k7wdA5D6fNmTdRTEKy9AWWa2ymPjujuJmh7ij+6OhlYfXZYFVFwimYn
UGjuiil0QDPDRduV7mQ6+2ZBbeGuGEvxOA2H16y9NgVoV5i8JBYdrXC/pAmbUi8w2TJD6KUPN/1t
P/G0zgsLq/BdgjkcyktTGE1JgzRbEX7uKXwREjWqvRy/QnzCBCn7m0Y4p6bui4r7yuycBJaae8cV
hlMqPr8NfKKzH3NhK4JrgUYedOnhew1Rn3nZCTzcW1nObWN1B2KTSAM8pXHowqsoWteVSAm/o3om
bma5XG/lK8ICYS2dG/ZGFSoXE2FSX4cKbT2DIYn8qQmjP1fMSA0B5HQxIppOTp9+1MDbo+Xms+R+
d0mKFMkXLWiP8Xyqa5u1xWYqWfOM2KFwHPPL4zzfzvfyZcvoZKBAb6kkDfEHjuLjM5zC1KLUccU+
RNb486tMyUGn1oiiWxn1+iyBT4U2qm6SAepPTtjuaey/t4SHdAm30aSgwVTQwJlIVFONUY5lkPTZ
s6muScieDIF6lA38puugSQxyrrXeefyGRcrl39qzx/T8jfKeOGUSKt1MCRWQfNCqpcbl53lU/X2h
N4170V9RkrVqCWbfmNPsQ2KqSlZQuKl1Ta3zwypWagHr7lIcMOeNEwVuxMTpd9Ff8ihTxSmaSbUs
rnfZHNIEQxgVnY4b4Q65UmE1IDJHbUdWViUe+Wh8Ne48ZNdibQL1EqnkcqrdUH1ykT7Hzf8ubxSz
bJRmcrFkbS9jSP/Oi+Kjfi7kUAc02ly01V5ku6k4oXnT0a6v3B+spLhoflt5UNwKrgq0h0iqmViC
aCoaVm74LyWGydiu/X+htv7U4Jaz8atqpWOHHNAaFUiZMGTqkEDZTTrJdeRIRm2ztrqWO1s+CIiE
URINYvoeYi2BPd5dPKmMRT+74brUrIoqP2XZrKL0iu2ozm/dqRJe3a0C7AbbNs/aAcpzqKdHYe5/
u2fbNXuXMH0fDKa8pqopoXaa62+B/yk5uTAU41Ow34C7EyFdCH2dGjg56mu2mp1KgYJOn2T4rBz0
ZRR5uQBK/Q4efG9klIoYWJKY1EwDEqzmvygOMFhF9eIJdIhG7/dIx5qe5wcJBu9Ov8vIoXkgNmgU
OKXn38CXyU0g0yd9Z0ER0HorS3qbdQ95i+tsvLVqzZ1eyfb0vUaFUDTFw8CnniWSJQh4/nZbFOuV
v7W0Dh48LdeP3za3UNto2s0uAlFm2iZ6CWrlISvOLcQ8dZY5krenLQZuTna9gxp0B0FxtnOhMOX3
c+HXSLz+qAgIC9khpBORFmky3sfItnvTCcCYuiUzo2+H4oos4cUt33XKS3ceUnx2dtuz61F8IlCi
WT2IRzn+YMwtsyMhvT6MIEzy2ALSOWO6Qh504Kq3zuDDdcFIkIgv2vaNAkwLq3bIiEUKfo2ZACeZ
CpNjzWxMLflOtfBgkAkNWjMBZQkQesoVkKgFB9PVyNp328zH/kWcATsPoC56ltEdecXUkvcA+N3l
3iIAx/BY1NKdKympE+llNbkXKOvNNIxSPSrZd271xSL2XK97o6k/DSBwx24vR+hCkOhnKgRt8bT3
8rvhEI2rwbeJAS6tZgiGy2i/BXACli+NtGHK+HL4vPo9FEdO81cXN58UpFJJ3sBQqYZWHkA/0nay
XV+d1cx4J9Ie6KYvnvIdzVSveSQygyhrcL/hzo6/AerH3p3Pz+g8+MwbeEX6pEROdxNH1Kyex/rN
XhCZKFBwpc8Q36aySvI73pCiGyGg4BscRT/P9nUEsP4wdlD1gNSX0DhblMcwP+K9yS/IIeVvzmXA
HCWb8C4V2n7caN1eNufmUR9GtECeq3Y35YH27wFIbzLH9uSwzYjgzr+yvRCZGx0hY7MiUmH67OEj
tvpkNVxFVLOcrbxUpu09CqIFdEvaNDAES+OieqTS22YE4h07iG47Tq1/PMV9H2kfZR/EH00Gpqvt
eC1uOKlg6Zg8pjDDReqR3SCypsA52/YORtQVwXnF4Axfq3eDx3Xy3nswORTSoqMhfRCrfJ+E4FNo
KpC6iiOkd24yfV2E8xVko940ZansiWrcN4Hzh4mOy+qTtj+uAXiAX6r72exMhzO/arMnjhZJh0lW
HO0BSKHdLVfHgZVt5z+Kl23TtXOpGWjwbiWe0Fz0haXjy48SjcmDwQQ+HZYHhjQE27aToLmgwwdf
WW35KGwgF0Q2iyE/ZP5ItnL5b7717W3K0Uhc8TtA2K6A4K6f55AlLP/w3Slh6WKfVP/3uoxrfETq
fOmuJ3JY+VPQOxW4uYP596jq9d7MOBOz3/PIzifvhbbKlRUZEEVQBeudhY9+vxeyAUmajzdg2AbK
3dwfXgNdON4LHBHbQOraBEOnufh/FXi7qbMAIhXfFE9z5o75xBEeTPs5xqX1LIM8Flh7DXJv1rfc
stVpe8VTI/1L9uz4nCSQAU9GFXg+uS0bhe1v3vIYvXNK1EciEtNHUTOf59EvMRsWxonZpcqv4dps
q4dBknNdwQVk8o+FTLonHLTJIVia9DZnO4FinD+B/Ct/omnEvCCvizNeQNu6BSAHByCEegctKJpl
2oRHWO4b/LO/rcUGuVt1fnpBBnFGWrM4q9kYDMd7fB5qJRWyvzZXK5y8cSpfMwp8qyh0IL5HZNiu
ROfVGCj+IhAAJ4qw/9t5nIvaN90spAupby/z0WhkB8+eow8E+wjsOF0KdkH9GgO0zKMej3l4/XIr
L34kewN1d8ziE0UHPv27WibRdCYVOKfFwlJT1ZLr432fbVowGZEUIcma/OodP+u9Gjo0xLplPPAK
/iIaWJj7rvibZ9cdg+N58/uoZE+T42cKBMuvzKyqxxa53VDxK9kmLvRLwoL9xxhtEdpjuzO45MW2
85PtzZOXoIBisR5M1FA3wyKNx10AniQJCMhRnmvmD/bVtFQCzI+qJl46bbZVU/7aE1qNVCrI2cCG
aIyQyqBI/y7m2wU/gU7L4XzLws6ThHAEKV/XoBkxB2cztbfmD5dSFm4nGC1WVmKlEP2pKJbRrVLf
ZhQ8LH+lKz4W9tvcf0mIMQbhAbYRpv3naEgCwKkiMBvdUByFcUWo90LNJzhdI6n2e31LHjsgauvg
DoaQKyyAcPemOfdXis3HtqD7iUAr5rAlzRlpLyHJnNdEEMmWWJHisMHK60eKDWJ4y7/ucJVlRCWX
WA0FYrV98mAnouJo3+HxVFm8c+1/lgts77rFQD9XBXUZbAAajIyldWDIjuFzJMl/99mpIR+X1qcA
smjuFtbrfDfYrOZW4e+qwx3CSVhy4qN7nnwUzMH+Z3Jez5DktyS5T5gZ/ZR0UXVSAHoOv1ttkl0L
/yL99ayykxAXK3ovF4ro6jUQj2q4/Ym1Z6Orm7E+wLQeKEXcDT7cefKzIPHVWzv+ZdHEWlfuFvzg
F1071Sql3lwYaqcTEPKWnUJgc7PnJFAUQKX2dPyG2/ZAmAYBqYOuANbpEoYg5QQZxS+4n7yC/v/7
ruDlYuv11TtvIP4LfqcdwXk8ev5CLMIC7Eqm/zyEKA638geYu9varcCC2C0wqgO5oQSpS9p9DLDC
G5bAaBsLbbcQEhmbtu4AF1BABjD4IaTn9emm5xxGx/XJ1WvSuVHtXhMjugKcPU5oe78O0Jw/56HP
PnZxLoOU9R9DodJ+I4DJC1CQFuy0u4VPKWNpWkMQSeK8rc9wRo0SdEWgJMtBYaI6Cc9qQX26fBj/
q89itAJFv95NR6LEGMMvYe8cOejfiIIg2rTytOUK7kDoQUh9fMNnAOxG6pyUw9Q9wg9TwBCmcnW3
uaQh3FaTXWHCBU0XGP7zltZpDacJnvJVC20ieyByN5cOomOjHh7l1CbvoEDqy/5UadX4NiFn4WcF
771uFLMbrUACbttbeImbfhl2RLA/rz0E8VtX8Rp94bbWaCIdNIq16Mzv1R9RmBiXap0AnoluH62W
WXlJMIJvsU+p682zDaq07SnlymFNGzavZyqA4vQOjGbDkUv34jLNYczyifsP8u9DWy/OOGXDsrfK
Xow6OxSWyic1V0nSFOLz9ayusstYJAPsMBzgr8xmwJSi5qDFvekf39Sl7UtP2ZV43YdFoeibnSCW
DKc5Qko8TEI7vafQZ9Worl9RdiiRi0YrBj7N6g9UxWM9nrByWYW+MuW0WtQEnjiYLTg2Ja3RzrU1
YqMypJ7L6xBB9s4VE7CWc8BGDLSLOirIblWvN9yw2qGEm6AXpSPPRC+kt6OzYCZxJI7ZvuwQUG4J
h9xONbdW3BbfOBUSJf21M2N4Mvh/tKqGyXYN8UCKdfUrZZ5edBBIBAQQPRvvB00UHp8vIhthjiw8
5owwWw+0+mbONaD5lp4QTC961hR8kcDmQVFk0p94F6KhvQhqWRaRqq6YMFMoGGVaFr+U3HVRNXMW
TuaX9FXptdT+q4CYlMRPD4h9uyocoDmvSlfR8pJaAihvYR/ozbKETDRcZxvOLOWXxjN+7ySjMVNo
7IRd8Err4np+3S30p1rxvdYhGgTmt1Wi3twaG1li9tg6kpDIctwtw+Rk04oLliGbfPz+Ce1UYRXc
Ka9l5lMfmQh8Jb1IjPOE2YZ/H0CDXXi/JeT8qFVA7/TYtZB04A7+crFVMsnRQrUOf24ajEa/3FKY
munRedL37HDrQtFWwmVzJOfVycb9F+UiR2S78nBCbzDv/xjmAW9ffud7UFaQOyGH7MliIdMjx1P3
r3I0DnmHR8Wf2aACeO8M6jyO5h63Abt2Xog0hNXfhUodh88l9IkdvNDF4qIWcwa+jCV2eOPXMbPb
CQtgzPlahbqcJpfyBdfqMqo+ZX6/J6tKWp78eSNsbLwVOIMhXS1O98bk9Gvbd70y8S84YGlt6mfd
77ChW5MNOF/7gxCIuynHOjfsU5BnPikJm65vwP6XYfsKREtNrHiZqfdPlgWOws2ckdniFroDyUh4
zKb6b0xCMfCyQLY40i/her/gWSDYVrirYII0uTM6u11OCIz1qwMxuNUYlsC8oprPDcG79G4fyIU0
Ofy0lR3bwQeKLOKb69LJ6X0ljl6UndRz785zmzTohmj/xKwQRlsMej5KGpd+UpgvM16iEZIEWD0r
FyuwE3Eqlj+VNGRGgzbKe9C5CoTpfUpElXGNv3vYKRm/gH8a557MRpXZkpvd4/KWoTPdb8fFqQ5e
4fRNiZIGlpu9n3G0grcdVnxnS6vpJpL48J9xCnMLBvyk8dNGdtvi5/f4G6G2OnMBxv+/QCY/u7Si
7IUcnQ6UtoGrO3As1C4a1zfp82un/CrApdr4JT5c7NfgbjaFJRoo7YDRvOtsQE7bq8eiZ0bJq1rH
4UNcig4O2Cmn6CvqCQeh+xy1H9TeWTZ55752CHb15PTpmdlIEE9TmS6myoR+G47Ykqj8IoJ8uPwn
AL1tdreuhp+ErprSSja6El8np/KPfQHTwi8tmMkeRpJ3W3u+RtLvgZX61Je3PpUiWQFcjU3zCbWL
NG7SEgei3uBPzzVS2xuicExM2UCETY57ptz0K/RpswkBGg0CuyA1gDdQ3rpDb7L9D4oJNTJmFL3d
NNt34klLLI2Tf+nX2qBzvwyWsfKv5zmVUYaCgbC3Gl2SqkJXx2KiAH3mvofdCnuzrfKxo72YkwUu
CtxzenJTMMil9uQPVsJGEssJGrKZNXnxhji2ZVkXkTxcCBTWefuzM6IIQyNxxYybvcgKSkgdvDWQ
N/MhOq36v/NPxltDd4PUXBEHVaUyxvb510SfwYRgldr750iQt4bO7hR11D06KSOv5BCevvffdkRH
S3R9Q43KFOlGiJLeyUt0gv9Ke/BJcm0aEamcIaFo69HxMSf2LRa+qAGM4+lk4KK2vgKfIcOdfYvi
5AT8ri4VNnNX/7ghzmAbuS6xsiQs5bOBVnY2c8oyjn1WmFEXv1+S7NTI7GrPXj/uZlD852cTf/Dq
FWMi2LHQfFStaGRpoj6j2iMserwK2aNzQ3c/2ki4+DiWCGIu0wOv6LHtmLxp389PIUKUHx8j8NXV
pocsGtiPc8s1yK+VPosPWAnt37xVdDFjjBsIKFMP1BDvEtiNRUWdKYbWt3/JW9Dd6OwqWvy6Q3nC
8gw/dx6tlBzzSkN+PHeLR3k8qTatpfXTW0thvVeSt6gq4BaLCl/yuVX6cTGmdUh5nwL0hPq7MKn8
xA2YmXI3SdfdxiLMDSLNIW+Da8Bbafap1ntKDbkO2x+VvthNKgzpTD6HwgiDtcqg/KtYqAmpAdFB
jLX4iqWVCEyp+7yF2k9CqixAngyelajFnvV4A4CEjqk4tfyP6BydSNtmVNgF3hR5ehBcb5BEngyg
eltGTH0RQqjkNUqbogsQC84SpflZoM7HAC/WEl4LGXKWTX5IoV/2Z36uWR2CewPw0ggNL75Q2Om1
a0eTOsf+iFI39mD5rFRy3zphcR+uECPt3mz1663VUy3zlnjt5q3YTvLJQ2zJmwBUKpv9KgBZ5wG7
ExytIL/xlWFshvOHM0sQhNzPLEJ+iAqzfR0akqg8jFH/p/CIuAaZ5jqJGbO1K9cqEkDeRM1n29nb
3qU5iZ+ZP4cckTwwpMRS0hWnCACQNuyWgR8I4xtQli/nRVH0WhDQAKTGjA3kIKsn0U2/marNP5dq
GD+YrGAivFhuwYacE+lMIOmjkhTZy2/pdlNDtH+PGdWEDkoFmyyF/qVffm0rYIJbb9UASZu6Ht7C
9KUozU2IZqtq33XiumQM5EBlAQ1T4BcmDRPEpSJZaO4kpok/M2NdM/GgC1CWoGrBQclS2uWd4ii2
EXnFyPiejSI1sHVTW3U0DLXneVxQucYEGRfau6Ku3gF0eN6/XBWHdXgEBJratQ/+VYQbSakMmKYO
jSaEsQ1bnQ5Juk9vLgUP1STfXVA/1uokZYiZWhoMmd3awyeCh40dZ0VrWW8OOsMnGjxbSYq4KZxN
HdQwi3NoEV8iUp6bcI7lssj+ApQIvsx6D4vjPK06N0D2MtohFpXpvGFzD1dNWAkjDiJLDYlaS974
iO8fFvzKKakxv2P3XfNI85//gjUBHHzOHixx9RdidGPX4PoIT1mKXaPlhB6Y7g5kB1E4ZtFy/fXB
0p/syLQevhC4splHyN6wm6uDO1hxSqVwLpDXum0VS4ilekPdA8OObUd3FAmK95eKUzWp8akMB4q1
xT4PbInH6weiHXMMAjVzTvDwdsmsRu36klMU95sXJGVxZTA3ll6i90ASPJOrnhhcLzi8cE1Diauw
Yhp6hCbLPrewN+5GNeW53FAsLPCu3GxPPYPYED6ixh1bHn6TixjQf1xpwNIa1/4NZtBTNd5kD7QD
lJZ1WvDGPyrnJipNNFyuT+OPoEyJGcmx7rzGZ913brmruiI1eVupPfzUfJJ7mElp5670nPYYnVVp
b67iMSVzrf1qmhO3o7mt65XOwVfyBwvvHX1iOCGZIqoXiCjoYKzoWZw09U7uiH/LXylgT1JBOsDy
uKIbRmPyeYkGFa1Pq0Y674nCIwGTftw3W97UcNv2lxgAbpdPbdgbu1sEdBddSc/xKQ0W59ufXa8n
K71BuEHcRjlQC6CYG6BmGeTgZAnNYzRi3NtBpGWlPj6bJXDJPNPZNTgeek0E17bXM660Pev+Es8n
Yhh5cFToX62KCJkDMUqF3puyIIbiAV5kvBzGqcy6WBYVhqtPoyd2FdbYlenBYRFnLtoYg4Su0SRB
+aMM3lupZoT9q0ZbnxkGoArabdMbgO9dh6QYX9VWqGwvqHEqR4/EKAD+IvETqp1LTzjSXiPjyr4O
Us2bh9H4lZMm0oWZOsQg3lm9E4cAsAQimyHriIx35gIU3sBNc9nydwx8Ruwun2DhkFU2mUSZ8TDT
YgI5UWfHf7sF9xURCL2Qxc0yroHQQB+TdYfShPD9g69WXFDuJSPuu1ARkgSwvAbBMi1YkNghiYfZ
Lv7kP9PgFKiEInv5sEzXfn8GjDLd8ZO8GtcqJtljQG/eZCXs+WsPIaKqWX0bJNzaDJn09wyXtz5A
SQMd0wSM93towsms9rY2zJhgZAA6NfA7PIzbqhggcVeXuWAP5eWD56TtXthW4g32n7VIelH9aDR2
ji+pskRKwUMddU0NWgwyLqQhRcO03bApAqfKIQaj+sqO8T2UwVlqR+jPQkxfAwNWAMaNJshClew7
acXomGteUaqaA/PiaIvddI8PRqOLYitmU8nEkwme2w1Gt2Nsbm3sah7Ur9+eIYJw3feKehMLEqs/
r7CD7vhw6QMcgmCrnvWvH1Is2OFEXs8rzktWsFOmaYn1ROIT3fF9ckXHgriiCIEW9qpzighPod0D
oHrni8I2Onve2EmdDxw2/Qa1+4AwOPda0b8dLdHYheEoHeBZMMundAubXix2L6OueISN8mW0zdhm
dGZRmFgtrXKHKTJ+Az+L3me4FrnS6rgIfLevqPzjWA5UTDDNb6RKfiF5/UdufnX0f9Q9AjG/cw5I
HVRwuvKGtAMbqIErAFSJr5wyT3rENRx53AqwExlgR95R6BRDF7PdGIcxN1LkmiIkcIFHJz0f3Nz2
le3xy8KUmZoG29Q5EPrPb59tFwftYWliLIqqrVMP2d0UHcSjFdR6bUehlLKEEIKaF20h+hTetdEv
J/DJYrv2fS/jFsxAVVhPXZhvvwvEcVsC0CrWSe7hgDRuHnyT3/aHKteLzTSSkgp0CpJTSE8dFi4X
JBGD7XYJN06tGY4/OVXgx9aVsFbPZoOxuYvKt8MLX6EL47cvIoY9KkVmWPgjX0UWlydHdODWc5tP
Fj2lBAeDXb3z+nhuhZZJCT6F80HovohH2p4BRLV55Pq+CcyhlgAG/Cl174/v26KSAFZIKdzoV//4
iJSjA8UmveqlgigGsyBUFgpdNF7hjICDPQ2qkIievLBuip3N4gWdyXqPvuj1zhszT1q90dNxYRES
4qW7e86mkksiLH8EA7v0URClMInPX0STeS6Ku64cB3HAnVNejfcjkUKWPgu1Y1DEJCs/M4qTxy53
HJeUMLlTOkf6XW+z1xtmsLEqQK0acwc0N3QAiuUOJxF/gsYqA8hmd9ThBO6UUJA/4lh1+hlC5GAw
DYbd0ctZ8ZTlX5rQ+Yzh5wcR5ImUORdiVolCpNskOOIIkrt1z+oGYy6rPAzwdT4bwRAOEts4uUwm
uEclEifLsPcVMNF9Np2wxGzJakzEUrYITcdphwnchW1q1NjEvdyVc5oHr6FDw5EfoA4L9Bl0hppX
lG19izr7VBTsehlFq75nge2+h9+vpLA1h+XSsluWpx8dvVU2SvVT8bV1EHaaY2AUalFLoM+LgVk7
Mr54JZ5mUroMNSX4F1xaqcq1nmYniLYrIs/exMvfjiV7GYZxsH4oCzcb5JUPcHjfDbzhw2JpM+jW
l60Jh8Q2ZYMJpjHpm7alvPM1UrFFGJYY0nb1xispAVYllir+3qfTim3QtBjnHAc6817Q61YSXQ4S
msnJDfUZq9D2NOb+KoSxF/5uflGzXVyKLSnTBBEpgc3EeO3nP/+glnBEmMPbeiOeegyEKDzkPURP
CN1R+Pl4JV00+++fY23+ydeklwiX6Luuv5r65S+ABQ9/OKDZkAOtO2E5Fl0eHHGw1oLB5NvqhkZt
ligzJcmo5ffQSBb451FlGRg+T5LbmONlJBmMiL5a1f3616CqANvjTfedE6U0Fbx6mofEFhsPSRHq
EWRGfXY7EhSJ/T0GJ0WI8dp8JprfdSoF1sa3cnoYRh1IuDUIx90vhJHAkjFcG2mjrAqs5Z2HoZom
r7/lUz0GUWyeA2i9BrTVO8O+YkX/OscDmEiwQgU2LawWwyf6cKY1B3wek9Pgtgzkr3suJ8YrkTQ/
cAIHF03xaX/erpwb1jnc3focxEcfqYVX7SRoDxILqfDmSLzMG57vzXMJG8/LvHNNQw/p44mmwMkJ
XYjzBIfV7GJlZZKL5NsmihyOwHV4zutoxcSftdaMlAb7MsLFhphvl3RGlMIVEcuCNZJcrsKdZUhD
IWm2IrWuSYYXhs2Nm5roFQSbctbo+eCAIocxhvUPp+b9MILcE8IhucHe8+uq6EBlqvOqLWWUCefH
UFZnhsRDnP8InFKKpvWH8a3nWrKeSKyp+ScvkPkcsme4JOnqbO6YrAyETOM4SUzsgQglEXmWNoT4
kY54ioypJDuZKfFkyQh+SzS2uBewvVxKHZ74om+/zPY21Gbx6AO6lcz8HkZisLIqEzV359JDwF4p
rIwO+HG+yC//vksjFtsBcJnKiinbGBci2TKRQ3Mlk0pHfBCCAGwqijgHowzvpcFDcL9EpCk0WCau
1wHl+cEQwG5Ft6tTmlEstKUHlL4cdahZyXfsCm9L7jUfDxFtUCIHkltFqHjq5hstnyJc6o3kudCO
ZmmSkHbuNYzZlccwrkIscIMimJ/wV4mBEIhd915qM0Ljv+3+7iYDFK95gBGuJavK4eVml1PLh/Gd
h0SfOJJmsFg2oo3X2sADnOs04NyeKL4NIqVwWYwhlaIpU5XgIi3KOF2/Miekx3VYU9jJswID9GI7
Ym4/EdzLia3idZkPcP+jnAo85ROMDFIUseIE4yvBWo/gQLx+vXmsr7l6avlZUmmvvY3A0uHLZbSJ
9Fk5x9mvWspOx6SErKi8Of/ZEC19RFQlN83KdFDX312tYV6nxY3lm0PUd6DRR5STR2GETg198dZA
Uy/vZuVtsX5Q89XxH6sDOyLu6sc4o2ObJz2JYAUMpUd7jVMC/8h3tv0vv+TmxVZ1AoWlIcIPFkp0
gE6EMCvoc2Da8QJaAbPAK2HEY9hwET97NJ/eioV8D4RkegFpQtl1ZU36drOYhMFowBVc7zMR7Lh1
lEj03qFdvVYj+m13+BOPg+bBXY6g+0PlLv7TUiLESVs7u4XnPoJqS3kCkE1HaiFT9FayNRinyAPo
zL1FyjNAaNRZr2IQfvLJkmRabobsxuZ4w4gnS2Tkyr7Iq4rmEovK/Cq/rbbApJzfPBxV4Ksw1JYR
U0I1+/t5/JjDHEjuZpKMTE0WJoXuLNmLyzxHP5FX7acEIOdTqZoUUcehboy75cUF8VPDW7fJ1oLJ
MA5yvgyG85Kn15MuSwwM6Mlv8gKLTM5bS6nGbzRjNPGWLuc/Hj1sYE3SqvN+OIR9UB2GGgleXMny
ZcQCzjjwoitX8ODx6OI6rEg3bY+FgeGv+HWqxmpe+UqIP2naI11jzQ6GufIvGbc2Im0V6FI+dn4D
DNbadaU9nJYPmLAIET2JxAtTba4LH5PyIEhyVZjAJhZqBzv/TzYOv8lrgN8cHHBKERgZOtTc0Ct8
GJk938PmBpg/mpYiNKWSiKBmCjSMMTq4RJ5HZay2ePX3TRBFZFM57J9wlqTYhmQlIYDE/wxOBU6G
FzFHRDI64WfMIfWV0QnJvx2P//RhdeCNDdny7L0kQfD+qXYjoXxYSciOJfFt2R7SGwd/Q7RxydDR
ytzjtwkuLXhIr3fgigVGqTcVrIEQCysJqo193Grj7oQgoJ1nvYTqYxcOA1zuA85ADI167FHS8HGm
4Lt7DdKYBSq7XmKUECxTCPuSEQJdlNCgRWZNvSHWypqTB82f/7HqjJV9mz7IbF14bDwzM3eMTLCL
IoBaepOFQmOWYTcVmw3tk0ZANFirStCxf6hQocvkaRKk+3MRsUT7lwze54+Fdojhsvbnw4m5Dd4D
I9FxgzWPWAJ4CpnIrgxoWP1asWWubdtWrfPKgv1E7ZuBY5wGyAsk/iECnpGWG3gPJXD+MxklNg/I
vyXt+gM5LLdQLSXs9TCzYxCSMomWaXlKNYokvyr+wQkid220QXyDPg4VHJZwrMAntt2zuLqh9pUO
yp8icFh3vfc7WXZCaXbM89Hr51Cp+1anXFnttBwGTtdUzIFzly9YrVqWBk+Dl/ifVlpxnYghNHfM
BgtGTtmMT5yKzng7Q25OSr3Gf8x0JbTzOYwWW2lhNx3QHqPSF+MRJBCuTwvxAFW+WGjpxMEQLP5B
vIR+UpaYI/5Lm4zOt61JGmOeDtZYomAt/cx7bizPAKIg262YAG7hEmh0cST45tPGaPmdUEGoV6on
aqAbbALVodFOJpUAZqXR1tBYgeu+w4QQNUkWESFy+j1reNFEarGbBS2eedUX0c5qsH/UyEUgMHb0
m4qOesbyySlZN1RrG+s0VeAbVQAL576OnaCUtwY8jAh+PQVtJx3CBFy4frQUfrSfRWZpulsYkZg8
aoEfphTKLOQ6NAtk9J3g6L4SL4nSMDRUSAOC/iH9DxW1uizm9hYbKXD8C8Bia+uBlmQ//wKID7AR
R33EaMj8S2AznCdoI1xmS37RfyQJFm+9rCPl8n3Wpwtial4HGHVlcV8MLBpOkASb+0siIS14qaJr
QdxCFO/uUOS8U8ejhzoDb83UzuIOVxIZLKxMRox6CSSRDJQq1uMQiQNxfjdf9AYjtxwyOZzH75qS
d/WaK1p30+qqSBHOznQEChxUu8XspiqvCKRH7JWZNFxYy8YSJhKwB9twKFX4PEcMbmbw18ZMcTZa
bNpQ0/CKticnr8eUJPwmovTzr1ulvydFK+XqBKA6bsEHHSiltrWWCPlQdhUJdkbZhEl2UANL2nKZ
S+36xEZK9NAaZmiXmA4r08IbDZmr91LSYAzFeXQII51N3k/xmQ2Dbz3v9va8OYTr6U4CcvafzWzU
Nb4WH46rMXqtc5zYlbQmbXlEf/NmbbKO965NIZDnAzG37hHQTxEiCONTef96oS1n5MwO+uMAxLx6
fJvRH7lwpbpeO9IPJ7aVZsgdHitvaf337jCkCdbffkv7CmeCnxV10RmOjXnN+7O5nMeZixyUcnHl
S9jqIoZ+hbWwHXxI5L9dRm2k/mkisBRAmL9OFdDEkhEmLhTSD3Fk/kIRQV1q2agdd8HyqEB187fA
EqlrXmBEuBgMoBQ9hy1X1khxy6JRrKTRSpCoo8EAiAs8OcY1qcs1sKuOIFbtC3FNXptPmliCYAQn
2MKhIMIvT9KWxUkMECrwFy47E6jfa/W04d5z1P18O2NJtjUYDHdhxr03G/MRKru8bBjwriafNuT5
hj5oyAkCY8nK/VHmtJ/AJ/O2DDYE5W80EyJ1oF7pBVqCDfTc+7zhENXga55NzwtSsTLl1MfLZnM5
tseOWokPiJNKpxAHMwyQeUcJYuaRQ4uFqbKwBSOrAq3Nsk+X2eMUqkW1v81sTrvoJwY4s9EFayef
8PgMXWAC1642nyCYcmqDBxJHNURiOm9F/zsixsuCF6lCzKtOALAn9rx83XVDwL7htU/1nEiIOvFO
K6b2AK7c18Iwa6eXg/IuvYa9Kj4sPThbHkH81/lMo/gjIN6Agq52fqQ3Y2bWj4S9aqbA2kPmonWh
UEWZd/6IvFHDxN+lPP7xJSWhbsUD6vM9EAW1Ey2i3EkbbEevhltxUYkwtZqwGaBqv7jczyOi0vCy
thHW1scceXc3MrkcfvF5kDC3w4CtvUn6RV0gGN3gbXUrbeE0lcFTFyjeYH5iR35glOf1VszJ8qOe
cnyTzFrRBXA+9cpI3MP05azAKUzLsiYqp7PPWc5yqdHiszAAVd4vvBMvYIwtBkwYqBHX01SvKxfP
FsgdbmOpij9dCwakdZrsWp5KcdAxkOZTjr8cnh940JdiHe/Y2iFfSzxc8q+XWiXMh3ryu75PFKyo
HiojDXpyN/heLcvbbFc6QotuJIhbc6kpKWOS9mfDpgIf+3MFD0MZKQeHgRCXaO3lpr7e36ydq2k2
uBH8A1UT5LPazeU2cmcGFTU0m/JuUXPL/365R1VpKxmi6Ku4BciXlS5dNy5Q73a9yYS8UWKVYF2s
u0POfxPU8QM6SXI6alY2AaD2ckN2zqeME43PQkkQPyWJnp6d8IIuvb+81YC4Y45dCrjoC6k4pCso
jTz6qwvyMciYuU8UWlW/fuuu18wGJW+WA5W2LgTSoE8INmM1SyOgZFGfh6jkX/a64Eyu1OQuCU/m
B3IvlkZBa8K/4ZacgEeaiE2A443zg3/sVcY5LM98dFkYoqddeJxKAPwP2kO57LRvS/LhxtdYWx5z
kMF8vZy8VCTT64BIRpb6Xhf+2U0tfFffOiTK6S+qDFUXT3Pks7qwrqq89uQXF0HB5rC8xlqRgZVX
HXL6QU7QlLS51rLQ6bzmReEjlb6tH5zAHW8fKa0Vkre09h61IKXVdi9SgZxBprYkw5ussyHRwKC7
tXhJFwjcKvrHFVmzZ4tLkZNrO1QiJczm+Jequmb3ZIW6RDEj4rwoHJDVRfnJNMSgfVpicNoRz5u7
bvMvPPWr3LlzdcfMjn+0rhIZxYld8Cs6/VIbkyMiM5/WXV7f7jA5clUIk7NhIVGniZPztzv9Q4OK
aJIsZPxw1H9a9cjWabJ5NaRy9ZOPrAQUpiP8mT3Q82I0XTRuV7XNtedZc9BPZBuF/chsLnm00j4b
Wk5/xvL77b9rVq9crLyBgGeUSA6z+XRIhI7qhTjZnr9EOXMG33NEs9+gvjaQqHmI2uAiTrWQ0JMf
0foyjK9yLJn4XkpWO5vLR33opqSGSCFt+ZgnE/op4DV9FAtpOcFM94/cdqXr8XeLuN4ZjALCVRKA
rdKoRdwCMQ5PORersgjSL0dYf0RPa1uvXgda+JTRXVqdbjKM2taXTsH3rKXdDlJPTyjTPlkVIgo4
l2QXxON1UOKMz/Cn2W0x+NMnQMMCJfRu4uw6TBJUF9KmCeUUselI1qKr5pEVhXbUeVn7Rc6n51EW
iam+1nspQbF5Cp/aIK6Q9uvZSt0QGArtUkIQ/cyIy70m3Z4LQ6KSAHeSwYwYfLLx/xM1dI3O5GQe
EayRZfyXyN8MVigxIX6ckX5mW/V69hki/tUcicqJAL+dyar+r3Mjs4WCBJsksu+veax7R4Wjq/cT
E0si6OM2FOs3Lnyda1YvaI1urlSdq6yLjiloSPcLaVySCHzoBeIhTIvMMfH0pqF0+PW1szhdhv9t
t3hDcF1EpVLFbwFqdZWHgVYCr78bVYqNWyC6jeGlVoMjaVt9qZP0dMNwPPBv2Id+V+vCFdygn1Tr
6F99Y4Dbpa0uJUPceNvIsboVTt+Z9cQyuwR3RNw9pCfHevLUfjRz+vRkhVPgjCDFV8VEXq/32tII
rPgS7CKQJt3O9pJuq6KJ0KyG3m4vPBmkbJCmq+4YtbJvE1ZwT3ALXduQFUbOhkwYpIw0bqSfHKKc
rgj/TYUHc8Pq0m5se5TRNKkDYGp7wklI5Yv7y/wmcCs0rh2M86ZWe2aTi2QrsXR+j0TouV9E/xjp
QaSJ2euvgsKCH8z5qU/8CnOR40SR+pgP+THfhi7fTuNmBSKwi6lKfa9mV6x26ZvGePIVoPJI2/lG
hCtZt7JSDRsXQMphiubZHSBLTRj57e3qPWYO7BxZT0pO5u/W0K3zj2IDoVgagXFzHzjcUSLaLUhV
i3b1pYuNjKrA7SUWA3eJ1CCry421ArUrCcOnbckoI0mW/2kFasXMbFE4j1Gi2IUwFwyNivEq+sJa
mpJRKKcV23LNCpnE19Bi5qujttLjJV0j5KnV/BxfjMexwH34opaZ+oTpYmyWkKiFds18Ef+HGlA8
9S+1qNtiaRUGr6xE76tevlXCVZchH5bxWB8TKehSXEEdT9sfLmciQXIrao+KJXV1WduVvbel0uGV
0+H5ZnVPmHI/d4/1ukgzvkcozWIN3mn4k7BfkLBb0tdZ8H174RLKjC5CT0tw+uyt8aJAZaNXAc9q
GJ5fTqgdcmRunb8e+SDkoCS3XVfyz4wl88ScxFMZtGS7S7vNeWw+dfs5M4QvKThwLPmlgEHyYAee
WGGI0Cxy/0xacvk0e0HAUQV/LLv2JTAdBCKMtnW7HJh5GptxtvklKYVlg+e8Yb7sK8tuQT0uSlHh
EP8qeZ3w7zEzVpESmuAXYZzvHIiuXU1mZYQmdLX6xBW7GggmCS+iqqypUzllwJ3/W6c0HIqeqYRt
GMK9EFZkeaGa33XP7lWdw5jPpt7cB4eurOrLcXUqljpYo5bzdqIeueh45BDNNBpOqXuufB+XqHbI
ZEmUPb+lv2XjUMYvmM7U17Qc6jSW4lGsYqp2s/Ht2/Q0PIvTiZZseaL7goXrKy3FG9VDFglAzx7M
NIOHqBZog80dUuYNQvGdqeFkUNW1LbDkDBj/IOFxUxELculqmbAXWE4nrC69D023svggqR3q4mrI
hP9DuRyh5Eaal66ZTMgnI84aSPKn115D8g3kwpYziz4WHBtIc3USyqF3lUgwzV/QSMnXymZZ9ZZ5
YodjNTBup46LogdL+m5BSaoRDkRVF0qdGqBRunkSrVXdtbziez/YfLgi6jTo0CfNMnonvd3m9Rq0
mjDHNvEl/KPWj2B6ACFwpgbjYVVC7aAo9cpH9kXvrQyot4DeZubqTbmW4Whibo9YoeQdOpeI6jGF
0CZwM8UhqsKYA+ex5S4vzudBCMwSg6uzpXQYPaG1uS41e2+FZgKl7IWrg61paLKrkeP8X7gq8SvF
uDIN2blFrD6YBe3CWYiPC87RAUJmZmRRot8dMOXSC2nZZkqk26BYbPpb8qh+2yYwZl9i+UVNBSXL
IDs8veCR3nZvTQCJwKMOn9loHQNzBHPVrrnp7iwiZy7JeP3sch/ZWRsxtEMuC/qV3xK6c3hD5eCT
Gt3F7mcuDNw7DxnA5P2P/lPF4dtY1yZKdOs5WnwnEqGOPTTs6eNvzJiv2xA1m0nzTI7fFGwn4rrw
+DIATaFxDqEpCzqYuR+j74UXzROq9aaCwkWYLuevIAR5EAgp56ZaRBreAnJg1X+lZ0MwRW1kRdKP
kiCqm2z5mAbhD7MsmdAyo7XDOvryuXfT90g9xD9DgnGKNySNd6OVv8p8w+oSOppnlAy2Rx7KXzdg
RVv5PYZx/TQ3rTZZZKKHtSTP35P0CVy2eM303nr8UglHIRQRaR283OjvRFJYC+3RsRtl8G6N0A2i
yLSjOmxHPDlu0REtm2AzCuogYEXFPFQQT5awgumhgsU5MiSL81jVm10dB5yWYygqngwA9KbpP6iT
2R4CT075+Gm3Qp86QN22nsQOpPOD8ZtDezz+EUq4C1DOIQpwU201T7E2TQfvG7rpton4KWzZnoXe
d/QhhF+RBM0ydG63HMHbqMSdbNYeVQnVOoD931AACREVBv9vd8iIDr0lzjuhkk19ktUoAIry4BSu
j+LxSIWIDNbZXsZAeTmD8Yc1SSa2pnj8Zf6P/aCXBn6njTShmstVaHmJeDd67IA/5aoxSIzQOnGk
tRmb/1dRZWU/3/H/J7HM5xfwElydmQLNfr4rmoEKO4/+y8CFqrEgFpw4rFrniHiKux/XUV+G4ZHx
VDLBCOjU67Yd4Tiqs8wcbdVrIsJDQLRsXuZbOuiC9D6bgi8RkJAuPN+iZG/B4XWiRkVYHrthtNEn
Z1hAEAr+gIuwQL1PCMminy/0Frf7QBSHJ4pABpKXm88LjwCscKb300EcCXaNziVqVCfsB/B7N9Oo
HGC0TgGKCvlZ45O8ouiCu+dP6i0yTgW77Ru2moCEefr+sgvOZne0TmLYuXIIwUyYy12pT1Lcb3wT
ln55WwWzSCjnNdta/yggUU7ja2hKs69YqmfZNDeUBxudIG6We4Y3VczAuy+5ZplTYX1W4NgQt8mG
jj0XKPqk3nwA4lsOaDf1Y7tRoSwvM5qJzOA574IqA5nnN6IYKro3yAo3a6QQJMh2YmpSht5/YQQW
sbbKk8EJL8DDiR9/kB9XI/qACnIdXEkRzrwjVsutPNKG3HS3oAUn0W1oxtIld0h8SoBeEAe+vzX4
1H5U/u/2Y+jJOaSmHY6AbcybkasDXg4BLFoLyLRdV03ayX4fq6UgsV9vKEcwxCzNhW7Xlz67NPTe
nLTg/k1pNhMc9EVTz7kIo7Sz31e4a3BnldUul9MhLgt2o6Qg1ry9sospUcOKaF4Ur81XN4ayV4o7
TlMo2rf5TBQLPvTLs/26w04g0Qt+pl+Pts1/9I476xP0l6LaAAlHfvOKHkP65eYUPnvgkSAvC++R
+cS+GcwPuaHOifdfnMmld++7vt8VweO2DvjbWrLO8xpH2S/a1PLZpWb7HsZ2J7fodDC/ngsw4uGI
I9QvJ8AA+bxRITSnLANQ0pEEJNE4nR6K0k2T3UyhcCqUVO+ySQSPTsp/ZHQF/M5SI9b0/qA+sm6d
rwRIiDSjEXh8FZ25755TFwphFQTsIXrHy/MWbk3RkKuAEmC8cTwbY1aCqc9BvYuzn6X1Nn1np/yt
ZrEMjxqXorgccGH5+04qmtEYivWKYKsM/SaTEChUkQJAo/Plz0I4WNmTGOxPiaNUQLnINnqmKxpo
eXcXbQ2utoS5bmCr90vEmdaKoA4F833MAu2ZVf8K+9WNhpfnSyKsAduwIgQv/euUAfmjKoveR+Mi
Tjo/yWMiPDhEGSKB+fPi6/4IB9ZFebTphocAYV5aFNYNfrY1DoOeXuhTtdU1bzMgeiP3LFLZDfda
Qper4xEm4tA7uADAhXo05U9gYDvu0ROaacD/xgB/T1ixfhpSTwSDeClEjzsUwPO0P5AkLezSRObn
xFx8ThwCto2S12FjMfgjrzutVVQqjE5xRPpDA417+iuUelgiHrN+DAeVWxT+7b7ht7nWOjFguY91
qLp0fTQuVMA2Vsgi9c8t0tBa+ARYiHfGh00RNDCZyFRsMBsPhpV+FCSWI7FW2yXI3NYlfAFNjghk
DJMF6yi0giWkrd8SK+TS+DiPY+LqAqk6FOpYKLG7FIyDWsyVJrd2Iwcr8h8hKtuWtL2+K6IKnkTU
LHuN6qT/7RZgW1VYmNL81FPxF0CX6bBm8AjxHWkUp4G1LrSPZTQa1yE8+IChyKbcTFjDDkGZa8sy
SBeQc/Nfbz+LTwkYxfp0CKgYxhLzhb/MMSZ/XesbAvEdVuKKqWHJWVlbMtN5NRNcHRouX6yD+klN
+bKm/xApCkaELTh4H1PVJLgka8ApGBHbvTPUkOeVVoOD8WB2h4INEObasPyqDKaAaQMdCkWByTPJ
2+JAcZQjPSqwnsowh4Rq4Zu7ogWsk70087Ae+iU62xUUQz3c1cv1H1j3wYM8u/92HieK0nbXpvMR
t6M1cyTk/y0HNe6wQ4Bk9jDkKj3NvSuoPF+6S4GHi5HrJp44NzGdbKrM50wYqS5xyDafPxYPgrfw
0+CwQa058BHffilHBfWgd0fOJsUxEmzoOP4vd/1S+2b3vgQMKblwes0b4PhN/3At5TSkd6Rbe2BW
r3Lyv2R6jUrLGSlfec00j8uCfl5C6f/k0AqvpTkdGYvCvr8oJ/9HJJfo19Jc+LXBKwJj/3EtktZn
u1v3IGVx0hlwh0N9yj7kOvWP64EL4VrS7pV33Ntzn2gYmRnV9PghUSVc/g0dKm/o82w9ylKhp3cv
IrU4LowJ7b5+vVXQciCPO6u2i2C1RoxBppLZjY9snHDZ1xDsAJB8K2rSal/zHZMRGdH9AH2fUHim
9eRlRutjp3BGXm37GMWxncMf0shC+LaLYuR2Oeqf3nbp8cokSJhmNTeh2z94y8q47n58VoqnktFI
/K0KEYvA1ZBgyR2neh4ysy/et08FVDg6Iqw27VqFF1jCxMm2ckd75wLuZxsxYGXDoeVbknIbz/Bi
PtVfuId1c6fg/VYTRy452tF8CMguTBbx0paYZbGtr//1GhQxFLkS5qagyFaOW/PhCq/EcmyflMXh
JqdjSfu6OJx1a6i6+bXcyWbQBTTx8MutXpUkzANoAflctCCqOOedmtxw0N54ojIlF6xYfQB4Z4Qb
shnPhvT8VjoZf8nt04pua7Cs2XOuRS6C10gegEpPJ6H5BPgC8+jzkAtljaN38pG6xm0Qm+uoSBJU
UsjUKeRYui7ZIoOWhWhtvoYv+MzTmEUrC+OCtcs6s5+zLlV3TInUzTr1T/WJcilBDBFkvAh+UB49
CxDIqw8YqpESNqhiflayMePNdAGcn9GDhRnFRizF9QzTxlDdB3c6EOH3ccwcA4CuhC9oG7qH/ZiA
op3tmETLHa0SgcSsY0l2nem22Q9lS+dCi2A/cepqnhptedXz+OGYS/Q9uUTAqBAPoTyecziBEXXg
PiSpnUtGWuhhySCf33dPMPIKwlwoUGv9QwqxZi0dPOUIUmEA+Si5nu7Vi4KPZ3+XTh30Jn8CexNB
YRU9l1ceROh69gMcvg8b7fm/alF/4Nm4yJtYm/ibyABIsY4Iyfp+c1wi/w8yyP/kG/24GGoh5uBE
rg4WpvSdghqDkBCUDzNOGcO+Xz9kFE15jsj8ZR2QkoJzzLiaQygOX+0nUdodyjkV6H8NFiqIJDIX
z8abXBNTYdH+d9O7UMib+iJEEnXrvBS3BRQwnlb/Wjr63BiZXjIFx4l+QkIAqz2p6mvcBiLxnsC0
XxmOiUygMsge4SPmGlTlh141FEKQNJeCQvb2uFoAFqubzj/QHSYxUgucCyThE5HvLtRln0hD5C9A
t0vhE0Y1WAQqmSBJ9RI3UB3TQQIPAkOd7iBBLAkGRl3/SJ7gKv8chkYu9qys+0AoCHpdp2J8F/Du
vIzxc8Qr8ZjKD418njbLtANRUNeMR2e02Pq0KtoE2njOUS9S7rTTDbl4HRCgYRMHBAs3YK8avUEq
ELXiEGZdWtg+MEPWELvPADnfaBaq4lNi0lk796eo4dpVRqcoLxUauhmQCRkxwmW3vPvHZcp/vKLt
5FKuMNSwRbwXTxH6nh/AN/RcI2Xt2X5Ybl5NH2/0dX+5jtZaPoUiknRCbt2QKfn0l3H1zCun7rvw
isEaXpTyRX9pcEy1CtNqWjQfnBmmc+oOUwB/SNNS3yqYjaH8CvTXzKUgZWonub2ZHqdVfUAx6BKO
ony8yOvCZ3dLqY/UObsWY6v/hpjeXZJK7P4wH9zMF5vc4RT+/cv0xTaO7iJ1Sohl/42HJPNRy98z
4QsF5fCi329mxtEXYqvOgBCR5OxVNdmih6sHo5v350qlbicgubeQyFPK/VRC4V39RSrCNUGzkFBb
UMNtNsA+PWpXehegB37ryeHCs8Gg6tPdvR0Hi9Vr++M9fAiHUImvQHcZASRucgw4pEU8U6RFvVMJ
NoRKqxfbmd7Fy+sxwFzzHKfMXn2Nj7yXoG+ya9mRGZfYzI1OYwjDZZulVDATBlbKyAT6cNsRDnZl
XlkZIyO4QF9/8OLhgyRXaGafFaX2jTf9UACiVpTCbgNEATe4FhAu4Y+UVOpjXjQTSbd6AfXMmEU6
o3i4IdnlckXKR+J0lL2QTb1TcdvNa3Plk36wXofl3wmLj7U43oX8q30w4IJiEHtq62kZiz5qoz9O
Ztgv8MP5YGif8fjwRmg94AcLQyMFf/2l6gSBcovWXtRuHVQz+Xc/qJNAJVqwAm+P2HZfIfnaVDPP
RsaXd/WILlx+zT0dJXfrEmep2QkDaeCkspOcKfWOm0M5wPdnrSUEC/Ncf55eUU3H7U1+LKyk7PGv
pAxHWADVT/H2Yp4a14FRK5ncALy3GygJR9RdZqRCfpdvkq9GF26AmNUoBBYmh0Gf7DunUBFZZRih
VszHA/xF2R4iAwEnkI4/L1jxBW0GfLVmR1NdEtasXPpaXNxdruURbrfFO8GHf4S3BQ3wVeY8AiQ5
RtK/vj2herZ27UoLUgn/YdV4rScjpYJKRXyM8J7qEdEKR/9t92iST1mSaa34zdDDT/wbuSNQZwxo
U8w2irTrZr/Vy/iCIt1mciRRs9yX8Nv01DC8Ie+/VNY8CuAhmdkIBq1kghd975hQldUF6hjQ6r11
mDtBF+a/s9CzYKYHL7B9r8uLJbYPUP/JZfC/2vXKZGqGrNh6M1AuAsJ3EFvudV81WHBqp+5tdp/G
GK7KlUolaYeWLdFMkE44NV6UGVM2GQaHNDOJ0hMAgxoVfwZaeZUPBEBoJw3AjzdpcKu9xS0yNBMy
uvOlAhLlQWOiGCGqlLbNiQg/+Bo+gTXD76s9r3BX9bsWlutruGTT4zIh/j7UM0MJNqhU8OBCP8Q4
Tk2GQxP6vhw8uep4V1xthxnSo3lXTIplQ7cvg+nlsjUJqwJuZd0iqnQCmh/ouNUTUTetnpQk5J6I
Pnk+J/ERvIcioMI6KLl7cOBRWqvJVlHBLApgN6ZEXjtIqVXuxU9UNfJ4l2E3Llb8QqpxWwK1Z9Pi
hv/BCHM6A101X55hWac4TyjVOhnHZVFP6ldzU0I9Ww7ICbcISPYUgwMrNzx4wOVaZbZkXo7+YZyI
eYIVYf8z6QcBTperPluyZ9Pn1nkfhscI347QDtC/rUbyD/mkvM2nCt8uqGDtI632pD0wIusUGHVH
fBVQpy3M76T5tTzkVy9XXUDyxAQiyODxFcFa70IxsuL9Wy/Vm5i0U7Ju3EY7pJ7FkDgHLlYKe8dk
O/kaSAPQuqrwCw2atzZ23s8vxU9LxUXQaShK6LvM6OtPdw0IbxEPY3f5f1+nFKxUN53No8YidZhY
6woR0prwIVjNa5P6DQI0FWjkN8r+6/kwINgJezQ3SJTCvhs84cfocMBXVG6cIQWoCnnjSOGrpNC0
D/twkiHXTb/UA9WNQwUQJOfGOADKRk7fDpW23wtWK/QR9tEZ4Z37m4JPFdhf4AIR8CsUEcOrO8PK
gaGLQqOCq+VxIcus5/7NrOOvX2TKNn1uw9foK0k3LyQ/ClfTUKsccxpFmSFpKIJY0cnNu1FBvLYD
mP93JUDCM+0yKmmP2aaHkMXDJasQpfrpYUZUFLLHZ0Inb0g253ba3EOu2Ta7AvW2/dTpsTjTQ4Us
T7Wrz67JjHXjzDEwgzJSHPAcsW8QZR3K5fMrET2JyVae04s33MFlNR1M4eUqfkCRBa3huJW03Ez9
MWbLJ5fvTjQayUHFbUxQfGs1d8DoYax6b6PH7Jn/49iywZxq/OlknMazN4bu4TXnpyeia2P72kyh
pp3Yn8yYQqdGI/zRCzQtfX8evckroKMs96jOPvm9MG4zMD7qM6fSGKHO5kqzfa4lgi6QZUgrn0rU
rmBwwJLBn7NCdv5bGOP7wIliqKwsXzAkzY1BFYRvvpX6311tvwDxQmY3uagKOJumnFDG6DE5IsNJ
Fl99ZG1ALeFy/YhTPVNG+Ri7POER9VUWdqqzQIF9ZntxXjpJvSO+N9zpC9vz8fJ4cWNlbi4cC7dQ
Fj88Tgpe09+8mDTrAsg2T4A+4CwL3AHBneV6UEdGEF0lebDgzbNciGkSLO3B4QkO6rWVtd/7WtC1
UOf2K1yO6qo6TG3/LlL71mnxAgE+XQz+A3Uqb6ugqP82Sqt/2zk4ScvZqu1xxhYK8IQdcy79TpYz
1N1OsixHjDVObV9nPoObQeP8U3Kh+pNxPmHirn589YbMzGQbnyFtzQFZ3G07DMMyhlrHrJAyeRmm
fl4W+kdXr/MSUs+YPksm8+NJkUpXVxrjkWkYKDNPu23ooVlpANsKGqTZyeeYAHHEbqhjOf72VzZv
8sas6/BMszmX9lCCp5AgABjNB62pO/Zk6ka0OfepLHNPXDyyxhhQ1YF9rOVhZlOUCy1zqg22++lB
7UAKVSeVTkjn009Ma0hSb9ZMmRb5wzOOies3VRrZH+q5ZcuFKMcUI9j5A98ziqlorknp2V5RIu+o
DJdljohTG2O7RTPrzKK43WSuP2VC6pSbVxXCW4lV9Ol50PpTiXOTOE8Fi3pc7GNGPqoT3LfKRLer
4h0kKvAXw0Gfm3vja+Ie/+WfV2meIPmUsSMMuK9ngvezywQ6Ycwpwr2Tkpsq5FnafXYcV9hQzx0G
mJLbk4rmL/DP0KWnMH89sCUnI7uW3Xpg8teUeipP95Rj2pFSaXTIH7U/MyhhOhSoNTq1cm1LeyB/
nrZpf8ERV+UESTR9GvchX9y1/jZElrNMaxyBiun188ggSl4iydofF/LI4l7X560m2AdS/ykSdM+h
ry9D0pO4zQJQ1B5Rv0NpoT39pIOrlHBpXXjBvtIIp0sTXLQrnhrPnigG+1Dd2GMvxpSd2C5BFLWv
ClYOg7Fu8BnO6QusLDQEEzUZpDNifQtMp3peo9KGUmjcQEOKUsHvjq8Jb19dtcO4xc7AJC4BHdu4
oA10zlP8WZ6Si4+NBmTcb2bGSSAxuBMOmFk9Xb+93T3J98P33Iyl5fFkDVO2TFFdDUZokGlhVof+
4QXOtpBZ3BmMJVJbPjtoo8DXU3e8FcPO/8Ue6GHGoTXFPJR6xDYi5GjFMHsisomqAGsR1fSuMIjb
snJnjQ1Z/RUbSdRtk5oKW3Z4IxzlrMFggSurJEu5ocys503CgXE08JN4X3HpSA5QwCrczuPi+gO6
TZowjZTt27ZjKtZkX76hDf/wJQpMVtMgHLQuh1fV6yNn5nfKGk2gmzbpoCbJQEzlKusQolgoLZ81
GIlGXtmeAhFJBcWo/K6bMzMxj/fwZL01fDpqk9Tt/WQuuJaXtahR6L9cg2Vg7xldSN3shFq5W3bG
KBQlg5oEaUMjKJ35YHcx7y8qRmC8fvQ7ZfsTVwz0R45VNsxjtXkv8zvRIwzf3NhjVbZ6GbJAQyzF
ycbSng7fYB8nmoXvVSqQzsIpLNlKtsEn9DB/TPyhJgIXlvBzukIE/N3UQP5Zex0lXInpyNhd2scn
eJkK4OfpS6OSvBzVs9Gwp8LhnH7vDFKnm84ImXV4ZqWbpXM+NBDiG2oaS8ZS93+ejfNGkezEC5ff
na1orSodYsXA40FuR03SOp5XIUAjBuCCN2yhoNjBV8j5JWdaf8S2YywTXbQXV8/r2lkNaX0lEurX
jOvGJqpGLHKK1gw/xIozmTpBUVP5lShCKd/CmTvxRd2bKLTvPcUavmEpaJojzNjkfDnRkp8tHU1y
Dp7e+xx4SHvR9Xe23IcJzWTrZKZzmVqMoeefHp+YPb/RHf+Un6p0w/fvfcuBcYLE5vW2f9RsvS6M
MAT9kt2nL82lSYmRx8QtWNgXhQCQD1uiZqakf+weL3VW/HAKNp2IcMC/fpnXH3GwortPuIP4IfEL
20Y+giHYJoRE28tUsWKr8Y2M6EVsUkKzkyB1tzruxZR9wIQxlpORcmo68se+Ao4z0CHCmlAWzSWK
F3vJrkcbXB91aHBblOeY7wN4u+TQhv9AXh6od3tk6nS5Pkqzybz+zpN080fjh2Nf0Oj8IkbGojo9
VLhsmgtuhT7yX98Bzqzb8iY6PJXlF66DvvbR3RwOwXqP3E8Toz/5Zoyu1cezOCN31Nq/0CJTk7RI
4ftl3+qaQe3+LCd2gqCllhPF8aZdMvLqf1/30FIK4kKgR4Xn/ghGKCFUvf/qZhEi3pz51cF63vQT
vUnf4W2AHGyi9h9atzQIFwFnZ7k3Af6hX81yQw6sBOk0kMoE4h/ruFEXm3d3KjukmhSFyn45Npi8
pzSFqglG9BSpA/uUJ41n/1KaEHhF1CgU0tSQtDTukvXWhowbp3ovQmEkfFIQjjlEvAIrlcEuaBFy
zdnlE/xu/sCnNDUhdamhVIhmHtqGirLidZkEsAvNlCQTDAYcgZUh8CRptGofteOZlqJjvd5qbCzQ
NtGpZm/M7H2mxKwbiLlFWofObZA946zs7ACp7U1uWATznQm/0oyyO0xH72dmakxhFihQHOiEbZkd
lg40OcC648IIup5btVkI52Fhj4lhm3rEKh2Iko7Ws7dqNDQ20dfazBqya2iXD/FAXTRH93CqYBVG
O/1NcTwIJKCHPS4hJR35t32vGrdhd+QZhq+racJPDhkLz64wSDV8p1MK0+YsZgBPuHESuB2OiSWv
WxnKW2EnQ9f+DyzOUrzvbdGWvW3UwNiOEHJjBhWip+rb4NeMl6f1tBm9msF2RhAnFH7urw8uPqMg
k+uPZBtjst1WkJNhgs64b4IkbdrXL/TkNiiED3NpmtcfrxBBh8qwcfmRXw7hrMQ40OPxnGe8dmzo
3YW695gEPCBJm7zh97IF4zC+83rf2E+o6SiAZHkXMRSznBIKItl1bHmpIg5T8qSqnxPK0C2K73En
sf3mTiH4sW5667aNeYnMVWZlG5cI6H8Oi5ShjIbj2FEsM6srgi4EGdAqidqJQ0Spcdvgpz9yoN1B
KsTnjhqJKMWVW/M8Vwx5Xtm58VHuELA1bqnPH+n2K9psbCj/8OVq2JnYHGYy3dyX0LmPZVI4xE6U
Ua0lh5A0f0XVn1TfJe4qfICqDINrTAEBE8WshY3OvF5eIxU7J6GnPdQyIn7Bf7lSHyG1cK0eljLO
57ULacJe0xPs+C2g0Ow99wG50lmtc3QdatrjwEDPO/GcBA0Cqj8dBDhgghIGzwDyChoDuQmL8Osw
n3qTRW5dtSvaPp4CNK+Pm2HPrCwU+xlsPVEEnwmp33npXwaaWDjvpuRtBsw2RetwPjf7yGZ4ZS8h
9IFBXe3IXcXKu66GdDp413dcvCiwP/Ro6+CYU5fJmLQgBlW/9yBS0Vm1SF02GQ6iQBf8BMbwYSxk
qbwXIao5lMDsiOt1Yfj/pxjwolTyzKD61rSX7OEVwPIXk+UiBy9l/gqjN492G7BWpQZWsJ2S9Ntd
c/6wfSUdUtC9/3t2/J6nHeILcJKWC/9ZrxJv9WXrgvvF4XHxFHcETewYMlpWrxtbjnKC73YSoHnG
nzkuYBt6I9Y11ypESb0OvD+/cz3Nbo1SKIWRcyKLwGMD7TosZ9iGu240b5qMr+ygcUQa37yT11Vv
WHoTIcpo0sMm6VxebT89jmgRKrfS9xaTkVSEtQK+0npTubCgzP88M6MefMl7jox5avThhcOa9+Jl
LwtN+nwKBpRpyJMPhAfjGmUoDyP8K0hVgMIPRMydi8WWs3fZhECnRhfJsPNNOD+WXVSz3GTbonJX
ZW39E6f7NJge7ZQT8OKXr/eegt6+iaGIbLngrX8puLhe6g5/RV8eZRwZMyqJXVA9+DFRdpTliCC2
IHQcHM7vHF7fhp6DJOlMxpbOBMGqDw3pCjGlDjubswFvTHs5X6kBENzf1GguxpBRt8doDf9juXpe
GZQpZdb4NrLTHOstNwRgO8J/7AUS+zzOeFXmH6GH1EdlF3hLmt/n5CyMSE3UZr7/Ey+PtMdAHhqY
akszEI1wJhQXsCiQPESOTNYqbLGrjbZPy1tBCnzfhSSn6nj32x59le2Zej44s/2a7l2rK7ydDMvM
zzG9A3WFGJ0tky1ijjbz2+pWy0RP0LJL44OmE2YCcPgpGIGuqD+a7kXZyxaMp7Zea17cOwYJRvpv
F8SW3HrhHGr8DC7XW04DAkekO5dxaL2hMiccQ+bCkSd4xfI6gtbASR7DVKx9h0UuBVMSxbqILSF+
MgnHhr9eP2SBJgyA1HRq2pObJsiSyodZEtRw3RZaLHsnuQ+M1F45i6fvQGtYw3h6puzIAXpdS4x4
YIjCSNCDCBDJdN4q2Y5wvqWvB+9IelKnOxAYwW7HfDBivbzl9FP9ce2q97wY4mon81gZoi3tpDgh
wPMvypQstgJU1npI8J8LBVstOV+NDeJXQt48gk4SdC+mhScPDepPz9BmO5S+8zfC+2XNdYjn0v8m
ziHJmq/rGQU2W2eAB59maBEw7HhrSvdcz1Vnqli+gjm1wW4HyVU6+RDGWyF9aHgC0Ql7L4c1Ib4s
AFl9xiCu5orhCb5P+W8kPg3NYLoq+qXtybmSj1N30K82CRBqmhGZMHtCEY4lFAzvTo4ld9TXVhlo
oBzVG3roi9YUsCHtNzCA11+MH4AiiaRhEFACOEER0wld3xpYmVfU1bdmeFHTvqrQIJPrDMnUZ3Ee
WH0AEdWBYLhLXMNhADDIc0AuPPKUZY9KVPqFnufQhL0h5B4Umepu4NQxyHuJ5pfUpkK/O9lnD2I8
e0WXScfoZSxHRSLjgMYv9Rv8uWRF/DZqOZM/fRxGUWUOWFKlPvBrrF3jTPnVm30LcHUktAbgbGuo
kiHsQ7kKDaF6f+u0a9E+gmPdM0ecVWnFmEhkjVQ6SK6xEqtRpyX8OQxdKtC39MKP9F31XMul7m1f
wQre0TenuqItxANzx+LgBvRQWI4ykToRoLF8cUetteaKARwzEXUJeWycKaTZSKdtTXfstgPXPEjM
k9iP1RokBIQ04KXlzACbF85nLA+ULrFy2hk04ojqUFnfSaF5x+upiMubOFD+7NSIOCjkA7ikTWwC
zJ8xdmQWGfs0s3gfnPCKfBWKG9Ba/qKI920Dy0qOB6hUYY1JImb1BIWkl3Eh7XGTRYjYtsmsD7WT
5QfmGYCgGeBAxa/9bTaUP7NINyIsk3FDhDQyNDatm/3PcduAUv2KwnH70gNtIr9bgcBXVzyI4kHF
sWyjXVk3nMyAH3AtZqJFhl57pOAdwiJkiKOowvzlBZ+qFBVS/sR3cqWZxyXKm5lff+kI5fhM/fWt
tp7Iz/eLHve04ri5ko6vGPuK+0Ggw5C0wqn818SHCm7y4wbPS1PyGi0zg7gcb6wFnqU0djE2LoQ2
bHjEv1xJXUZotB4nH4eDG6sBQYkxYy9gAYgGAUMXMfAXMEyzbwjtrqIQkNIGvQKo+hYGKK4cb3d/
UXtgMkbMoMo713523D8t0aWrrmnqQ0AbIrYoyMhcDs8o3wWeSWoUdghs9uetw8XgdgYnTYEnwCjX
eoApmM/O/eYExH2Vz/awWYoTT5bdRbnNB2JuAArGDnO1aATDHFcTGTG9BbQQZVT+ox7Jc8KAA3wo
YrQfo4Q/9BbOrpem88kLbfRpBE//dF3+xZDOLtq27ai1JRll2UF9nCTW6DlzwTfLYHtIdnaevGWF
f7kMY/huADmqJhA689/5PJvtan2Upasr2sVFmnLvQD3dtopPZsXEVsX8TZ/lS6cC/Vm35LEQCJbm
wW6nys14r7d7bOod1RghWrwFK0tA8H3el+mNqoKrafRfAmeO6ztX6zIh94uQ4/zpJAaN6RmlCwmD
oHJR1E9rR1KjbHv1GO8QvWKsp+vYaRWRCiAVKPm0DXPTa/nX07jmGyP4aiQbEM4y+hv8XJ6AFBIb
AQiBDwL2y0NZ1s3N/EyyAmAkVqAXJyz+MRfEdetHYgcSTVIYaLey95vr3KbBGyFPF/HQGqBCZj5c
4oVnsnXLt6RKs1rC76mlneTMH5I0FhUNI+4z3v6kpCPo97wENi9f+zUyydxxC6PFPnVgk9C8UJNj
1gMJr5jVa/3MJ9tOjB+LM5GjZArcC6u0wsD046gdb7xuvHRodA4X3N9+GM9VZAgA4P8xHer4x+z1
btb2sPohfljcf+OrCkUaaI9Sau1JSHAQK1MFlCbHmTHTSwJciKhem5huow6w1AnMa6MDspOC5Llm
RS4VT4tdO+r/aRYCy+qaowSswj5tFEr9nvFdc6mstwQCpLFQAWV6FtyHb8bjwt6y7EmgV21xABu3
yC/ovWPt0tYkOgtf2uGi96COjXkna+XW5CejjuTLHiWI6j1gOpjh0NVrrN9JLkU5tSJwqWmyUJOY
SIBn8enXMc8Dk0q8o3PN1BFZMgxHfaRytpJawOk2AYfnV9w4lBcH8jglbhJX92nO5AW5hnci5TXf
SYtuQ4efE/ApaGNqrLUfMGLC4Pdu9qLoDpDgU9426dUQrn3URqe2ktKWuNXcyXEGmG6IVIHAy1e9
s9FeOX6DFtAw94+76LsNqtRmE5epRf3lT+dQNBubBnRoWWM+r1GzURcgFyjXaPBiiFtTsHLWBbQZ
Q3tdesBg6TL2mArx36pFxCHl2r1c74XAejD78Mj1aGfEa01bwezjboLuOPoUHKvGrclCuqZMXbFh
mENyX6ndbQ29VnO8sGKHPNayvnQb/6S+TXIjDKhsezHp7OWqnWdDWULvMTCWiuA6rEHK7hLc1Alc
NZao6jlt8wJkqv4kot7Fnpgl1vgxVC9Ti9ibGIe2x5Lxi01zWLZ8e7SzEIKJpheAX8AHj15ty+7g
GZsz3OTgvSOLA3BMqN7OvsOcKoEIKKKCERP8TediXJapsTbUTqsnDv1eONMaQwB8Sk980tkPVO9S
JycMVAXfBfpV7rvt7kXBrziyVWzL0csr4pl9sB0VilxdRYhOvR/g8B0QE6YmHsENwJz88z/iW2MU
WdYaBsqhN3Db8AfuqL0xQ4kjVqhn2oEtwbhBOF55yooATossc01+UJl4wpuGZLW4w4DCCddNMzEY
SIY0nj3fAwn6SAlDgL4iOSU7mEyi0i7CzSQtlefAe2I5N+gxAmv3IExUPfzn9KndcrDbC25Wf/Qs
prPFKX1Y/uXv1p7r8t6Rb6RNvx8uJBB5OtM5ZPf5FJambD3w1+dVY4qNnGXuaRsC9sk45ldQXZAp
/hIZ8jWc+Qr1dmXBW7hUjOoI3jyBZWrOy5ATE+dt+2bMn71Zn8DzMWt/UHvoS5fS6MFHdZoz51Hg
5IOO3nb9vDwcjAYHIk+kQ5CDH4cFfOgaGLsUxzQX2npD5VYf2YTWuoF8oKuPKDPw5A9BDkdx+Lq0
V0HcWwdukwn0PrkoXbrkR6YdWEFnPQ+P2EyU9onkI+5Jl7NgpJx5V8JishX5rCZlSDMdNy0vq+0c
eS2K5ghyPo4woKNh6MtRwMtOJFRpWhzynAKgPBMR8RtwhjviTLqp72g4giDqVDMb3WYfJX8IOLK+
lqfx+yGWo2Jd8fbYq+scjSMyrTqFpyH2TnVsnd2CStfE9kjcuYmQ971fe1WDjZGvqYQIxQIQ8ewp
Gpi2LvTvt4W3HEWRX8IXKDK0PFA/JfP+wrwJcJZ/PcSy32oWa7rG2ITWcVFO2xGxo0Q52uUHvrr8
8xkBhANouSonS8Z/lNqafmEdoZJJXcEUqjZ1O9eKszutCV66WMW6QPcSnFthgZ9DSFU1ZrhyTm9K
qPFP8nIb6kqm4DGIu4A+r1dKGBSQzScpovfmiwNRwtgm8jLz0iO0Ue4uf2ph0E7ZCUzhVY+91k0q
kHI0RHIE00PG3XkO4tSuHBDMeT2hgFdyEjCutjhllhXY8hYABiX57KQU6qzPtM4cmrNP1dvfMWJQ
Nd2thTSiaTrYXw9H4xOvK//8y5DrrVmnBfIQcPKbY3tXmG0+vikg4NJpdI8qiyxXVxZ3ArGChWrR
8X1aEQ+POYM3jJdB34OZt0BTGg2JhdYaOUUyl3EDw80IUheTuzupL7gGvQFy5yKubFPhzJTjTi75
QSxxtLmQaEZpM+NkoDkrvAB0ahgeLTHZeGnTp9125TUKqclZf7sukLeDupGuNP4cOYQEAvw5P2fr
IZ6vXFJwEPorTn7bBCP/e/dZlMfsF12JDc9E4RxeCBH5mZLxlnRITY+M3DeZWJ/hB0ZsC0wavwtT
hDi0ld4uPWw/qCTfKpbA8PK2CidgOwIgvQ/TF7FmTqbFpTz0isPavwjIPjWXBZGVZS6ztXIMF4iq
EklHiduD2Ij5gLqx5NwQoTNgOK4pf4nLw6ecFXxd2EkIIDNwIbe9kLq7oZK8t7hCmtJ0mC7L5o2Q
ZHVfSFKvL1pXmLSp8bBtGh3Dbr3YXIqlNIJA3XuwhLdLKJv+Lp7PxziZUgpQy00YxuPW86UUlVYs
8yRhXcElUJB6lZar33wNUDv0WN1NnY5E0e3ec4nBSwjyBIIi4SEAW284S3dUV+HkTZke4ni/SwZ5
0829sdy7hYOd5uHSHGdc0eiTSZ2vhOWi1OvnLpsQ/aQ4kD86Mbl1LxOpTUguwwGl9sQTXskRT+g6
wNIL//AkFX/5g8Uipxv8a37IN2MfggI6DKLmH9/eAVpAbV38/rMdZhCsruqnrYG/K9wbazfddZfP
if3Zr2eUG7p1YMaVA6exDnE4uDMrKnxfM26EfghIPhxStfWsWX0IvU3WgJV0QTVtXdhxhORzUbqH
1jsq8fFBDLAhWl9asDjyuWo+6H3HQGABT1s1KC/we8DEkLUCNZWs6Pd7jKaessydr65C7N3g0sh0
wTqQ4qwFw0JcNasOJz6QLUhnvkKpMr7AK2zA2Nubf3DYeD/OH/bGhwBd0qZrlrWGsRWYyo8LL+Th
NT2LqBrRB6UDp4Q3Zxod2WtfGV2SU9xwT/6NWuTdi8ExYzLDm8N2LkuBhqCLN1AruX6gdW+1eApu
536z05Ho9v2y7ctsS4/rMdszn+c+bHHf5LHPt+bw+OlhQkjH9EyqiC3AqqsfV/EwGWYANViJUPb8
XvpPF3WAIa8tGdYlkeY4cil5kMtFNAWeTIWI/xc0Y0OO4scMPmTRro9IDp5kJKWBL9lXDpzRbmQl
elkxGQvCIuNUFgTaR8SSxuDdN8Hd8TfqHTeCRa41Pbc8MYVkCQiX2jUvnJXnWR6u1BwV5SGHajlE
Mvz+n8wBButeysgxsjBKYDNx50YWT5gW9MYF1X6rdaDw4UO+LDQ4u0S+SGH9I/P8ejrxLbb81GVA
HRyzDGWGEVyT00XG7mlvudSOmQWfSS9YonAuvklE6GQcbY19Hr5ZEuiPNbjpeJmtKZemVzAVRVM1
ngJwY2OaQztDcvWqLk4gfP1uQcUXCpg3aQo5nWtT9CKu0PerVFF+3FDDO4M97/H3AxUConcW/EVb
ija9TxFJgjZ2FenFUWMdnGqNdo5c5KteYfkMoWdJly56X3XGkRI6gtP+C6aHeuhK6IEfkjebG8Wf
5kWR3/lnm/16BBacJE1s6G2g5mxxCdAkCuV6P841jPs0M9YXBo+PFb0MT/8/BLCLejy3IomWxZOT
90QHT3zm/btDkqJJ77oaPhG5XTZ5GofXwLVkPOXKvI83mZpeVYsSmilI8SHjmlQiGpfmDIgksqRy
p4mxhv+auG3nfh38N1PS7C5H4h2VUGjrVYv92vUIjaiR+u+Yep586lKyem6MbxyiogC/EhGoxmZS
8Uo06LqUB+s3kwf2pSGQYhRB+U6MDEhhj4hd3F8xmiU+trfvCl7y8+8KWLbsPpmwmmeVt47c83GQ
EH/TBGnmLnT6nMPZyoElMAQ2I2SbXkq/KQ/UTYlncFl0GPYyQqCCDpTtnT0kPE2DNkOnMs/7myCY
1SVzRzGseRRZ7CQmA+ydXRWw80zFou+0YpckzpJ+wgBDxRPiZOrYeeNnEX/a88Ktjmm54CePen2u
6uaytiWgQ56tGhBqeMD/oq1MDix06P5hxmw0KHuQBi31eY6evfieX8u1UHaep1B6pyiMSQJKgWDK
64OsprKXmKm1CxAz5vH/6NUfaVZxjXKpe6QUH7hD/K91KmHMLiSQWAiR55OQkXRuALSCxAyCkHCF
VsMEq0KqT5yoiGytg33ckTph57Cr0hp0JbsRnefTVS8v8H4223CHJMHSAOoqED1u8svY1qazx6gM
m/Wi0+Nwzp/XxNmn8JEuC/L2vwo1WvXKW8TqRUW0RsQOnAvgrsi7LL1XBOSYXMlBXj1c/pF7ij21
IO6gAE5FLoPzJfjTTzeBpAOvMUbBruxXAkIgm3vr8O8REH7v3Yl50LW+T5yntiyBxhbhM3lXfPnN
wjE7tQh/rUCA7NFLfsTcDQzCO2Y097sZ8YYve398t7RxH987xWZXHi+C9B9owSwfwTBsdHfVkO6H
cStCNlksoai4qJqnqbYuph6WdVe9GYzEd4Avj0c4wB72+O8zveuqR1iss8EtGjNBOI1ba5eIr0RP
7LCnYTE55UoifkzRIAzqMVNS4NoPnOs3fxynfMWHBa7Gl13FtSMn7OybzKZYxTkKbfRY9kWPpbSQ
amk9uBKE2OhWw6H2jZAzDjjHU2yDFqRPUr23+UL1LXTk8/P2es29Fq2IRlARdaW12dRN/kBpdBUb
0rrPXLLr3ozNyYH9JH9XdfvKVuoAiMhmJM6X4/F1L7FKuwEVWsWP/WDSC/J3g2Jgw2gD1F3KFsl7
JeU83pFYek1yP2nG7+kuwvmkdOqA4GIXWte7WpC8WtXkfTMI7y3dAFIA2olbsL2w0nYtQCxlGyoz
XY2RS6d72YpcIKwTPfACZoyUstYU48Sjrs6wGgcj1e1xvM2K1RsNtHMmNeH2avoZ2PrcDFehf/rP
phE4+mFljhc178bPYqshrToT4QVo0Sme9x+KU0CYpHEzSA9xnsjcVIm0WOkcJmckr37cnYpkjw+c
wrvyE0QbJWEAkPF3Y/itSgjL9GDEltS+b5kt2EGbENy8lYLTufqbw6FkCkmvUbYKKzFRIaOUpMHq
1WHC2iwyAhUI9IMiFDilNqUbgVfylmPOxeZQkDgxNXsaluhNC1MdX+NrNQDqq2Eo3iRCdLV44Dtm
wvbJx/KHtHXWexhASGNf+Fp8bf6isDeX3DPE5kO7YAQcFuqHCfevaYcaAj0+oOJnjIQbcW0V3EFx
+1tmR9++kyb6+IECFLgDSXqvbkLOiJmu2vxA+FfR3PLjHgPII3WU3YkirUrn5cj56uXTT+hkMtnb
UV6cP9Jz6WPZ+c7DO41ktC0RmxYc17pUIBeWKM5M0d+vK8SMaNkRa6xVQykL6JLfoz9A4tfP5k1Y
aB/27uNXt9JI7J1aolITBiWJ5rrv9UqsMyDEETx2haRmizcNAqEjS2Ffvjvb313BGFgbS3SLV8Gn
jjxKwBE7lQCNdCTtU/eA+vUuPgL+edAjyuPRVJQooLJfClvOeFsYnGl+utPRCi2SOIaYBnKVxiyZ
ZEcNcHQr+YLZPWW46GELonundzgBo8KCumCKaxwpWQxX7KaeSDd6BVTWphFEgSCX9zQ3DNdbcQSC
u0MZu9mlDNvbzyCgBCGMLamPudaMg1G9kfFZBR9RXfDtbee5DpM7P73RbryRozzHfpgy8jk5iyHx
xtueJm8uQAE4AFKAVqLjb5hu0q5fPeoC5j9iEGw8eCY7kFAl/I/pc8SK2Mv0SGNUfCRsq5mKFdmG
f4uhuPMpwoA3sv2AScEX/lHRTM2+XBRCc/sWlc9KmbIikr500qBLapmKGnogh+fSrcGS8Orx0Uqs
4xQILlb0SlbGk1TK9EF9X3HTZ9ynxdzoG3XxDRrRErepMVnchRCmkp0mXHBuCjCexkJO2OpinryU
wWIJkBY9BlSzgKRgDszQpVJMBverrLib+PHAckW4oFxW9lJRFAGo5AAOYeVBd2nw8xwc09tth1IL
1Pu4xW1L7uJNJCer2SsPp4AVlKkAZcq+dINmcdNW4BO/WUmQXmNhvnKRRuusRU0r5QXSQfnLsuMJ
CR0ijbJmRsJgbkwqtLLHzWRAM1rBxXGK8wbodgbbRtRrRUsyh1zeG9b9SWiouWOsotGZE/dF5ZP1
VoakgMLt5a5Vad8LROXRCRNZ7/EcFXjGZJU1aMGnqXWtduZOSfAkIsgaickvY6SffsSgz/CC6iOM
iZQ0RBCAwZmUdThoyp9e/eC27hjAtJdjOuqOfTFT+XwbwSBB47q1zn/T9yAcH/FlLXEcXWS1emLa
oG6447GtsJIn6QfyhiCiJjcNz/WyaTiIb9bXzJx2Nf0NdWVDThIcE4p2ztJW2RHLsJHth2flu2r7
eXu+muvd02FonhmjHGHbdBpXGg5QRzqJE2CXz821Sd02RVl29a4vG9rPjJpm3KgkLUfcbJZqqQGw
p3lFj+PWKur2VVQx2pbam3kv1wayR6AC9NrwL1wescy4cT9j9gKlfop6U+rcu3mFhInwWZmpbZ/Z
DmpaABuFpHaCVzc87dNz9n0e9dhC5ePsvRxKHn5oiCuClDPvRK/HxWzJ2KoMHj+x88BZskWSoD2B
LDTokkV9gNDv1vjGOKACMLdFxIFmNe35a2/oR17M3GstMUVGT4HS4hBGcxfWCN4Bk/2LV+nzzeU0
vq9lIk1yiBP24tnnpWXw5sKHvOrOmI94L3L0RFGI28rPGYCDzAKx8Vhv5qDGI/ov3TRyzouys+xj
AQHfWSbly+ZxCxY+Mp9CQUyQuv81wE4A1+/36VQmkd7t7Ib3uubDytR5vI79XOmZ5kOdICWXhLTv
LXN4psubry8Ngd6Kegybh5HT+3EZ2Ww1jy4L9W6CMC1wRyMYIzhlBL4pvyxmeCBas5PsX/V6qM0s
qZ/b/C1iSvm3MPNffr+CUNsrZ1J13OZ07eWbmqnDO/yKI5F2WXlj5PFbdAGMJhpTQyM7PkVaNDfq
ih6uzsIHckzU9ohvd1E2RhDs4CxaTm+8Gatg//W5uL2up7enRIKk8ieBk2fsOA24c9FeN2uJLyz2
9XA1IHNISg+THGUPh0TT1qjtByTw2q9ipCCaaRYWNrX0+U8CslLJ3MtF2Y/oqmGiRG6mFcUMxAfm
qZ+5f8JJGmG//Jm7U9oJpAn2y64cYATu41nAU3br5zrCWVBwrKr21799vVi5Ic7aB+X1ywJ55ao2
bohFzml2lHOmRNZgWWtWLlQrpjoXTRynzEVCAruB7v/Q/uTDlga8tj012DiOdLpUeYVCR/q7J/Jk
N55ikjZNMNEPIqAYf7MeDbcJnX9B1ezmY27cDkAdtwBQoeLpKXOD4lrweDWcvgHc2SFT7NsjXyZN
bKkpHFJTFNo4RfMtDQYLbK5kFsKw+xytF++nTWF5e5kU44EIz+9GsBM/li3lNjdfyCY5/VuLPYne
vsRcLcmr19WZdzzFOGZnLdvP9koKqLaReh2NwPbMOHZs8UNOpWXJb6Lbmj7oBs5Dm7VOlfZ/iCu9
A4awrKuLrDMQXqdvjyAxWnJ35LatN7sUDxpLibegmqO4NTQmZ/Jd/Vu5/Gp71xx5tygvrBXr5b9c
JgTLX3NLzHEhEPtAAXQgCVHJJbvpazDNUVsbk5pD9bo5C1zOGKGgJrAATrrotq1wvhw6tJyu9Hx/
DRmYARxHejW0jn5jpE6KpyMLUMdvb0GBfpIJMoSUYwnHUwhtAzAU4BiiJViwAhlqkVyH4JmF5eDA
n+l5ZtjMsDWMGtPW85G6Iai5HcU3J0gBJiJHxcu/9eQp+He6dMYFnWDaU4HPkXscDrPPkPMPzivz
RJpJMGwzotOwUzxvptkYnPLGrE+uczldGpBtbhXTtXGpLOJ+rVsCkQriBAT+7/Tzs2x0W7lDFZT1
+Ik3eL4VbE2nc3qTb62KlfDqxmP+xXOXurl8nkDxp2bNyKkEFdy8btgU5ntRGmLu0twMhSB1r+Iy
4q4d96hotmIdrIl6RaPzkGCu3Fg412NldY8c5y6GLiMCthTJPdTwcY3UhC+zEq7qe6y/1mDdw9+n
U3lHk6EJ+RxS8fSdq6l/5AM9gJZFOjHUx+URCzuLJPCKCwQ7dPzHnMMGWfTvOA+N299ooLqezcml
KNCwGWRXn1kmafVVHzSOWxze/0IbowmT+d23NfZc4xZBaKjLSGRx51Iq/hphXbfMaQdvkbMq4H8O
zuQ59oxtDcCO2IsF8/DbHGYfJ7WEuH6e12eaK0oGZcOwi52LOTznMbVOZGhydMrmVOP7hSMWHh7a
mAYh6r16uC/YX2ZGhDLlW90PVDuEATLJrHfAwQg0mYEbB9VzGJnpYVlZ2Z6wUHQV9JYRDWRifvD3
kQ7pzvai92b+zTslDDYEyx1Ul5WhWLYrgGzy8AyZzkDg4nlrGKyjH1AXdfVyw8jT95r/yhVwkien
VviTEyhvRO9LRRBQElGX9WNUfjfWAMGc0Hc93EklmIGocU0+Vj3nz91Dt02ExRJxMGmp08s4pEet
xAh1/buIEaw3xEe2qWP5xsUVG0vjLedBDxhBesN9P+jK6x89BYODXT+rrNyqKjLF87TYSxTP4AJk
FbWFSxY/Kx5dDDpmxpLWj7vQKTixqyGog6L5Say2TLNKzKm/fqZzhnhO3ARZf/hLGKNHMXBrhhzS
O6wyRXiyXt3hyl0SIrm6gz1GAChdSboBmWUYYIKaC1lCUJgDvQ01kaKkNgK9x57yeb5xv0/Fz2ir
qliSj+A/D19fCRY5Fy/pmiXkOBVuKuMuD3y+bPZ1xDf7gwjoNsK6eSzrjfJ/ZvezihSKntp9J+1E
/a9OFg+cnynUIfMk+yJiy7QVvrIUQOEPWkOe1ms+dCCVui0L3W2zRBr+aKvVME0HUr0ATOEH2EJq
uigmXiwxKT88mCbE7s327dgrwQDGKhvDdB/Sg/cA+0RneP4Khnlx6sh0+3W46TXNGsebDI6gFkRO
WVJ83LDDwfbE0meeLp8ij6o5Skre4Tm/86pURq6jydXPRs2ST8n2fP0nVaGDEekSASPhLqrjTnCT
yNLTmJo3WrIgSTLpzUnu7dKLkX5KUnNif7MDUGe5FFouAxX2TlUzREi1AfY1lIm/vcKluPcyaQIt
ggqVYMfbGlG8WVzemvcCbP0B5PNdbmVeizi3QZjuCuG43CVIakIiKJIUvt0i4cDdP4VZOBQMZ9MP
F5i0EwyQEWb5guTSRYnDPzz9C2wJjcUygQMEXH3NhhKwg15aXlqq+jDYpEdn48W9TPCDHV2m7eH+
1uBbsvHNtdM9/glEw/5b/NKrUlzuRZQeEra3tuu49RmEydH8bHrWidDfFT/j2fP8NbMkkFCKuy79
ZAx+FM67PYwRSi3zTI2v7JcsDbUqhAg2G7jqNeYExt131V7eZ8LZ2hmPayAGkd01kqWNSkB+Si5V
ubUR83XXotbLaOsyD+SZXhvNoc2gAvmJHnk/uAHdCSdkNyNN4PSobusLw9YUqs/rJ1QDIJeNNqgb
dq0C3ZCyqyE3j8FqXu/fT4ut3R8QnGH6twDuAA5Oc/DnlRSa/uOz528zn8tDjiJ2PLUmIrOXc9yZ
42mcuRkDOZQopXcfXhp/pU1XhmromdX0579e3PDIgpDqPHBWWpsMSt6EnXFLfOZEjrpXs7cgd2l5
73/+OyyoBypybDwdCz08TkfFi01YnYjAVcMRc8HkIQQs9Cn14QNDIspDjXnTJEq3LT665UUx6kAq
WaUHy4eiV/PSQXaQ6O6QsjhVS/iEh1UjJrcmxtqwGQHqLGvNps3YkhgH3d1t2rf9gqj1TWn/Orrb
O5zXRHVRuWssHPtRKzU37ZRgGc7UemrmfWZA4QIQOQtndFh2lL0KdjbVJbDD7Cb1khG5+0/SRFX/
k9vaXh4sbUjPlWYqAjF2KA3sHngzaxTb/94H1gJRq1QRSOf8COe2YXG1ANLP42A6R3VeMCAfLg+j
4T7Rp5PWEjAWyVqtcJLN+bOTxnYmbg22Ey4YEyuQCkkgH1bq6X8bvfwBixdLtggjp+Y+HMpHuoco
pRAH8H/hl1BfhEYBgPdOJKSxhJe4AxsAjbUmS3XS4Rb3nQ1S2rESaqNq8Ww2v0PbeptNtfauMqOs
78lFWG54Bo041oyyujlj2f5tYrCQjdzxY4xlHrX/af+Rl4kM3j+h/CnhZCFiXGj7R6JNz+E8llX+
iB8UDFxBBHq19DW0/tbc1urPA8NoTxvU2s/QvkHXBEYObveXTr9TBmUmyA7J3vMxjj/AjfV+Z5Yo
hGz1xQ5Igeet0y8J3GpoGXQlJoStNdmFDyUjv1LPDVtNtvaK3nJ6GbD6glglT7TuXzODn8FLu4WQ
gYoArCMT+nilYfESpZpHlwqDFpWlL+lhEVEdIkrEUKPmDdeJn3GzPdMix8qZjuJ5aQN8E2qe9Z+S
i2MKFaT0S1OY9OzB1Ao8hctX9XQXVf9lRIcglxVVrRrFuLWfWR/MUtdR5liMa2E0mBp2qB2zhBoP
IHbpFsGQUua6hGqTz+iMIaxcTW5hKm8RnvwKcBjyNv0baqG3VQN9IM1jwlXVbY3lbybLbbJocwGR
PcWv/uq0u/UyLdIa8noq//0CUtF43mz9awuW3L0BJnwiYQvqeKbxTz0WrLW07kl4TfGRlO+JpNwP
s+kPFSTTjjv574Jh9Uts7zKwInTMRPLC75C+toQ9dMeuuxKBmWNt9ob3uS6tBi3KFjMm9p8U85cM
ZjcnM5IVjHoBzkPqlaoCd8BILuXH+JbPtVlBsGzF0AQMGQcsRz2aqY/pY+H4hqn7kavPfQNSQi0G
6lKHDKKiPkl2ZY0zRJpp5zMpJUvf6XDOK5/4Yb9T6bE+wA+x1FfUOqTCFmx8kAcD3nQQuWu61b9X
8RoUQWqNIYAVugVaiG4ReHJma6xQkUV35setga5q3xCxxW9ygbEBdskZGCjkbDn0RyrM7LPYAQMs
WfgKEtpibbsAeVIYTcY0wp4bhLSmdZyYNTOadDhNh7xNcB+pghsrbNPBf2++b2/+4++2UpooIbkR
kNSdf+O0ql4lqAEL3chQyyj1C9lffc5I+s6O4Up9GZZ4cuNbwTsp0giGxByYLsSyb/EUlsCum3lV
xO0NdClKmShPC0evdlLEi8rCXBzFm66tG+bBbwAaM59LdvB6MNq1A64YQH0TXiTDDEzFkEvLgdZW
iJUiILPSzadBDhOP6II4JWT9xFVqX76rG1ZQgc7Or4boYt93jGEvAbRwoktgHJcjaFX2u8MvFmc7
dF7Ru0jrj7PKulCY2Q0CRdn5Bl2msi2x+MsJLb67ADDE29lkxhWpY8RTmnpmPkX4m+7GN+t/pNlV
gnVCqXMpLqcMeoam2zcNHk9mgWql08ZVoG/8/ude0wQMjCvKKP+FlS6gRS/EwHP3Jimb4DJ6rqUw
DmK1NLcFfkljT9coTUEd66aD0uTidc0kUp28FWJGgdz0y1K2vBatpOMSHlELRh2ZU6bXGAuKnVHR
yyZ1u7gEOoPzFi2zzBM+3mHhqbyZayn6YCDZatNeZ3Fz8EExAE54OfURQuHOiOVT62C/2X5RJtAC
F35ah0AOxXCKQDPLSHBsvBjha2LhRiYw0QIn22L/qCB41JKYAi+OKgwN1djskBUoHU9+f5gDQEK5
Q3HSdnMYBW4fp5TS6HhriV1aW+sgpwUSInl1TZAOWde7FdfuW2X97/RbtC4RFes1mFiVTLAroLwu
e7R31SZXtsHPlQYYfMDIFKCA0ipg41uydGn2dWPp//w91+pNJrh46gid46ATInG/LlHR1kjNNU0s
AExivXu9q6+FfXpKS+NWedz4F3JpCAMOKTV38J+GV86A4qXN6jWlkCY0IcdFdLoyfynA/KPvYVUR
v6s2oU8hawWNdE0B6PBvq33jNnrNUhQGrD0XpIMzo/ySefoCN+M2zGrBZZlzN1fUJTK5LK9X8fu8
VMNTmHnGlIbIgcDN70wa/ssmOlhahuzREsZNhauWrZ/0S/5b2mL01e4KXDUgqOGJhiIvf0d6PSUV
g2iyS9xp4CgTVgGBSk1Zg3CSFZ4xgXC0kdj3JNH1NvMec8JSwDhNRilA3ZCXZsV4wOT3KSfkpHq5
oG3oApEuJ4tJ9nf2S6DZh9N9TqjxLLOrWV42plnndmIZ8Ow2MPuilo5QErNVqwu0O7p7abp5pNx1
+ZQNfrPBOAuOAqGnyR8JPlVwbE39taa66HKnfihdiB6P33QiZv+pS4rDWiuM9wwmHYGsVIEXGYX5
V35cvMNrlMe1JPRVR+9ZPtQMCAfI2S3kQJa31vavpr3CiPYQUWQRHPCrlX1ceqGKTOUVLsKB0jDD
IJHIGh8JcGzbKogwl3GLOEh+8w5YZXM5wh9EqPLOvrWx6yCCMtdKLFY2c7iLb0lH1toKz9foqP0x
E3Eg/BbdID3TCZQWbMdRhWqg5mNJVBdIQYVbeiczOHBp49uQ98haOiik/a7SGblvoTqri+wgsD0v
/O4XCR559IAYZ8r77iDuwwkw5+1t7FmniVAQ2OtRKNL7y+5dx8qWf0zZ2JSZ6Ba28XDBFq/jOTtU
r3PtOF6BMNocIp7xxdPXPxkwppptNh7BPdrwjM1fXJPeD3MJaQCfuOZusMgf1u73qymgfMpgS3yX
nEHNHj2tDSEzduZe6o302vaMDURkvjUZIzkdEttFeUkA3i50FW5pudgxyGirTHaxYGPDzbiXDp+k
AgI6kSb6RFkNrlc45dKQmCYIh3AWtIG/GwSQoMJjzqVV35xdkUn4D4Kq3z5OF9udZdvXJsuDsaZN
69bMrYlINujH66pnmMfwPUCHCrcUIg7yYp4Vy/TKPjc7itCpowDsk/Irs+ORKhUQ1g6+/pe7LCY2
tTB4nPbWDmMg7/I1UDfpTcTpC9VZOkQAoSqlTlag2P35XcOHjGS2N3OwuOURNgva+aUGp648M/D1
JPFAytBd1ARTCXj1TdlkKjYyNSxoVTRNXbh2xZ5YhWT6y8YcaEDj29mgyt4EB7cjiUewlTeIejk1
CP/QeJTPKLqb1QIUIclr55d7416YjTmR6iv5RLe/sYq6IoWS9sR+WOqG2m7E8tz3w9bQxyUebrr6
dOBsazjywB0bYwFLeL7HuB74tj0SlCk6yTL+jt8uvKhFB0c5eN6ePaez4wPe/POhzO2ing2P7jZg
pXh2cx67I5u5/7YkwwLL9Wx6zSAHlv0LROMm81Ucb1JTSh7Fki5MVm99M7x6UxbLa1qzWKUZPfFC
UwSA/KMagwvbxgDA2rpvhbP/GiTIpq7KfdZHCUKpVuEE5QQCCO4zml1JozZ5AywCxj4fakSvKWIs
ZhjmGYEovwRm/ar6jmFZT7oEX7ukJAcKVxvFKFR+6v0oQHuxe0xQyLmUQN8RvApDxVNuLEqRbvpR
LyeWEXXyZKV90rslc7I9V8uPLUf40G47votkaBPe6pmNCeIC2yVP2vmvg3na3neuViKFC1XFA3uw
D3Gem2NKa6E5bNiW7ecsfjYAEt4lKmuh2XRf4SABr20Kg2csbRAeFpzjrvGg2AZEN4dv/FyYtkQL
IQkPdPLaoagizlb/EfuZ3GQhVRYioAO27JHcW8bdHOKRatTCE+Ycvcg/y8aI/dSlKzmoOa1Irei7
nf1YvoU+4liH5m6oFe0Jow2VuTDxV/4Qc550Z27+fDDr93laBf/XiYhNFkllcXl/nx0475yp9sWw
uBhr4abw8mg/0MQx3lqVG0I9n4WfcpObUs0wXByz3jft2hYrsIq1oyuU2hF0kv93pEykXOyp1YVf
nCNQW/21Z2LTH8LakbhNquyT+ztgH22f9CpuultWfFeRgJb8aG1icEXD0dW3GDPtKcyZrIDl8I25
MNtltM2ZytKvdaLXd7OsbvLrOOZCjcpe3jnwtl8AZBjm9cFMkIo0EiOvLwQ7q06Pg+jCS8h52vyr
nQ9ENTWQDnNYUexNCrIHJyGwoyuHHRyM5wBGT4e2hUvlBjQC1+FofEcns4pef71FnGsFPOBVIE83
EyQUHT0MRB+6Q2NJoqK5Ete1ZkWCumoP3eIvKvnksRrU6JsMlUtPyB4oABCnRCEdzsSIoDzUf4pR
WIs3JLbVzHkO4a+Tooa192TKd3WLsKp2hSfB9QchT7U7Gwr5YzleESNRFXuStNpGKcZsj48eQzsa
VgZNlWnr5wwyMW2DxLF+mwAgzvVWD+eytPtHtmxOqQN72gJPBM26Ar99OK8hB2ltlQcFGgltwqR+
/XmIlt06BcvufT1TnL35KvDNJ+hGrzo7ZWPcee+9KaEWs96w5t4Lw/ZmvXVi8A0yqajM3d5GYnTo
RIPFAjeBE9v/kMcFYTogO242yJi70PFCZV5AaGp0Vkgw/yVuy0g2yqh464PAmfmZSM2RtpSBAfPn
i+sWofHcDkeFTEkCraFBYcqXcjYMpNN1E7TK2FDFvUWw/knosXQwJM79Rai+Z62IbBIeCCSglBZD
6E6k2knPp1qj1f18LoV9MaAQtx4ME3AnXbtP9v7MXQlew1+06pGTxtHc5pNl0+TRk+SR54WldcvR
hTyuWfeY6S25Iz0sVf5qvdmRBVvX1oAcIUWf0HAOqEtuGWI7ic4gGBHLiz8T6b+UitqiUOG80LFB
J5OhxuTVeA9ihrxbOkd4q2+loKMDR2fwlANAaEXsxpLkxi4rp8BFXzN1A01aD7F+mOVY2HrtCVAJ
RJBfvVA9c8SdU8zVLp2naiR4laAOGVGsgLRt93p/Pxv9A+lkTnvIZ/kTeFxKG/ENV+A2DtT+Wbcl
zNX6Qfu9IgPnJ8SFHmqGZ+MrwcEkkqKpkWX3bxhyImOG43ZFcfm52IRNKGYJgXpa3HylJ79+Xf5b
yy7d/IJixFhfGk9SOAKFNVVi4KKdpMkHGjE+kgiDPriMyt0+laQrN3fY8APLxjp1zxtedpz7U0BQ
TAsVtEVeme8ZRkRgc9Fg2MoWEd/SzC6mw/nXLuM7MICtIHuwNCp4JmvgLI9bde45NoyoCC/Htmnb
E50Y9kWIBn/sWl0lNzDLpQKne3QuRfsiTNkKzEwiw4BzpA3jpV+aSnejReWG30DL1hSWrjscCA4p
WXlPW6wirEbETyt9ivtUN5cZAAHJ8+V7oJdSPkPdSCyG0SVDu9uf4lCT6PYApvai3TqryF2WZcQ8
qvcpv4Yd+NT9kXGodE+WABUiFshWpPokmZHBLdwu/6k1dOg4NZxR8NHmV9IB8VWsI7sCIH5PtTpQ
G3j/xCcXHzMdYpcwnkzLgt7mrybq+d6lM61lF03HuaHwtntIaz3beP3bZMAGG0MNnq/4U3Bk0XKM
yc+FUfz4yGXVt3MA13Gg4ZI3a65QmOeEX/XwLhroI+BwBVBqvCW8weyLDzHe8g76lcN9awkY7ACd
B6P/6y9t8cPpAmUi6XLPDvb7NU2Fe8YfD0BCxLS2CqdFtKgqtWTuP5eDO3W/p4boUmKspLc9KCj+
dMly0ne5FZBvOj2kuDqhvIGQHAfI4V9DLg05oluFVIkJsGN6CQlOvO/l6BXwLX+b/KMWcdzyyv2H
+AMSlMFVIfMhVBEM3tgsLmQONRqYOQ3kH7cjSEyyO+/pP9Xkxnj5PJbxCfGMgZwq6XUl3ZISPcAj
VplVjRjo0j64nkA6OZTqMWi/ustpZJCFxxsqFmAFLfIclEf6Umb4UY52yjcepSL7HesAR6Mjsw52
yzd5YN+l7X6AMCvUXxi9PUcE/4Ieo5K7AHbGGamgaYvKIuAVi/IcM6tkvd3dYpU5eVMTRPU7e+Xa
ltKIcDBOozsR6bbSkEQB5iy2gKTawXogntom2EOtAN23a8SAlEN3/Iu7E1Cl8f2c0BmBw44PQYjR
lZlWDGMgs48r6xRumTRsyRGTPdNYJqh+bh756Bsj4C1QN+G/qO4pH1Dvub474ywxCajR7Q+0Ytkp
oYG+Cmn2JLCiFH9u2lzxX6khT11tMH5YnO19ZyS34/xrjccN9GfUcyR7DPJUfI1wH2kkvfQS3jEj
Gqzc5oII3XrkfKYK1ENjM/+MROGVgEA4u5wEDeToqcKgkj1679VccU52oYMWCC3fOv+kTZqr/CQJ
dNOK4gwYidXvWLR2yQijm4kXej7z3F4NxeXJnbGBZyyVa/nhWMsOvWC4F9hw4Swoq2s7jgLHD7KH
nV3hSXwCw8kG+SRAO434em7iEdXVKS4MGI7eSWYkxcGqKSJIQjIszWm08tkzPpf6lWIZd1i/EDZn
u4HOgJU3F/T1A6Y4PxC/UNBLSQZlXWmBMDTZC3DrKAIYxiI6EwqAYZYXOtOuL1TjZlQfviayKb7+
0kbLJoPgBylVaYkf5bem8kwfMbJq7MT6b7kq7LxwCSvtA0yMry/paDt7PFo2EnEuEuPmLxLyHojo
8ofkYuEhpy0zKBmLFowKxbBfdmCiIdOZApAvsOCnC3HawRJnxu5bkZlfqUJkGhYJlEJMIVJ5AyP+
JdJoRnBNAu+4PYChlW8W1GtuBv+7RNcFb2VkGo9+fFjtEUV0qgNdTjO5VzHZdjBTdIvhZ9Gp64Ma
qx4tssMD2ibvcZQW/AISh4TDr2GUmbxoucSMPtc1GkFsQ5CMhUVxmKTb/NkGFy1N80oXBUDdpMfe
+vf9C4WlY8j4p8MlN9aG0qOB0HRRb4OsyYPMfBDWvlAyh4mrpq8NKDQJmCUWZdvIWUN9TWS7mAFc
gHpZrn4GDhfBXBPKKp3RxJKhCJjFASC7pAoXYhbS2QS2L/+mh+nooQOt/9y1pzhkZjO0FoqcYFa/
WFX+m9tbYrLmxBbcz/vgniZ0mLiUspXD4MgrB0qoQYLDf8vbHUrSUJST7/FrkLn1eSljCQm6hI72
1/5jk2mg09KPQXYP6jBgYw2rqOLxFgX3JFEevMFmBZGKQAooNsAlwklV5sawrRKncdZ7Y4sFo0s/
+ZsYHS6v1eRnMV+8+bwzSwxBGa98xYrsb4LPcSMLaVyYTqPyP1l8mjTo7q+GtUYWBRIYrpF50hmn
26zWek4y9BupyH8GHPGqlOiLaVem61IK7EihbGWlcCa545FqgbHNHL/r3G2x5hn/oNfz+LiYb89G
TMypOX7dqDDqE14yBNfshrFuWBbf2xZTWZQgC+JboSKxvDEjMMHaLbvdQUz3N3LexCkzUK8I5Cvi
KxAplld9ZcP44uMapLw7EpMMpqnKAL7lP4btqHXz9aX41PNNL2uZSleSIIQYQj+GWEmdetkJ1rmw
/xM0Oar5iJwVuDvEWe7k+MoSsxGKrTz/OmgqgCRTcWrAKndiqtQZATJd7jAT5009jAxkPRwNM3JC
RlQaBr7MNLBuTWTHm2nbm4NoxBmFK7cHRNw16TS6Lb7xPKxqeh6MQo6Fy4L503CaqP0BSxCiTKhC
tZDd1md7i1Fh/9sEmUEYt1tbWNK2DGDHU30/FXFNjZE7xUCaEWLSgnWakR0X5zLKSE/j1l21iSWB
kAkoplNXL7pk/wON5D0SWQhueOVwwn82mKrYbQ2aQzjaQmQF4K/vLmi/B0nP5OcgotBMU9yi//GQ
IQx7jmak1IoD3J5GrUYFpVRMuG6PeEl97/PYVGw8mrffZBKz5eSVk9+ak+5yaexh5IbMrSAWbUx6
B8cGMMLSaEDc2G71pdbZtJ8huuQ5GOj+oH3cGBMeOdWimM19cOuCu4GBDMwD+0JOndzW0zIYbjIt
Df289XetToj0CFMYLCko+GC1Y8xLIpD77iC5qNaa2AQukx+3NFmHBL8VK2PUk9raAm9EaTZ0Cdkt
SdsLqdl0nBXhlTymjzZ63iJA2G03993/FcZp/TW0efYFttQq7JybfDBuIYv4nALL0agUX4y/bPMT
vN/9ciUPTDWUi1gjOGOmm07xFPxjtWN3MAvQsHjqWPXumuDsBNhagMcP38F1GNwkv3Z5ZCKZt09C
2E0J6fY3Vsyeq/0H9PlNbpxIAuFxlxdj5JyZoiQGmw3lnBsffxvx+DO1rQD4skwxukA2SQYUW/1W
j8EBQhrqTMQPZAy1sI0hqtVkQYy3VjKDx0jTvqsngMAQPduqRDQQJGQYOZmPd0CIunRh2ikq7iu7
cozjz2tUT5BiPl53dvOiKuX/9H3d1Q8UG1lncztltbIOEeAED7niilbKcDGvOQ9lY//pkObIMrU6
H/kLkCKIvmOOK1n3oDJ98ebbXmc0laR9WtwZoGoJJLSStfRgya+nFORKYg68nbfeXc3G7Ek+rgWR
ygBPV3ccQLUfVpRkyY0g08bT1BJTh6yU0FKH1HOWttZGkGC9LlHQROrRjMNydhuqtZOcLXIIbbVZ
CK7vPK/JKGgd0wTzfTq0R0zc83BqtAvzb2pJNAx+e7LgdCiWxZ2lRMyLr2HRBwyDB7DtVlXPHzjy
rDxJBWieWRXCiKzC3ewPWHktH0z9eAVIV2NjSpNZZpnlWiv2v0XcpoWjXKdVWhdUVAPiUPiH7sbH
cyL1F0xBrIc9Q+8I2cThHeZB76Tnhma+FjEIM8VPuheLCIbce8isVmDgLPizQOhFiTh38Z8bz5aY
3pp9ldLSttTogBt8WFAQ+5SoYUBHHp3Tk1PP67tcry5mTKeKe/HGkPUhL644rNL4n8O1aQYC7FvE
fpMj7WQL62pnO2mjswQaNdfPfApIeATDvCf4bcWsL4i29mK9RQEl+HBQhzBMqNRkuJtPdP679aqf
MifxqiEVvSrn6GTf139jxAqo+67upPlTiRJwU//HQ3ru1z9MpyLn2jBnD0af1DpNBl71g0U0Tft/
eyt3oyg+uPIiuEs6cyeQU/ieli0djWLA6RfeNmk7SF/UbS8oVGuuM2cuW5nqQgbAHmaMsCuWJ7JV
kvlXwvMKYkxaMWqFlaM2X4QnUIsUjswapPNQU9xAoie7iUuHHCLUvNo/gfoRIdfeJm/FjtsdQsHQ
F7+y74ut+ZDf/DZVbjIlDBBuNe7vz1s/dzpHMLCPuHD3CVdKkR8wbnOIG5IMgeaEEQXKxn/NXaeP
Nv9aps0pZLPv7gvu76VaV7wTYTNE/m7bpIBJzcfeoZe4uuGxyMa2DBj2SPzH/P5ldpJFVRfNsPX5
ZoaGikussxiwhmh5fIez4RVwdj9QJpGFQt5BHUMjTU44VyOG49rLRNdwL3rzalCrHBeDlA9tB7Ez
PV/EPOnjX0b3jGx6On23O5/PJKx8Ajg+s+w6b3GA/VSMIiD8ge2lFQrlE3dBWGAjOGSJAW4xCHVh
33Y0wAfQAJCv/LAv4zkANvkPkw1eyMrUIjM7JKKNZALHGa/D5MPjBdYatEPJLIqYiwetq5igU3El
PO9BMnlgOtLKVDITWaAQPJFbwTyggfXTXf0cU2jarM6V/tAZwg+pCktvlNgpJW4Kp2DMjf0O/FWm
KnpG9FlCMlj+HbEogb7/zsJN2sN5suEDFxxPJBe6ZLNK0borM4zxpz9d7ptZP5MN9OI0do0dQtfy
5lkO7goRx3gZ3/QlCJ65mQ3cYPpQy6UrFH7GSPxivd3WBgrex3O2q7ujIF/x4tvL7/dMaA/kO8QY
+lwVarx8xeD6du8PeQf4PVo9aRvcD6A1YVYIagp+qY7GoAwyqo9D0HA2QebGRm2uLGEnF+o6vIYe
XRMnhERTpdTjMq87T7hb1iO01kLPuPbTVM14yGf7l6GU0QMd75kGEjY9y5FhUTPM5f+2/TsTWwkj
TsexFnCZ4/e+kD/pr7fxm+vnpVNkeVK/my6dWp7KCAjb2Yx9D2iCn9JVCfhZSesdjDZDQTNYV3xJ
sZlfBt1ZZKwWmDBAADTlbv+WbRgQEXL8BHG485HV+5Qb4BMCV3vVi7e/yf90i+PUDWtM/GKLODDi
D2UY3dKUCSfWB5zv+WW0IJTM8r34MWlO3ZAUr9ysG5bvHh9v/TPlZmxtu7pk/yYGnVcwdFQQYG9h
uVPlFehtLGzOM19MOzO7/Xu/iV7Qqtq7Oy9lvLbYMQqaFYaJqQE4yZew6d5CjP9XlSUVo8QQExme
EM0k5V9eGS5nHwCTDftxx0Y2bhDDv8HSeTcZDjjJI98C69dyfY47mn0SCxlXpienOiWwmxykxju4
Nq/7rGWHijEiMq8Mgo/jIIyHv+tL1gfU12roPlDVUBTKFnUwbransDzigxvtC59n3A+MC6cR9yra
EY5zhuCYC2gQzfqFiKGGJ036vKeKgPzzbt94Yx9WpvYPxRM4jAdfY4X0ZEMDhCaItgYU6zoloDTj
zNzCac7PR/d8GuMHeErhxUpgCrOT6+nW9/Wk3B2D0eSBx6fntaz+lDkViEDXAs6MzCxPWX8ud12b
OowIdbWrzskl74UP32ihFXpwssdOKu3cm4/7POYPtRw7Myqu1KpNJBKoMoCR2y/dJYeZ5ZBxATIk
IGmqp1X0DpIkCeCC2ypLX6UGOVS71s6mIAp/+fuS5lPeDP3cJdEuMp94DGFl7F76Nxcxkkv4nLDW
O8FnX1aO2VucerigYx/TdMhusOehqgNBty2vdDhIcKKTpW6O30wQq6mffm5JBWxd9PBKUxU0oolc
9IX8jEY7AM5nqXrpWGWUMlJxk4ytTyJhhbnt8LuEuAt3n3RtmIhxIpzygD8LRSGPoPbIxSC7ANuF
A/7T97Acvx+YU/8y3uPDJjMkrRwLKKJoXBt/gzE2VR20hzk7ib5VAo6DMNf17S7lo6cr+6tiWjLs
p8rxEusVJ4ipFBY/6YYrq/veiMyTsm1FJ0UFILYWVwI34Uo0Mp6WoppvPSr2okFfhJsGWVGWSo5+
1L3+61pU77nQzkmTnjM1nEP182RnLTgOD8x41upwcPJnSObTnjTVrWv5NZtzY9RaLbF5AWBoG3vZ
ElT4KnUV2Zk+++uTIx+FRhH45o002FDsC96YpnnjbVQiULpq7fSuikRUiY2o0dclqbFq7Dc7vWs0
+ro/nsZaZHG7HKuTw/7AyDROuJ7KXKh5nd40+bB6x7MLkKYJjy8TTpDrBK2gj8doL0jouLVsukSK
pmk1qaal1Yqfm/AEduZ7TlZjoFshVy9kd0G9Ahk+nfsve78lgF44rn6EvRtjmyYI7FX235ufIKKp
wy8kYDeuNnPcGMLrBSEhLSJAUqSmrO5SKRfduo/x8tPhoZ5/NENsFSwCtB+BFT51V/oVpqFdvZ2S
O9gJVE52UXJ6AZECAPrSpv2Tuhzxp9FUkbDtv3ZixuXdd8fE5EnSwdkM2zUWolD27rTwQ0VrvKN8
NKrCtkYdTGEIsxHALM5VBgCEWqrIp/yHLCWcosy4aQkj44Dn/1+pok0u670QHTfwnwwvWIDkladG
qkh2j3HwiSVrV+RKY6MoiyR0tnXgPCJCG6OvvG/zDIlAiUJ5sE9Cs8DzRnpWfcHX1KaXKERmgtep
AdcIycADVv+J1YQKNDdzQL411CnONgSRe0MKodJ0OSiW/McAG7X4FHuhEL4I7uRLjaOcU1WK385g
PAs5KajdJ/sF91LvbHRrmjA9R4M5PhOVN71B/3LO64rS9DvIMFiwSBZ7EYAS0VU+OMyHgJ/LZeUW
buCZ+UourxHEycjezzeJvw3kkHdb+1j0R3fV43o9Ox/4F3CfXL4C7PgdIUb+hFEPEky9sQNLOy59
HSshSX74G3Uwt2ogs8tCXQYmUNd/FTQ7LN2vt7+OwLuCFow0k88ku2a3aRbI7f3c9Xn3qVZ7ws7R
b7iGBxJGKhdBjYffyw7u9rILcQNsD3Q9MrqaGWTvXE2oH0TmwRPLMTWNeOKEn2tu1Yx8hrPqMWGj
Jwgyq6pi0chGROKaOQfOy6cUmwdAmeIQyAv5nz+S6r6S5cdVMTt4dHtUDuu0ou5mcP9r7S1nMtWR
GYNoB4lGEVxLyDJIp195jblw3kWy0vaVixVELBaBx6iIDsQgx/gy4er3Eq1ppz7gYzQuIHAOzRuT
WUMpRBgwawctLLSu2a9kD8b3TRdeeZao4qxiFIaaT38iJ0FUxr7Uu6sOIjiZco9h0/kCXlgdSvCf
Cz+puJ3PSii/ioPp4vPkbPL9isKzLCa7+we3o9Rv4XQ0ORAUXd5qcr+2okMhsCU8T8KUAvxUfSyu
lqkwXg6tmFSqe02xEhU5XmkQA0gPqLPIWZhDu46grxXOXTIEAyXWMslKZUza5ofds7urE5RReK1o
OTEWHe6v82Ya+A9WQLeYB3j7sIZkM3G3lmnGpeHIBLAAgfUVFHovQFa4ldNyywtq/fKgujCyA6l7
PQyuyjh29sexPwi0jGbOKZ0YLZf8ey75eu8y6XJXwHgcpbe9h3OdyQGbRryj+JbuRr+pnIpnrsfH
nXHYCVU1bY2RlhCPj4DPyJivwG/6NcoxqsT0jdbzebPo4Ztc5IzpCXOEbp+b7SQvZCIKKmSjgPtQ
fsPl+LKEke3BH6Nclp9QZJG6GvJmi99izQhRg9Na3fe3SaK1yKFR53hcCmVKtQne/v4kR1fKTVU5
HhS9YDsGfu/Xy4+qs4eJ38T+Ly8ntYiX4/jD0c0tmBKGhAWL3ZUvLST6/cDlPxtLdD1627RofdZZ
ebFmjg5l72tL2iwo40Pyx3arf5d2vDWmqJ5T+AiklS1kLdG3lgtmG97sHxPLpz1POElVvODYySKQ
mBC0E5AxrBWxS0DQAHhcmjmda3n73KS2ixrGYxpU07AQEPoApBNOzF9soz2U2Ny0kZPajOgKu9Wy
jyMje+/CKiuEnGU5RbKxX7o2kcBeU1BbvIg6B+17rO5pyYQxwjax9y7vN3l7sn7zZZw983+nSPSK
kOUmRhclGdZo7KXX6hN7FOuSAAaJkkbLVx54DoCIKctos1XM6DP0+KOsvl+OzJn4jdYaNE6HihES
0qHIgx3YTojaXMbvDJNPeaXISBFeS9/I1dKhIhPiEujtcZmsIVTDrFNvN0C2zTbyDUzdCBNh7GoW
3BrLNvlMy463js0xVpLiiE5oGkbGPb5Or53yf8djUY6GhiKDi/H+zxtBAq2RoKh0+UClxZ2Mhc5X
MmaUdJJKSEUcqrmO0sN456DfOFY/FNRp8W2j0mDfUDJ5oMpJhk49vguSfBpVqRjbCkXuAKMuBptQ
tyn8ewfMy0EAFd+QE0r/A8TGBzGwjk+XNbsUlwkWmX5LQdUyxdNAREaMuHT3qg2UMQpWDGRoRtoP
W2EzE+bW5FvXs5OUKRyXP0TSUu/T6UV4zz86LVAS3N5RRnHdMHRLfu9h9v52Ln+cUUcXMg/J64wF
Qrfk49+FCWu/Zfz1wk91rcw0P2ghPYOzGew5ezm+uUzti5aDMvHivOhYeVfk1zM3hduwQtNWVXqH
S8Qy8R9Phx65dWo4abxc1XQXIb7BsyceheSY2fbGGg4CQjdU7yzyRDp8cf4iCrt30Fc5Tz8UTv7F
pGgblCsUE7CYUMcLaCgf57GAEVAspxBY3cPXyvqy4FsgDQNdtX83zIiqJVMPzQ8JGr0hJh7QEsj6
tJl21tz9jfiWXB7l5gG1yPRcRVIj5+IAVF0ASTPue/LiCnnO1Tn3/IFttyaCrMc/npPNMR6F2vBO
OWABlOEiqwfirPpi+queV2XPlzFp/WtU/JwNHIA5RjErygvDR8mtP5/o2snYJFSnGzxIb3kcYnzo
eS8L82rbIG+XUA1IOy6kPolrWOTwTJRwwoZNwMNH1KDDCly9nQqkgAaKGASUXn3eOSs+ZJGgllh+
EW6t6NhUygDsO4irBQED0oSjRsofl5BqWzd+a4nq/C1hxDkRw9Ijfz5jTUdtG9Rj2lI1qLsqaq4r
whzKiLimwL2CcOUWR8aSxRaam0L3fzbFXExeWSyN4fCP3a6Xya/w0uFGxXZT6fglP86N9raJSMT4
CS5RU7cPYc6gd6SMhUa+uBL06njZsbDYFbp9DStqujf8I1p6ZrCPjV3Hg7wZZiJtkkJqHxySAjaX
G9KZ7gkvR1VNxpHPeGl7LUUsKirEc0NhOG2Gs3htWip/wV6jlKXUwswtNWtUZnevB9bZICGmSgaU
3mQHoZqSbbONjoakRcdQ6aWUB8IuSSoROf0OoX2mqw+kEGXCIq3zzmHokkBffjy/Xdh4V8bT/zRS
xIXWhPZwN6ptvXE+zxDE6wsYt/d3NXUbpvcXVxsJLEN+MsNmLUPHj7cSXuUy4OrSH47JJeV5JBy2
5O7+i42Lei6uPBzX1BW+ZaDBfCCNhJT6dvXSBQ50NhVVEg66ZViyLbaBa0YmdCFU7FQMR+Kh9bmE
3Obv/Vd7TuiSQPdhlo+Ivau7JyGjYa4k3q4InhhUBVZ27YdmsiKd+2OqfY0b9QN0I+HoQODJEdMP
UuOLJYTtb1uQ+XH6vPKQOvmXQFf8xu5yMTs+oMT1iQTE0hOVkSLe369wcZj2s4e8YuLnyBt+HE2A
Z/5hLWBVr19zqZLxzNVcS1ZTjMnhnPZhVrzL4JZVuYi4aZvo8MoBmBKwhFAFeIltvFh6nYCYLBEi
YHWg3sp1FPfjE89DaaiUCcpILfQfvsiWA68DAOfqZ8wvHb+r0DHTYkEAZH0uNlvde66SkL/HyI6X
Ckd/Fz7wxTEF/DQ1Vu7WV+w+boRVUcclrF5D0HOf8AotsJiyKBiH8m6Kq9NLOvYp7BI1zKCDV2P6
DXgH0JiKoFB02gHNzzsIU6zcgOxgI03D7j7kC6GtiGTIDQ4M4ksIVMhIxrqUIdRYYtr708K94RQi
INcqV6BIPXbHrr985Noew6slsdfUdMsb6hI1Y7ATP1AnyKA5Ukj/MDlmC8vPMn0LescHUdE9OzqR
/F7PNUjcEUPyyKOwebiYY3m2N5rxfVLNSzGbTm9ExLuvTjXtLXQXP950P9REJoufqpAXEQAUDHc0
7e3MWm61c4AXqTT/upgVgQXxhEJ3gJePUQ+WDhmzPCqD8C6j6o0DWWvj8EVVqtYEfUUrWLaxtCkT
/27DXcGYk7N1RNrPqGf2OnTEXw8AHN+MeHwMCX7j3fId65y5KFUWPAm6wMDG4a6YP25/D7Xl1kbR
FCKoBtVWiWngl1SfQGZnwS3bzFd2WM+MJKPPCJ0KB0zqC+EhX080UaYbMVztSLOFWiChIQDM2ekK
dCcMidiM6Dgez043OuPcejIsmgpk3NZUwTIyCi9haXDq/XPvvc3+X6zJNXQefXKOjSFCTRwsCyn4
DO3b00OYJ80KFznaRi5+cp9ddAInDPex7BNYpVnUeboz/GVSR9cSsuDRxiamTEmm0KmDmAQEMewB
gFcajlgbXVswaTYgjgPJC2Hl8/blLWKRpc/i2JPzmNC4djiiCcgL/PdEX2M9NdYfrwr8xVK2YUsK
dxGeEZMEpdUS/qWBJpZOYKaqf4s+bMvvEE4SDIJS7EIUjZFJfDDG9qzyLsG5ghCfX2aapHMXIlbC
TGKvlm904vYgCl1njiDJADYL6fkx+6RZNA/flZEnUr33XnmrdPxYq3b+urycdi5C5TEnY2x0J1Mc
QTBcelgq8aCCZf2tPzGa4Vb16moj/EDewx7QpYLfGtXRJXZxKAM9M5a8y9fMYuE/RnBPsIu1/4vG
IMax5P1kM/noIGMRnz71oU3AJX3K0KI25uDpPDOCS8qT8xeTDqMuReyPqGaF7A1LkqgztNkqbFsa
LPaMSsUVfGMzsGYNExhTlyzynGMYJm6oZ10XvweG9uUwnLHYClwut2EP9CKOU/euUCH38CqRCmul
LrBQ6T8uwAM8923nReIy6w7Va3N66tH1aht8LM6uqPnuBvEbydhDoe+ma306SHC6YTIaG8jhx1wE
Q2RANMJmQLr7Mda6IXZ0HoReNtJKpMgYfTKZgEvmuay6BfWRPVo1P4GzxBYq1YEbccEVu9L2Wqie
Dzy5f4MpaltO+RTV7n0b12CMIkjIvNNklr38qaN4+C9sOPJunc+6CT0/1LQA7nX7kgeaekD7wv+t
t116LzbOvUfnVqXZOCpwiNqrwSnsv/zHra2E08zSEujQI40MKy9sInzTbEyLw0bdJ+XEVMUozXph
qG/3U3Qfg0MRjyvbnLTL8YW+f2r1n+4uUueNejyDnlPXgWALiiu8Tjvjd2wA/Q7zVkP0D0TYkExZ
XKzM+07krbu0yUSod1qGtyOd85l3LN5KbUptedJV8AK6DjqC2I5JqChwFsrASdZIj51xpHhd+0vI
mvAOFTrO8T8Oj3gYKjctdLK+QuU7wxTslQTHf6PsnYpBzqQda+9Fth/2EqdW7cmZreD2Mo4WghFY
Ii+bMMQDmmDxWJ6oT1wgIcLV2u45wrbYz9kNe30hww7TMrE7XAXm/2tPD6keI6JCtWTQQ0z2hAIu
rKpo2LD0CFxAJrafeRCzC16KdfHXKmWw/nlbJ4KwD2jMT6RRnY7z985zfSLH+KjzHOMkYeA3CMld
+aXYqBaeVkcWM90+Gja5Q0ZVUGCrdoObUAwC3etodlddLzm12xmQ6O+AZ1vk0Cx5ijnB2vXFcbXy
vzzaVFRYFlc1w4pD6+ljbQjXpN7/KkpJgt9kSrNadjMuI9rBKi3qN0GFPJEnNEPBi1wf3XmHTe2f
pFuwsllUFqoPDwdHdCE5TE6J5WBklqv72vhwYorhQBJ7g7Td9GnjE3qiV9+bGN+mbeOaXSo5ygw2
PMG7dfX0hUU8ba1CmIpN2itXLkDjx/cWcY3tP12M0fchdez3CI4D/yTcrcaGj0eR59KiM8+qX3MZ
FFNkrWxNRRlwEAYY1i95qYmKEq6+tjVZH2ONygEmI8BVLO4chtCr4KEvftCajQkpsbP/Ja/Xp1XB
PI9yhD66EIhqZiB6BQJBps/055rP7/QMSRmcM1VQaUGaRKKy6Fbf+W8vimWQSAGLyz6h02jL7tJi
gBx7iiiF1Ng5RdoX3dDaQ1+gwNjFCn5UCWTBzxXD/sM3hWiwZG2yxoBJ7km/sfXIsHuSeOMdzrIX
bqrNKOlbwPouXszPUerv/PCja0leAGK/UNJFDbUU6bo4ZsZGtPxFzh8qwMyKhbxAc7wz/VPVBzr/
zbDKXqm1OQi06uMfnCKVWBL0pgJtvow2s2HGxZoCURj4vt/Cp7IV1s9Ca4RMlzUweSQeS5ZrsOkQ
iS497akM5j2gnZrQ93uJm1vYdCzCvHzNRYfSBRZskhELnfh7+ltmROoM/vuxDyG4lNICj2ULU6r/
yvm7mPhbZvQaSPAZkfOy9JBohSqfsQD96aRU0RCu8/OpkwsQk565nJU2B/6NqPARBJYm74YaLguk
1rm8jmQXKck1tnKMDObQ38EVsaZWRvh7QYvUM9DQ2yrlzTSoa241/4gLSGCcjMTa8Nqw/dR7eSXl
PHRBBlIL498O/Zi2JraUHFuswbiv4sIu3OEIEJzDHdijtaHIKy3NbxbtcrpGjQ972avPZxNQ1r7y
m1widh2c3h71aBKKxV9lCtj8ktmtrPU0SSByYFK0EGWC6qx6oCq9KfXz+udTftU/tyAxAu9TWacd
mBQwkwpV9P7YdeJu0cYgEcRe8D6iMhulvFDIX8uqiseMl7vEkBFDG6+OuQOI+gXVZh8iCq4AbHVo
f4Ha2aksSq9tR3fYHRL61oavuO+qc6ubTA9wVlTJtvpOqQNJwZYup6A3edjTNA9vBgfSrYU6CLwK
32aFfAZ7XQUOR6baf67gQ1u3dpiggxSEDl+/T4v5yz7BrBY2K8ftbqYqi7BEZpV22m3C4mAmXuKC
mV/nkdJLs30aZVuXhGR9uh+8ex+3JZ0+ZtzLXMl8ekxVbAW0K5pDH1pQdzWZw1f01N2dF0V7inG1
HjwDStyYO3aGHD94mVMz9v2m6LV1Yvrvr9J6vYLN+qw8rnBa8xK9CUFsYD0PQFvRzK7DQEDDtpn9
mRexMTszQVTDJe0wWrZ5/i84yh4R2iNCOu2xqEPAnBx4LM+h7vv5IIksauBlxsoccWU3wvf+UkE6
l6+BGMvXe+CJw2WlbS7taZa0yvHwKYpcQQUsSMahY2sSrcMkzKFZ3GJZA6S92ud1t7+AfF6Yya+t
5leOjumQX/E4OV0y6gJb8iYnZMrFwx0vyKJmlGM6KT8cZNY4j39yQC+vaRFYSTO+mSyRy/+VFe5L
wdvoFGCpzCeautPJJWY0kipIHwvS9mB2hsw78LAqsKfusGUug3k99K05ZqFPwRU0Ocl98nJoiKLb
lzYri0yD/TfZgKtqwh9VSBUnx4k2ghWj9sdwgmGVD+26ezQqgo9tidUAtFiJUGj6mxzZCfjLFEGx
+3sKRn1xpAGEVv4JeBFxkr9LhSwYbpX4eW4v/pp/Pxgm6gHqr0bNnQu3g30oHcRBxuIqQzEFF7IE
g2SI6ALEMWvjcjlknlnjz/kTbeKyxHXXe5CkWKmlzHewJNoQY5IXySlaiHwk0N3I/t2ImIDGgHfE
9bo+J6SDS/sJN557ttDpDAyB1h81thx+joyB09/+u7ulMJPo+/LpUBsO7wUBSgEGq/t3usPw+/h1
XpBzTy5o5M9nv4Gh4aT+AP777pAANDwguMbfFALeYrEZCqfA0uebImX1iZr3DyWIQNuQC9JhzBrK
VAVfOs+gmuuLni/D5EH1xplbx/VzsxqdQRHpLwMTsqVDuisLMWLG4knRQhO2gg9Q3WJRlrs8WONH
qG43qQWRLRPymvi7UBFlB4rpC+KBklrZ9QuC3LZ+P6oCG5Scjc54FgAJh3ernZeS+1rz0ac11YER
TEMds/APL+I8Ain0jqg78ZnQvDbFZ6lengWvjn6lQyxC6UpbkFIQ89L1MgovfIzm1ElAobbaJEIG
H1z7W5SoYmd0fZaCMwTlZ5/bl8cIS10Djox8XK+rb4gmyqJ346ixeKs9scQYdr0665ruBSHNOOuG
+Z0jsS5zON8hxVFNswx/vqtrG8RmDHvUrvZAoNrv+I3wFyu5B5SEJNL1/YuNOLri3winrMUIGl3U
qgvoda+Wfee8GifE8+aPEkiBXnxUQBRxIvYluDrAkc/ksuCCbGLn7WOL162JSmP1AQWzPPwdlMaA
eawHzjKKoJttQWsbuBmzejfDWJSKiKPOYFTARQ/ZgRtaz+apZzSF4DXMbNb6xEaX8NdlrqZ1tee9
R+3AghOUFK4xvv494XI5nlcWn5db15kHaSRo45ts/6qpjrMX0Ja8CQiG1SWwVVPSeK3v4a4uU621
H4exXbM6KTnpcW9/9lFtkbm/mSB8x9fi3Ajs5IeUhKKJYc4Kx3ONoHRIRraml5VcRUn6TDtj2F06
T19r7GBz0s0imkk2DE0FAWgfbW3f2wZTRAF/YUIp5IxgVjoQtC7X4/d5bCIdJJxWGKPeN1uvhLwb
BpuzJu/l553VgSLaQ9yJMIDseKNsfTsChxmQSf3/Uw0jpc5YAJBEN1pKdUY1Eh9n+AeDy9iv4MFp
I/gOkKnQz94qj+WPkK2kEQGshjIdHysqNtl/wrjuE9+oXe0+aqLXZwdA4MbruYAWkI2GSu4XDpu4
LUhLgNuWCWM8gXDAdoRvejqI+GrVMsGZYlhvyMEjIW8ABIyMs1PZcyCFzXRoIJ9kj77C1HARRA7I
aS3iwPnqcYYbpkHMmCHWhp8F0iSzuya0e9a/3EVSPTOY6qOY0ZPvtE31U4wrNqUZel1mio0JxGKW
OAHXKlIrEtArv26pZBxh2O10To+ityvyXvdMZ1FhVTD3WDrL7zSIzQDH2/NiS4ETPUf9c3V3izGx
gJn10H2Blpoo73c04a6qnLdvNbMVmnCGwgFKe18dfs4IRj/RRWikwBc5ttDvwQp4NL1wOqiIgBIJ
ALXIcX7J6ogr2qWnw3RHAHI8D1yWVfBoGfm9ntfPrIcOgHUCP0tAmMH3S6+j+zYkeBxDKcu+2AO8
ghXyc3Ssv0RJcow2M2hXIqVtEoY0d47rnatCUVxHew17WmvcCTitxSKHUgm8BLzA4eR0hXo/FFIU
7kxIa6cLGRYam22aH6e/oq/hMXDipwQesMDfoP+ywTTSjwJq5EflBvnr+iD4FKofCMjpvOzF/VLZ
7vg5AZA6HUahUvkrjAanLGn2vmdnADSLIenvgzXiV7ls28X0ZE9HTEdcH+wuTrUnmOl9ptE/ys3x
d+vL/A5xFR4ANGTrPKYMSs+YMlLzH5+owfQLcv5ELExqB2cYHAQdjJeuNDuTeB3veejJHlczkW0h
DYBtu5de1RPYd5rxqttuX0mSZY0w6/TBOqOqYR6zGZXj//BpNWHbbnzwFH7VmXHf1QnnMqYWjlA5
aaNP973Ng+W06syLGgVS2GRcmfuY8ONzC9YsPNbrMg5NHXV+cb4IO1Cg6KzEqvT5a+hZ/cSi1iAC
W7UBi+4wXKyf7LPDLw645ccep8uIavxx4kfvsQrPwtRen/9pZ5YBkK+laTV8kRmlbFFB2T0bpNBA
towoyy48Cn3LEY5hloia5iu/DFAKRoj1+xkdltVPqiUZkF275OE/Ci9BiYG5f+TD4wAt7mB8v4IA
YJXCmRCilzUBb9oQe5za2DLjPESORgx5xgvhsbjdWMiuYgpCWaWnfHncnTwx/kaNjCpJ6YDjVfkc
R56ahaNDN6P34tROBTIBFjuFTVLWJHJ6qpKsWe/wySir3NYOYY/zEd9dJuVDeIUoXt+x3TiMF6l6
JiGZgOWpMNc4TOtsZOgrui6/M295zhqTfDDHO4bS7MNrIG9Kta0PUxRtQxfTL3/UXJ32BgogV0qP
CTvDJUW+yeyxvd7A/ka/JQbVB7owWyebFippu7lHHcMliE6UoEve1uLRfXojTZ6IEZLzE908huaq
BfyFUiXhwNC7EuqQ64h7degbGfvgnE0AkgbPVUxnUEVh0YTFfXWBG3xRCff3BGB5ncI/rADoqYce
jAuyUUslUY2cuWdZ71scqqPy3m3NCMbFEnY8XlrIiDERBZOzMxMQ0w0c2HMQ4+NJDrtYaZ7DJf4n
Cta41PEOvd0jxJBMwFPvSFBm2tOCthcGZZEMALt6lwMu++RMRDfr47x0ix4Ck1mljVgyFJQQg82V
Y27QKAizuT1jPrIM6Jo0UZhwECIKXrB/soP1089NoMnh4lujUHwdAMJrYnqRcVECUuElgLatTuwe
+m7D4mOniL5fAtr/6AuRcjlfxQhS3iaKW5HexxuZWif7cykC7udeibinTS6Y9d8vjuVD+e70Z5sj
Gtsaci+diyY4j3suosB3aQm7dsV2vACfg+Ixzcqk+HT4ZPl8P0qb4i5fQp/ikkbaubCZ/vEbpp+e
KuAZt89IBIg9FLz9O7V8cDNF7i1tL6ZgmSSzsStLuQvTxJlERAcUGpH6IQ5XSzowAX22GkfPLQlv
Z7aKdxbj+W6exj2NrUJA+tGGhra6RziDxeoJ9kHi7fJl2aojaGdcka/Pd6ZgOykshJufzWnq67xv
EQiwsDBX1mWsuKpSB67FwV4YYjm1NLxlw1Lv9ZF+lBicD1k31Qj8mHLX9hkxKUadWpUzqHhq6e5b
OnNPBekqeRVjmm5u3xZGpQJkUReH5qA7m0E7qGANqDvwGL+vxrl+Yyis516uOVa26Zg3ZvMV/mI4
W9vSXLi+6l+bueNgnhaZEPXcg8K85HQagHoBwIRXdZbNj9vg4cX23/UjxTIOfGm1UJTBBbvio6ts
djA/Uym2Og9fT58h7bnH5Oc24ed8sMLd2tOk5CRNeXhToikYRTXL3jPanatWNhlmAo+YEPvSpto2
JT4Mee0HH+spf7H8nb/NguCAhVz45eKLnHW417ChcaMVaPRiXhKNerzwfOXRbA03avXsrFh7umDe
o9zDrwXTt+PCRsvVPpvjTy9d/Nq8wtaUSHCwN+HXHTPqItJQkeeS3PpVTgKkj9G8b6t8qBZaXJ2D
VDKcyAJUgdWEdNWpFu5OwClV97L7PC11j8dWsEjgpQ4MyEZRZye6HLF8dFXSqFFk0LeDZ3vhvYWP
DrEZXgEsSQUA0vJs6BEqot1hURqC4Qt/kXjsg40uRj7H7uUU2/cG9CzAdIfeO4XeicqdN4aphkQX
/VEyAm6L9lbkovdhrzBln2Qu726K5rdjn9XA3Wn3xDQ15d+of/8jfAGLpfm5SanU+w8/kZwHmywg
LGEO2QlLbjZsFho7tJpE18CvRo/NOx1oQwD50SLz3lXfLhX1N98SoqRDBttme+uximQ+X+c0WEyu
wIqhkhBc4aABkqLm0Vio8t2ML7gNLyt+VyvXBYN03sludynCqaDPAXcsx5tiIeKqrn4NmglwyAmQ
WKfy7ZVVV/QJnKZm/zvRZDTuvmxcKQ4tHWiqXoMcLqzzjkB86l6+5XgXIiNII3hmvYCmHBXEuQ7I
AoamC1mwGZ3X6ALaVD58K5jH8Ykxn+DYeMkGlNgmsOswibQ22+AOzGMmRwWRiE0AG3jpWAp05saF
BqDW4OUnEDyJkEcDsmd3wcBAAkyoT2hfm4OiB5NlpOZdMGrIiuOCFoaXthktOzjOqS+LoVSUo7M1
l6KHcG6hYm7yQaYJr3mlCcO6meP866wPNlq3DeOxjvug/AbWHX69lLvpE0dHwDODyTdjKS/nbiRm
Okv6GQuM4MowAfIpO1ees85uBTm8ZV0oxhzHi4Yva8kga3JxL97bbwjvNX9XB+DsCk9LFZDPESdf
+cdHTBVeOMEWX95WXL9GIhdE1j66fMvxwt442f90U/ZDBsHshymwSOmKgv3OSLUXhL/D08jTALGh
nY4E66J2bD/w0oePqjPHb7x8xI1jopF0gG1getU5Jdh6SJKq4TOf4GJvtGJgmw0HZiCtrPdjP7Aw
jGdu+hVxf7ZWwMGTx9MNJFmYoeDjK8XXMaiKRxztzxWr2UM6iOshWjNdBJg+8uYopVCXfuYwi/RL
6Q7cYWo8CIsQNru36ZI+7sl12RKgidcvP7n0kGALU4nNXFwhEtkNn+fLbbs9ifzmJC38jUsWyqsr
4hCWRsAfz0Tz9IILduzXk+4+fIYJ19wO/VnALAA5hYVWMQVnUTjRJFe1Z4UV4Jji+rkGXX7YRb2B
ShKPv2qecJPOSq+915WdHDGqkNZBqt3DToNQo5QEw4SgFzjDrgOgar1JN93WHAQ91dfcNBlBYP24
BMCwT31qdyBc9ZZnOKepR+nsE1SDI8q+k+KNECG0q66odu01pecpUJ3nEBQuKXCz5EyJF28bX4C4
UmprtSyBwb6mWTHXa4C5PVvnx9jzUL+0okYxm1MP4+vfAGdSzpcmX56hpemUQkFwjOV193eIpGbt
mGzfiA3kgJr8M41XQJGGn74fOrwnF1i+ZqHK2PbMN0wce/QlHlfnCplqN5tglUUYyOgqwGOJgDxw
gTuTGFsBqW/Lw3v5AbazBsFMdLYJhCcge9sWjyqkAFuklhlCog2DSTtQZeLEwXabCntsMQ5SfNmw
QyX2ki/nMb7AGn37CKYef7jsSQV6cB/oGVRyuaURnJrvQql8p7e0ZadQ3yTozmDHxkEWQDy5ZWTb
JArnU4bz32F2is047E6XdjrqigZQsAN58hmASrcxrkW+gYE84U77UqVd5UA7zsLZmE/AL5HXSo2a
iERtNaSkzHChHWY4WnBL9zwtBxYfeIqiPwOI53iORwXuZZ1IytiAO2vPU793LtAlzljVlde7bYRw
fE8vhL6bPUjceRONQkkSMa9sYXUdXhbEp77WC+ZGv6qF1s195X/6ZOBasvsiN2+wMV8Cn+6pbshg
sclGeOwzHIHW1LPDln8OlTI/wcT+g0G0m9WuRDwC2ixQhIqjledDnHvdbbVIyc75ZkRRr5ZJKOzl
lUIxLKl17FZmRqpfPPCHhz6O2vCyjcpFz85RNqak5SJwle0sEQm03pCIX2ruDjztu3eaxbA2P9gV
cQq2mEVKaH+HXZnvb6eBvz3N6RdNU94ZcZBZFcVG+pQPEaBIcLUtOlIIRtbHSfdXEB0e2FdOvou6
BEx++qD4mbuuO7qM6VRLgDMC4bN9omJfU0+a9hyOkrklZQSQ+lFCWI4tWfZAPveymNDb/yzNrIzQ
uAPrOwdx5JYoSpFM+WQhoe4q9z1MUj5Wv6onEijcNu4lSd+4TIVk0vwqEPZ3UteS5KzqFqF0Juck
kVQ8/cQRPHnsLOHmlkbpIAV3zKYg52T3TO2q/X+Qq2yoECt6vTCNY2sk1HvNbXm762Xb+2nJLU3Z
zgT0DZrf+rzZaO9p68Q/1Luodjv9foByxUWb3zg3jX3uk8TRZzJRlhsGCICz0CIzalAy0oi509hq
MBO6K11Wl09AQ1NYQM2k6SO3kljxSY8v+/Xtb578qnmX/5xaLy5MZgiSue7bMm4qrkKGDVv428B3
EspE/NqBzS4enHaMi7yqomtW/pYGa0qVbBY8Edno/+VY2c4U9RrqrcSYsj5QsIMpasVlDwVE14BU
yKfl9r0AyPJJ5V+WiIuBbE7dIEDPj7O3FBdOWHez3ZUP/dWwpjjoasKbDnC6TIeaGg3dNYTFnVXe
Pz8HseQmU6hmbAJurnAAYhedzt5sMoemQJ2ZywufI033geTB5D285FDydZL7wPoiZk/vbOVixZvF
UFGajcPZD2I7ysL4UrcY1Zu6K7Kmk5yDmJK5VojkzjcdMsww1YwGntmSyUMA0lVQEJkmgnEjcIAr
oSfD5R5kkywANGiyRIT/S/5FGzl2v1DOcsAx/Ez2a91wuqPHwFqOcsYAiyeUR+EfAp+iAiv4T4bQ
MPNzLG+oqlwLvqpYDcWVIhqHJcJkrEG2/dIXRxOETuP1XPDha3oDhK1sTFoGcno583leFlIweLV3
f/K7dCzZ5idBendcovFC04MSoYM3HHp9aFeR4512GsgDFqAEPSeaz8HOcK0n0LLu5ZyXGY45WA0b
GJlNggMmT9sXuKDWHHLBXtosyq744FG21Hr2uW2p8P9B+B0HQrLh1IaBodbR++y8VY/B4TVVGrEl
P9/lDDvFPZ73qVhhZVuV8arPAZw2K6S9uQa9SPWXUCuHzU7dBEkKxezg4ziqdcrbXcQlLSjO7L+X
4ungszeTYB9LEwXFK/nyY8gO7ilzq7qxR1jEPLbPLxw/3fEwuaycCRbXmlmFOKi+QTpBi5PRTZdN
h76xemyFgFS3OKwYQUr1HPljpFVJYoZdQSJacLG1b+6g91vV8ZQKU/9TLRMdgN/g/G7nFflaRagA
rvXw06TqO+0llFFYkon0RP77bh6zen4LoGH+2MvAL30pHwFLOesQ1P+wJxZ3FzzfND8w4eghxrPf
pkhXB9/heeuPb/IV0WFjQK2Li7zeiuCgnLUAxZb3VJiS2zPpJYc4JOzIXM2w1il3It27EhWHYvSq
8iWkLfytpfJPM0XE6aAe111fWBLo0k0prZB+JtZSA2BAAZkjsozVEyA0VbIycO3KKYxGLGkO8+15
WjGeL2u7xLu28CdW9WlvB/EXr6XLtc3GTuUt6jbWA5VSGReqqXvViXRI9XTu2c8ujWittsGT+19R
HgxxUTsrsrArp3C6irRyVnq2yHjQBMgP5zpp2KK7amttewIK0CGco82/nB2V08opal7ZlDxNJyTf
PRy68ggH7pNcBguKIr6qzHi4pmtaEmL1SKbpp7iNCRiWDcs+nUkEdgao64flMlo7uHK/BiqcnY7r
rHiWV+wAb4UamIEoH2alOaBkC09tR5OGtf9StK/avZbYG2qdu4sUwUX0luuK6YZLrV3jdGEajdi9
sL2puVrdyHqpRvj5onQtpPR+PtGdc3zCdZVBh835wAfs4+pe/1IqVXOaLbpnJKo7q31nK5feC3Tj
Een2IBXCAS0qlIlUQoGYZ3Qxa/QLzJ3ef/nPCfWy9WV3MDpCRWcoKF1iNboRt+WsQ/RFLOgKt461
7PxC9Yct9AulHcZI53Lo59TvHI0GiV9shQMo4eJO4lkgnFta43zG6BAWy8uyt37wBwkvNrHeOv9+
IG9NZdGIwRD5eaz8suFLPE4tzccsYfoe21poIYj1ColYxV69gMLn4PfD5mz5vq3TA3DwC0pH4XIC
l/kURKZoqOWqeWh8H2NQ4qIjErEIzfiVKUwM7dAuR9gm8wyJAegvXePNzFjlo9tgmjV2Vwz3DOjX
JRv6RWTir5xXd7pwoeYAeuKmLSm53kJkoL0e+k0RR3CZpGmnYQgzxb5nEGA+S7bmlQtHhMshmWg7
BzZKcmWck6hkCFxPXztWkyVnhZvA5/cCTKS3FmfA1L2xymsd5z19bTXn9x5bAaYIWoS8JKXzoS6P
hxlebOzph4h5bF5g0w0dfFIx5vM2YUpTtEKJ+TqRb44bQ0jv07HgdYRnluuhn3jFXfGGuztma+W+
wuKD4eq1hLlcrcWGdKe7pZu2faiSELrkMsFYgaZfXNde5/nDK2H5sBLkBQayRcqhaFhnaGeykZ+B
admaXu5eEFDD2zEhIM8ie2vTdzQbKQUS0p85A4TzotxUFihJdXFdkM1kMLd9/M2uRFk16STZCy5X
s72SFsur52xz3LYTcWXU68ulKG5YkB6F8aANrM8tpDFfw9+37+5qeqKFfxR7EwiHmPa4TjAxgqNm
zgNI7d0Fby+5BOA8jkpuLlKBugyJeqiaegrx2hiaUAQwqfd5mdhBpkUu4+aC9zTq2QenIG0qj4qs
ix6hl9pntm8N0wzxq3JSqxjwso2qvuUMj0esooa+XsnVcm6souJX+9ys4cME1TyTh48JwFYD7RcP
PwdO8uhr5aSF7/LgOh75prHUfLk8r2CfpqCrDsOcr/jW55cdzb45Rwpf7T1Mbh4nTBKAVgHIYGqi
WWWeXFT7a6UWbaoR91ZKuPJzUm2wqXiho1/IXzoWDrNKqhS+L5VKtYabgFbCwQlcjTfTNHp86nIa
l8fJMFXRN0opFj44Lw5n61JQ0lOEP11E1ssVElNbbiXJPvKgP0RB1pZxM6Y2xWPULWsBe6CJ+bqt
nW1sOWroarzE1kKeNPA3G/U2qkJm3Rvz7C3z23XA1wbrx9BWfsqbozGtl0RSXwiCIpkkqe/jMxLw
/wR8IcW0c490xScbiPuj9rqlRPolvrDVeP5+nhTJ+qQtLFd6bqXJcJNVLDVvry3awdsWWCLJIZA9
p4b+asRWZTyf9ntPvGpoq2IJYPeDKaY5qKoSeDNx6RwZXpDkGmPNdvovbA91DROLMeJXGd0AIB7Q
2RJVLuiryGQRrilZLzC0/oi1RMQzf77gZ7GcYaJmtkfsOhxlRsDUyg2e0YTpqNNevvU7B3Q6YwOI
62Ex+wYEv+OS5MusFfl5En7Om6kZx5Ys7Uwy6Hz94IPNkvfsgYcoiBJvtE9V4rUudX1Ot1A0N9h+
H/GRx6iYGvxo+cneWXldCbPbPF6HMYLZevD5OdMEjuroOhRxpsUNYt3GWX0T/PeoHQWTSZ4OH6m5
NtTe/mzL6vjkxajYQ1nTQSmgxXbCwmLn8+jTfYu5BDxnoaWRy/9QzjVWfzKcJuWKk7xinmU361/5
DKZrFibM9PHkgATNceicw2zgOO4ARYYX3X/WxDVjq+Nl36TQOcdyyM4vPUZxbPVvFU9b90Mqo18n
V6lSlN89vOA5gziR4hUTrsMdfcxfIXkOTercK2L/KstjImVsxF5jDv/2Uis+ejnSKIsG4uAXT/3M
5kUwzXZAr+J52JTe/vX7Ax3j3JGnc39baB1J3bGoMWABrz8w8p1HO6roSWdTyr1dRlnxwRBvNNA3
MPKjN0LXAl1evd93Y/aj4CYdhYKR2P5XnjBlmFeeHUCh+iMDEBq4yTslwcnE5/XZMO+YAhzPnBDH
+IPiCf1STM1Q/wWtqq6iFsFRaye3+PGdyF8a3AqHnBrbC3017k2d6OZYwF/g1BPO2uS/L76lDppc
SupYqGFVbSRGpKlrjlqAsz1mdin7D2Ij/7ZQg6hY3I08c4P/3QitJ/JTjpKoMnG7Fi+8kWazxcQW
z3kdisG9auXf+/SnlPoJjaJ5CTByvvD0rSFur89SLeZVLkIjh9ERchts5TUwYS2seHCPSSnn8sHJ
As38tZPS98BNb0Y0s2ZjHRhyQU1fZFk/m0jWsQbcZnmtKzWnugIZIE/9tfd+5Lb/xGA6LVzaSr0g
dRRNxnVv5zLdAzvvonowTDiJJp42QSLlE36PpMx7jzqcCsqQX528lte0DKtf6H+ZQoFhPTjR/bhW
MmMVUCZcXqEFEjvEpO4m/J7di4BIDcFHqY1tICTRX5fEqjos4/gi5qc+V2RB8cZw1xf9WUKL/9QE
eEpdy9Yxd6U1aE/FyI51kreoxrm9P6RSG4W0ROZLfTz7ryGpiWhahmtJ9cmegmfuC6hB1AcoKHPu
ZvTJn+wFzENkB5KtZIvUn1bBibPazRql+l7lmJahokFSmP5ZFnqlNvZ5mEP+SqRwdnXvIvDLHLeC
9QFJF7+T1+CFCnh9Ow0WSZrM7RUZA5KXT3I2xYST+ahP6eoMdgKRJN5Ezg4lI4Yvxy4mEjK9/Nxq
NrD4ITkUm58r0njGQdDu0/P7dHmLspujcggSuRDROAfOxamZoTyhTohGysAlK3+PWEyHLZli2G3r
lobscM0Oj/e7h+5aBfuETUnaM/ec6/csYwjawDNFaKpItGTXgUxy+1mOlQ0vYNYF8+ucDG7dyfjf
1U2lrPtfHr04N9EgTx1ecsDS0sttJpvimSo25GaopW/iTjD5T2vSDWWA44/B4TIJrmJ99winVuqU
y18TA39YdthdNto3Ej51Y/+iwDFHQ5ft7IRasqkSNuhjyM5nvaG3goCPOw2V98Bdvj2NhvLVZaAp
nZaF86rXuVEbRTfUXFukCz3wSnq1hgrTyIpmhEw2OvEotsc1S0Us0FZ/WXuZZxDUTVOXIHNBbYer
4VTUg9u12TfLk40y6YR0gA6KVXIvU62jzSyyRZLpUdW/ZVkDlWoD0BMmD5Yx8ygydTH3OhTVdWyu
4X7jXDQUy0e57jI1yHH6laFTuBsjNVO8wMvfCKxJzcKVQCZxESh79hB+hn9sHJFZnYyBBLnDGiVp
Pzu28lKMgEACIUDsr0A8KLEyp6yyP9CpP0KwTvctYLYqv6n3AzE4o3T0tWgFPrxfzsYD1XueWrqq
wneNCMC9f7KYM2rPLOc/sTfuSTXH6F0N3XewNzxDdY9Me8JEPKliVx0KQzFWTC8KQ0X+J5fNzDSD
gyzyMgDCVlhkO/q3XFL2nnvJmhR+o0WGS6QHh7n7IW8jtoYSmPftOxbW2ektqXXtKlJeYqxbjOYV
9pmjrOQizECvGs+QgzX04/ZlspvcBhj6gylnJvtEaabjbVx3xLVRcanJ4FfHLMLl7qQozSpkiyrc
eDlkBzz0tKmgQWUuirFZeiHiKWTvkatg3p/9S3iskwjV5tFdsoMQ8vg9QrJdYMupHcaMbKNAnShP
XBU56zR6NL3XTtHn+u1hwjUdT8uI24WBYXYGsjwl3y+JnUcgK5iFTWilONk0znEvQKiKFncFBZDL
owf/7jla9R4VjNQWT194zElK0kxF/Ai5xv+RB+zWvZpunYYpDRr8WoSyMKPjL0/xoyqhJlnbBuIU
P3bGV74eCvTBkbPoFnJ+YzlnrXvaEUDKO+b1ah60iipkEzFlG8IUlk7KZT08iMMaK3qcgXDa6px+
jMl/NNYd+c0yVF5G2SeBu+h2nqgLnhcsqCOKIBJWBOMiyIBZiO3QYT/lewnbLO1JWNVge2U5fErf
1RdudRngX8nn0ZQZo4+z+HHgYsNROw0SKNsbXkbSXOWL149WB73ee1yD3Tt4vlFsSrRSYxHyjott
4tMYmg1q+/mSVXMoDvpSOpg92Nh8ybyFFdwVoetDRN9xYxe6hJIixwoNVnCbbj7JM7MJwLora6cr
s2AP/68m5sJx7VolNcCw/Hf2fnOYCT0dcO3y6fRK6AxJv2KyUsEd4UC15lRWJfMOH7vpuX07q52E
kH1wm+PSpPmVMipE6u1VuDFoiisR/p4xqfyohNJULcwrlGtu9OcHepllGkorwLjTYnCI8FiJqVSR
kOLoVDvJ9IFI773XcSwQLHoH1XjQgW8j4nHHYhRS7PcbcIGkeGyXykuWZATBBg96pA2Rdcrf3FJw
o+r3yfSzjTdkPXoFaHxM9SVLDi9rAj57PlSGFljsLK+I7jukTnvhJdR2yrHbFz25cESAoEhKVwEB
Lm/wQYZ8fyq6NVvunXEX4Mz9XMYtTR3mtziSdH7TCKPW/wTVBFmVn6iNxRoPsvESH3W57pOaZ1I7
AZvuz9YU7buDMO+eUhQITSBFBpZ6bh8I7Y86Ad6S+ApSHFy7tzzu7PRllKXi/85vYzz9IjAERvcS
jlbAJkiv8J+GZtjZJ3uRgqvFIgE4ik46Wt03CP4y+8XeAZJczBhMVj1Y5dltjmNCcZWT3VCaL+cO
5Ox9UNSdRvCpx6Iw4+rmvI5RkRrr9EhA7IiZuerVDsUqzdMWgkgAvMeJRpqtBx8pdgM9NelWT1oH
3ahYiDMCfXj2s8GfKaUZFZ8u9qWgp5+BLOlQo+rpyNBYfb5swzTFoGVwayPovekV6mPRvN4a/Qz5
OyBIAdTCHjAgDpTLE6XN8KFoF2KMzeJCFrX1lBl+n27FIrnOU7qb/KQYwMsQRX7BvCBGrAwrsOT7
SmTyDQPCYVygSQCnDUklmPM+Z+bKmdswGwgomIYr8Smrpt3AqQYRfPktUq4SY/XZfYi9mWU5feYJ
VqbaUThDobs4wnWJ2OoObDX8zzNIVOqkqvFafopTkE/YM9WOXCwUQI0adVPaLr4BOyCKAqfpk1vS
YxYIvtVCFdAJYIxWqz+TDrngR9OlwkGKs7zb3vAffnMVEE10HfwmAkAdfV6pLAMkGdcHH8y9453N
sUxyRSeuyqddtgz10wbIUWUsopEkfFIBeGUEMkuON2SD8CNHbX5OZmMV/gXcKRwb6NDrogO8dINB
Sw/wKPTt5kkYPL4QUExnEXqMFXJL14ITrIGihYqmwN6PE3Nc+7rSUEfoluTc4XnzJvzaOTYqoqL5
2UosdBNDGZFwuBp4WMq8dYh8sO8v72GvgrpbpHuNhCaHpmRGVCbQP/gaHZMjruObMhCIDLHgFl37
1lcuwEJHjxVWc/U3fHMVkGuEmnIlNBabZDGKKcw42HcpsYNA0Si/pWOmqeD7ONyaBJpjU9jQXgt4
B9P7fwnpBfNSA6sYFblhn5PmQpkwduS47pKiEHFmlsIl1iIy+a8UrQF5TR1MJGLa8WJCIFRSXDGh
CGx//zhHD8JQNZ6Nm+jjyboMkzlEXZYblzBegcn4tddbDx5v/WtYljlLencJnFcoMSYrG/jrQnHS
tf9lY23PqyZC5iFWN8ajgOZLudjUIJiB8shEwG4TdXHA2DmsrsRySlqxm/bj+0xaJjyIFtADRryw
STo3YKGymov49QT7bnV+FUOujSRwHb5Sa+7Je60FRExlsOH1ygysa/OHM9ODbL32gTTy90ruxEbw
TyN2eSfVuf1MFYbTZOoRF1/VY5flGyiVwa5F1bexhrGopxkmJQO35aLx9ihj+ySDYLbJU4fEzxvS
zekPwEeR0Le07XTFBQ6+AgPQjUNJt4K8S0hpXeCQrX0WGUmGJBKOO2ctRNMVyeqMZC+e9DqQKzaS
scr09HJrM7zL0GmzcdTclrOtYw7OmqL+YcZ9OdGzTeAPQHMZkZ8jkGKELHigBXee1SqYKhJjRteW
cVrQeYviOhNLegp4n2/yOkcnYFgtqVrmQ503NSjyxaBBhIwik+nHJOwEEYtEGxpv3WJRzAOOGakQ
tbS9YA7MfDydREY/ijlz1jEFz0hRDO5ZfhZY0DrLSg7baA4YlyorLx6AS+onJQHJ23Wl7legDjxC
0eu67hXvnhy/yDtQI7kBZSZZCyjGSR/V66weg4YFvEvnXrFmpRG1XEkL3aRb5QCB+LEwGNwvDTlF
PWvmKaSK3TM6TJdP/iDvQ2MsFfEKVolkPFyS5v5qVmVzqdEBX8jnmIEZqFk+X6WKWkxW5605Zgne
3SxyUxOQdJNET5DzVKi1fXwwhmMgjUxzFFIREzVJMxr7XxcgxUd8kx+TJENl2GTVeq917qawV7lt
YqBVRNo5LCBieOtZuv2/rGGNwucoNxnPJUGMgiF3MhnC4CBDdZArHoWcUJhGSYChKbJN48t6qBgF
HPAHG9JIj0G7PHiTIV0xNcwrSiZPLdkVQwzR/XQUy+Dzzn9DXtPIeEGtsup3T9t+En6sQb/MUwS9
nngWxJDQ/ZK4etpdzN27KATKAJw0OutLj1MgplW59WgQmBUhx/ns0UILVzLUJnjqHAWGm2EV5zN8
36qIxVxgTSuX0/22AfujvNbni/pID2cjlCuV6uy1MGGyEuWLDC1jcFSFM15pDd1CE2MEEEHcHvI5
SrSFt45hEkFknAb8WMr38jPrSLHv2PhqWyb8xJ8QC+u5pC/8dGneYEp4C8SXkf+IRzxENj0ChnZs
d5UK5EDygKAVq4Zc+68dwCbtLcBGr6O/7P7JJG8a7KEYtRolodVxLSDEfNAUHYWGJerPvvkejTJT
b2GJU9iZ2LbNApZJFvHpIR+xYQvzmE8fd19PP/0C72j520pwr7NpTlquqDx05Big9BKmWCZW2/e/
f3lYZgZK28+gnqZDiuwCHSplcMRegOP0ctbmOZWvY0H7R5nqQD6LnRkxxt3eMUt2D0H9OzHNcEpd
wQmT20nKZ46qsLYrRmrmqbWuCeiDmTnNItn+qa1KrYd0bLfaOGnbJG7+Pwv1FBCT5e/ldDL9zdPX
XTuIg8JQ1BuCm5h9EI3VCTQ5JRU0SnWhh1E3O5vbOGAjEU8Wuw13KPrCcNwH9xJA6+bfMK74zVKb
7HK1rrWsitfnlCZuGaU9RgDOSFO0c/G9VQdGgmwnp2oeZZ4YrF6BhGZcPOKhPlOY6NkDBvwP9h/+
aD7ybV3Zl8wFWjdeQmzPKoSvkU1VIkoQe2gdCghQ6tZuXFUIB72ghOXJ79qhdm1g+0V+QT4cQaEU
TwM1QAUPQjm9TUS5dyUwbY8YnJThmg4VBqPixFrHoVPCYFAMmXo8IIlpD4AegJpKU2wyb/FcZj1Z
L6BVKvqIPvgyvXEhqRHpu7qG5Da/sj30sUJq1D+HV8c+P8sJZY+nDDWUA+kN3aVvM1y5Rhds23xr
1aB3NV/GprDC+TKLvWbBYAYyO8HZXVyjhoBR0ac0koJaGr3FqSQY20PT4gswYqaD5JLYU3ioQ3ee
JemNOO+S0Ze2tc76urHw8mKeqzZfcIfBYjH/+mHUzZvEDXkgWEt2pxHQhr7rbGKUpItUbjbMISCD
2NqBvYmhE2k6hXv8EYYFmkpux6x+psIW5ep5ieZaiFiNv16gXmKYtP4XqTpf8785X1WeyfmlD0qy
+rD8yNq5QkH4Qso2uHg++NfmMbt+00RyzND19CHye8jWwT4izEL48v3Q1qE7grz2NeZcj6tdBAex
+P5qtqse17MyrVQCYTNFYvHKn033P4zOwP7uKHirvt6OwZq+ONiL9J83k8RHnU8IVVxMzUQnaXev
49w7X0BxnK70TIvovRFmKZl+7shiVlIQClz8tbzNbFg/Fz5L2WD23Zvytq1Mg9+1CPRbTK78WN3C
ArrpLzcDoqS5RnmgdAsJLiFtnkoQlVWN6Lz2tRw6ERFg5+P8gNejo1mKUkn7ilOSsojrCv9+f5TJ
7+n5mAdyX3yyhBDeYy1yS7ppPCGpcAX/GUaLjHmnUe5Js5LNp3FSr7JenPwJ+vJeGqwNLzfR4XZa
rxN07c3f0RNPsCfeCU3FMX5N2ahQpKVhOo1kDt0Morok4yB2N13wQ39TrmU/e8aQ96ewyJppeyqE
bbgM6iCiEicoFHur76gt8v6NIhzM0Lt+C7QZkkCKucsnqStraZavILdsxBntxo7GaSWBCJOl/tWk
SvztLBsMnlzmL4QwIWSknDJT5AV0Wh8HX8bGlP0SD724yg1t7yFELCX5MGM4ZiyXy8gkehthm5Oe
cfmQTCpdvrCfeOTWJJRnlkHuId248IWRdpkqQl+SnDAQkEK1saxqqbacDRkfpbppHO+MvwgTSLoC
6VBfPkwuvv56HX5qlf2g0Fudtt7kJyvXzpAD25QN1mJykZo0oJ+r4wS6nLlXy3ugL9N50y+iy9lu
AHmN4JBmtf21bRbS2T0Rq78ipKfhdMXFnbDN+COnsiipFOVpV3FggsiM5Y8VAOJ2xNSaymnDYJAR
VfCHwOztB1xR4nLUvEIed/JLLX0Lg5JN2W1qxP0aYcabvmWArKsZPL9RnvLPwO0c7qIvWkBxfILS
XiMw00wqoCoSIOlu8eOUuD3MgNRZv9HVJpF/mFw8Xt+MBTFBWJzJMCCy38vj5WxozYWT7ZGI2wvV
DZ3NwdI8b0C55T4iGV6OvZhFKEflqJNNq84vG1y6W5oAN0S3VAgYs+tUHoSg9JnJ3q9jT1CUU2hf
k3FIxeqTYEs09TtHUEsLFo01b38Ck9fhYiDpO9eawvyp3GZnh5WXkbC2l3/nYFH4X7doIv/7WvXq
t+EM2zI90dUnewULfCgrcGmvfWp12aMTEAKIzrbKWLgxTPlIWe2qakkid1kKDioVCTvr9oUZPvEX
y83Wr3EkmbZy5+YEvkQZtb9HngkPNU79fJzMd3oEnpvtTKJLiyTlDZWl5QwTxPDbXo55VegFLGCi
SEij0ze0GIpvGzwlZoopfBxNjbC9g4sg7LIlMlaaHzD5+3EIE7veZaTN/bwYtGsxvsfkrBwvoiSg
PONUx7+59gFGxtV0zDNcIAN+uUXrLhBNGKTfMXdDd8Ic1U6TWTNsrzNhEu595SdJGCVl8cizJ3u6
kbKmmd7/yJekzqsQmvBdhfkRqZsZQ6UFVQ0BQw3/c+b7gYzp444QHLOHFqDYsaNPgF+alXZWIcSA
bJ44+ozusXANlMplGCn/Rkr7Sufdj1FOReg4FPy6QvIhu3KeEREybXm9Inf78nG77kcHYbrr/gMq
/c5xcSxcNkP4ho2F4O4hNByIv+LEM5oJ+3nayppDPiHomMuKNzW9Xutant+TrZo95G0P0posAPst
ml+sx9PwaMnoZL/iaiutD56uLVTBJIc+qnajFJl2oR3MOYoSaKvAkiofecM/3c7jhIea33yYVlKj
ynkhKaiqcub1NFj7KlbWdLNuX5ZZs+yNfGkSTRPgO8jonGN4ribQM1tCyIBjs1e9w0AF2Re3TABk
eXbLQQ/Oxh93EsWEecmvRSWffu/aOxS+ZvFhTl0SqBWfD1qpH1ovFrzIGfaFBQrjU2CuRzIn/432
t7jMMB7ynNFTFWzaslQYxMbzOHF5zGaIdeFeCf+Sh1CUhY7bKv98856+c3FMu48YRIImYwGW4OY8
0OdlWMB+QA/2iANFgbSzivDf40OTEYx4wJF2NBQ4mTjj3xf5ze3gIy0JbOOU5eQdozpQax7FefAC
os3X5rycD3dfwY+YVvCj+SiSTLv370JYBgSbmBf4feYmyNf772nR5+TaefI6m40sVZbrBUhW3hX1
clWKbV6TckU9/FWtyrPsolVl5KcPGOzCTHSJ0EEPOR2uGHrhNISVCxmMVJ8rEqWWqM1wqpClvogc
UqYJmuROCycoxUx91Kxd14EMkgdCR7sBKXsvE/W2ONxRddKTJedfrbHXpEGsiiMtKhNBXU5Fc+qP
YImKVjH4c8OHDNR4a51n0yMLbcaQRGVWsW7PcNOULqY1XIC2C2VQnb4vWAuRLCJvYUKk0AqUUPvp
gHRABt5ah/o+fW5ueP1PmRnGRAGSrSLan3bxQpU9JOIcfOgPRac9bJ4OYNoGFKienbd19fL+88DI
+OcXXvkq4QMvxfingsHSRAHxg+ErZ5TylIAlWJD0WDOmT0JtV1QkAOquEjKoHzWbn3cZcUWrKrEJ
tEqht51w89AEvLfabuvaM7Sa8vwR97kmt662NLwS6IHQeTav4w2lM5YRlZM0ekoLPSpBtm5j7x4Y
7tW7B+KtG3w4sJGBF6UZ/mtoey15bvPlxYKuiQgr7Dcgy2etVpmHCmiXdyIx9etoJ31DI0DHkzbR
iuLQGrkQjdVEMe285kA7vpPVmTcx2ICAsCu+CJvLEngvbACM1R3R3ky4l8tp7EffmAEtSVlWk289
QbEaSmjfN96muWToZbJYWe7aTId9TzeTyYCkP4Zpju2MkzcqdcQeOm5C05jZ9hsdfSuLZAXkgHt+
E249pZtNMFDiEt+XE2wz0WgOFSh2qbFgRmx9I1gJdS9hqqJFmlSaXdaTlhc6kMUNhs5ZAm7qifDP
JBsEmIFipEKMU6SROL6l5wbcAH9mv2hmIoDWvBctDix7pzgoFCLYs3ZL3l4E7gt6tzjrbCnXpQKw
kGl3NXN1yZOny7D5CoJP9Xbvz+CCsLln6XMTwswnQS+8/GtHGrV8jjHx4fnBKO+jgM1Y+1phSke2
PZqVIQV3zsT4xFRXFcOMnqMSAsKI5JOUfdEXKniiUtC9cwSQ75u3bezIDNDfpvJ5hQoadCGSQqFJ
5TiVV2y1Jq00OQoaU9WwgSMmG6HEJ47gIGngO7fItZZO4WrWxy4Dk501/2UnO5GHX/MI4IorIoRT
DUDjbK+DqR9D0v3CAM+UE8mm2wnnBTlQ/6X1YAaKN/dNrsTxwBX/KX7+2C4rw+L5KEz3sii79VhN
E3kzQ4LyYDy9ctLawsnU6Ym5qanv4joCMcI4Vu7ZyVe6zYtBvwnFs4hFQV43I5cSu4sNe+YxuTQp
i7b8eTox14SDp4zeezWuS1aJ6q7ZDPytFsllEiUhOhf+o8czzyPNkhM7hRf0BmP6UwcH+usLHA0I
rOoUQO2qDyP+u6iIrplNdMM1KLu6U+qVrDUCcAmodmDWWpOPSS7M772GI9iHiB2dqDjLjtoWR4MJ
30PyhOAxEY+yqMO85bZP9EQmoBmaAzpy/rc0oUpluux07XxJMavBIP512mF0Bvx0n4MKhU02LNf5
t+INsKLNHgGYqujcbmuGNIxTj33BtEoD6TrvZ+irI9SciAO96NZQQV9xucdGPzk45R+bwNT0QEuX
qxNZtj9lu6ysX/XH+4slRuWNudOKPMU/vwhVCDsO2hijE3FazzrkdjP6etOgIPjBbh7V6zIARNO7
I24PfK6YvHP8Tts/1loqLkVH82V5tuafe8NqxQWz0JzRjdtS7bvhVEQ5E9SIQst+R/waJB2Cppz6
vwDUIRBuGGabKYnp5GtUqjFiSviB7xFeEm3TnjX6lfe5CmULT8GSALbN7cGWamasbw0nqmTjUlda
MT1G5SB4Ce4sZLcbLGB/iie6NUTopWAK/MMSEaIH1Y+kk/EH2hHfmR0CphFfscWjpemgOw+p7fAX
ed3C9pL1YX56sGnkUacBhMbAonroQCtonF/t6Dq0Q1DPhDieZURoVuttlyA8B0u4cL+WvhaV1C4K
i5EDXR5eKJ7BdO+bHxwqq8LSdQ5XC11Q8PjaKPK++C/+2DPK9RvBTDnlsYXkRfHGuufTh6tRevWX
W6m5+6Q40Wn3yE4i0MLPKcY7fvxIY4woZDmQUKIN1xhP0VGu4+wEQjT/V8OAeZLdIU3ecyuG6s3e
j1rp/tEIPd+wOF60mjJTGCFiN2UmcRBOyvxgw8yAL6CLEtgiDkTnXgex463MgqcPW9JMKnhhkjAD
Fm1Tu5+EwuGrNW5gAYl06afVg8qLGACKw/73StHjRFeLhWpRXmjGJSx6i9hJMbT8rRrB8SHu2juV
Yc6PyXSHqt/+lrjoS1sESYGYX/OuAkzuGY+HswBfiHw8Fhox1Idx07WhNf9nmGvuetfV1Xizx0d/
UFqdgH5tpgjiThorevX8kBMcFOeMTZbyPH4n6zX55gHR6nkrEuX6V0a/7qBtpSM3aVm4bK7QAuv2
o2FmBYl3aDxsS/8YhUId4MQt+zfCRRoxt8AUDTgAYmRUPb/uSnnmiaaaAoK4cDOc9uPp7KhSZxWj
WtUII2sy3mwcWF3AR6TI+hnnsTVZml9LlhXaa+WLFrc30QW755UeLd4o9T+qMavMTaFxaXu2qha/
M/682oydWNnGMwdf1AF07IBy+V/LMUa/ihlvBLod8hvBEWEtNm2d8vIhkIKfqf80Jdur5CqYEMys
Tamh8y383nALCDK35cXpqhalqeZR8sW51sDxmJ41KqJbt3Tg6fyivqqCgmAhhDDmdI8vQIMO4nA9
oLY/QwqTO/AL/Gvm6xnf333DN6aOz2zblpgMhsvh2Q/WPmN1BIgjmB/KFfLrGO+ErvYp3RRUkRqf
rGyRGcDx5Bpx/vmETTiIsbr2ZZQP+C4cYxmeP5vcfU23V7i01peMKrPXHPeUdbK/+HHHFwIAiLGh
A9QxdEWtwRKaCAeU+EyQ1ZGqKF3l13CDYCkqwv76lLuJ01T2Es9jHlzuDjs+6p6kcnDaO7D1+oV4
79hvI6ZMuHvMHeSt+wL3ULl3TI+K5QdO3JqwMERtG53CSuey20wSOOElr/CldAf5pBJcLnGmfYKK
wmHdiVqiySnaahOXvKftLvHThXGP9JrySlm+my2Blmhhw589SIIpbYpevPa9s5ZEpyA4zYfRrrz2
b29vLEzPFXROtxgqy6obej9nDbA6Hi8PgWtq9n5Q671Lx7JKNMnuJSQNd6hiJ6xeFLFUkTSB4cOY
YXIxz/RtV9jlVnqaD2hLAom3vg6AcOdrYj/T+hyLUCiLpkeuPkNhd4t1UZuVrMddmhBiAq1qm+bb
VC1rM9TPB6FNdp5evqdfhEA7Hg8ZcoB91NNq3FlrfqkMLNX0dKxEF7Q7Ttxx7DLKLtUSxvk5h+CD
puscWpWfZf3ieJzThfE98d28wCyGkG2bVYVNRSPYZ1V+ma53tZCtpYi3u3xYvCysKH3THTqYzMIi
6KiEwIJ6dLcbUqGNvmuu4aHx6jIrzhjEkr7Iv5YAFOvp9A0fX1eUHAvCUNF6BG/GA1oA8D9XZdP0
+DcyRXbU7U+EpjCNBTiiN3RySgExU7AVS39EaOjD+oBBLnkm/VTg7F1DK/+Qstj3T3dbWAc2waTN
XJnJV6GzJNwmwThIlFgtq9pDisIxooL5TJNQJDWDsoL8xtNHrrkoQvj+QkQYynzAD978PggGRqM5
RRmsHocN7QVdHPhjjOwPt3rkoJVHo6paNVMpxqEvOgXRuG6AjaZTLVBuxHK1AHrZGSJiak99ldrG
2Gz5gYxBx8o/269VG/XrR5jZmzxdpXDyCqu6dGMFyROT0RE9HfQU/YI7KJSbKYOxbNFDuhQYYrZL
nCxjK+FasKRQuVMeeGPvX1i0qfe7ViKWAl/Uc4bsZPtdTkrFyaVXGOaJyThFJcCQ553glL60ZL1U
Hix7gkOdsKKw7V8zzoN4iLUquAB0e7yjXueg7OjHtBNswvbgidwMnCroTtupHoxm2oEqYydpK/N6
XzHcrxCGR759Z1fyCwkbrVMcGPElBGmFF9Mkzg3IbMj6Xrxw5CESrJiIDFne/F0gDzBque+uhW0k
XxBwPEVfQYjEoCao+ik9xC3KXICbO7nou/kM60jH5puyckAcpOET0EqsnbJ6LrWRDDtrUdRWJJo+
d283rp2fgqLSa59aJHQgMlUkY9ZvLg/maVg5rXSwUmiLzyB//H4AORpxovoLNy8YzL2p2GzHT54K
47LQ6nF6XJWHD+l0Vv84kJDW/qNXObNUDcVNTwZnDPHt4OhkUqmMdKU9vStrV4mrcqRnB7RA8SWo
OrS3FlvMnFXAPlipVuGwjQepivtmYXwOxTOyf5+234Z/LX0s96PR56bNwGDo2jwpa4zCWdq0Pdvw
JMMrJMeWcuaxSvNyTvXEgkfx3PUVrpliJuAYya4pF5GNTjgFKeCpcUdhv4N6WlfJFGR576nHp99d
EsWc/oYWcXXMmWYPVfg0HaMcFRMypEfnL0bmMUCfhIcLtfIaXQbnh5hO73cLHzE3TcEXm8CfjspN
t64H2X8gMw0OuTgtPYq5etH6elFK0xOWXqgXxzd5kPOTsuKTutr6Iq06UBpUmQRD10GaaP2S6Z+z
woUEcHR+Ub8+0AoTtTWTIj1MGcCmJwZyJvRKXU+NrmLfunaIr2EnGbgEe4nY/K0vEZSHKBXz3cGZ
zmIjCc4gBznv2pjZol4G4N7rPn3gSpL8Rqs8wMtGs2ja4IiKyejlbTp752MQYnWSwv1HlLNlGBam
imvEb1DhcDZVEKyNhe5CC9p/7nea7PGiNBa9RejangKmjAZslxlYbtAyqTqxbS5GveaiF7xrBuDO
LnBcwB3k0mIEb9MWHiFdy+7WGHqjTufoRV8aS3+aNCDsB79nSEPYaubQbc5o1q7TtWgM109+V+X9
Wo6JwqhPFMvUJZlRhHRy36GVZQxMBs+7qA6gv6ugArCcIWDjc9avQcDMLOLNHq48VF3rYzkPP6sO
SiYpOSBOR3SWZju3z4pjhxzrUp5ZoNnjchibIc7nxJFjrM9R70e1nB5CYdbAOAeb6zt5rQSFOi5M
bC3nCER81vwChFk2UpCeqlSB9xzWE1pkqhBJROJC0dOLhEDv3a3yKwsT1ouZ457CWd13f0aWHAJH
RK6PoYz7yfnejSvxUWoPRO+yXWuYXJGJWUDj97+qNc5XoKafgIID16DSH1eeRJajnyeeoGH7NXN7
BIwtvQGvrKjyUsfuPBuYJ++ZXxh4oI3chlQtKR7pjQxtnaBg5uufqHlPPRqC0R8J/nkiPl0mllY/
6drFmm2Asmo/n4R29erHZsaMjkw6XJX0yV0OGmegz60quV4VFngPTF69Q+jCyyz9gsb48GSXulaC
WbS2YTf7SFqY8ZSC43XVRJLsDd8eDWxqUQEhqy29gHZkPDIvzAdwOKgRFaQjuLETadjTChasbhtb
M7GYuOwNw0RP6WwqSPZO1f+iHxx7VezmWjdxxfb9+82RkVPZ8mJ0ct6F83k0MqBaRnA2KKdZBx5g
FCZT2H0KLBYE1pLaV3P6YfT7/MKr37fvMBauNpskW/xJ0gly0BMxjaXlnPVdkRgtogygNUJb9KfK
wOAV8ZywdfkKbMBDPCYqDD7i6EKPArdXev3dTjHnOhOWsb2EXf/4tVbBQa1gE69A9tmWtS11wo8H
5P1NUvnHQCywOwRiGOcqle4ORxdQmi3GbeYi6BRhnmbu1yKA4HdYaHSdUZQHnBiXZuX0aoNUHK8X
Nu/VzvkfW+i3ISZueY57ttB0dcujrexJD/7qbr6lyvTWN1LGmxgMIFMgqWQQQb3+pwUlxmyp6/2d
Ownr6rDbKgktoIVV4dGOWqIMpzMbbKRBcW85n8GieRcYI5X6sRjPVgRaknPmZFt2vu9Fb0wrWu/C
fhoB+gs7ZOBZ/e9fVR/32pxm3Lms9/mOD9zeCybi4Bf8xUtY8R40gm7pDhJNNEa86zrbH7jWSjio
ieigNAh5YuZNvV5jJiY1d96hz9UVVNp4GFy8dkqHEmOL4He7/fpW78oKAhvVOgSxNMprQgZLXgbT
NPvbIk4CBr61cWfK5GfQqmVyMLoaoJYlEvga8i5lxAo3dAbzD4bKUnK/VMGYiMPvcJFT+PaQCv1R
+lOt1Rt7bLDysb4xP/34EixPm1C9ZMEqW4DC9ILRoJdgcoeY3X7wMHYtXS1bmMTxDwHwdZCqbw8U
yTCTe4jHCw+6lSjiYAfWNIYXj9JfrWsoZ4XJZT9L9JZuRDOnP+nN1sQZuukBq13By3+xvZA9P13+
ejDERNm3WPM3pMRzAGbIJS8ZTHG4HWyV63SXa0uTWFVP68SG6BWkz0cg7DLTu1BpMhUGvQU8NmGK
1SukQbzZy8a4pQQNSnICLW9RfVP8264n7lonwOysxn15K7iMHZyZrX6QB18d2L+eBjMZic+YmB3c
ahrxhR7a3z1ruhkQ7El55QZzPZwXwYYaiDum35nkp1w+90B8DHv6CZBBa9gMD2MnTcfulSfftRTO
ZKz9khe+MIN/fbpAdvRbenjQT5Q9+S+9gYtz89IdCTtjPY12+4ni244xtg0G7QtJxhZ4YjkEWaAZ
+IF6gsnevYW9wrOFN82o8ASz2HbR+Y1Ar58ZSIEcKsB4M5LplDteIO1HPVJ7DsgYpZbJE1nh2XIJ
B8XaLXXLlhcUaKp35Ui3uUHksMOzu/6PELf/UUPNnAwj2YAiN6++/hxfdnAra29MPg0082ouB9HY
gYZxwhksk7nkG7npXDr/m4nqmiGeuJSKJ24YPJUhLwWGY8pKCbcjzzGMEpQID6ChgvjbWhTS7rAy
7XtrayMayIINY55WvM9rDQOB82FFm33Ras28qpPEXUajDsUtPPAzkwbZNfn95epYOQNEwoEN2hK0
3bJYqdBSUm8bhQ4ZRMTbCoqimwKcheoMELiqRsG/G1wCw4LYSS8msa0IJMADdBJ0aNnMt6Flge3E
6gtwS+4zNU8owuOr5ul6OH+0k3m/MYf8dW1SBtME5YuN9i4iWUCqwXXi045R+6wTIwudnr3W0kQh
M9XyFo2FotbUtMgRydwq+iWyXIRDh89ewjNKrcDaucscq9EtR1eCpWet0FBrfC52CKE/UtI1E1oA
D2D7CBk3/Mzyk+jsu77s9kw9/op3pi0tUfetTXw7ruV6s/iY+T0xO2xC6seoFu2IegYZGZ1XAbLY
tk9oclwYKEn/+KSLRo4MQLKt1JoOcrwuafugiSvfdAsijPxStIt8x01cnDIHIc1yPBHncPC0F92/
Yv4n4vB3ZG3Q/UkoWjXJUUvFhqBV79OerSs4u5WxPKJ4G2nLOG5MfIQ30kC3rGmARpA9IJ69dYve
S/mqFJVMm+EyTUY+wIB54NwrMGeWvY0SvtdBmuse6UJ5RUZvq2oapxG8/JQdys2R4y21RLc/ai9x
LVuuxDss+HsYQiYdEqXSAZTN9Fzc2r0ns7GGy5nyAMj3SmV/5Rv9tOXk1J6BK+WgGyk0rrZ+/qft
h2t77tioFhp1kE/HzmvzIDeY+N7/XvBTwnfJ1rtS3iJX1Us3MUTXG2EAb57DBWRjf9tb93eOr2Jz
nULeLygG337vtlwJ8wgGcaDcBpb67jMpZz6fTaLsMHCG3vrH+4BNXHmC1Vp/vRGb3Gz+lJLI6cmt
12FIWEagpQFyYmjjfIFrkwwXV41jDsQ/c7bGIJwSskhRkpQz4lEeSHX3rbqhOgT5eYrDnedE5TLI
RC70tN5mg9hqjAO/92Dz57KKA/rsci7I6ZY5NZAEze2pw8gEqkogVV9eH2c9Lh1BCCU+BIMZlItR
uslrl06t1g2Ieqf/bR95S4tDTq2uBPy0btklsl8CNrIFGt5xCJxSzqlbPXzoAmPwbrsGTv6xa3Ea
N8qL/j3oHVmy6I4dsQZ4UF7wz8eMcjCyBhPyFLxokwMmDl1zLiNbS+Fh4VFIyVA4oLcmQ1xYOMHz
/OSty5tOsYUEUVzymmVBq0uRrfhYyXCOUR+U2CZtw9h6lJX/uP710iVJeZUadroTGnT8RyL0YX2a
3Y0+ckTHtLcQnolJnzAgMnJByLHqnFFXznPC7EJbBwrTw7XzgT7iKhB3RYNlrMALZfXJCVtIAt2Q
RF0bBZzVnl6QbhU3yesa1R7HTbWuQIVvfYDE+TaAjK5RGjyOqERLRdXsKmGSAMR3ix26pwjYrRJL
fImSlZtNctCCJxXDiyFdeR3DfK0CT8ngoPIi3qIu4Bnsi0ViHmzseM+YJ4EuwCIod4Uq96GmXTTy
FOnQeqGXe0cEh29Kb4CIp7fetR0+EzEVUxtvnDB6wl14A4RTKL+1nBk845n/rpWvzaYzxruaGolk
dHc2/58tJgWnHbm0uz5xmQjV+cwDsg41ywAqUq1E0GuXABlO0JLR1IsfbiDWWWkC6IFWFPKUmuRH
M+SEqJh/PwzK8gkulqZqRWoI2CXH/ki+IXLGwyEd17QOr/Y+N2G95dumOabjPXlMH5Z/IyAewXUT
FBJdp4U8bebzPNh8yo3dNNH0Ye8tHCqI0QS8fB7znhP3g/Kg1i9rWPDO3wI2xy392G0AN3T3rB9x
F7MJASCki4M2J7JX94u9Gny7hzx7JfU7OPcFst05X5MRFhAg7RfT7dz0+l4XxnWNQUOfPdC6vlYk
wFe2ti8kKdQCjrimHQs/QVoLpTle+GoSHwX7JJvXX31/HQNFS1RIVJ2Fhr58GjHF5E7q/PkKrw96
Cx4CZvOZIHdg4hEbvd8eSjInAnWMtiAaVipCUQA2ma6MYhyoyIslPM9GRAKufc4B1FfSUELTEWYs
wOvDx+vQd6rkD0M3JcFzmVjjE3RWOZ2ROJ4FftxQYqXy0ftASxZhs0JRWwdzay/8gw1DdQ3/6EvP
Z7+3Jg+KuHD9uUtrDQ9FRRo4ngFumtr6Q/F+1bbEQQV87fx73k2Z0wM4HT5RfQVP0As17rmk4qCH
JAdIfpnSCBcUQFcEWKzKwVXg8kXENkfwwmDaz8AVfG9tNFvy7xrDj8FERigZaMvG2ADMWxD9QyEB
DZDcjOdlnr15X6BLP//x8CY7hmMUqNvKSMlP3IVH4NMuUBU3ZRjnNTTlydqCiYMv8dBiPUeKaGXR
uXaXqQm7fGJGS7Hz6s+F6kcmo18+eZMpEHfw0lFS2ShmnrsRa4/nmaVpJP6EzYNCNk31O3N2w6Sk
157mRrGlnNDH2uOvGkxegkHgNevcPivVCqm6E/3SjD/KqH/9c5wcH813Leei0tMhxgEePZBLIA/O
TjXC11knjNAjao82CjbHxgd9CbB0OTSXIRfXcpZqQJ6o9lG1Vjx7vWJE3c4WO4Yppfy4fIi+UmM5
qQCSTSMVUXkrZTCc8K+51vWGlp8xtPTfK8BpCZ4pW5bTN+f0sD5u/XiogYSKhqP2aqVqvXM/r0ZK
uemgD56Cb0WyKJL0gHRtxRyUok2bfh1t9ad6bTTqHzal54eVXqpUrf60HCbu1dXznfej5TLXg3CN
lQBkv6rdC6MyNawMaNNDroLrYaqY0NasW73JyPdNcUz+qEgekw+w57ogzpKYc647CnFZDW1aL79t
HXDf4cTkLCIpMalXIqLA9G7ExEWBrgwk6722OTBkCNOMnCT1HjTzNE5UEtQyfIUcLaz62xpriP5r
nDWsfKt9sMY5s8tn1UvFLf8m+xC5K6CKKhU652voGvNUK9JprPOnTFIc50HpHBleOHRf6vbP+arE
+wqbb98liJkko+wlGXGRhbJY5FLnU0E6isBJeOAO2rEWFPnxBSYxBigiJA8WVGzj8xEPna7SuFhk
SIKYmqq1HVmJ/FIg7xeDTvja84Rc8q5EDAFFxHpjBC8u5JMFAPP9uYLun1eC5cDDtJ4y1jGaDf2i
0iqGuFTxeKuCsqY6jylvmVxJhFqBGWavDKRMiMK3n33St/SOre+RxkApfnwGI7SIxb6tluoulr6m
XHRDymofEsnS0t+yPWsewf++XUnF6oYRbxIHJ3UyGQJXNETGTqkLxViZkND1aqqXyBn4BOE1AHAb
8saprvWYG55niFiqfoiYnQSOUptygCtCzQk8nYkG1AlUr1IjdrcB3LF7HDlmcVrVmNEf0wsQQO+V
BHq+OV88n54Q70m84JrVo7gQOT083mmxsEWhM/rKzLINT0wSAKnposQwgwCtY1UnuNkRMqVcytWL
YLV8KavyDqfcQBpcnaTBY96VygVRGILs5rNXnr6lmfEQ1nJyroZVRqHwuSoHxjJs67/pHtH4LAVl
TBa40h0DvBTx9W36jakrSlMd3zKRGCHUhKTQuxaYz/t26JSZ0UlF/7FlAjPcsOXe7f18liOk4HmO
moNHQWGLxBf5DL705kgvGXmLSPGI06r0iuVwa5G3ztNb2qvd/+bHWuvJCNIstu8pWvzuaM56XZLR
uTuGpad7ID2y4+ZiNXzlvWKqk8gZ/LEb0j2urCwehrzb1gJ7QbFOBb1euz+T1WDXPi4ILjiJcC1H
miKGe6WpVVXUedcaTf3yfuOaPDZzGtRaU7ZkufjryPHDMtweJuXn+m1VEygfON4SiG1x9ofJRtyE
bNI/8hre2K/3gEzBxBcmeH+kuFvVkvkjhH58SsuGmlfFunQghtOanrbDQ3jByHQZAOLJ81A/39J9
h6TtBd1zZfzk0q+G68qCCz/2YuMmWu0Ilrq9IEs6YcQvIowHifm3/prhNzACvQ7RARsCCG1YcLRK
mp9EvFGuFUrBnnjOkWdmQDxKo6Kk1EA8aFg2QKiuSD6Y1CzARQrOP0uh2cdTWrbgVYJ0HliX2JLJ
2rQp69Qmagr1D0PU1BbG6AqUJwMOSHxDMf4zVUtzPqNWtT/KwjakKn34ndxoxWUmkzHWObJQ6VMi
HSUVJLrgM8h6WWRtAxz95/oRZWfovDAWMAfZRwN31oZherad3Jv254JL2os6+tc+HDYOWCICcvL1
aeuBArLGAVtUkFUjjeka5sLvvJW+/+8b/jXqMLB8VHka+ljzk46LTfn2YxLnDaYL+zxp4bdbfjsC
dhqBuzrhILoegQh6ZT/g1L1IupBASqVwnRF2fah87SVAl51OAbl4S4JQxWkT45E6bNGC6H+pp/Ro
0Ad676yk8GYKB8za6MvzRWiS7dQSfgOusp2+yXzy0cOu7ywmzzOEllnkNOA2P7r9J5wTpn5tvYQp
6Q7iBOqnYWcAJGlzYEV1hsCRBih3nRhh7K9K8eOIYLt2iimi60OBi4U9Bfo0Jedatzm3+fx1yP8M
Z0Z2KaFuL1FTsciMrwza5Ylkv91NBW3UeLwjV3oZqNbH2iy8sUt7iSNf/aT65KhzADqZGFr1cX2g
XsQNPs5ir48MuoIgouGlY0fjTbX0RprsCbxWzkM1pJ6TejciihrJ3jcWRMd87wnsnQ6IrPxsYzaD
N7uE3/dB465ZwOPEAMZiMNjlbT0PX1MG8E4Uo47vsa65Cgdbt5oyh/Cp/VCN3prM0JC/pUodM6Qk
+SWddn87xUEguf4wThw39vn45L9er9r1/ecQGpFKmA9aaHDyTOehnjmhdVam2r/bIFcoA+vCpv5y
sFjmAoNudI9WuzOSJdEMC6X0PXnl1M2/7MiBSetQWrW4qP3gT/cOeA20Uk4/DnhP/lH8QMS2JAXm
Al/D0eAAbL/9IcAuTDoEXZYoX5iC1DBDnrZ2cjSh6CtWFSY5PkoYFuUnKC34fO+gsZMoFCGRVwFO
T5N3D2t4f5tRcMAxE6R6FW0rXgFeSQXV31jL6aZAw/Ju/6vB+mf7F6KQ58V5XjUepU0LYmUrhFy2
zIcb2M0p9vGMq/psNpDOlq+9Rhtd2ttEEwQ3Ns8vhiCfBxa8PTyAXVyRqCFhM0Fgj+o5iAbAK/D4
Bybxpw2HoKhwPv45bQDUHDheTs58PAIDU7zlTN3/awnNf8pkvKiKvVeAQTO6pgaY4/vPoyWM/9ki
YMeY41j5JS8FI+OSPqZ349xFeIfGE330fesE7AX37EnT9nrqfh2zLjNmy4780JrzTcfz5xKCEWRn
cCFEuUQ22yekYDSbn7oajVksNCSPPbB8X2yFCqKKBMesN0RoGLu/nj93HVUV9+0omkuUd7SBxBqz
YLQe9u8Tu5SwXBa+21pQHmH1hCwLe7EFhkMPTJUxQ9tR43gpvHCd8y7DtSQ+lE8XxZBRGyw23GgL
jscSZD9PX89IpuJdrg5okRI3+5WCJIkWwVBXZ6aJh+T3k6ydwLvOx3EPaODZYHKIxKqO7VzK6HnI
4s5M893I46wWXJnFr4G2JiaV49lkFpp5VANp4ghWca6/iKaaIjolvSURCRU+PqtLM1+RaSnXEJ6m
KhFeihnx8YnRbUN3m2+p/XTIpKOYd0eZbwe3Q5qaokvDTgi+uSQW3BbWsaxTV8So3Wq5kLd9vzLi
/KKWCDT8l4kQRLz8lE775+lkSz1IdAU2ebNjalFWXsSVVvQVhuNW6LJqILlSPcVW1fqOgsRzuRow
Co42d5g2tw9LwUugtwpbfha/oE7URhRFfxFRjugr8UKTPHU5TXDVg2tiK5B/yWphTFHmX7lF2rzm
4SK3AZ5f6ecTZSlUhFXJE9XRYG7pOD5Jm2bgIvMVQBVdADoAymWOaUq3mLu0NqTdDhBnLB/VQTPn
I/2lIZ75mtxvRuEa8juXh4V3Im/zNeVWnD7x47r90Bj4F+Rw16rSl0/1HqnsCNOoFbu5a/MZP71i
uAEtlmr6l+gi8bL98tvVsfEni7STHAF5MTX4l0w+nHX3Qci4QKrugwVzxTvIovwvgsn67bGsHHvr
FaV010LERzh1HtuGUdeRPqq+VXfG9Rd8nC7kyXQnjWguweGOIe6BfUc50dMAvyaRgXe5FZInyBYs
vUaJpWe98W30tfT/hy6WMnf4uxeSfp2u2ldSJ9FpiJN9w89OiHTtl8x4d3kGRf5Kj8OWHdf7D9Qm
M4zJX5eGOMbkaAzIWU3AZly22WtyK2fw1T7mVGZvlg4Yul12KaW0B5KsY0KxzNzKG+U2gmUQBbHc
CV43PEUzxX0T3FNC/IY+trBfHlcXqwxNmDdB7shJwVJBj1M4paF91cdhvG06FIp5QxIwvtbWePRC
wUS7xDbEy+3pEDRgDn1HZaZOiV1EwCUu5oVPXoONWHQ30BxK1sW329Xfx9ZJFQCeWO9TJhjnLDw3
rmOs67RvD/+daZ/1dMcnc6Jz6Ya+BS6hSRaHwgWhD4pNHIk2fbfj2gowyRj7aAFcpX1Ro6GOK9Fe
Jwd+B3O+wBpubbRDO6Dt7I6QuhNRQFOFgzA86MS3rxSFXobm86ieLnD37wGKfwKv5B0rbY3jS08S
fPb+cXe1fM4HFOU8GchAf2iRYlcUgFfEubAG4diFkq69Q8S+qSTiNVn0rWP4rbG/DPuzKICY9L2v
KCjk9TIZStO8JXrGQ8kgRej7TohN0/BX3BelR541E3TVs4N5nAjKj5pvCSSezO+AwtU4ThhbG9aS
JMYjlnWqXKSDuyv837d4pOvXqTNPra+KhMufrk56krzPxj30P3MmyTDzbXfRDi5t8m352mSaSklm
V8GGz1reJemFQejNJvPrb12H3kYyzzkTns/uJu08tUfQ1dxdrLz95JCqskrO7PVfKtaqycFgoScb
SoG8BtoLHMTbCPj6lv1fXVXzu7Yz4F65tfIdioC+AMrl873byxggVsQMbb9xlci3/eErCj/nbep1
ki8okYBVmwrnsy1Qkt6ktRgIQwT15/nThBpxtqnGWXYL4ADs+G7rdi6YyH+TgpEPwhhJJBd/uNMd
avXQJdkXF/eAK56KZSCmzFuDpu4qyq6gNNykDR9CQkhVkg7BoM0OlOE0CNwRgeZZ9Js6X6cuUviP
VjC7SOZA0267MLYDBDKGEQaCOcXnHkZrrU3V3btqoguMxRDclAaWDbPBbRFTbB+63/zcjtvZ4qiu
X+kqPLNVb5MyaZKAnpLmJJABkJukfpJADeqJz/hxchsZKIRVe97IgwZS6UKVQcE8yEtWUnB959va
GAu+50EedApBYhIZ7BKhDqO9MjTaec8s2kqz9ZgpY91Jt7GfA3NgZU6Pzt5SLH8krTxWqlhthwZW
zCjMnNCCYiMt45Y1mmuDHNP0wU5iRNc8iOK5bbxDo+9rPNP3JEQrAxAQ8FoVLLmFqTQhTmkrgrGL
IrnEqzyklS8gyaN+FkiKO1Uqw04M2EKYJNxVQNfURbOTxrMdKohBQ6DP12Div18Uyb0neCAaJa9F
nnVpXYYmlCKTBwfqTONooGsngXvQgy81OitEsIOcuxUcBxbuEEDEzP27taWjthDBDXZy0V31hWck
5N0xaFGTF9CPzrrYSUchV0Q5AquOrHVf8KILsr+frfiOZFkQ/CV3AaqX5ah5iEZnlSRA3JPgWt4m
j4RgLHRZiWoGROa6h8Q6ZSbA7PVJYWLEnTLAb5dHP/SF+Fmm+JfdEJQXTS0hsCa00w+LN40CH1Nl
3TafVbfrpzHOOWKqRTei1GrdRrM8v9t0z7ee0qSrW9BhBgXoiO3qG22rw21cFvBIQAe5gco7qCTo
stSJCdUYJ9zxl4xgrc3Q6djEJmEJciNym1l3QKg8DahwfOd2LUdZksZpFzPKEZj2mhR0c9Irsw9A
6jDnyPDovvZVag0f0GcO97IPXvx3kAAn3xK7x6TCVAJVjnZAzk/Fx0OJnwLYqgQ4y/Qgh7hhbzxp
7xKmvzf0ar2vyajiguOQfGSzw1le8H9+ArbUMZ34Aw7Ep/REFzN8zpmmzsGRU2x9U89//cwHPg9B
HmeigwllS+wBM0jEkM24IB8CBsX46bMQoQpMCmHPcRj8mg/U8CkqXPdOlfHTeBHzIXwoTOl9i8zL
8k+daNr8tNd9DYE2ybgPEEzPmRQgFysnD/tl7nqPfPvEOYG/Z9gkuWz0Bc+awfImHhVHLDt1apa8
c1Z5APCl04j1As6bo5NMTfK8n75rsVY1q+ODLlHQWWdsjUYB0ouFDsjyrTM2sNGaQXtDB0TzCVjR
tsXmQV7N0SEwJ2bfRgZO5QwxrgYJQ+CN97uRB3R9AVxJgxuo6SdDM4BRKjM3TBKDq4YuF3AmE0wv
+Vl1+tHlVWWaJuXJbHHItdf/neq5Y6Y/LhJL3s6nLn87w3q+SiuRUf4UCjFewZot5hNzl7cyiHcI
THvJQIfiijduyOITM7Rf4TNlxo5OAKThg49PmRbf5PCQeMhgA3PRvDgPvMBQpOxjf+8BG7TRpBsc
dvhOod4uykl4eIuozdSZvpbdxAz4VHYw3bII/d7tA5hpXgf7FJGgUYPc0LFDZKVHzwOlvof3Y5ou
rcG5cqwvMbn5fWHCnh6t5+z7YY/tje/+kwBtdF1fzfqxwtJLNMGmPVOowhsOBrtZl8L8FCwRvqsK
uU27mOU6omYt3/vAYGXsT6eN9LlTiREnZjzkuS9FoM7GKbcCvxZRAXl5eow3Epe8E+CKrxf6Rxic
B8bou0Hii6yV6lzS5fTbV70MsqsshywZOBszZYzOhGodPijHFSaFI3J8rXCYQRLYvA1ry4JN1zn8
54mRkhkfsLqSJBzmTRdvLwHAIU+p8DIsNSV+ad4YrTshcyRmFhKI16WbOssCo8hiSmxgs/cvIKxa
dYNh/v7vJiry0KMqzziB95QYgkp0Xob/AKq5ImOBVJxXKuzSNPPyogLzbxbbXNz/5ceC+2A+IxQn
b/C+KwcoIW/sTweyddKgyzg/Iz+hIZ1giMxaL2JCl8cWyKrblPS/5q2csy8Uk3UXVT9+bTMbUON8
ed/bGPY43ZOQkQVpAq6CwOovvwvG97TBBHzJcaXiG5/+26jkVY33IxZ0xrgC0IgetO7PM7++8Et0
XG+vEJ2iQFk100Uzn2zF5Xy2bwC/Ckcs1HnsHEMNKkS/V1NyOMVTfgKVCsAv6I5joE0sVNx+Q0e0
CiJk+2iPe6QYv2jMYIUdGVGABo4Zzp/YDn4YcKZf73uoVPs94Bl2gwnSj48kvS489YFck+RLWPxy
PCmUmcDXSIV8Pge6629UEhAZY9E3OVcvj2Gwpgh0KfEpdkvgm2N+CScJgbEYe7a6ZibM40D0MPQ7
HyCO5EmB7iwC3uds2UN9ZPuAblNeExi+3no+odZKfS840aCaBHI2OJsXfuOa1AjK3eL7Oz3lc6iU
SkxNDOmcLW/PqTjqKjUpg0zGjaDCKhHxVPClU2Xp8IJ5ejpbienefb7nsCeXIq1yjNNirzr/pch3
8Z0zwWJdIte8fxGs1Q1I5LCF4QF3vYeKFwYQp0+V36KtYak2LbGi60IWDR87VNePGtlr7bfc2N8u
jguC7XMdWxi+msIZtPqnQGswuBVNxj7Ny6f3g00wJ245cfnj3cDgpRWBPH9NH8FzcpOsYhhDiE4q
yUxRwt8WIgf74BEqztr9kk/ZYqAnURsdWjlg+igYvzRhnEuwMioSr3eRGvjuCistbMBjbGR6U8f4
DkpgGKr4hnkkvHEYr+V2yf1p+TeyhtFSvpkrvkUXWIHwSqyBig4GYFx4WmeCbdgmfquUc/c0oMGk
yew/jtFbu6lN9wFJN5u1Aha9omiNjvuQr7pHL2IVIss1ErQ57277bPKubZGz4r5zQa5uquv4NfWu
CTYUdZBBsk/QJ9FdZth6yHFCTtuxmhmvVvM/Bm/ZOERwvoHa2Gl7uiIi/0w7bOAH9zAJleMv4DIY
vdS4O2hR5cIJw/LmspsXR7CJyyFGyR1QHdRxbJYlhFEsEfw7vWLQLBX5YIxk857NekY5hNXkRjt0
8GE28Ql/44ZiFD//qazmAVhSj0S2+R+wmZPRLGeWTXxth+3eXXwAoo7r0M3zPF+hSDpfEN/E/96g
e93cx0JEkgmSQY5fjm7dSHpA5yPeImmrDCTAbR5aG01pnMGiSFE859oUEDHH0D7mva4U3C8S//zj
CXfGHUADEoLV9uPBCjRm1iwFOjxoRxt4rvB/JvZo5Efkip4s3tLnn0OKaPHI4iU+Pwsn9CDVwrkv
tEQMYLb/If/gj/FFj0kBQwyOTlL7NweoiHEyeNrQXPjGfpSu5IZs32XmdUufgUTzyGUjed4NuJ4B
daEbx+iu1esm97i6RlcCfH0bbACBKVgbA2FMdjeza/aM5Vzn0xx2+kZBtSy1BtOJ2o6lJUmHDomx
ySFKxho0UjLfWEIQOmOaeQ2XxtDqdXcO05dvUZci9WiOFdpeqX+03kyayZfuDcYELL33SV/tZyjZ
VtUxQTobCiURQ8t3+81gLCKe79BIcA6Y/9S5b6diTNsL638umffDrJEz++8QsBeouW18Yo1kCGsm
kc9rxZ7Bw8IDCpCI+fFXMvzJN4/TS6ezFI8ZBY2xnfzWZDG8U4x5nJm4ZxHFFSijOxClz1wCvtQF
DiEpXelcXxkTuITjpzxw6+j9RwGSV+Vh6S6NymV/LO5p1oQHt9TqatDGrfsq1MJElGggIJpGK5BR
pc9q08FUyG8+NrkV7msb1uGGUy1nDuFHrxwCcGxIx24SebuLw86PJt6fI3PNmV5iekS/NXms/S3C
7Jeecn2Boe1rDTtMob+6wY27SkoJ6/VVFprUSM6P+PM1vl2zS7IL3szt9MLV2qruBnNASJjl+Qlm
mMfR5/rI3ST9WTfb8zn+yKJaBI5HdmLpWiOdbMG0iLikoNdOan93b7fB6cDcZ++J+90biIvFPSAO
UTJ2UNNxqYw+uwl/vU6yB7rXHeT1o0yYXc8xRO6ztXWd3UMxEO4afqUXx5eOV5BKMuuQhfnrk3Qf
M1pRogkVOTF4Dbzso+RACu5uTVrjX6NuAbwgD02uSlrGMqPcRz2M8neSKVS6A3y5OI6egq9/XHCE
uk+pBVFiRDf0YOtIUDg2xUKHRC2EiQooNGP/sWlYnj/ARqTipso8TBbijcCyXR5vMD4RBnR5qv5u
m4VQ0zrkCGZTmq9Uw2s6qehV+iezvqnGY7eS+y8h6W8GPSCXyOh1XJgVpzaYh5m9TkRAt/1OYD74
rtNmZOVxCOPTJqE2otN4eXzZlXeKvBWes61wWewSsnKuEN7m/x4WxyoG044EIIG+5xpZJms5p4Xs
oNPb9FE736p6rhQ2jt3/Tii+BLzfLLGOcXGVR7050e22lT9YmQmSB8g/QQgVnJzj/lnI0XZBxFqY
vnOHwIWt9lrawYs7j2BWWuN21EFVuYl3OOSFnOTh7z7bGvS51g3auL4zDLi1t21V2SJUQvdjngA/
dfLJvQdJkrllEBYBiJ5Dk1rm03YZpN5H81EUtsvPqOBnHz4/dyHevcseIXzFH3Gac4WjPXFU1RDH
RygvNRlfx7WM0sY2xTY4rgP0bDF41sp8DFuqdxt4kwqkUChUoxzPm6wrAt9SAnaqrwZwfsdItsNk
XXuMXy7LoYQkACqNcejOOpzo6mguSFQrahFtbaoGNPDGYcjBK1bviVsWnwqRhf7ilKv+aqa9D+PI
HegDTdEdJ5ghfmpD+TD98jFjN01WsVRgoZXz4T/MztkDd87Aik7oZLl0S6SzPr2NNh/W7pRjGAaf
LJqE5G30lKeLfTnsxDdUI8DCl8JcX9UEMBpY3y5id6S2JCMKjn46uzN8eOo2nZsaeumauuePAf2c
V6f7E/JxQmQn1skis7649UsyGesJIOebZPTPKChFn0dtQZQx/Ike8MvT/AW1xyl4GN0LcqBVS9aP
JuPdi1lJrE6drxuFZMrsyUirKebQOfwBxqdkOhIE4dHf+H6zgVOGpnF/MXpueEJksJpB1Yiniagr
7kHt0/SF2mMmcX8rWY5XVHhoNiN9B0CYqTxSgCFHfWp7n59o4veke3EQKsOPDwA/JsXcz/URh6mB
Mz2iHaCsZZ3thGJWWbcc7jkDQUNAVAlgviKFgomd49KqUeHA9a4pY9U4iJja/CSNP/O5lg1LUcn5
qBFwpgFsXhVOkVcjpVlXLIbZ9X4B3F5tsMETsV6ZjqY1jdxjkuxsbsqJvpTt2tJTlWo3JWwQN9SR
GCDeVVerXP/a9LyBeLcYDt5vp0gScuCAaBYvPcr2pbDqz9GZlrfwl9Iz0iCUpTmQhhEhoIBKeXk9
tXQHsWhm23OwTDq5cV0T5DBT12dO+x1ipX5+zv20ImviyxcENl01iVzhKs6vQ95MHX+pxHblxlBU
YPuFja3EAmW0t5vmvz/OnpfCXy/7rQ6xgCDJJ75MdjYG+7HhMnBInTv5xG7jQu6c/k79Lvbt/xRv
H6QKPvbfMWgJ1i8ogd3JeV3Tix8TEePXtGYTfChpFv7hgV4AWmBYf7IgTlRqrU/HUdIGKv9BI8TB
SzBqVYPrzcU6g6VpgrJB59d/qOk4kR4lAN2/7BJlcai+q/d3mZgxVADZdl7nrcLPO4+BMSDjbD63
fMmfg02IlozR7RqU/XNrneoNZ4K2GUgrdxjrka8niFjdW0gpF8gjO/fPMP3B4w5iG2YpuMobqNxw
5oqcoxdOZrQmG5MEujz/KuJUyPpSObmewGODRZo05kS/rj3jVxH1deDjxGXSsXpHUXYhktPqS9TN
at3f9giJTtNuh+kFkS+cNNw+svwWKLOannwTvP1e8QtTTr7NPMj3sA0cSAhhFkwTj17lVGYf8vWa
+TXiIKgwZCAqEHnofd/x6wE/S8ZSQpwV6q37VYxLa7fD9THwVlIh6GpvOGMUrp9dLEmMEiJFjUmQ
kIPN9lGeOsSx1JMdYp2oJllZb3+wF+LnSIGhQ5lDkFYfH3CzctZlnPLEk6653mFEHYkCAogWlBXG
V7mRofejp8WjHeHdibIEgejWEEF3O9uPSoRafCY9ztvr9dKZedp1I5/zu1DmFaloTC2ifGMwiqLv
IDT0JYWAOlbs2yViH/mkP+9YKjs399+HmTNobK6mOrUr7DjA6mhdxKHh/vaReE6lCA4ud0J2R9iJ
h5MobZwia8/7liFMg0ayfjlSsIaRizcf0Z/aaYi174uxOFZPA7zXwtAeSLRMTxabAeA+bQrc+caK
29RXXArraiZM9IiOlMII1xXwJpK1EsK+w98NP/P+x2Vo2LXniXAZN+4CRi7zSLGRRzASHuxSIm/8
V7GaB2dSOW+X9iFJFDpwnLVJRLkmeK3+A7VlB3tfWCsAsAL5FJgtIPj/OoIXEDRLOTwVjGeIaZuD
xELN+lAD4BQXUR9MpC3SSog+h+Rs+k6DBktyg1+zuYJQhkwYX5KcLB4XwvHMz1XdKmjMxLEiRvZ8
qENJ3RNURsd9KOUc6b+3ee8MFO9dFjIPFOV1E9l7yzjK9yTVN7O3YMzIHkpvJP950BGLbyJDPoho
LT2fO2i/N+G55kWyyRD2MaAhf8hF5mDikNEFu2s/fB5S9Hk/MDHOLGsVdXy5YqQmYWfiYyK2TwqG
0GtCmhodfB0hc9phY5j3BjPRq0RtA3pe1osMYNLDb2GKAvIYC+QqYFQYWWJyRc00zelOEPkpaczR
wafQubsQpN6nV9xOaggfQtyY/DUBNDOf2bZhmLYrdRgVMdiL+bPRO1adzduxYVHwsaKPLvTw12+I
YJYWaA7IvMp+LHFsAkG04IIFzaJyf/NaY1JiBtw5nEkS9nE+QwS1i65OwNFq4Qasu6f+tBVMZXh0
MMFXSu5WfQr77HBfTQeODDmkbe/crVy8BJqjHZ0pkH2Ule6U4YpiTbFWFYcqGojjd+XpGnJpUPwC
eGBLceb+p5Ix/CdFvLXJb7iolBJx4i9LiNs6Y0WqG5NLxOHMCPZpMO+OoyWT0qQIQgEmt2NmRUUK
D9AD/HsrWDr35Iwixsq1ddeVg+1hXnq/p9Xpxf8EM8rg9+0QIXgaBg3YJa82tZBWDt6x95nxDYPM
+Vz3iBE0ouL2vsiTV8n9aYogW03UmkO5tH5YwF6CY1ga0ocVTxYSdza4iXl2zFaVR0ZtmTDzLSDE
5ycQWKKdo6lPcaQd9olCcrHaHLZ4yjnZ/muyRVYWR+R+bn2CKF5fdqa9vGaHX4qnLbuB/1VKWlWJ
IFnVrYKprXCpFj7hVYJPdaYT8Vq6MlOBt7LSlJjtzq+5yLCJXXRsCJKVK92whCPJEZPgOtT7iH/M
lVeScjTCjA3LZY5VyZNs+6x3G8rF77L+0LkqQKxKxDJhSunDQFGDKaP7oxi38uJ8tnnkM7ONXd8B
U264QjdiDbBMexNkD8QoAW8fJifniC8LCone7n1q/WymP6yIMWriOD8IoGyCIEhzfbLxGCueYSQI
WX+fMHy9OYM9HR3vy4daYHRQtZyw0QIwUiCyGUhc83XfZ6igAQ7jH0LOSEsaigTnNRiA8JqsPate
qgjxfpaJhzgr6guPb+eSzkIuvcqV4odmEN1PC4xzY/ylaU+j5cmO8o8V3F/rp6q8NNXOTxJ+ISyK
22axDmNL+itzyX+amBLXssENXzxsbaGUWLsvVoGDk37PPp7W4MrkSz/gV2d/t59YybE0gWgoeaZL
1204nKZyh7rvP3SqbYyQ9jFIQpsUFe2Ogn9ekyruBEB0gaZgQSCNiZsoOU3Pch9/d7XdVvT6peHT
SKU/4gL5RlUwJtcGgd16ZeF+9aK1/eAyloyqpJzMIbQ3b/RpyIVSJi0Su/3iXuZVPCdlMWsXasqx
YsJKLTESEOSMvsCzBDhPPl8NkG84O1bYfhv/ZAa0rohL5EAEpR6KlWlufRgCCl+/e7ads0ksKi7f
ZULpPTWEcaNN8YFb1B3Z/M/XQGQedn093oUgCfV9LpmDi6zl6syv5yZ3yOutyYWVRpWPCOg5e7to
Yyhw+mSDxSHnhHhdd0fZkdoUbwh8XFtsvwhF643YKpH2DLmTYvJ+gxO0FXfWwFkS6mxWqGndZfa3
4H0w12aYaURh9qBzd2XKUONbjoR8S9awLZAN5lvaMuNnjKj+CZemQuEqD86lqQjPkc+QDbPZzcH6
pZvguNbdLDAmu53zRtDjRwvrj5rpG6svLBFMlDhkRB0zOSTunKkIVa8BKoIQwE5ESeZehhRIFxNj
T1D06Mj7k0XnaUQ3v2VYo8S1gE6ydR+XUvkw5Y8AucQVFP1Au44hKcAv0PQ5P2dD9iXTsiX2awM8
iRZgHB93fGoH6ZYR+HSNL0Yp44omlQIILrvRTlP0GE4F7zgs3OQ+W7mNU8ewcsBG/4S9j4cLIaij
mRxD5dDqobhH0w9o+lnkuR3XXZIvcvCuAXrBheUSLIdZ+0/G39Y3qjfJ7wh2hTTYDMSuKze0Ut79
MpizO2Um3rVD5kSg6hG52e6ShILuWYkfVhWWOJlYO20QmCpYAwtdAnn2u1LP79t4FfrcfED2AYFk
wsYi3NIOltbCuhsI3CWPfAPfAyNOwFSVqk/bcyuo05nlsD8f5eMfIY/g+Es2ys6OlrSbQV1fjIVv
kxMB3W94BitcXoY/AfCJ8Kj3C4WYwzJnwT2G7p/OWxPdXgq4ai+4BFm7EZA0pjl1l3brkSEW/Vyq
aLeFaSGz7S6Pug9XNMHlwRTMD1n7AZ/4819vpxAZGtFLyY+CXV692R26tA34HzmpvHGwa/1Em2Rj
tqp4zPxKEgVew2v+Ai0ryKHTkm1MM0WXd1mP5SEWuMHsxTyYZYuCbIcTqertu0qCTMF6J3NTOS6m
q9Ey8PxHiHG2QC90YA8UHloZna13DQjp0jVt4ARQkb4ujDGiFb8AesQdG5UDQogtS+r8kY4nN6pE
dx0QYOl9NqHvBUW261yyWes1hU5/XMpfixurKchxc1F0ndOCNy1Tj+ZM7RSd/sui6y8Y/i0QJ886
cU9xs+z72arn08xjFeJSzBpvqZWqpiyCnCuiL4q4M61ZGFrl/t0Ht0HIi2N7HB6ZUms4qz0eoVS1
zgrBlUnB6pOgZQe7jWwQmjohUFI4O3wCt6Vi2en7XDb1I9R+qaeyxp/W/tnBVNpj+/59PqAxkgva
hR3koxYowffKrc0+gZndlxuTbKYpQur+bs9TcP6/2cQOib4imANBrhwXXtVtlwLth5PLgp/CqYZV
mgQzyfszj5O9iRgqas3bAMMmV0s3g+mqgFB56NM0pglDt5/25H/bYSXfl3hUvErEe3PxNAlFOWy1
DhX1iJ6tjpBpLWw8DfgfSkUXbHskVX6uByJRfKCgX9apUsrSemHNAG5aDNVMTnu9U1k3LcJnj74A
c4JTBgSwbwYOcm0tmC2nm1LiErOqybYQV1AY9Wxo5dRLbKUw7nJXPljwXQ+YRiXL//yK4QxnVhCv
rAwXAmbApiKEviycv2i5EXpChYnpcwDVlkizB9G0pPizXOjYJmZypq4/mcJW2twJ85U0+COWj780
EtFqARFG4t5vjuOz1p2hubtuMDvespJtZtm0hcoWSRLGi8w0NiRE2E2nG0YnqNI1O3kFH2JbbPK+
zvhUQRS6BgBlFeT1gY2qxG4HXFdfPTGXhDTW89fI73GGhmaCrLdc8KZXK0t4VbYddviP/SecP29G
ZowyZ0PeTdohZKn60Kfvec3t9iJ4+OlDWRDfINPtOA/bsvGsiGBZxQXR0FBmc6tyVngD63FLWsP6
MsCEQRlBa7idkUiA3BV2Ri1xVu7utkculhzuvGiXon36sBdVRY2b9mI2OgdzeBJT/9iCpEdTsp2L
GmPgwsH9E8QIzica0iRV5H4ixptNTuyQ1fctJiLWeNBsRYPS3Ta51+ARiim0wCgKnh8xNL280vL8
Dxbs3fOxLE6zXpgMOymkMXYjk/eSX2i+z0kymavmHbH1wM1r2ds7OHM2+7gpX6lwtPwye7870MOB
94XYWRK50+FNVgD1PTMxCqHAeoJWVkuR5EJB5oJfo8FLhBPNGh1eI3zH1Uz0qxWKi+cmoT0tX1v+
iaPhh68Q+xVHlGwgmJiSwwF/p1KUsutF8T1ZSz5EQWngnwwar1oTgo8iR6KhnS99GPt6oUpymQmx
Q1FwxgLAZR89nOIqDeelguPhoiVwn+wg2yUr2iOuV43T7RmxDzhLDbj7x/4ioYlY7EWRD8YmJElf
UAMEq1C4uby//fPJjXs641qFGWPfwVSx2X1UziK1dR4vo1hzXtq+qw1Cvppt12zAbHHLgeMYthgn
oW73L6T3hTvXByhlgMsrTduBikZyckSEZxiUbFdJFjZA670+g+lpP+mQT7v/QZMBSZeLT5a4jODp
jAtipS54pnVcHGKX0aqdtJxnwqcj+As/7Yj7dyCK/QqOaP/S89EJiaA64VKV0s/UJU0/rGfgh/Z7
u/bgIm+IUkw+ilIidyB9o+YD5xVd3mtGtIy8HcR0/I6QrRxyXqtfOQUSHtUtBnhruoWGOpohy2c0
ymtTtauCklnU6lSMuGcQO76l7Uf9rNJJsbC4ivUsnzR+Qn9LgT7e9Rt4Q3Hg3jEROIGvCGE0uLvc
Hqr3S/BUuIvKE5mloJFpmge8FrhSZQ7UDMLWz/lgBV7FILm3NUIfYqjfdy2A/xgECyuZuQN75gms
3yzBCZBhtfPAyc2CDcgR5jknXjDEzDJrPX5AQWrgc/fqZig/vRd9DkEX9LYEXzBSDvAyeMH/3hhJ
mCH14mb1WTeStTanB6mkLU9vIZYWypZ0q3pdi1V9H1VEZVx+SzF/rYZRZaaQU+sYmAUb20V5sE2g
dXnQp4d5m/L26KSHCTftTty042G4ozxwGnMbIcasYJcP3XvBGNfiJeiTAci0ykwV9ECt3mueyEBq
/GtS5CoCO/0s6i9KBRlhI+5wyNvy0qB2aHhECZi1SADgX007DdVKfTHDPYS94aexTXIjCii3eCN5
n10v4/iazDY0lvGoZ8J5I7+I1AK9CcPmmGKIznc99iVHOWmn56XQw/b1M5EJMZrs4Utr52yFoaHw
lRYZRepXeD4+kCtK2bp0/mO8JEPBp566KI+JW5qoDUi0bmHJz3AEZlTgesV9+WL1VGQHftHoysje
rzEpqmA+SUMRFTJADHETXIsLdWRWF07FNpkboSPS9k22n94InNZaqrvbd9uQCgncRnWWGRvUfPXm
twCBvPJvYl7ZI8N2z3T0d5UgqjFiaB1Hm0PcUE6Hka5dsQ1PeIoBIrcuJbLZSKhfbsQ7Wx+Lft5b
Bh6SezBPTWQrvv+l97ailu6jrrFS7EjLTYce+2jN/BuM7+w1YTSeNSgKpvg0YKFUOgl/zklRmigP
ulDy8rBfewcI1z7yqshtg8TOTv3/OjmMVv+zAdoz9sVzxUemjwwT25N7SOVlQukRkYKBK7xB5Swd
9oiIztnedtdrMVDaJdwYgjNKtRX0LamtQDv7UOwXXjc3rDYVEt2MfBXKdzq9y8Lh1qTCjxoC9OKM
0ORYShNE6IfZtthqHSBFK7I/xSh15jHJEWRdZmIH6ZJE/P8ssII5xC0MhXAh+91SxR/inW6chyT3
RnLJ3nkYC847Y+SJWIlqSng9UnGE2Jru6mJnmCJae3/kJIiOMekV+1fVDvqEasus/ogjiyLMxaNG
Mt4+mJvQM47xUv/AAvp4bKsP1fWI5lMz3KVUWNoNcgYvRAnVcSuf+YRC4I0HaydVTAj+J3GtHL9V
mqCPBg8AAiNpet9sgK+LJfT4UnMn70UFEzFyQ1gMHGbzGm08mYntXP3VUFkT4gGEjNlwax11x32R
zur7f3O/+adrGG8tELXPFntUG9/7n/bApJamhllbjDTxZW/xTEKswsG62PeFRAnVObRmLPOkNbga
nLcABAZjDS4GPP167FZvxUCB1NJxvLkVxdiPMy3bkd9UN8Q4kBfHBRDgr2h4ugynPB/6yZFhhwbI
e5Dei/U2Vp1ghD1dpprP6oJ/IjOSqVVqsBirbNGzI5mYne3d7SU1DupKElpU9bflTUDcSdzfiwu8
ISnwygwJrFQIn3HpGnWjLFwK9in4GePiopnBzhaCLf46VkN1eXpj/TkK7oozcx4PGDDuxVY4ccna
lmH3iuHQFpAjJALhbOIQOV8YSqn2HdUS8F1WfN/MFYmHRf/nEKzzmgZhTvawyDotB7TTY/KggIG2
qnulHXZRL4fL7FhuXW6rZERniRTv45j0Z6IVHth7xSXb3vW7qsV3KNxEVmYY2c+o8zc2v4xiFvbi
0v5rWZJOEy70MtbI4qLl44YwusJR3uaBdtgpawvkmxUfmuS4gx4qb49j3qSA7+g0nfiS26JpNhvc
tstOAerrelzcBJ/fvS4jQTXjKmSc/ToWspID9jhzMZPs2u6r2553qP4r4yAN/+BDRNQggNJrEB3h
0ngdcF2s1cF6s1qg9w2SC25sctmy/QkejpH1uKHNfV0MZifmuHrigrh1dZA+zNgCYfnXtLK0OidY
skmaPz3tY7cJkf/i2B2LaywsZn93uMQKH2J9zHaWUcrhHPMAEBsz054E98VskBh3P4ax1sfn/cPV
qM8TZJCpihxYK6OWSMSSxxOMGtAIm31RygKrQpdWTepO+7oDEVwcqbTQS7RMp4L6q0fmTQt2tHS5
Ku3tMIuAwXrjlk2RBjUcMZiaZUGuEFO0g4pXQfKzNM075eWuyj+tHEA7Wr/9hEhEbdjTUfbFzUtm
0NQh+ZlotDduBaYnG5CFjLVDNuszRdzsYi0cHNh/C1z3abqVzUe0VztIFhm3/J8q2Mlu1gzxJTHh
iYGl5vk+23NUHG7XtdU1EN9WynI6LhuifPMX8HZffdIagJEvPYXpRsBIGbR9dxfaeDo0R6XsgC9G
8vS5F00mDDK1ucYcicMCZofGED4hsnB9SGWX3mDc7W93aMrQ4wIcIadvuP8dhS9pKbZ/WSIM2Oo2
kinLyMiEywKYIVi77iu55Xrv1Y95EYok3tM0qeeobQ9Ndb7ax5C16tUgW0nRXZ66AzdbDQvdLf2n
9INtl0Wspmg7sR8vXhK61JZorTZK3XTJQ0yTZM3xl6mzw+BPhQXmPveZ11LJrbTk2MgCcwH2n1CI
yRjWwFGNODqDp6qINtrV7KgoA+RJs9JHoDPEnjkmxBTlRqf/LkHGRqCPWXOk1TaJcFy66zsDOvH4
kIj/dDuXLQlRd3jZqpbECPTv2lMZriX0OAqgISgmhQEno4kbYAYO/KZvmoeasIyoV0W/A517hxPP
zN0qtPT9yxm2wSRioDP23xfbp2n+u5mtcmiki3OdbzF2dARzmgBH4SLGgLW/O12pK/EjIOCnclgq
Jm+bOeuj3orroqqicuiVo1tzqe+PrMYicImVysqJIoMy6aU3bk+d2oXVsdALQ8mFeru8eaqc0S55
JrX0m8K4sLH1/54/sRUxKFD5lcPgmtOjIwyMiLH9vJEl7bjFuxHNX9tN9vuJG6mpZHLT+ATHrq2D
02JjdJUP4EJA9OGOAmLj5O1GGnPPKakuroQ/lbiwt2Hw2iyKmQWBW0OYgHJxdeKzKQ5tU0cA8tP6
BGT2/6qjiWYzMlI7Gik1kQJZDmiLD+GOvtGRgMt/LMkYFV9MUNoJX24vqz7+91WGFwQhzuUO9YUb
HmqFx5hkb8fPR6vHQXQ96/vvZEv5mUZpWW+ekf1bahywK8Em15qKrvCVzHER4TefU/3RvP+rPBPb
gflcDMdezolG7wZ+YBoeWt5FkXHD0qY6qaKu2HdJX7c6fGf3UH2yul2FyfbyiE3zavtOwHXyjL2N
jnAt9fbghXAoDUAlefgVuvH2d9uNkclxqVBxNcxh2cFFfNu0N5vs3ojurj+ZtP6/zTBMo7e7mdE9
84Y0Y1iOlP1s5d2T5jw1yWL52YjoeOX6mAm8bXn5ummxVHlufY2GtWcfqJIwnBln8VqpBkeeOuvg
d3twO+JuLItXhqHIzTiGJPG2e1iM1ui1Pr5OWWOVVu1kMx27DTFjsFd9E0q0jjZUE8oeIJge30OP
wXQlRazEjfrklbI4n2j0Ik/LHhArX9GujRJ4iFek9Ip6xan9NMhqGhLx79NZvIkoK2uLaafX5nh4
vzKeKpWG6BRsLGRCYi0ru6pSxr/g36iCLaEMgYiNtDXCmBOPAARparpbKwPDk7jar3+9v+S9EuoT
aZnosrI4AxulSpavHpvUgxd3JGTayKXpfNBXD4HBamoDgv77udzUoHTSUe7OFce/+Gb0jFKtGJh7
xOgYmTYrLOHs4rD17gprboZrBS9wrDK2MYM17iinpTWIBINykfNIDkIS5WX9tZRstLtA/Ibd4fjq
/leew7GKVRSI9OkL/kyPPUXGvDlwX31WXk3Gc1IIF4DaFuNLu8NqM0OcX+xT9w9Huxj7z7NfRYbY
mPhsnbTy6eollMpM/zJTYbrLQwVZ9/y+xrAV938e2Hf9SJQEnhPh3D5qg13wQELbMLg9xBufRfMm
cbSWpaHh3F7nG/9q7oeEBmdv/1IubBaFfpOU4+GAuPLUiPNc0WvbG0vbZXIUHmmJqX+iwvUkFH7V
aS1t5Zzc97+beRrazM8eXMdQpO/36r0z+m3QyjvRdahTvRFTa0NczLaw5mjiUEvDNyOV4NXZqi4e
YaN+NL6cO47gA/59wkB8t+hNzRxTFq2on7PtqvnQegD0Q9C66phe+d9VXQodlclIBJ7lX2KUOFkR
FNHw+KcWtpsIFjlCU5PBrGGWiDx2hS0cMLE4pnoR0cZlfVL3Wg3TU2tHHjnWnvhNUlU7QvINpipC
rx9CiwNYIG+KOg/UnmXnsfMXr1Hr8xLZU4BK9sNclCLn2DJVTgzSBN/GiDlB7J0UELBwtYUhtYOp
QSI0PyMgp2LoGDkUdDYQVkCBWKlBln+amJhrGWcOxC9TwGrDtcRR631qlRMnz5/iIEzHSLrlFO6J
JYljGDPG0txCqFjuX4PnFJH+3qnf+YzmKVuL0PfGaj1F01wKg/IcaTCHY71FT4KVSaXXWLuFfhMd
NIDAOxQrr/DQ2+66IVrCqLbh7bmpBMWCXK3AgEM6w4WSdw54BRzOWTULkveKwbUXts0vsY1ELpWP
EZ4r+YYfzrp12RMYo7IfwU4gIZj/QU0Vu6kO9uQGIaEmevMsfFbXYGVLRlBxyCOSLAcKtTuLou/e
8fq8uCEUkt1f+qebKPXstJHegVk0/1QLfSbWO1F49xhBhEoXrMIA8N7tm2IAXucxb+Su6Md1+cIm
IG5ng5IwDKovCi+KDJnpUS3Ntv0zQ/qYzmr5y8kgtr2Fp/gYhKCE0aG5RWou286uo3DawrS0Rlyp
0GZkgjBqQ0uXU6SKZUcDCCqY+NeN2DhC6td1xzKvl2t2ea337LkjSwY4JXumaww68uwe6JplGq47
wwFLvEhxNc0rpfKn/u/nV8TZx47YrSKZqT0rFrNNBHuvkRlZ5wb3+3AeErQEuuRUFY0qDPEfnrPH
46MCoKAe1bNUuwjFs/o8EJLr2VI1Q56WM4+tL+6RHcDb5+P6IryAJi7Xh2qQEpEMzmEPtGJddNET
PxO1A0K3wVZptpq8Lj9KhFM1RROCyozslsfffpew77ThrezXSGCu3qOikiTU/I77QfpmS4x2R2jB
YJCBKj9/lsz4riQU9ICsfmd3fz4QJ8r6AaEfIz2iqBdvcB6DuGMvelCrmZP3cMJg/TAEO60SO2xB
DoHprRrJPp+3ptgzi4HCTGdSYl6FMDTqu0NCXurFN9XDn5R66Fn9XkXcvfCd6+fRDh7o6QYl3BvU
mD404Q1TZuen8yf9wUeUR+CX+0S5sU+ZOk9rB/YDj2s/1020j0TP6k8RypQMfCeZsDZH818k9GtM
yuxktTXRbahK8a7qK1J6wZ9bmjXJHevvsBR5kBUO9uwrgXRhX2weHdOsFfnmBiwImVipJXHwuqL5
ssKhjmgie22hFsLUbR5nIg7eJdL+M8ODcK23JPQAd/V9MRwoPXGLaMizxPQhPj5Eon5i5qu1N8O4
qxq+k69n2p8PtBihHNYcnTLL9w6ee7ZEKLj/94QbYClfbfJGdAQ5mknngPZ9mtC14lexEak3rpT/
PF2ycc2Gvh0b72MdSkK4JZml7FF8qoeNLoQz58D2zDG0rlRtKR4MdrwQ0A65/H9m3ZIqnap5GOrr
mEMtMgMaM+n7dwuaEVbbIgbjjm5xuQe49lB706NE7cksuo7lhCpbt4aUCTdqfIozLNej0JaGL+4j
xxxCk2+QbnmJy3g5ZsTAsVfIiQMXwpv8JV3Ia/0w2cWRYwEPKqFG+JVolxlIRdZqYb79IO9E+XpL
kCmQ4zTd6O8OcpYz5nhmFS7VtqEFLWUWweT9Tcke2PDv+jZJCapAsS+LynvBeul81g1E2vSbYywu
C6KIJFBzk5RGmLMoe98pDn9MHeUJmD9/A1x8wPgGLbDc0j1TQoeXPrjsMXUFCemnW/ChseOERYp8
b3byRBVlgEDnyXgwmhiLhK2owxMqtOZp20XmaWnoMdfCOA3qxnTNQcxgUHL1rHR4U69B0D2ZnNLC
j16KiJ4CDpb6D31h8B1mCnCrrr9HFBaRsN7aPYAgDfh40DhJCZ+i07pTQxzfEejyIL/9+EpLzdhX
jaVUoe4UCMc2yjJiwO3N38HAUlwPQ7YGYbG1UAaO+fPDmAyUPd6Uf5CeiVB3klFzX6TZy7HzEkLy
HMONAXD6u64/7AbQHt7B6MV/ZA6aej+XN/x+0j+/3lITyW42lFyW5zvrz7GNtwDRDySFlVYhbts2
0RIUC/pu4Cn6VLCg9XpKt5YAl+YevlUSlGJyYdBkgk4eRNf3gLcPqhzhQ0CiFv1ucZ6WooGx23IE
OjHYIzDukt0SZTrXLn1RajtbkcGkdJRVBsJi4zMvU4unMI3mWNJ0xLlgHrSXcv9pLmnAKdiJ3iPh
ZDdZ1uan8XAnLqdzk+vgC4L6LcsLIJ6UC7u9nhIXEYNMBGSWS6VVTsKvP71b9q4P0SEgWQZl5NoZ
JkhqTyo1iGEbBfuwlHAd4t/ocTpkFXvQ0HQIcnhpX2kKWQ0wcsFgaA03Vc24DhEZQaqwgGs9e5jq
K1Yk96pnOkvNS3fUtYw57TcLRF+TqmjGCEnK4QuDr7XVl1t3teg6LzEsigMey6izrFvXC6ma5dAX
44mS+MvQwQzLIJOciUNgcWyEz2bAwBjY4SqpeLCUWJDNCWEPzxhRa3dHN0IaV4zW3KGHkxH7eAJO
ZkjQtMUY5SRMFpIQNexjCEu+7C/y2FA/yWUBRmgESRO2+DRToIftrHg7a5zZqgHDbUqqwWcGl4GF
3XkZK42g1iNSIW7ZNGw2ytBkcnzqyjhpWwZQPKfGRNTYUw0xR/hjvNPk2i9SbjCpFCQufjcN7lvx
2MYUCqZdjlP3r+khjTytMVQcLUoj7c85RTP50c597Z4zxXCgSqB0E7+Vejqh1cjfvmfH7IXSkup4
y5YN8NO0uYGazo3IR1imaoQFn8zEgcBRQUs63Rsey/9+pl6/4euOkw8XQskTM8yrCnRKztPXPNIL
BcQSs/WSHSuWJJpoU+vy/B0pKvb8S1dXUQvQEm6fJ8gTNknAirhRKvX9xHrjyUp1ykf9ToiASCHk
+sm+qzxuIxKys2eHWQtHsD+dyZu0rooTVu/JyYXAgBKU0GOJZPo66B6SXWFgGuFWIFi1smveZYeX
SyVXc3bWB9LF9NpNBnzviVfbN4NZiuNw8O7fRiixyfFcGHYSnyEgPNyTCUsaH3GQfecBWrnG46Uy
qstxZzeNrITeHhz70Wi/lMxuK25cnNRi/5BWLNppl1LFCFrfc1Kz1Idh11G361Xcc7eUhnEWv0PW
PeltdYS332WYa97fFkzUW09epSCSk9vgJJxjPGgwSVdT8n7/UdMjIicFJVTG+TIwZBvjzKvZu3SR
L186nBQmvSCp1Zm/2AjvqKk2/YMvxG7W+PToipahr2XJ1+hFIFfv3iUHdhbIB0mSI5mDGN2WHa+S
B6roCGqb7DYgPAKrIBYi4F+uk9uezXd8M6YsUAhiq2wgDzTZg8p1uix9hfOpiiWpRSPG0iGnvMxd
d8A8hdMrPIpYI4QVKcRNB9UJvbAzfsOqKRaXU5blYWgsggUYFTGoAT7iSQWCQ5jmDeOLiv/tHKvc
BWiYvNwIAwTnhH0MVKENBRquekMHWySaXkJtNNSISvVHeGIUJHjtBRPc6C7TY+WsjEZFCJRQPrrr
s1/f247zXDiNgzKd0ClxgdYPttL0fxEoOsZyz3VGL8kAnFJUFN109fU3fDdS8+LQi/fpEZn2tc/o
NAv7cvtZFWDKAr533y428tc4+C5k5dL4Z/Kx5KXla+PcatgHMxD0HMCv7Vm61rCRr5eNjGCbfKve
mNCuXsa0s2zgvHCsvosAzwSisiZMf3QVREhUkT4UW+YDLVKsNBxzuQKhlj/bSNtwX3ukZO13HXeu
7KpArIuWlDqwK/tjeLHMSPFt0VKBO/4EVhkdfyQAtFTJzQve0RP3EUOJ51srcUs2VkdrJeU9NHzk
YdGphLv0k+4qL7PhWLEgtZxeG1grxJxxzP6hvBSRaYq99a2tpsx/AC2vicY4m0C1IuJMWJWcNbqu
hlVNQxE0ukcxk1qQUXyr/qKoXnj9MnCTSjjZLJt2gyFskurEDlosL+1sIg8xfr4IiJIkLgmlamsh
F+3/8b2kbN8f9wft/e4TJO5xhP0/E/YNx2COOI2Bef7bxinM5fhsIqL5o1ateYPsQAKYP/Yxf39z
9trAH9AoE7H7d/qqmgOQTn5XMIPAPq4xYfGdfPom0ROS2gM6tv0MjFo+J+wlBi/ypzanW1Wx6Blu
JpPVI553A7rPi69pko4Gni+pst8sQY3lhgVYhlyZkWUt2r2QPkrHPXgPEsvIvF6wZtcOkc/7ocCg
07say5ZUtvdd0jAyQ+o2DAaLjUZDb1+/aeMvccSCX6o90cVX8rMldgD5qeS5BtPX+VLN4AjvMp1E
EN7vfftQ1EvCQJfJ5+G8/qOtWlpYNIHispVnzPL0Rkzp/anbHpYIQWizeKG3IY+8GrTAk32MiU9a
55qYV+QCezXA3e/fny15WTdCAuGGm4PX9nMajiUeCv8QSWxlkjnwQB4xGBl/kIdyv8+Uids0VCfE
c2qU4BxkCjJBigU08qeAuXNsG1Tae8IsyH5QZ+QTUGBYwFLa5AfEe9Hlj8ayrQwiCy4HQSrYjVAT
efIJ3q7spIGsORsdR9acpoRxo2sSiga+foEEUOjtL9shSAzKAI6id3PKhaxkFeckWx9irpXa5wt2
ll4P2fGhSX1hfMIgCEI79Ibv4CBbCLW0tQ8myLvJZ27Fm/W95uOpLxnyJnMdZhi/MNIXFXbwlxa2
/jZofZ4ZGrr4vjXHwrrkYBgM+ypi6u2XI85xi7iFExo/I4xjIFjneKnbCJEU1bZE3CKWiaQwTsfn
owCNOESvsZNz7OQ4P/b1P5A317DUbMcjbDSB7MCWA7GBDhLDxfw2TwsJ24qHazsUM+aOsmVDvTiQ
nPwk/Ruj+TsK0fVD3hOKJOWPagI99StF5tPwBHkIrVTOTPE3s+JUL8RJ55xPmB7aPcfvSuRDS23Y
i3yI6/NGfVFzWsjNtSOi9kqOqvS8gcwtK4iG5bYWXiRoRoT8fROrZgbbvXs7O7yVm4sovDU8odDg
E5J/REDP8LFelsbHCZyP3NMoL0JO52XPIpZEHJl0Hg803mcfIGvZLJj3SBMYtvPWN9w1VeUoWzSy
cMgBU2y5xl5JQbkqziN2Rx21w87yb5gjbjbDoHeu+VfOvMRce4tiZ3saKhM76yn5c/D738Oqi2Bq
26o+2FSdzVw6+iaDSlncGeNtEApIs0A2GvHE0sgFPe0Gs/RyrXSL/VlKtyiirySqCTAvoqc2SHKX
Fa6HFxueHdhbJ5Nuw7yip0i9JwPWI2yygkLxyBREuu3eTJNAoZEv6nbX6sjyVXu1t2Z76I7yJMzt
6MHC+iyy169huUngdIJ/mk0Z1ggHbsxpdlOXyk2fnjlfPApFQ+MOHeOEzkb6c19UaCm9IesuSpV+
xDGJXf4Ww55a9Auk1kFE58IwSyde3WBzzTFfnOgC2dciAHqSCrarqRlWYPi8F7DPKeMXjbnX4oLG
tEyPdrz687QVmwFR3tJ3nV5RE15q9hEvDiFak65YLs+M/Tko1CKt3G+a1OMjtMkK6R0D01/5i2HE
cM2Hdas8WHWAH0QB078tSd8fRChhOdGwfp7U3VSUbwI6549Mj1pviSHaHmiXJ0+IeTH/iuMivxw/
xYoPyHiq363cXwU21mJK4esm5viSaXwgxvPo/ThNzTE8BzJo9YjzdDAfgKu/0wmeoHtEuSdzWnut
+D8zZNbRKhdwfwoHJeDmvMhvHbCq4Y6wztyP/lrvr2sSJsf9NMpTwAIMHNQfZbbBgAB7BoqApU3j
9mNZAnUScErzJCvVYunZp/vpVE/yRcMetM4PPnBExuKqnS7KyG5/GhHrIds2fTPZ/JrptoIQ8wuG
yXN/cLDEBkaCqdBJs9RudOZQhOLlDUT9whtjIV1EgS/X/adHByVx7CKPv5rFTr0+a0/wZUpMbbgb
DOMCvpxeUsVJnHA3cScDkLD4Eiq3F0uK/J2E0KH7uokqpSWenxYNNxcdqDs1OZv0rKC4VE3b2Stc
3LZ3JBTJAaC/NAhiXJkdi1C0oPBLzHpJ7ayYobZ2gZXVYc/6MIY/LFsHAc6GwOnIzmayypByVJOW
HVqrf4gOR/0NYOvAtk6uZ+4cmD7aEcpV3SjaWjbAxbQzTNp51hbJ8UiY84XodA8sSDX/WqzXVt1K
aBOPARDIjND2ERnPE2fXvRUoylrvWpeAm+m6Je5x5Xlx52EGx/hOgN88zzHrDmT1bbkH3+YwlELG
C9m5SWEc6S1tXqv0pf/l3s2LS8GhnpCrQyBsNLPzVREqvps9qSFKu3Q16QzcWHGm++Vg9XxClbqs
oP+wg5dPtMwzs/z6InNhfr/HoZ87mQvAehtUXPDoXw/4jU0pOIDyWGhJkqFRk2m2Ykl1Rm16Xdsh
ddsidnw0P+s8Q1Xob+Cb12Z3eqvMHKPvj5VcuE9GSyNE4PPBWLR17jIryBQVJGf5r1jmT7fD0/b/
BAJmHkBAkbTunkXf6jGSFc1nh1YB+t6O26OFdA4j0Wu5ik5pWfyNlCWIPFMc28rEx3yXuch9Zpl0
5kSbqZimwxU9821AKN6O9KY/glrBnuyKf2xufDT38ThNBCSWJb3v4eD7VNmQdamn5dfQ2FUoST6I
wyuxKKUXgOAkK5t4zUmX4YPSIFAH9kxJmnfCW9L+EXejdNKpyGqV606mXGivwnT7FHIZ2q9uqpHQ
M5p8xvuThpZnCiyAgvmsZ5RDRqf+TfCDqAN6msLtZ9qTBpWuREXtx+vBJ4UdPR2oIcCEZ2xW3lhZ
TocrqamHoiY1jN/DjngFeZ0FipXum4cUWhjnvR34jmkXkHOgClfPO8kdMDPWu4DXNZKe2fnGgPsu
wCgCsJz6eymTP4QJECbwjWxYMQ5/j4rJsmECPAWgVnZb2Ey0EDjkV6pdjTxtu9lBGSksOkqcxBRi
XJshhmgCAsmFurlQ1Vk2cuXhoue0BI46t3qbFmQQ/9/X/eApsXPAUYENQhx+QjcOOeoDmHNEwRzs
8Vhj4ekSF+hcmQ/q0FJcqLI9/zAVoQh4ewSgso4M0B1Toq/+hOYCm62UtK3fNGeXkUeZPacpKBtu
K2syf8HkYDB4+u1TWvEgv/IiXeq920MaYOImIvZ7jfeVGU9M6fhaxdO+eBTnTyenBWrkGP38Ks35
BT7VdOcH6UkrvjfaY/DTiONrsA5EsTFDgVInJBYqbBf/nnrnMpP617oYNSomGn8PM09Ly4BfIcsZ
GExY9mGpMCk+ETGTSF92SY+qYxrRCiu1Ys7xjS7tpcg1PY14CTd+Ei8IfkcB0ZvNtXzs19KGiAsL
ezNOYRZzhqR8zmuIGgogOT91qrWMzXXqyx/1VMuQXmzGT9WxHkPP/Z1il+/CyMHK9VatVAt0yxTe
npQs/W2zEbwq28PsZJ4M5bCGwhcIIXX4ABifmhn8Y9NYvgrT2IlsGjC+U54n0XSd93sQX3cqKGkA
PcSLBRMZ8AN8qGOL0poHNu+JkJXnEjvKaLO9b3yjEBMCKshwcFki1g/BzE8vOnbbyj0Xz0BWuKUT
N/h53bxz+VJ7j2cQFvv61OqHvEnV/rReRrqFcdJRrQNrI4ASo1B5i8ukVdxdzYHNsw/hCvJrcIPE
reF+pZMszQ99/LrUbgSwH7GpOAFNq+19Sw2oqeF7X9ACwfJQet7Y67Tk7lxmSDyf35avUVgBo+Wf
c9MWl+ohYSP2cKQzP9iThNArRKb7ih4kh1TtHAwSXrMj5EcUw2SLzyT+isFIw2aV1/MHTR1xHUx3
gRFHQVedwbKpGCeX0YySNZHV0wZ1DhqMuafY1hg02NTsVgdIJWLuFtRULMGwYl1+5mu/DHcKwcRC
jVEJuh96ic1kmfbU7VImK2S3n6wluSAaWi+G/jMJ+aMg97j+55y+voOPr3yO2//lqmarezJwkgDT
2Y15YpRc26RjD3YRfORfQgDeFZatbYJOxf8JPShxZg6GoKKtfq+XoPaB+AfNtgWqdQ/QyTDhirde
ry5KIqtRb0MvUZvoolrO4i1bqvTHYXaaS898+0EI8xu0MlCauCQ0Lohq/HfALEkNLk5Ew6/LjVt+
2upjByQYUMH4Cd8pqi9tY6CP3AczMsFOcLOIkjNUQHu7/fvFOl41lDBhNSDxBcIIQAbB5c12uhBX
h6A2KJ7Mlbn1OrzTm5k0NfaSNlviQCCncPhV2ulvc52u8rlMH7gIlAAT4ra/wD93ZUWFIYe9iqPM
Njizzg4godasnOXtWufkScpcB2OdcgwjIO92COvi4hzDhmcTJ1t9/hGiAwi82rlHcrHH6GupUUWS
NIgicQA/HBwLxo4pk35MZW27SJco679fw3Ty9RHywgPVnFAp6o6pbU+fG+tk5zvXZeLmh/7HWf30
T5SDroBsgSYFe61SslYioZ5fNT4o0agSW8imDAq7MaNZuKvbr67wngRT444snzbiHl7q37ievA9K
d8ZnW/7TSSNmTF+89tTaN3m2/ZA0iFH2FNLtuZCG5pA1NspuN3hONwj3h4PKrWhPV7RfeF9V7tuf
oPDZyzc15Q1UZR+fidI7hPj53DwMyHgfJLsM9MZrdxe8SGIYP+Yg6niJwwaQBdItg140/LrMK5tf
sq2rFB+bZYihNO8Gl5qJUi2ClBNaHVDJ/tF3galwKsO/dhVDUzXf8xKrP4KJah/CpiOCSP/Gnpd1
kFSTfuCVOqrKuEvDf34qA7RWPx35k1cGrv2BXrwCojdoBEkrpBS1H+O4CYDUCiflduVEGS2caGXX
fQpLNW85y9AWqZiovEYHoTubsCDJqom+GZ9lYwrqX3vMSXkVz+PstpyfsakYqr+LS808A3S4vYvM
8++Sn091itIW7ZKDdw4otOF1h5Mw3qsUNcL92v0yplnuB90NOrZDS8o45F4AwiEKWjX4gio/h9Tr
KVbnKFKAYsuPWs9c6ZRsU7rmf8G0HgzfcfdhBAmDPyqs6YwIQNYd7g5ICpH9W5/uWH3auBTBCUK+
RrU5F9PWXh81cGn4JOsMWILXt8ebYfUdqTIfABkhJNTjy0VOr5pXn1Hz+PNWTxstDcOt9WGrl/z/
JDrHMVlCAXArX+bYgrqTNfg/jfVAe1ESdd+/VfSlAG4imn1esezvW4Zh4/ZYJjsVvOd1nN/l3Az+
mzAh8+FR7iMR5/kt10B4rcuNegkbtQ/2dMbVO1t5SWgh/qZ48JnZlJhpAjgM+5Mx4oftQvVGk4Fl
kpISQrK3JuMYb2Z7TteC2qQAOi3tG5VMTrPfCOjmLWVQtFhPUevzEm3884ox6ejqCczjW4oL8Jl9
lTLgcUUUq3s6rrGQis/v5nfK1dlVySLsGtKXGYUBkN6uBBfdLsaNSIQzr/eLigH0a2oevAAHmQTw
hVgh8RAwj/x1BeVcPKcSSakTcXfF5C/+idXxGwY9pcC1K4B3DT1qFIv/R36SWQmTPkhbVHpZgJ5k
GqVXBONSFbRvEFwMxiBuX+VLU4vdUZtNwEVvb5muFzC6BpbmCDfU8w+eE5pq3sO6GEaUZ87BbEjR
SqRpFWS/M80WC3lsdnsuTlyt0/3Vca9HZ2bTNHYI+HPya8Ht6YdxobVlEG/ETtOjmS9/Ft/x9aPD
jISGcoYS6llQjH7RRTuaW0/toDdKyzCxvDtcbQT7TRi5O/NoJOR/x3mvIbxXQNXUpZzGEUBlAkfv
V/DF5M7k1TE/ht5ihm8U+eGwS+CfMdgS/8OXyuYcm530F7DevvR8SD1UyI1oidIcCcp5W7eX4bE/
r/VRO9wOxxuse0hHtetF1in889iN5JMUItfx4SNb53Sh/IrNDJ7p/u3hyLnc1Ekc/CCSAeNMosXa
etHywuhqN6TrmNHd1lMtCMfLFvUAqZKryEfiROxEQ1xxxC8ySVbnvBEE16jUZ+XwZ+4oHA0gfF6O
gr5LrEgA13aCfwKitf2hHQpI89JA5827tRjuDnLTka8VilTx7/GheBZr6IzkvgwiWYDUOFyTMwQw
6Z6A3wZLslZFA7EVIAw31h2J/1O197iGQuz9JZqzutJem0S6f3c3xwmmnGFuXGOKc5cBbtQNQ3Ej
oG0WeyZcokrXWCNxuMTEQXUzPLRSOB9mGiQ+9vt2X0js0+gP6zxdlOWPGEcyGlqMWSHimDcU8xa0
rrwY1uQ00vSEWpdfentD/dsAnHCLoDilAd6lETAdDm9YdkheSrr9htz1VVpOyB+Mlbmi0ZHInZYt
QyRKrtN2PJESCPsFVhpY18VPYMPny9fyjkrmhBLUioKgT35b0wxIy1MnpQRuKZZ3oX1bfT/NBI9I
Qn+yWY0rN5ogJQ/I2MSskzs5oQd8hTRi1cdHDUUN9pIW7T2BDa6lIsNPfXIVNFcS/qH7XwctLg7O
bXXjtLQ1o9vvsNoqWN19DJ0TiZEvZndy8PA8gpYeL6Y5rV83yRi5YSr7eWXDzTz5XT5sbCfFbfvW
BGsvLmwjGN1YkRk3ih081L6pwWSwDo8u7nofKKqN7Ung4C8ilz3BZF45VfA9PLwLDfd5oKJGR/ng
KcZOjjsi5lwXkArcy28hM93m4fMUnY31kJ03DCRX8p3y+pl9pcFW5NfBMEtrLb/dmAI4P6DAPgq0
vL5wroMT8hLnS+VZwSiXPoDPFgdXVbOVIIaeQjCfcHXybLTeybzZyYg1sE/+D2ZXhi7Cy13vmH/C
R7lkUd1d/YiOG5PYFEbEYjHhGsn8bSyOpOM5aMPzyrxwtrOVM47sQSGvhot9Ild7NwmZV4hzhs1/
ZudLZdGz3QWijhXX25GM8NO/DKW/9pEfsiR+ERQkXbPlIgKRC1At2ybXSHCgal/bhBdEBAmRnsXn
z+8hov8WXms44jWW686mW5H//cc4TaHYuEAgYFU9JmvBFCjBl5HHq3PkFEjxC3zvjeDgY66RYyFU
fnWxuszNQalYFrlhe1Itp9GfA2Cd9+sxs380ExzN72yh+lT2xgZ4UaG8o5FOU9HuHKaNi2FPv/Kf
yQXkHIbuB1BghmhiTGH6/a8kKm1iMLbtmjrLH6+8lpGPB4O9ifzqOPu4XY1dNMc8c2niS8l9sARv
nsc3+rGZY07M4HGc+ya/a5e503qdeXY9B1x+0qlmrJL+zt/1Kp9qAshMVQ+B8m2Qewpqat+lapxl
NhIkYWa37sf5mBBn40NnzAj8qNDXSlwUi4wiQkk3a5Din0bW/SXdMQa5C14VQEGbnufQ3s4DPVA8
ihVZfIWORYdr7BLctDeSU4FZEPXP7t7ABq2hjCm2EBN4N6SxLIViqsA1yDJBRXy6TLiHuQuvJhJ5
jkmTwh1evkjDfpyDLbIeHXes5u2M9OVeDTSNuWzIj0oqhUUoEv5Et9aCeIHa4AlFQNfhu07HW+jA
BTeMFI77FhGZ5E6Y5bcCaRpmg3O0x8f5SESxw+g+71f/hlpxiBvHweme7W6SpX5L6QDOvCWhlzwN
pKWXvHfXGkPDwxw4dkDlAkH9PhoyAv4XeUFRBohg1svcqOrtDHBHJ1EZfIY5VIj1ldrJcYp3jv8K
kn85BtpC8BJgBC9lVtzsHdeUcD0VoKB2QNYPBOrpbvNa+mp/1mXW2rjlMbeLKbLhEm0Y68GhDIrK
YJJTkYb16YqhRfDcuQ05fQ+1rCj56Ogde/XesfL64WHcFgtPEDCtY1OAC7PZ36hEevzYa9wZGRgl
pk8VVOOAlgtSP7QKfQ/h831S5YRbCdkpR6l/ujnUffDHlkgBvbV1B0rR/HPmkLiXdcfG15Ectslc
m0R0ivk1EzkAl1SxEM3R1/s6QaHnN2cZwtZ4o1NaPp4OH0E/geL/M5oRSltZJVt78exU4PfbsQxg
G74vamgOFFIy41nHZO3ZO2bA8F4YrQfpynderto2BsRJXfxE2V2wqhPWTIDpozE3LIsdGiNxhL9p
QeymfhcXtkGvPR8vheSsyKkJuS4LgkX7Io8KwWXLS+yzhXkY3JgGicplAgRHlhYsdrpMxTwwkiVY
hQ+g1KEF8+j51NlmVtbK0rro9xi10A+AdkJ6LsukGAp7JdXPDs+HDj0z3TeMv3RDzLdalGDDaYcA
tWYguY2e5xMgoOO87x/YzReljXJxFF/D6efVzrHMne0x100namaIUl/5LdMNG3R82JuA2tQ4I7Pk
kDV+jbDSvxwbRNtN2IfQE2TVgYQh46w/Oy20GzR6W2i87R+GYzSH7gEIi+VAPBitQuuVSAPg3l48
Aay0GDHHjfgw7DhDvcsCJQ87YORjbnUuoTTp+56HocJqdUOq0pT+BAxiCr8BbaEUjfrKS0hNP9Fu
pluYvczRDy2KtgNxAmCcVn3qHbjOKP8xHJTTVkZDml5R0Nax8/v+Wv09dcb0yooRXSLB+GxWKjFv
9Sq83hqXpFJ4gWpulo6AD5NMcPyqx6OZtCOEVSjmdd0USLRISUg3XRXy1EWLw6h9ITnm+SgWh0Hm
u4w+5zYBX3P8KQRVkeQq/1qSuI5B7UUM5iJSxobVn9HWdBbdhaFP3zRKOzprq5h2CWN2dKt444TD
KJqvoscZw8yb8fG/jp9A73N1oh1SKonq6QdaOcskVDFTL1f8tNuLW2VgIYPtM8A6fFmXgeH+HCO4
cnxTXnSElOI8TDeVzurbi95goRjNvy/Ei3b9FdTI0P7oZ3WIBQrBlF+yQI+9LQPoNU3G4e3LtohH
KbG1gaGMo7XsU2bTfGkDzoeMjGxXJlqHabKD7bycb9rbOgkQvt9Q7bobX9asFkE1LHz6iwGqS3pR
ZHnpV49gca6ZMduWzH9WYQ+7MAcXABFKeHEsks/LpNDffWxxScDLlF7XEozNshMBW3hoZQG3+OfD
dPC751mhASN4mPOxD+fWPm5FSWQmkM1YPVEviRH/ZNrMACaH3FchshupL4MbQCD2OmFbMQER/HVr
13pdqlAipaFmusjb5h74YSc8m5Q98/gKQSxmcz1aLX+mFsVRN/1Uu2HSRDuOoCOHYi3Xqj0dDyUQ
NvCbjLTZSn0sJNaI2kKi2HnyfL937dvVD06cHDX1y6MFrdQC5Ol84Gq4dMwsAjwl5/2pvL9iU28S
aAO1fD16OMTMiCF7wXWkyEhXADY7aT0S7Bgb/qsHiUW1PjErpbid02hY+og6+icYnDs9aRDMc0jP
hkpcc4HlGsn4w8Ld1NUQEwBeLa3nMXzFrzJLWjyIHnrgcvFxNVgLaDoITsej8SvvF4En7UclAmvd
aNpFAKFMb6lpT+/TzQzE++SEBeTCt6tkH5DBKGx7/pDzw6dSf6YPyDsVBUUcwVGjv9HxIpyZMgxR
yhhzhgN7yWU9TMyX/vyDkI5SR6mBRy5Vv+FVKodMR0wu2lt3m2bv8A2JrOyHjjffpEHVMbb+D3Ou
Gdx+eOCE7ihcW/aR60srrGUr5Kg+WA7ysYwW5FsvueMbMXe7xRmsVfZ0BQ98OorGg9kIgo2hyqqr
y0N2ABdNYmdQkxUgVn3jMt/ZP03yTHXvAbjyZagy64JThIv7YC26b/Icxkdw7ScO30pQ5PnAaCry
NJCPzhth3tZBjbXI9hsLJW/qG3aJIm5181CobW1+006dXwzWSwzyGX5MQCWPLH4hTURADKjSM8h4
wNmp7ww5eeKmSwCYwabgiWF6+rRA56GiY3KmGJkxESvnXsHxdV+n4CONtUZ7Idk7Q7rJ5vt7N6m8
b8X7Bn55+iTXv1fag2+aqH3isIZa/csnwdrx/fbA5+JxjUlrY0zzfD48Kuh3m+h2TZLNh+E9b6B7
06czIyttSDvfAIQesqR4HictbPoHJYu2AcElK6nkZIrC11/Fvv8TaRAvNMqZeJSPfrF+SKWdhQRs
5UJPsyE/CURd30kJs093Nh3gUVoSJ/F/rzl4ZM9FPuqLvWVmJ1hCG6uKS0mHkP6q4t+UWCJM/xOf
PMowVj/QemoJ4LFigfKNp8C9HYGcQEjzZ5hJKxfyB5/sxT2JTAmr/k3mfCBWff1yHx3Mo1oz7h7O
aKRPFXlP87RId201JF4V+KEv+rbJw6VYs8yR7xLoXmapthbb5S4B9jLJD1RivP9AFg8rc2t1V8/4
TrG7mJZ6dVhwn+AQBZwfzz+ImudUlITMMhoYe+qpmDUZayy+ZNig6V8Li9oRZQg8Hw1ppVjZ2U1M
VKBYhNrdG77oYnGpYD3m1dj4fPbuflrAT0TzLpbenZpq3WbOGWFMXcs7NAWFcFuxf/LbyW/P0syD
jpLV7JfH07HuxXPhITgIda9g3oGl6rQXRrKf2i+9jCYVQXYNZ8LShAevKJnoa5eNP7s987MZOddQ
ADoYInHmuU8XHcIY/76CqBFLhxguQZjBRz4wFSp8uTn3i/NL/v4BRorg77F1L2SAX3ESNyqQe0wj
vxj3hBbdAZoHW6yHEqF9Xi4hkn1ExiiID7lYC7s/WGFG/0hXlvzyJAsMNPangoUd9BQExkHerSHi
GagJhbWSRTlhXqscB3BHJKNgCOGeuLT2E/xbJuicu2jmzX14YS+MlBv/evSh8ptou7wZs7jcO4Qa
2nvW7tkMXdBAe56Gp9vLv1zrDb7F7LdSkYqVbLBlM5gkBJsjzr0oqiQ0YkLeq9fosqz9BSQ0wCtN
Gnfla2Y7V8/l5oKmhFfOWnyy5muqUnIpGt8fBXzahI97ESNH29LHC4s5BTl3PqprofTrYZ9QZpAR
U0ZTFKKgXRvlZtQvo9h8eUN7TrxeYTsvv687FGbJoC05kH4gQHinEEeSl4hlMXtfmjRNpc8w0dAm
CqEnAz82Kr3uofIRJYfaW2Oep1Ev0zpvRiuz/z24+IUxfrqNzkIopgYkTPqDKgxtr6CKZz7M0zDQ
gQeMUyNnuT5FfDAWtQZ2190i4C1R2oEM6oeolWG8EKoeWq6WKSs/Za2sdn0qpM4w+NfVD+zMgdrL
52YycQkv5r90bwSrR4UTfCMYbQHuB3Eqh5ihcMCDzhSA8zXt8B1O7gQh00Q69/3pijj//4AqT5/i
Dpwt5Jr1dF6PU0bbJGv3CFkk98NGRZqoAaW/9b3X8nIpzgmi1l0kw+nVao8JPYmkaVIADrvU83NI
cek80xLHprmhCcmSoynE8RQepHrBGeYaJhBLqj5GvPnA5PrHOT2DJrjDGOk1hDRWSisfLkCcBlkE
cQMbBO8uP7ctjXMLdT8b2jnIVsWGvppuRbbsTgs8EmRT2xxK569Al2WqUOMNQRGqu5mOi9fwwTim
N37hO9+mG69XDm5DxDw6hYHFjK/CwfXogqa3mXPcPtBk0+XiwGvxeO/KPeAe4Nf6baz0W9/cFlYf
npywD5wYoXr9AJ2b2anIJZH4uJgl2WPo1UEGOn3dLFk4j0biH9sqFvzPAJLhhxHgPplPtvjVOOuk
DQc6o7aLPSK4zT360M/sOzCdIEM67YeDO4sM+M4POJ4AfERcbzAKGsqED7ov2Q4W9AJV3tBIfjDI
20lCiLy4fDc9sybLNYqqe3Z/mq4N/qN1lM4RJenwk/0swAHcPoLM4RheZ7VfuBmAtlv41wW3ZV8x
mVc7p9TQDk7I8DIArLDre6UqESnVTi0EnhH+ZUBl9RXsT3F8Rgv49JNy2SNleVACS0tC5CN1fbxT
icHzayBInb7KpTrrBJ+vAFgh2fQ+T3Xxn+Ep4WMTnhXrGCxv6ugfzlCLCO+EipdzFoXS3g9z/qoW
/7WICpI82sKPRQZ4jKZAZBNHHoZ9kqQDI2rgHd/9N24Le6yM0phwg9LDWQL3D6QWw+/ZZSgZxsyI
/Oc8jetKLSHQDngMo3G0Ac2yb5sSAl9vwjuOhWnQyXj6ZY0I15Qdt8hW2pugQex0m8z4l9QhHVNm
7B3KCdWqoz4S0BY1SlRThfkVMDNFOnofimo3x13nMeh180cohsQUa/g38TLEPZ3By3HKJXegeoRz
jN3NBYouXIMNqmA4UN7AJ4jyk6Rd8MPBpSV9kQijT9P7bVjOZwflVAO2nIgMfAPBfLW6AavupOkc
/mOqRTP1exTij623+v2nkBg3XFHL83hqhCXdIsWpICqtzpFOmvunZgJQckfH8ffFAuCd9eDuSLg3
gvZPbI6BX0HrXhCMwyrteO5d5IZ47OAqREEoxBqSq6xTBNUi1VwA1ccN/LgmL1/8HEh+cs7ohfSX
vYvfEVFoCB58guKLWwUewM/BEdudtBgyltKu6fCREf4Z2VpfbNFf3vDIHeVgand+zgmUmYAJ1mpd
sUGYCB0m/+JAwTpVXQ9TMfR+/NajxjEJkyeU/bCw1eA3VkpzXJqzHs3qHfqL4KwA25HlgFgmoeah
rANRtnWxScoRcvQvo0uicpGo/UsPnU4dzNGcZ7zklIoQ9uOvpNvvxKW08dMOyIwqkgsGVkU9m0S+
m0To0r22mwH00XUbcVQ+KlbZPTyXsDd7DhlpllnNR2HZP41dMRWAbtaIULvz58UPdiodQMMoxZ20
Pn4jAoh5MkzHxFHKHdICm56B+Gkoe+4ZL4dPd1BOegOdOdjmuMcR0CzKxpc+ApYItvMuYzFza1Vz
kjyYtwJz4zx8vyfKffs2sdiI/VSEHFtshh7+HMwG8jOBUlULMThTl2hG75RcxoPC+MEy1z84XSc3
Y9HmzInZf2DJDV2/G7XaEtMlqp57Vr9qwhDOvEhZoCWwq3bXzgW16gKeroOCmqdZhP7UOQYKStEA
LsfgugKeieL2VAON5ZnBYiDNjDMXFTYj3evd4PMvzNumIzAMlrwNI5jyQ6nOwpqzMjj2pYSJdDxy
tMEa3wV/GAIToddWoBuhymtKSSgE+OI/TcQ4Ra+QhWuSvBA0dfrIxEHnKKlB5oV8/5cotOYfCAI7
zIiK8Lw43W/FYs3jwqF+Z5A3MWCT7+40zqW+AYvDyVr8qnsj4OdLbK58BxVCxLKjy/2CwoIlm1KB
eIWQWsJLX+ObRjn19Y58VvFOJwFtU4tMbSp5H25t5XwmQOxF0TlySpYG4UHFS4MordsdyuhAg+UG
J3IIpyEg8TOZXbg3SP86L4aoku/Nw37J82VJKYDfBaTHl0iSPGwCiHzgHtQJQ7eX+SZVdZ/9s4hT
ryuSa5/lIB+gSncsTQVgRtdOGFL508EpxQaMqG5OcYFX4ZWItax/A5PnW0dr1Vrfkkkm6dzg2rbb
xq8YoFqmLAwhj6Zxhg9mPF2JR5ZPy7t25rp/KWz7uBRUXeXv4ZVoy7SbSfhPoeo7Zn4uZJ36ezwm
/cwZRRezb1MDcruHbRa2oscreTMujY8C0RdFumi+TGoav7M7COd+JR24mMYCP7eWaR+6RnQ8Qijm
wKQJSE8vAX8GmoGQisnc5k6xRL0WcY/zd2W05FCI5AdZ43kEeLwkHeFjRnEJOQF0EhpLZkjdVc0K
U2rY9cLZkvORvkuGH16SlnmeZwyTXJep71Evta5dyIPlvQTMPP3VSiJ2tgPCYlqRxnDl+STereF/
W+/oMki2y/OMrbM40928Tqyh/4U7eDytdld4DajW60NHaR33CLyTKRcyexGluqkUC6504UcElKLN
bEWKfGuwe8j9UgbX2aBam3ExNrnPU//qDzN1EN7/dthMAP5cE5ZwdZy94tqrMwHbIKR3uErVCBdO
0Qx7/lkM5/DjkZjgNhGe0nuAPfRVnfsV3P43UiO+VHKZhmQJDyGyYqn1N5HC01/Mf7AzKnDgjwAM
IXCFDsuEa+zcsj+xs59HzEoBM/4YBCRVuacOLpNZ9yVryl273L6d9H9iP6lnbCsL4Hf4ZGT4phFa
qSDrgIx1SDNftpeQcDwPEHTXnX45DLa66O4/kvmg/2NsWyQo4ZrZJI7efrPAxze33mg77aQBIrN5
QoPSzw4uGwPWJjSkEFA68axcPIu8I5Rh4DGXAAQAOLuzhfWIljLScXZxZDcroXowpBlt3wy54O8o
gcli+COSxxNP2HWm3ZMyay+7+dbOftkmkdDLQjr23+vGldfXl9fdZtgrM/XjQsuj0wZGS3kNqJ5l
WqH5j0reRtXiajppUKpt60FksHCZHQhz17A4SrtF6aCkBvuBOc8EHVcpNBZzPbF4/DyR13MdXxTi
cyCPdO7adnsRsRqu3BYhxCOlKD/phKzSuF04mYmo4qLQk9afPpTxgdP0BoQJucdAPzzk7qzMFjuQ
fcWS9+LmT8xB8aPqB19wdfIU/6OhZvqz+ANFbmSgGHXKYRDDdh54Ig9eWsnmbENuhCC8AoLKldBk
mtVkeOjDw95tMvOSS1XuGRiLyPMnMtAGs7jJD02GHAwXmNbeAMNB69Z6o6HZiROee+m8a+ttLIKn
H8rfw/EnnLi8znte700by0cWvv0kJQaqo+6eIvK1IHHiEsgQkPJk1dhmCDp8/gWR09pheGGfvkms
g6S2lHkA9PuB7/TQBvHeGKI3r5dg/BLwHuZmZgCMj0f1MrbWuJRXwO6AytEZmeiqz5e8JQ/UlRQt
upWHNsWL1/IbMM8f9z74wMSWwR+btqzxQFtIiUaSz3WNY5MvX/v7xBbCiJ+KLBAiTDjOPWLupuQa
W9VwFMbsbnfY/Ihc/jIkP6/see8ZzMludZqlLt1Skl29Iojk0oTVJUK+KR2A1GKe4OwefjdQ4sW9
9dRjqYP6eNEB2nlqB13lGkIVlW13Eu2czpyf0AoA334xVoH1xriyNYgjq9qXr73fVZQneHTw5fI8
95fCxPDiFUM545Wax/Sxee9THPcJ6nQVS38JsN+6BXk/y8e7+5fWEEwGewtpdAI4u4RwEn4CJBWv
bSPKhIgr8x8SYnetWtBxBqCc71O17CtguZGVx24zh8Bx/jwuuDVU5ZFPtlBG2Qhy+9CGVMdADLyE
DYWnOzK49zR4ZD3W3dy5s91NKSrpbw2NGHwVpavaJqjqyXpjNrQlWFFysElJH0v3VHecknrbGxLL
qiFahExqrgoHb2y19LwXXBOwdl8mYyCzZpFm8dD90I6NUrYjf5USK/ddfbws1HkyZPvharU9pWn1
O1Q+GvnztAbXHlutqkM8rSxwO31QV7Zqa19lTK3saNuqK9neGbQ17PFHRdNBXmhYPAkrM8W6oURL
7K4v1XfgesPJPDngVIpoAZPTx7MMIhxLID3UoDvWmkYJzsYoLP15SQQQ9Ro/L4tm4HcVNj2xBmga
2YuQvzM9XcDUBAInLFF7k4ghWA8BhKwr+boiURMbhtluM5XYmBu2CMGMmlHHvh253iQ972n5b7Jr
tAdan+766wFZ0sI/yVrWLMoNMj6MXURCQK+twj6OImakhkbcIQlXB0OjMru5miG6tO2SneYXt2Zz
VVtkSqXOWTvHRoWq0PeKd5p+MpkQTeNsT2gnwnYvXohNJYfwdPGa4l0EiWXCnn8fCi5HRjD9RoYS
X/iRXXQFBen9HYKoyZcQesqakIC9EN9pqgsBsDk0ToM5viKvcQoxTqSR4Uhjr8FOuYII8mhm3aqE
7gwBTvsumeUZfWOZcTMt9nAk/YN1CaO0gxeF4VO8LuXItPzzmrkTXZEhIqFLwsHCZIpVcxLkByoY
ioQS1m85yQ5NncszCyyeHMxsdF6ixmV+SGsuCJq5fosIc412NTAN1aLU1ol8SnQpj7QH/CHE6mnj
Ih8DxQzxW14UzHPS9Nt5ZXIaB2HnANmCghkjj0+bj9iOpcSG77gMTeH1dty7rBM1mHpwyQ4CNwBx
JROEfIbbrnpLaKoz4ZMTYslS7AHddlolIKS2o1CEKZLiyV9YneWQa3d3Gk3H/r0IgH52qjvxG3da
x15tdmOFa0UOC0a9NKceWKFEozdW3GJ4tBTX89VxsprUbaTm9cKCQde9vfcol5tPlv56CSbwAFvc
PeZxt5ajE8uh8B3Fky3dFO9EMUKFZyMTYwNxBrtfNvLKR0m6CKmXtrIZ+VR1WK6s+yxXlPBu+zs9
1CGyKR51YM6cFfxIcxph32H6S0qp4FzboAybEtIyZwDnNiH/jZY31d9TimShUK7GzCDPRvPp59QB
RIzMzKRWae8g0DWf2kP/AecXf+OCgBiibuf1Xw3HP3W/7BIu/xUcYWmmj7JO52ryV5s4voMsvYCO
byCgHT7GnMGYoqgx+GMFQ0dWyN6eA/9a9kbHtgGbWiSUxub+cNMYPHhmalEc2aAEN8iFJz6EePY4
rrzMf+3H9EnNu2JhPvurIo5nPShrVjSSpHpazruOtHF9dDobIIHGxgSmVSA18qUoq/3NWu1gsYtV
rRMNnOauYRvwGLzeXSquqDvoDJka2x6Z7VM7qMY2F07/R4BQp3jKkRh/xWRTDB3renQ2sLSOIw9X
7QLEZvDByEqTR/9WsGr0xYqjeANekG8aLamneQlwYRKrEu9z4hA3nxyIiJ/AxFWGUCEzVbM+//kk
tfATZNafdFmFtTdmP1QXA7Yx1nTfqv8k+aeIdjlm5uGWUqBpP3oSamMC2kvJxf1YeDwpoohnxh52
14CTwDN01tZ4SwYb4CQkvxCvFY7vwLOdxBbdk0pVPURBhHrVA2TuWDyBNIzHKtDRDXLltXirKdFx
wnyLzcVEytdBbs45vlQ+Ma7XdnBh/OgYKXl9ZY6qUoj6L6Rx9wKwbKt94gBE5uHzcxac5rBfT6gV
xGsaD3FelMJ9vZ1AJi4Cnz50adS3PRqznXhtdyyXqHAeXS+ABsBBOAkYzgVrol7pl/rpW9GnhTZz
yMJ7TJhgrqn1LWaum/NKNgrghbvRPeJ8CAKCX9h/uKDMbHKdO4ZHDexnEu+M3ndAh5/tuJ/xT+e5
UXsGW03MAGKH//MiQXPJxcYGWtGRUa9uax/wyohb6BE+QyxV0UioKapKH6tLMGpRLygOuVDQkrYQ
E5TVXhgHoN3sl+UeMiick+QbKU4nRseQ8B6+hXgt7oiKLzjZy/CbV+k2mmj+urkC/o6UWLHPe5VE
2bD4tucn2uNJYJqlQwR0e8loWnTAi2gm9CieKqnfVlj4V74E2KWJWcIHd2vpb5EmkVC46ZQM8bkp
Sq/5kAfS/40NNecHfBpJvVmn8pCio/D9SbNwTE3OqiZj5RD25AlxgXvb0AburBOjEOoatVCUr61D
TYgVulHholplslY6ScKnc+it8I8/TGdR+Nt50LxN8Ztk5OkSfFWG++KSA/kEz1hRVYTdn0JtF1TL
6+iiswplY3PkvUNNf1HebFVE/VSUGdot/e3XqUir5eD9fMEmdpCciMboFi5sOwhsr4tsAhIGdTVF
Gfw1DGxe7X1tBOwkgOcChhEelBYTiEe8rvpI6CGYdNbCQcd0QcQYU8X923v7usgo97Uc+laodQ0K
NKkrldorjQ74rh65WMPS810gt5cJWN2FUcomEOCJUIKLc76jNNpEBt+R3W5s6NT8q3vIX1B4rxiw
8XRUmyUUerE8aMs6bSPq6E9hpZwPN/iLWy69vq0TKlyZCgUzf63dS6M/WhJzfRFlaktKsDwSVEz2
IjGXxDWptchZGvcsvdztH36UQ74VWKBgRoFduY0U9rRzgJiGuKjKng+hyLYkxEobkJmlaqNvO5tx
t0o+Iwx1Tiz+sTp0iGXMV+nSh9rJ8HWdbMDQV1kbWc1FDU7EpotPUD9XnZRwbbSEETXMdBr1+yBN
mczroKSGN9pWUXjt7ZksxKFJoUAMC+gjdGUsGspDWetqe+yS89/1MvlJM82jvetJrZELUCwoQgQj
O9SbNT9OQqqqRZfFOAA6rsktRZwwiW1B8OYKe41NPwoPf6Cu/WD10VY5c2Skxm//hO3C/EuagyRk
ipNkqu3jPfK/7COjTNLRfPLcjxvpc5HH6xj145IV9RHcSW7q2tATk96KGOORHj8DoZOL0OtzaNCG
s8DAYfr2MSF5JHNXoDTm6WSQr+POrVgSJux+YPy+v0e4++xTB48orlN5I8v48U6Sr1uAGs8yIjhu
ScAGRSMhAMHJfmLzP7H+CUBuabLCJyWq6UExCgPIRKyKtO8yCgxMYcJnwB2JB8eGH9pKEXMyvyAC
nccISEvClsJI0B6FNMBdl+7LPWHlcjp6Ok2WCclj1vPGshNTrUXTw3sB+1gzgnwO/3OctDorUMpy
/8CAZCoSOoVwpsZ0k/rA2eXjWM+fzUgIaRbZ0sfixPvT+6I3m5P82F5ut1u/TcjFNXidZ24ZnJyJ
lCk+pfWxV3szy/W2PVFSfsPeWfn982js29Cf468uzbE5jDss0xULkTKxbYAPc1UKuEdhPZLUBJiK
X2brrYnUfK1XYqNhH9ActG/MY6GcRLcUCj1HDE+6RphJXsmN2K02UAOJjbisZqtwtfHeK9cx/R35
S913urptmNSD4ucEjyQq/EQ+88cxnMCutenArSaerC6x9vgZqOLgN72pkmWY2ajRDJFPk+mf4ggY
0tjGhe64AHHWQoh0R0EH5DlOXHl5SRYPjKbJH1HZ8mPuAWVB42wgq6vIRtetD6SPjA/1A145h60v
P6d1uJ7Z9vlccsq6lqdu7NDYk3CsIHb+f2pvsEv9vYFkSsvYrmTtnB6dWtijYgnU0fiiBi368po9
MnuD0aOPZlceLhV4Nh2QMRppg2J8H5ekiH0gnUoTw/eO++bV2VbiVAcd55fLeeDmAonAEhsH/MlJ
AbgVO7UpEoWzI1vhXu0UlHKCb9DQmrVTiq6kYXMA4Y4H2Dp8bEr5N6Y6QdoJ98LvF5GOAeGcWP0w
bHvsJrBPL51hZfxRFq9ckFnX6LFxEIfijzQvGFZBAp7iRRt2Uu/WxEasM8v2/m+XkehAnWS3yfJ/
zxCaYv0CH+AzXv45IbtAoremg+ZWJLxBPr5yiQ70BR2VtxQ2CmRI+kOE4gBdOc8bgcNrwhS3Yxod
8w51WgX77+Q6cUxmp8vGOWjF/P6Fi2mR8fbCFlf+ahjEO6HdV9hxhJwiDrX0yiC6kHD9WVJ46goj
rqYmYMhdF28sUOP9nZYoYUdeFO/bRRjcv9iVsqFVy8Q8NOum8oW7gsciZ8dnn66MtR8JOxPSW3Sc
05dHG8CRDfLZmlI0jUtybA4IkqZv+VTk1YYZrZcG+pLDODGFshXKbMlWm2/bAJotyqluwGonTAav
0k2oTZMg3Q3Q8m+HjzH0xJpBZkXaq24gNjIgno3uV8zEW0RO4FYUsEgewWcRIZd3V/8p8LF04FTX
AYCJm9vnR4Eu/Z04Pnm0Uhz7pXlGI079l3Pg1KOveUH2OBRLc/pTbPqW73bAEyRX7Vs+XyOa8SWa
DQhlSOlzMpS1c12Z6lKtCkhq+vdzJ++z6tphDWXD4afIrvVae6JtZ9uzjdrP/vV5jbE62bYJrW7D
PYBJhBtaKAQ8keeBEvkLY0Rz8KDfDwSvN8Is5MiwmbwE7l4rpNSUI2qeOz+AQLCc0Gha1YdVJ7ZU
YrQdcbrrT+b0imVQKZJ9AUX3cpqv5RjGgRIlSS7z6U3K8mba0jQQw+AaXX9LI/jSqveEz9NeoZZ0
53IqEqTAwfAGImgDuASxyl4xVHwDE82rn/E1OxxSoQEZSXNQQep15Qs9pFCmAnQ7PphdMbdQMszA
zZTOV9HZLnwczwzlfvaxHMSjf4b+7ea+M0anfsRN78p3YlT5ihy1PVH4d1zG84bz58sImS2pPid+
Wr9lcEnTwwhxAFzt7S1huhru7Yp4wUNDsfg/NjJduZn2AlZz7CQORnXzDsTzS6johZEt37V3HmrI
+h1arWWiqUhUHnKx1HeyZFpbVkvH3Uv/bJgUKXZQTK5ZSQCVhyXYjMLTdCx+nBvZQ3jyIIbK8cE9
In1cO1UaF2zQztT6cECnk1l3raseleB0rsSGPBu/SKLe1SL9rrgY3lAQd4fqFEWWxQWYtxdljCuL
ZdwLMjGx3n1FaZyT38b+Q2sBX7Cc6xcbngK5r/TwaMOHyDrcnAXmaqHScZFZDj0+03st3+boggaK
dVpxOZkyqlCevSOQ+FE8bU6kHnRvR3fB7mMxvhjneaImQkjVmtGRQjhx192U+AJQWV76h9lbnx9Q
7qCApE99U4n80zceLI+Y+BqpBbE53ZHhVcjgVGjD4OJthBGmqpHVXguvoXzRHj5ydTjxNxbyZ2Ef
1HgjbrmvmmV3hNpOX+X0IwNim+/MvEPqvBhc1MEYsjmSdV+orx9LK1F6ib7GNN2kIrfsWzjXRFrJ
wYF/19LX5V94jOdpTMM84iAWwicAM1fcYq+cUWmGqE62anmzEWk6scLTVrSEiiSvIjkkNV1rL4aF
j8TK+9yPD/0yTkkTRwRDxiTT2w0xPNiucJPoYczNcuzoRAZvhnywDJhMM4ysnWscXkOZEovdZeUC
5IuccvEFvBnYxm0rNcFL3lXeJHinaT77eN2VoKn7+FhSB2zF6DQSiQAhKSGwhk4DTCbEE/A5jOZ0
8B8KiLZcbrTfMk77AGD42u5m8Y9rQDNyhcm2aS29+TguAvONscV5UGwy5PFGdLLyrU41NZ5nGRXY
8ByHI82z3cgX5kf9bglCfc/jak6wRtA2NdYbuL7M+iR0JeYo59i1GFYZg/pCs9cBq5HEJVitHNzi
pW4CWGYog02zOdh9fYpRyS+ZmDrDdNTlo7wtlfNovgyljWFUJk/s2mfOL+3PRif50W6F7uKhbgR0
1hgfQWoPxawxRG4Khn5zMdqhnz3I5xvfKQJh7bCywccMLEHJVeqinmbskrrN7mjI0cVylU5egmXR
nbjd4kOVJA4EVw+eRb0zt0VZClB2q6ttw4F6ZnS/lDGSY8lL4vEgnu2Fg5XdZjJuTtKTBQCY8ssG
RC+rPCnOIeXZzww271LLjJje28J5eAgGwkXvL3qILNGSPqI+gq2RroQ5qe+KOwfELz7Qg1bcUJ5q
huP2pdylJTQkgv99Ea1q/HUWV1ZJYxZwzFAsebzVG/EGe/UVQpV5dBwNMgiMvgVxkbyp39jVtl35
i7wUyGHefrPOGb33QnoHg4CU2iSMMhr6aXLgSOiyBTRfyc6ZP8DnXdF+RD42oerqW8EY/JLhdxF8
H4wepK8D3LTCcUtaDpXTTdFnBzOF4ZdRsZJ0rn3qILIspSPzDhd3eSjVMPPGVUw7ptI9EVu9yq27
h008iExrr67qptoDXRt63wHbLmRDHuZGTqmWg1Kv02KOjcKILUb0kbco6j/x3SRfaXLwG6WUERDb
9OnQRsXinE0kg1qnTX32PT/2QUG9oB25wZ3hcOedcdNnYLL2ZNcMnl0TLYFbeDwGexcTYMH1UezU
Utr+ZCtrE8ZeSQsHsj7DLAeLAxnG/mNp/ljExsWCqtvdfyNpdVySbDKZ+pChx22OCJbUe265A3SK
k8ZXn10e5zNURQuPycbulHwbcTseezoovcfSIi/3Ra7xFueofG8QCohL+4ln71rla2Q1MDDjlz8r
LFy00W69ifmY8tbJ9eVCy+c0PVZsj/j+91IkI9yOHtBIZQcIAKzi5293FqOByg8wypJZuXz62KYF
2EYGwUGQ8p+dcmgOl1YLe2yU0QdqSg+Ln5olvQC9xcEnT13JP8DYEn4PSe5yR8svw0Fydac3nKDw
YxQgSpAAuYBbSaQ+fpIT/hiuFasKHsOxbsjPE4oAiVjb6rebEvm9RaXe7URnCJO66uT+d4NLfdJw
VLtmhte0LX/1Mx+ec0esmogN5XcK8weT5TZS6eQmWaUyu7BnX54sVKWtTlemWipeWZLjIfATgNSa
aaXrc3KvaF3tWarfLf+oGOMOySg9eVZtfjvwucwTS626ek/6z2v027Ddgn1lYh6ytEHrO0+A/Ehm
n+V2Vrl9jkEWIrnL7gs9j9JzuPZ/QiIDIYoWn98bQ3waAwAHaVM+AWgHCJx1DHUcn9IRmytDQHQx
URFSjvDBNBbWkwE/CT7wmxXfA2Jq8pxNwxbWZuOUzOCMEISMFktB5OzTj4XMLYTEf9XZqyRrsG1p
0mW1tcaQoW6pC6W4jE0uLOUfMYNLxnPSZqaPzvUFOd7CMtbbBWmt5QXTdH5ZDS5tq6WIpuWl8CFr
KDdchLAIw8hrhBhrYpqVgqG84xQOK81UwYkiR7QPzCxxwLr+67mHClSDl0jBe+c5Gh2zjHLtwPeY
UEvf830GjQUEzVxCd8ubo2Z2c0V3ddkzw2w2eL8yimZNw5eL3/U7ZFSEXFONeRSvcF/UJlC+/OL7
mPC6FnEuLISebPisvq4/7FciGcdqNw38cM0hxGzHIeOHtzULSSfCQg+LU0TDkSRcPr8vvmxAxoaH
2/Tyi6StkqeXe7SR9SJY07ykijDXMNb/RnpvQGOWgBE4EwqAJonTiJ0W51kDBwrum90ogBE+8265
JTKmzZngH0GXyizBSIS/FPHorvDqNG4jxd1Wgfaa1Dp8vJNrFHYeSxTvLMwnk2ZYAedmzLtpEv35
OrflPvMY66+a/g5ifi/aPMqQXxQNXo9EWrdLv7Txo5HPe8hmI1gO79Wnrd55cWaCndxonG/+eYwb
7PIF7SMPny9MnpCStWyVNRIRU1ElCKO0bG4dEfnNT3WWncbMOXs9uaZY8HxlG7XXs38gOM5WboQ3
Y3/ULPr6++sOXamb0mDfyHmSnj9KxDL7GVaolbSpJO9nqsGuN5shph1XLigZ10XqKLjOXcXFIge1
SPOAn5fhtSLKi+zU3WRqJPWZUkYu+A+JPpeTPz1Z8uXMxhAsh7IwP3qO348wmTc2wNaP03gfG0cD
vj/1WJCTvVaN4L5f4qCOzs8N+daLfdHoaFJBDVgGwe8YsUlWavHFgiufHIOYX+uLx2XKEAakXehB
r7Oghy6bcKKDvepU/aSgwzx57tszbQ/e+iDpTRYciNbyhbxGo+yMCJXGyFy6KhlyfKurcFG9pMq9
nL3e0KEVtA4ZuaYUbn8AfBgyy9F7drEHq1E2V0KdTak7aFtt+VfhyuFbMP1NxefNOQN/uiVb6dC4
N9HsDPHPWO9fsLVCkNr2c/9wtbZuy2INh9zENOyD/CCxxkZRJxVZib5mxK4hvauP8qf1s2l/3xYC
9AOkkDFnGzcEqOfppIIFdSSG1rJJK8IZhwdUFZnmsh1uzKwV4vJZ5oHnsaA5hYrvccuG3hYo209V
JmqcPQwYGFAy4m89ajPdGR3dVQdqvgLCEQ1pDL3ybxrn2etLTsS606SKmmdcXn9qXOgFCnsGTpio
QSpjvyqrPJZicgOzGtToVoFEp+AH4k5ax7QRmcliMcUl2Xhzb4yntwdod6c9jb9BtvLn7jBySAda
Sgx2dDNm269VX47y2+TzW6fntC3ndwsT/56ewpeRp7zsenlG0PDD3bHHm60uw8DzAqkb5cLxlWWl
cBlMSPMiCKQc08R7SpX+XeQwCpyTLKQIbMGNcZsX2DK4wSdXia7XhfeOkL8sS52BLoDkDMTHiy+z
3cY4A/Q3sQmeR8ykggny1fz7MAJjXJ3GH+KJ0Xh3E3KgLUL3bZPMaTQ44ZVkM0Rl6tRH848Im22i
qGoGiP0oRQouw+qdCxrVlrfNZZM6JAf8ApVZS+tFSZCBtmzFwW8fDPRA1uX9G4fVokE+u6dhu8XW
LPYnf8T6WWXs0tczD4m9466MObSGlot/JhcT+dF5vzSYNwAxVgv/PQc5oQIg/xrX8QaZmZ6hWf1i
jfFB+on1aVNDFqtspxUXm0EKLn3ED4qQxxBirL2v12ueGxBjXXl0ELf0pwO6ijHsJlge3hqQ1vof
XYSbc/PYEyoroVH0nCY+wOwmiIYyQ8flIbkeCcsZIvO+8lLuSXpP91dGyHzkke8D9SlqjC0rOYXK
LBpqoENozgHu77WyVLYRlzx4HYB5ksHk0N39Nhrf7fF4fPm1MbKYtF9RCp2GcFxYIftz5j8evjMC
h+e5HLsQ54o5PbU0WUDkxbEwcJVFG9R7MOM8ZBQ3vTBOxI1QjkPrhKI8rIc2jqZER5rmu5B629Uk
rzyTl+dxBJmR1bnbOLnmUXos/s7M8JokIutAVck39csjj/eL1aYUH3F+W4YllOuP2eCwPgph7OwU
7ZYKIVagP/rdZXQIiCxo6NiohzeBxmxqNrBrXx51eUfNqgomjSy5bB1mbCm8zbh+xK4vToljtgnh
vTgt4ISCaz06Po5HabWjIpqx9JiqsK6lUZmlyOfi2gB4niSNn9VhAwwrJulC2RvAyksQ0Y7BtEei
pjWxbnFZNuI2F8e0TG3talYpcJ2vWmdTVrHFdy65rIfuqgZq7ze5J9BuFi/SqOUFkXz3pN4a7FzU
nBVhWRKWFqXzgQQCorGXb5878e/tmVMmzUPH1GxFOGn9hJj6XtwPbSK14YzsLfmatTy1iXzUcG7t
sVvMRhAU6wNvZikq1dHDO7Z8r2pMTYH3bXIQSkHvi6xmLnizGj4JgmUgCcrHwYMJ/hqydFkYG/ym
aoZKARjRN334ayeZk2lUBTav1SlMgUayS7wToxroN7PKRQPrc2ioRpofUaYEZxrd56DV91ojqIv0
6n1L0UKGFClJ8psQh3N6RKUBcqQheTnFq8aI7DWEGsOIQlQ/P7+8X8j2lOkJHOQTuXIv1XTEHGoK
K29U+9DW/RFC09rp7dLfTguV9AeuR0APqf1hMOtxNNS8cIGbZKMCGTDNwcnr2j+oE7sP8jWR0YfI
0ndRpQGcgaB1IV1/ZXNltbqcWmwmoiEJf5d5An6wJOft+ZEHfIowBk1EHsAnhVnnHi0RM9yI/YbY
tKYqCwfHaTWLS9Ff2dOGIXbVei4EFmiQiQe58Ggq4LsvDfhYTSAO+HE66Z6ZEAQsiGttgSyB5sxt
k0La5da0KLbpW+TpEcfinFGytT1dYEOkheeIDe0nfWSA9y4Wezy9NyuV0r2LZ6uty0Qc91UyP02p
359lxH1pA5r9rp7OwyfeTpjL4FNf80wbTpTFZKQ5D9t4RWu+QLRyo2rdl6fo0qj4s8XNl16Ws3Mg
wt91Jr5pzGTHu2/dnKsU1o5f2EGaOtgrBqgduGEe5dPXjxAXbkaAFJc+HZptm4lJEAIiL2X0wWX6
LAvxqijpZYKcvyhYoYiZzEhNpv5GhEutURN/ccG4s/rnNYbnIOq3+4BWiOddjXSxtn69MgsGcjnb
cE092/jNSYSMRBmvKimc51d/7aXHQP1NnLr0XSMO2O96GUaNK0LA+/w4o060jEB4/PbWFTiaTqlE
Zb/euD30TRw8NU2PrXnAm+De0ygK9/S4eBmwZmajgYLJb2PpPrEwu1C/5YZT2LEVFE5xKUnVC32K
CnaeskUzyOwcZl9sXIRjHkeClbLeF5xxiM4otLrv5lUHGZrQdc9mLeMKa/AP0XW7+u628QatSnxU
INIjy/L4tGa4A3lbKvdLhS1BF1FPimbX0HLqRLvOGhzFDz5HMzWlWjEtcv8q63gqdLnIZv1f2Zuk
y9rpBkhQnhX3jyh+c+vw2/EEgNHQet5rX135X1JyLPN75EqecCWJj52VYw51g1VT0FZy46kR5Fta
PRUZexsgjLBG9nIaD1e/Zv9KQH1pafgdS63CJszFXBk8ikaHbBarxqme/zA0gdTMdWDvvpw4Pjm5
7EvaRDQfObI5oIRC+R8a4jjKc/nnSofwkZK7Ys4YPHfQhz1lYwx72FneLbDeU2d1TKzRY8qwxJJ9
1jDeyRyZ5y0N3ckYTrWYN5AQADu1jc7L2GC2cvMP4ODbUgoA1+hotoNTiuvp38Zi28K8rmbuyV+H
U2RiFqorZ4wTyEnSgX+JrqoCAF0ArsCeBOdTtQlJWYMkiHKQTJ47DOcFXIjHd/AnJMshwykn0h7t
beFlZdsh1TLces8BYihGCw2ordyNqd4MZvmw1I8OCKolyMonnqO6QDGcBFlsK4j8gPBbhDit7OFK
kiibjBuxndhrVigQSlYlOt9KzoMxcpFBcQ8tW2/5YsSZd5HdhW5qfuE8XGZLaVNSNawAW2ra5ikK
q09drfUVdcwg8p520ll88Ub3lYsLND2MbRge7fk89ZkNu5GcuwCfEexdBIR3W0zVq4TinCcGD6d+
LqLwE0rAkkQvKr3AnVtciQExJKO3KU3sVKR8vrPe61wjPFjdH8Q6sTIDWRZSii3u96+NX7Kg+EEI
JF4MYa2+zNSxW6aiTVY2u83qvdUxtPz4L9QOrqNvezXOd4WMdLbwegf+7sFPshLyuJLWB6/Br3ee
Rz1ZF4ifkwNMcXZV1DCHsQ5z/BTV4GdwvoSUW2vlAHvDGRe1BJz5pWkvxJTX5OjNSP2EX5Qr8Gtr
mLFKNXdoDLTg0P3y/ZlQacJTN7cz3ZBk7dCY1ghF0c5a2LPCgtqZlIZedvN0hXV8Gl2Bzy5fecQq
9pqoL3l00tsvJOek6Ax4lmvKB//fpal9mYUqF9KbGdA2TP/0W4OWyacID357ba7to89xQJL2oGn3
AVDwpwFEA4S7TcjbjpYhVkD1Tw9ID7fcd5kmxIXR2culC8HKIuXUZrrlcmwsmfm1YtDuSYroY2Rn
i/pgjMs5SnHxGj5uqT0fzMZ/YToh1adJJSSsXx1BiBvYlLbpiOPTE2IB3E+4zEvtm8Xo1eywcOO7
tbQbYCpBjSGsHMwrYci1dpqmsTnmyjCqxjKmXgiZgG7NvLAbFngrydcwm4oNYsCdfRdg2f3qy/T1
+kBu/xs2hZplPsAyt2uRLWFAXd5SqJgg40k8JQ2GgEuFAjGkDuBwXqrdud1ukVwD4n5T5gR9eSZU
JCTpKnLtMY8tWut/bwJBuqMj0LLbpicC5qiSu9hoCnKu/ThyLMeR3NHJB0Dq7mc1d8TR0YZAlwRq
dxXi9dwkv/OvqO9upHuJTNr/CKFZKHMPCOjjf/UaEDvlQtauVbbXi2FXw19ByKfj//Q5WxyEFF5z
e93fNmee9ILbykNmOwFxyQlJ1Tlrm5+horwsdJZecNk+mVuELMvsorP2Q3d1fYLfNWAS8p0fiK1M
3tiAtGMiEI6J1S2LsRFlb6rEsQYDFWzalBxCo4wmTqlvTbt/XwdpZJBJcRTtgj+DMOPD0Km52EEr
zhWlNoVHcFMXgR/Y+bexJwTxdNcG6i7xKy/OZocVrDmkx8FTte/+6BlexKbjFxrRJva7k1HzbCpI
lEHOgpZ+SYYn5DlyP32T6HtQ3eUTpy6zwo2Mlw0fqctmZWH8FmAeQZbjWhARMcHvi3xFy24z/6tM
Oio46E8esIm1VtC+CikXUewi8D5wfvpQM0FfNhXRqhVHEcUxnVE5lh9sEmOUFpPZDE5QBTQE+mUi
pQGSeuYCTyLJVFo2SqldqPfR8i/GHhUEjfrUsAg/KbdgAFv9b2SHAFdbfQo3NCxbHtlUe1Goih5K
eqO92B7vILWj5o1DNIIidygUyiG063am7YqjNEuvFXwKXjk8+QKQ35Ox3NYvx3CxdtXeDG+esUHO
2y9S9fTkhxYdxrARclmXshb1e4gkugLLwVnLLV40ADSVOQY3rc/lG3PvPWcXcUNYH7nIeIebDsrn
rZni+tfxKW4VSgXKV4sAd8CacQQZueMenbl3Mh9lsdLYDWMu3TVWAmJk/ZFgv4xZQUFmmGkuNN3X
3EP7HBebTgEMIzhucacvZKNlQNm08B7zK1NL/hB3Ew+MMrk6v8+b00rQi4wx0iv0TRpKjQ6BDrxz
d1ygsxdDQxu6+jtGIk4zt5X8+ago0vnKwCR3fI18S1BTukJlo6pr6c4BbD+QHGJH8TQdFIt9Z4YB
jAFxZSmALxWhMUJAMBoYdQ4Qsc23cf8jn5+5oSgZfbnH9yzxFMumNZ+SlxaXq+gArKfjoloZo8ew
e5NZpwgmr5OyWDUT5y5j7wiIshL6HxojQ3Qk9Pq/YYHx9qgmvVs4vX8wu5UhD9xMnb1yg0A+rCmi
r89LtQ5UGYRx/za4o4FvsIRQVCIHdGCa4nfTeD+/ZVR1rYfpTCfX7smzdp7O56COQc2aplldsB+n
reGF4NrCfR+7DP73/lxZf35yn9M5Au5IxLQNUMV4W/pkk91Pj5E3YkRPGUPVlhhJMnZEKZk6eNvu
efvRmXEKMjTWRvD+XZA8o6adv+bcf1FYoOmwZ0Kab5Vy+XkVilDmjRmafyKSgWLJnADUiG2VY88t
GB8B870xXIA4czaTJsmoF8Sk0/Q9bB0etL5CMWS4orfO60ImarbsLBhtb1PLH0/8h3s/HFWTo9w6
cQ/XsCr9YCZZFEhkAiJstcUI6NUD9zyBYTEG3mSpaIlvjdl4AyKPI9wAc3g/jNDPpzpKzPn6Ru+p
4SS839nYh2/1UgMUhMKD74JapNpzZsGemizSsktDuLRAkb7MhD0CAt6FgwRX3xo59oW04e89JtsJ
h36RVcaGIcT/YeNsYCTnJUkPmohMXvYSaCrI4OLFLQUeRW9a86EZ0U37Zmn604Tk0RsAC5nunvF3
PctloObVFYB1YIGQu+aDKWPLoBGPs4Iz4NQRj6FaSHQe8VaBVHBO9E4qkOZYMIPImoxW/ComFlGF
mMAddwKqkN38uZAp0SB3EIA2YStBnAgF95oXKhjDjrJhhLoNmQ/3SvMYd43ZCcVowyve/LPOr/1H
qrUKqpFawhKumyRTTcEQVwW+8NRb8ScLiroTW6pCZFGhwMEMv7HPtgQbVsfJVPndTFFKrs4GJ7+h
qwmV/msG1xdFMG7L8K+tEQAVgSfFpdluJBQSPuwrVg2z22SCBy4v7LiCQ+IokGIspXgNBzpv0nYI
3ILzFVwH3Tf4/7cDz1R2/DUS11hlbP3zLo9PP0kO3wjcMAZhrj2RKp5bxUCLSfW3hrLLODUX0c4H
JkpqpSjCg+njNsJO7/qslg6hj+/K6RcaC/RqDwqEQ2jvrSVAURKqxUHazIpg9YGuhS0v+Jfdh34i
e3nshbv2jnbzm/sjxT4/dLApMNr0Php8wsQrViKYV27xGBakRGNvPESGVL1UXe0B8HfpDa3s3KeY
vslkpOJ+eplJF+epb0HL853TF0PCmnLBLUO1sbDQJs8vEti2Pc2hkgElWxvRwTVHHCvtzxqvaQU/
iwjulHuMbvWLqrj8AjJFI/PUyFQkagzMYfPWXUAOim+ymzVHYlLBBX1H2PRrL638CPSNQo9Npkvv
SxsXiFujh7+BRTaXLnIrb7z0Lew9fFajhUTv5BW5jE2StSDBRbVa/fHZW3praaRzlptKzn5V3pWT
uNS4cmI/PHWTlv/vkFR/rBPMNPTcbxM1gmFSNXVaJsRfCCtO1Dl67aMN+0XOj6XgHPX3/blBekw9
aPkhTVp8O2VOjPYS9gRhCvDgpYv7Ejm8ZmN3mtMBnexhxR58JL3VLZbG9iLdn8UKJ01+z8iY8og6
yCAeCm3ltnBTpTaIK8s9Ep7WKZTKM/7BhKrb6daQl5QdzUDsCnsLcyTxhvY9f3TIAVcwqScDW5CQ
sHfAjNcg3pbleNKPac8TJxUzVV62qOKrW6mOccnkgmAoEtNLIJMoZIN/vV1CBI8cPUI5fUIaiVbq
XeHjdhQuG9xX8Y2OpgVCrNHeeoppsElFh9wAJFD3l2yuTrvP/fe2OuB8Pj/YeZDmKL3xoKXcyyiH
+lv7Feg7s+saOq7zCWYuwsDd7A/x/Mv3OyZGgJ2xYtHePSGZq53X2GT/wEbl88fVH9w4Fv1+REOa
x9gfLrlKAZe/epsilQxZvbZz37QMWU+JUWHsoOOxjlr34YQOAIk1UzZHjYs5amjJf8YNEHIUpBMB
IckiJO87TvJXqNq26cxAvbhdlcMueHMYmHkM0nnZhhvIgIrNwgExlTkrPJW/xy6vJ9CslD9t22vR
ytUDUqNyNZUA1dUa0FqOYG3nSuH9md0HEWBNDwHZAUqRsNmdERfwGP7khlS5Yj3RYAK+FhFYKBlJ
QJTLEH7NTsc8CdNcmMpeEJ/ZcoAnXGWm0zJ+9r74NWZrqw9nBvL0cOGXf4/5ZB5rGz8Dy5GBNlVH
23e2RMvlNWxQ5NtcaeWqlxU113BKCyyvs9tz4AtMPGgR/EDV7vND1D66Oa3sf2fUKSPGQgVe1KLM
tPk1PjCoKf+jFU+Df5jwE1lkdq+0KUg8kXe11JAWk0lgGl4HmAYKO1Ox6AqgTBkUnqtFki53/RnP
ABNe0O6GQevfDHcZl5WKxQ3dNfrCFgBTrobBSkHJ+qc7GXrlnP/+boL8wbCAbF2jFoRvDf2qpx6V
LA6Mj68gAhZtYNy38SigtsVOVyGsmOGHjKchmgkfPvgXROwx9Iu60oR5+ABgrRNP3qeecBJKcd2g
b/uZnSpgGL2t0LMQ+bKsJ/0tXXe/plwx6MRLrXJ/0PBViQKRql+hQHZd6A4NW3IA5soQx+JW1FkN
9z/hULFwEE8ECKkL9wnO9r1gqPLXnZUDlYpxScCHgPcVHSmSwFPkFQcEwBxiSOLjaKjwKS3lEqfN
chkBkPRdttYswVLAsN2QQjQHGEKNb92lvl5DKuUKBefa+SPUYKnpjcfKBNJVMVbORMtkmOoM4ufU
AC0LhwTQAygmDmkvhwxRA+EyLXi2F6SbJdqiA32Y2BiuwCrd/AP4xEPxBReR6vyKOwMZ5aYXX3oI
e9QssfK9gX3Vy+ZExUpZZ3TYWbPa4uV7mwKbPPLitFNqVBGEsBh+/Od68peZURbUxV8z/JVWXSeQ
UQlNEY76RJbwe6SDIGhV+6V9M+whmQ+sjVk4u9N0bQZLL1PlIqIoVsPDjqMmtg4rv49Pja1DsIFx
6Xzzn0pUyBM+tY4Y7caPoPsSjbCkLy4iKcIebhG99jgAj+zrmR+m4Z5+tjGZksg6fJpmfMRSqkil
AUjvUclwHjHxRCV+DAcVba7KcHDEV6i7rQv8T9sntzb179rQDHWvBvlx/FMWugPykfQB8t6SCQtf
vn1Zv8431aO/Wp2IPjbz3q61vYcIRJTyiiQIgq2YGillQnLjZn0SlM9hHFYbJtGzDETyyVIdViCI
ZyKzVK6Ery/YO63rIP+HyfFn3J/uD1hDwCM0tAmUbP6dXyJijE2Yp/hYyGci+GXjrPfTbatt0D46
V0c1/CGncjNcp4RUVDcuAO9qyatyXb5sEd3uP3jX9lbgMhWaty4UWPBHy2IP/CdTT5c3b4YIs0CL
NQJXXhyTuJdbKMtoQNpL6RBGS2OIquc2+h7ST0IbZumPxZCCyfWpBgrY3o7jk8SEIjY79BzIoVzG
ZHNdLjTPJnWVHAj/6x5LoSBzoiB+sNQtFk83GEF1PhbtKPV11IVHok/aFLzbLw/qDPPI9bKoOATz
GbfVSeAOCT53AIxK3IqlfaFQO4o9Ky46DWTFQCSj5j2LH/H4PBoSz/kplU6KhiI/g0NsY8KZkK4J
fx5zI+WVIBd0779AnxAqQfghqiXQkAVjqhIpcfL4jvQ9Wjm1Fg75d+mwiBn8i48U2SzcoCnAVE11
EXa8yKh7Dut01PZKaZsw9EooU03nY+Qhl3tKdHPV8EgkL6XEuOIq+/iP209vknKjw7ZJF4AFntQ4
3p05CYVb1B4ZUEAzk+mbk/osp928X5FeLITdblZYrXVHULChm4PjZeGCO9GB840pfPcC8jmctvt8
hbpym/Xok8z0O1jalJt521dOSuF5th7lWT7eJAaA5t1oVBbsXy2vgYjvGc413YpyWivs4c7ha+K2
8Ec8PupVN8vMnVi6TDqJOlaQMJOk+drWZ1ZzEYLPDUblybT/8oYO/TYBhf4INLTxKwMXrzs7kxMe
pTUcPSi/tzBSIWHLywVJfdlXODIzS3D5oeO7xu1ZRZL0yGh+Z27aKOM7lq+AC05e759x5gFPBxgs
YbHz8NMQEksMPiUmjNd1QibpZ3HJBUIlrqfFHqi7HNywXtZ4mjBd0qce4zi8dsRsMySEGjyUVy99
oLDsJ05wPZSHbh2XImbFi+l2U/dmhs55Q8I+DKKnsMCDP61gELz7CNmGx9VNIy87b1oqL8yb7L5+
1jjv6D4PnFBh7zkPtT/YBoyhyO1yjqpXl83EW/3B3JCylVbYewjd5WEsfGM8y4fwfm40xX1Kvw4U
VX/pkFTGG9ZS5pThAvBGgnLYwdAw6MZn1RGhbuItiXpE0x4/4WjsCg15t1cml1xnIVWLk/k7jtgI
/05wbLiHH81ZV3nwk2Bl4njMl8ECSU3MDeHfYQJ249oQdBgSv8+m+COQDvwpkjChX1+FaktE/SXh
LvsEmWW/cPs/ohABKvE6zLjxebr2nieLi9EgYDY79U8aC6HOX99CqrYcFjK5kxNWj2j6TM0dFwgq
4fniBXymfVY/IYVjqFXX8XASukJ3kdjFkmTlk+1uAIv4jV+xP9Rryvg5oRtUiEx6jUgDyfRpl7Zj
baBQWqVSdWylIkXjeoo2ChDtxumr1vIT6IgqqSHmXlOrO1s0gJLdThut6U1cngBMOswdU+1SdYt7
qd9c0Hn8Zv6zaxnKoPp6cJ5ODSKn1NnSDeo6GUshsA0ka+7yC2T/JhyhPr0d8/k7LWaAXl2nAa7+
D0N2uEptT7+7vVnBRhCt2Sx5eqHrXI00zv3UwUd1AfxDWi2ovO8QE/4fDYefaZc8tOOUMVHv7wy+
pLfKGPVY2CeTcvneaeSVafwSr/jOgY04ailfV17u4h0LKlsepGAq9YVQ1UIPb7TZ5T4x/7B1VsZ+
DqwHGJWzt7n7i5N6xCbqmsZpnYSTt8UVEvFAqv/OsIF3+U3sfCTxwg2SSlYOXFm3NYWYx1dRhdHw
hIKCO24pK1wfXD2ecti2mD+4fwYTNEqiSmWHOq+B2Q6SilZcJPYliwoLZPKGuBzRS1OJt2QtOiX8
5+nqMmXhFBiAA/64KhXkXSaKLL7qGPtK60FZNtJl7EatwAiRV+9op243opyt9AR3kQ64kC3z2RZy
9bm21MPZbLWFyNbKenkkQHlyZmJrWqOr8HiCZhQz5je0dGb6/rR1oXNT4NlzAQXVfK52z0s9p3zQ
kYcosDKxMb7EZzrNam047IYeAm62TKrQ/1TrSVK8/eIWOXvKPTvPD6htwTV8cmKgH202rxxXrtHo
ZQ0Jls+G6NzDv0SPr2B9dMtAX/0BLz+UG3AFYQWYxALONIeV7diVdqASFN5HRFJsj/4ADv4Q//6G
hoJkdcxw2Nb1Hip1x9arV+PeQRmw7bHeVbOallgxlfHPBGrgYAVaxGKYtclHQX+lHK5YTTtCvDtQ
WDzlZS0nCSSRypLVKKeCBU6Bv31nXr1CG6vqO9r0YDQyxheUt9+xUy6r6PIfVojTUM7AYSjJAEzH
s4lAjAKRGIa4AZJfHM9zPWVLjkwoyG/GW7DBkC+5EJfFWz7SY/VLHfa0l06IIjil2EmdrsaIQtqr
tnmTOwjaYhUbbDU28yZu60FufNOFvD494Iur/HRraGotOjEoIM1S015ZsaLXT9k9T8x75UPllGWx
kpSlF7Qv/jrohvA4j0gFPcls13uLk8WfrU2iSwwGzWigYBujWSuJA16BWI5R8G8wE4bID9sl6RU3
fswMjEelyGD4e4OHHpF+zf6aEaECQo83baujHfM66tYzWf3dyAdcNQHWt252CqIPj62TjWyg3mCY
UgBXeiyr7BB32ZWFw3C1RecwCvfxMifQgDpUe8u65Oq+DR65yZE9xvwm0R1kscKpjyKOPav7cERo
EN/lPhKQCAPS4NlOe6l3i92KPNFVQo39HUhe1A3ZCYDLtDss0is7yyT5wHMXmuXfV+UoAhgFJcak
+pv1Teeo4bGSekzKy+PWrFQOSIZ1rW97y+ruIJlHK6Qv/SR/SrwfqJQSlq223IF7s77Xy4tMOBe5
XEI8JKNuPsQ5xP5Rb8W9mSpwaH2ilwHm2NfMwVZpPJVAm7y5zZu+EL+I/MkvXZ1yawrv2YHcooo/
QcD3IUePE5N8aIGJveHJxmOlzTMaAfI3aCillYJweS2m8JEiQJ5NCn0IKcrzrAj9as07n00ATBYZ
QFTVuF9PKSeTgjpJeBmf6f0o0LDK3VyOVym+4TIok6LOF40332Yz/2WmNqSwALswH56R/QXZOiRX
ibaRqRxNJyjopLBjqdO2P98CLDM6gvI3DoMA18oWNtw6UxWQXucFvJ9p13xlDbJ7rtzs5xibk+xW
D0BCPzlfTqjf/dV66razXVX02/y9g86sl8qxWc9PozxH3FpMizddq11w1DLD2ld1RTKDeuilecYa
Ug+xyrPCzVYrdXWhyQWZkXagRWAPIpTvXBkD4TaPuMPug8Tk6Yw3XvI1sj2Vy6KjMnpyGEdIPasF
mTB2eBM4Mj+nknnq7oF0ixcS9TKwS1+WC4jX8ckTFfNqxPL6dTmb537qGSpnUfK1FmVEgsdv0YVk
vbb0ME3kFICRIS6+1xkX8oSsuVMXSZsWwie45nCZHgTH9/UnfidBL6vHQVM7I98ANGgnaMQtO5ka
yXxjB8zXsFN13Hwe7b75teBKquxLkBUw42hUljsxmAxCQ/RFg4A1qwSvq3ZiSACzHx3xl/TH2Zeo
S3YFFBtutWJH9Sqp+6R9fG/7UblkypY7hcnGuSuNrf00Smw12Trf3X5ktf1k/jNxyrGe7eTNMKKs
aCX156ylf6ONA6bzllj7jc5M6hMAMCVjJKP/Ch18x4OsKQpxLMNHJxrlc+Z7uGJXX5pSQfzEL6va
v5FGbOEJf93sRG0OC4OjrcirMBicK6GB4NN22szgcUIzQeIfMWELnslSerHdpQi6o1mvojuUlXt3
bN7B12fPFDQLZO5tQsMVW1gYc3VVIiqYA+hLlNz79728K8U8uSnWSogeM8BjHKOETi/Guhzt/m7e
SWBnDqdThTXnftW9ci6yYDPTwK6Sh6HjrMdrtEeDsXPRXDqUnlu8tPc8SGCYjYQySEXo4SYA+rf0
CIO6NQBjy9XvCyo+8MF/rH0yOJzClXs2+PYEegP9bPg2G8rO84r4I2BAPVXlQ7YC7QVFHpDJTMWX
g4NmgfO/hna89naiuhi4++xdRAZpZU1Q5II76DJzZmDDAVxN3EPmHUkRHIu51V8UX59Mb6l4lDae
c6KtLYJuPQZMSNj+0yunfjtIhWJ4K4Hnc9sPBzD9AQ5OoHiPNtQk0NYsC3oK4NLt4rVX3QP+QxCf
bWl0BEPO773dQdnhzxXsRVvH48p3Y2EpDiDYNtj9Cigg8068zVilGYA6ylJlXXRiFjYutqNYAAY8
hRm+Tvd7+A/Jx7YzgMQ5ZxQXOQM+isThSgdVAui3AxTYAwy0VnQeLUOKscoDFObbcWskNMKAEsHh
tyBZw6dgvAt+p2KqRS5meXF4w87sXnVfmfw+tKtaWq9uCxm376SsLWUwq1k8NkGs/txHNWrWLy3E
f8uBq4FoBQd5DAqfJW9MiOxFzdItkLSqMfPSOvAxlEIGpYJ2fRlw7AmE6UwUHu5MBmIk3E+VyyAv
c/vrp2AIw2hZkjxRDA7L4hFYFzz6sjVHi6ZDpfL6maZo2Z6yXEQoSHzaUMp3wcLDJZOUveqau5m8
vFCSGjOlt9fToeIKebd6t6B4XbFdJRuq3oCHRWh890EAcmJv+Z4F1DMTQ6xjzEH7j61MTrUPfUIN
NOf7bzvQ8eqeDx87UrUXHWqGIr+tOfvOczyxWaDi3gNTpWGQtzWf1pbVuhQFnm/WPg1fZBEo3HO7
sMXt1rM+0R09WT7h/wyTrzGBcNRkZXneKZmY4iXxNTpmNoz3J4qtepowoswgSnGjQ+N75dNk+MLo
AYRS40jLs9cJuyPKa+9qUy5gRON/rZYF4Ga0I+Ak31PcgAMOGQvXuXlcsQwbnpILUSAAj2MpE0m2
T4oGwgU7xELEOJSadcOaI7iFjrIG4NaHShLlrdSYWfflPRCTYpnS89c5qD6k+0/qCSmWq/KlkQ6e
mNBI690Z3518hGCyLNyF00CDhoN5L6w1atoTELMJlXJai5xqTnEgzTgy+0S9glo+8VrJXX6Y36Ti
hH3PbTFjVjI4PuaoKj2enNJfZMrugk9IzslthZODD6w4p83Ffofo2Z3K2dSo6M6rf+h9cH0pAKwq
t/yN1m+qSO/VvnAp1IRWh0eZ9xvTXqiARHQJGU0YH+aNJlWwwoPnoS6zvv+mGQMK2zyW0aPO7blV
pSSeNd9VBlN+o7BOb7LhqpVuiz3fl47gT0K8J/72PS8bbXr5GvncOIuUAt2mxY7W/6zAxg6DJ6kn
1GHnQ7TdHyKF0X7BPuXxwl1lzct1zDRtED4TWAzWkzUBIKofXQn+Cd6fw/7eWEOssUP/vm9BMWJu
9RDkq2ulzweRGx71OnUMtZcRA9fBTMTC7Xy8rcfZjvPFR2J1pftQvSLQ5A5fDdkehdVDufDH7F1Z
k+b5+yKqZrF7HpcYViear0KoxOLDpr2sMb9edzmpq9OtRmcu8EIhZLPCGxN11lvfYlRE9NJ1SBxu
xzNmxjr/WZ90Gqyqj2qP93FBRx08mQ6D6z3kNJDly85by56BTVnY2r8xTz/JdB9OmFUSv2zsUN7/
BFBgSmYftSnC/3ktuKKM5fQUvxHIlghFj1+Lcrotj2vbmXtJOrMepuZBsknsXdaAZTa7iK9W9HkH
pIupMKZTqncGpS2GCn9wcuVZASrQd0k//6CqGVruPyt73qea4gm2AaBsNw1si2wUe54bqH7dXg2C
p2B9Bks7IL2i/uz50rUJEGURziNztxAEZpARDAanM4qryT36TqGxCAcoCV4ML3j1R3Qdd7rDAMtO
NV18jaQPD7J5+YWizmL3K9YThYfkWk7+lYweZB6h2lobQR/a+iw9mlQRi9kw/lD5lgZdFSrf39Fd
4G3B8/pqIQti37hpAFrDtt86U0xpOmSGGz5buDPAqPlitgsPCiqK7RtXEkwX0i55npacpBkE3mB/
Nrq2yuC9T/8X2IJVWFP3dmM9jGcpXR7UC0E8EMMWCrcMaoEd7pfFXOpzENjmu/9xsYzxABfM82zG
0Jrl+JXpAKCbiPnlHegDHRLBIGwkcX+lYUQUdCf/QOVqObrCTNUpTNCICa7G8NuNQ/TqyHqB7fBg
Z20HUxb/0jAH0QFyNJ7M79nwVAyZPl+VgiFwIfHA/TME6tu9rm17tsXk4pGe9XjtQGEofGRgAuAq
rHN673yojunuZjR4uwC7wruGlJgvTKDtBbMUPLFMTO27FtnxQldxWjb8pbVLQ//Ex0rEjwfZPPZ2
YvfAtYI5556xGWSfPV5iq0FHpJKHhx61NU8qanjyCm4/vhve+vQCC8okkTdqLj4nQmbmRgH4YzqN
9y3MgcvnsCTYaymFmCEVeU7Gha7bWphTYRYv8zxTZ+vL+fzvx2XSE/pJH7TX/zJlamDvJpkAFi2t
D/pUxTattE6rgyZF1HFdsgTJbGP6O4REw7tyXs3gAkhZAWbjuLCmaEaQrrPVBjdsnQNWBIXVIcnq
cIweQ6KioDRe1xXCyxDAqhVBsQfxpMFQ1T51zYGJRp7P5cdahDwIcTnLauUTUnkeg+xbYVjSF2Xl
Ic1yn5iqvI/sSlgu5z4EGCokp3QZuiz1qUcCTd7/0elsG1/l4HliSKa7R5s6YEa0GfurV+9zRMK3
Ikx0pXACj3xrDz2hZ2hgBej6oAMIujtQTfCeFTdz8nlOLrBk6aZKHNqq44naujU8r7tuR5MKdNNi
yFXsudb/ycRBIezNVhQhv2l4Pf/JHv5PY47xrZAIzc/6CHBif9wDLaiexyq/M+yQk1jeGAPc7rGJ
NgSdXrEdXtp9nm/LZpR0a3Fdmibns+9OWy1nqR2ihjl8E6CkzcVXJtmem9z3H3z4td8usbUwWLz0
a/pSMVkxZ/HHkWVrJKOMKAQtlRGgDqmImq/njYet3RHAgVxmZrvAlPypGlPObxZGqyFaPdAJzKS2
LkFj+5cpwdU1E4I0Bee/f3TsMbU1MJKg6mQGwO9qNRv7N7C2U/36yJws3pLVtK2y+xa5Tk2uXSGi
tj9ZzyPIIkJXoZfaRR2fE2l2RDXTmL2aOHTsViViyF7/wHLaoKgGLsjTXje+iADpWWbc9oNk+1Db
QZtR8ndP53kmcEEvbyjS/HM/7OiEOjk53p4eFYVZw5NmHo9J8YyeeXn5hmvchs60UB41KltK/70J
EdQH3LykapQjV/ifODFxuKPIF1HFjZXNDkRXBexg1BGIyYm0lGlFb4LdpKtY15rNwgwnD7oaby3r
Vufg6/dHDHlF52hn2Zb+z4EvSh4t12VbkbZCXIw3xVLFpbsIinAs9powcNvl0+h89WCcTJV8lYUX
yiumuwHq2EM+iu37GNSTLFLDNKQORN1IVJ5zyceRDFzubcu6D9Qd7x02q56FytVv4loH37dzpMAG
WAJiz7FqDiGAM29wSib0U0MAEB3hpZJagogVt0n14OUQTXESBEGA98N49gtNqK5bcD8TAOUWrJ32
eTGf1n827wpfrifThDFutaDC7fGWxyhCrvOCBvx2dVItveIXawYQeyHnnb13GyPIp/gUlDBFGaa4
BcOqhrVXMz4XQ+UR40MbZKejhqV6bRv9v5f60LARpV1Yb6mZ64YPmqLkh17XCjGt8CBWBmy1kV0/
btBSkS9hPshmN0AjI68FG8WSgy1P2qsnO+zPXDVZYtneygkWwqcbTw0ezdwaLWkQsb4BjVSoy9KV
IWbWL+HR9OtoPIaF00B7/VGadPPiToIAteQvbJ53ZI2sElKMM7T1F0okmOpnrPw1MJsFVSAlhzMc
PHy5KTQK0fkmGq6Nzof3OIB9xDzJZ80nVRbzqD/DGxfkxuMU+wwZ2jjhwsZt4C60oCWs7jzTtCJx
Wrjdjf81NBvY8JzjC7cENNhmxO54fCoNnDoXqyWGet4RDrRD492VFkfJ4RaMaudvDOoaAr9J/x5e
K6bQUvdyUkEDQBOOatNprWA4T7naQ3DozGeeL0d1U7xUfuN+HgH4MDE4JqFyYjoYDR+4d401330z
dnG78o2HSEv71AXcNGQW5CniN3JJrlYLJaO5R3LEWrUAfjKw7jJIDyCQWNJPEFSKdh+vmfHcalr7
MYxbIE3NlJyubzV4rTdBfqQLGHQjXYOdxDJo4O8L/2ZzSKSpUvAQDUTEHPQHHfF7AsPeK6uj0uCO
z/tn65cfCleYmG1OWm6Oz5sfF9EWtJ/7Tb2sT9e93qa9X5T7hvXuIutddF26v/SHUhNMq6A4/s+G
RKEYTziCuLo/mqcClZg3O368StYi+g9o7aWuolXwkDKtoSa/b+ZmNhYKUI/CKWkDZnzcCD5XMY6w
8zXg7E+1a7Pn4ArcK2t64mLbaZs2RgQSv+oJNsYkOTIjPaZCqXAcBBrBrECWmp+GmGNrv5gY1Wmc
pgMOhTNATxjOLrx4NO1LuLuH9t6WWSQuWJpsuSUYUDg5BbpC8QD2Ig5DuxDPPIGRrOWrEItMWOT9
v76heDdcE0Rw3gO1Da8JvOksysS+YF3obw1mMg2jWj38ebSjD5u1gyGu0dPntlEgfAOonI8zhoD8
RiF1rpV2cH3xVJ8f30nELg0snwA9NbZohMRQvh+0pygOnilwhZxQpv/WXtgCe1j+FpIs/UfZgAwl
Zwd6Db+UGCpKOKwKeGSnBHlF6e+yxd4dtsEKZ1pqQgA1lJ/u7OlNHO4E/pbI2biZGanehl8qyap8
aA1Whzmv/TdFwspjGz5XxPPA2YvhDUnnsqJQ3dmQOzSTlvbJrTgSNepDES4RRsIAaRTIPwmlDx1J
z11F79wHkSA7Ve9us4rSC6RhuLLHXTYcuKYw4gdTXKcMFYqPF71R3CfahRCCWXonpLp+kOEOpKxJ
UPEGniDCuIgAygQN8HPTQ0ArzKTVZH7uE82ncDt6vz3JCXyXgRyBdB48JbLc4fcHddVHRqaYTFO0
qZE1egpi3J6v5lmN7gqR12/wqH36BxhWk1Ijj432q+s464KaipJ059uiI8TTNFB2pXIrKH0a8pFi
kD0Ptn3u2LUxKhA5MVc2Py2cymMKx4JIo4duK57TqpGyhfKL7s4di1C7LwSWgpj1DS4ZqrIcBQx+
O+MhjEKs0qF7w18RYoCZsQRECbNrahrx5bgs+uvAiKIWmdWYQ7BjdX0CHZAeWGFel1YN9qNcBey9
KSINnFF+XFCiJZrhMNcK7CE8YkSIUsTtdNdqZ5xLy1a4cpFhpHr+IzOCNkAVgY5Yy/czqt9/0F5J
0WLf2Ovkud67cpBb4orIsZPXwsu81AooYnPxYtkwPUuhUZRBgmOxJo3nP6/94ErObwEWy34+cqH3
ilduct3mNGpX/7NkhG4ZJ/WN/hG0fHkTsCe9UNJgJXxQTS8GYPtVI16qk1YvgM/KmG65s6dj6Mb5
RYpFy5h+Y7K09X1kvHFpaJH5clE+0rkQfWUHqwHJL4iAW+I5ESRrib9ZKcIaZBVJycAm9xs1EdUz
s4T+VdxNbhAD96P0TuQc3eJT7S2NU6exSwA9z3xTxdw0PvI4MjBbjRSY2ZCEIpOjsIu8YJ2tHJJr
rLx9PWfSOyQ0Dx5Ii2XmdJI96rkkLcmI3zKqnwHuCNcN4jHXXsP6DohnkSZzjJigXA6k9Ff6V1Ta
N3fa6NW3EtJTJTy6NtKlrZccORS6VLxLhKqj6rCIIbpxvda2qXmKn7HfkQ5Ks3ySSl7J+mrfo52M
LnSV0/g+c3AavnZ5GTaq4TV3pZvsX0tGEfD6x116JaHv8dE4MeXVZ75fvjray5LeQocG7VsbnFKQ
JhHqK5RGWcM11azI8UDJgN4dTKD8O8CC+pN/1ny9gbShHu+sYKO3c90xx4h9YNYmQJBlvnCHkMKF
e9e3Ue1LbLmtqFUEBqYMo7pb45MEKqiGGXbObMkJvIF/h51UGgmZz8tl3LkgmKVYtroS4IKr7XlY
VgfGL0C1+u1j8DGV5wf4Ah13T1jfjVfijwcHp7NA8vFUYaTuSqzcWgOuxE0vUypwgMAwJKvXf4q1
phJJlYE5iRn8wPBTE2ZyaTe7oOnfE/Z+2GuiYLmTCeky4ID199t3yu1HoQlGl/4OgE90+bQw3Id+
E9nGnhgM20uiBwTmcgfJt2aS2NvEtDC0+yh7RrUef59PgMNRmyEwph9hfimzu07xsJP9isZJUKKW
WbNckqtPu62zqkdzdTmi9SrOxRMpN3WYskGiWjdpc0Gou67GJCsjosUJB1xGzAKflzqA0jfUo3z3
Id1I1eAHpzbwej6MMuvEzWENjf4iEuFwXMTRSIqbWEeh96V6srW04Z2LBmk2dtd5D6dMRCc0fkqK
nrnNTs0DUQ6x/H7fCvqz9YUZjiWUt7NPFv++zT2FIQQrzhhaE+/Qkwu9irsQxGHSIRVTZ3YYU0GP
PpHWmRpIu2sUloZw2FEWAFLoT73Pa7eZvf0n3c3P0UbBBFQyQyirCUBX4eEn6nZOS/d6a5wOnUUd
YSPRTnrAnvTzQfQ5tc5V1HsyPOHwqKXKBcvHr48aNt/yV1kbhG1pzdI27m0o0Lxf8b3LMoiTGy1v
yWv+rKJak9Eq3LtrL+kgTGZo8Z8rYGP7S/rIes19vIiYSqlQshU1Mb8i5M5JAkYGj3IYUnD0dzcO
cym8yccjo++PBbIjXs5vGYhJRt/pmpk1f3coVmOGI9SRlH6qIkHXqcC+6eb8v+wMvq9ABpyl9lGW
CjhTgGtqPBuQzkMoMRFzV6TK989mvggrQWD86/xTO1ClfJwto86JBZEFVguIaovT6JW+R5b5AGwv
0wzSe+9daTQctsNAmA0B+ibRThRZtQ9Z7Vne//QRo6UvdDOpsmvGME7la9pO+cRaPZBCzS6igDB2
U3wdFwOVNQg3ksfdp59pe53TxVLp648LzRmnwnoWFydZiZgfcTYxQoYO0z+o5W1FV/ALnJTvIk87
INcY5tHUjOuTwGnytJelE72rzOJHF6ahptXn/s4YltBEYcoWheOIHV7bR/bqhau/Ov84RqDzlBh6
7U4kYRKlQlhu24I5LjiB+x9yH8t0kPBStgLa8pr6lTeGVen9B/B4Gqh1bZcnC6Fxk3eco0S1kfYG
oQhjUFraPPYdFmYudJM2tA+dQy/tALRzxFBgj3J/g62IUpO0QHRv6oc4/P9hjqEbP1/OB0T0uApK
QHtWn/g6E+UlD8TUBA/BJ8EVv6KX9gcOZplukcocdXf7XYU+jflYxMeBBLiYD7en3awPJbJK+WvJ
QYofMFbmth7wQQgOXM+vRA+WrKPaTXNkibHoLTDrsiVtwLOYUCNUbGo+5TIzuuJdP6sotOsu+ZWL
kzrlr8jnOt2ivqavx8ok8+pMu5fHZ0QrS6xJgke9JVscE3BhlXmi+fNw5jx2iRdPL6xzJ6tv+f2Y
m54Fl4OgZAheKZZYkkWTM93iYxViTker4kX6wEmLqo3VPMw5CvOVSxJZiaWbzwrEz+89D2vv1zTV
7fXhdP3lnyn/8l8qkoo/oePV0pb2GyCRl/QxcAwR1Ucze8dudDa0P1S+We1pd1V/VqwEUQWZpegI
7Zy3P8Ky26iLGO+bBfYKhbN7PN8DrZzJC7TAihcc/5Sc2htfX6XzJqERaQNm1jQqj5ddnCJ+U9gw
MUpHMa0nVtmTdQAOoqzefUeyQvbdX2XU+zPT9brIBI4ictMMXHmVsCknselrFDQ/99i3aeLcLdvE
6v/LknVi/Yuk1/TIEnU4YDiY3sks/g+oTIwTRBP8CZ3jCzz7nGdCjDMsUDR+2G16HeOkV81nMwwd
sxPS12ld7v8FLzQkrNOtvr30swam6vdVnSrwRuLdJ1derKUTVoYAw7lXtt8LXpYZY+9LtICnNzS5
47Sj/os8nfd2gBosWllH/1dqyueR3S0o7BX78W5ap5jliNGOe9A4aTzH3TXJ2tnj5gfwK+PcowTb
fhz5i1J60t9cuGj2mouJ1ZhbrFaIrd1Uaul0ZOvx2dh7pFqlC6QJ2+d0CriQYAdYlYNOszhO0J5/
zSWIjms9l9Il91n3a8m8UEDDmgyPaaI29NEOJHvx6kvEFeV8P7nKXVjfBCEY99vWWVGGbe6X9Wnj
HZp4dIxFm8meNiDQVpm6Jw659PGx9xWyZ4DCsIET06UY/RYUFubHOL7BxB5aKexkturtJlLWiOC6
gmfIoJZaKW95VH1jLGIfli3f+hZi7ZeQQd909dTeG8z7fvord/RVMItJeTqupzpYcrgl2KM2Yyey
72Y5iOQK4gf0lLxyNqy6AdhaA8f3jSuQ1rOL6YKU3QcdnAuvTKG6HqOsnIZaB3eA3+cX5c910Ho1
g8A7WrYbnrfFcbOpAjzcPiyDFgsBS2Zq4o0/b3DDUgCT4lMABOxWt0fYhc4p1vbIZn/k33oeMzLg
5b0tOFUWqeyhOFn3zVZmWMH1/Cr0P83TjA0VOYi7KT3GzkrlU7NoZoTSyUXVusTZW3hBD5Sxa7St
rSRdeRvnOXo+ToQwSYgAZ3tBB2xrcpenzw1K8yvOo/coh8dLxcb2nw9SYEbQbc3wDPF2E5S+Y1Mc
0c+8Y9Fzr2NLmRsp3ALWPhm3j3tYaff5TBXeCUDsZjhPQ03LpWSGxoOnZ7Xe7od9xE6AbkKCMZH2
qB4twNi5U2vfZlvIHr1HaA5LKAb8v0NVFFac77+MUaVpRhngx19Fd6FMlVWsf23vQXmQ+AR1eczb
0Y8kFupR4VjZhitgyQE6oxy32mxltSBgTFFl17c5Zo0FKmPUqDm5Wt2v5LyXC3cIb1idsKp0yxHS
XOL9ChsOPazA5GvxpToPQF2ezJV+xhNF8Bp6LTWA49iWGmPdq2QfWTJ7M0tSR7P1g8iw1FL6THY3
bJb0vt5wsV6LElsW8IPDNjkNZ/VWPHg2QKnQ31faJ465R2TAO2yMwvzLhAD2a/mjBOncmAhy2S6O
cThXiOhxHAQKIPPoZXwz1GDSxPh935ipPwUBrzR2/WM9caI7Juy1ojB+j88FHxx9YIhVPLtws2oq
MkLnRz+0Y7c4SRydtOPVXeqZt0wmYRtm4zY2VdhWiLJyx5AUFLglmjPCc1JGx9ugiOGS3Naogkqd
nQqPwFXzSEUY9vXeBgTN12WAG6nEVVgs04M7l6caE6VsZ7eSQgNnSfz+uMSEsJMdao+xfsgQ8rMi
rClCOrJpBMsqOsatKJdYWIWvhBKj7z0EVfh0V2i0pJPoXEByC+MHoWM6m5j0nZpkUfSKQ7JCxzuS
KB8q6Iuntamp27JrAjCf7qROhMuuhnyUbCXFRPVygbZTUdFoKbZMz4Gly0UoffQXif+6ChzPCckx
LjXBK33Fyhb87S6saFBQAgdgTjrNoUBoXBdEA2+e73UK1QRofvmV/4NXv99PCfHUv6xirs4IGnYX
Ec/oiSTp5dQ7l6QPnNUteS2bcmqrhbZz3I9Q1WuAQAUBRiPRSwBOEsb6k/CnLKpOvIN12bJpPiqr
Tj+jKwDMTWlQ0tZA8Ow3qY+EmbSe5x/hVSRbStA892nHDAEpFG57RDOrVkZP1qaLtj60MqPL9sq3
Ub8rYPbB0I/5EmOGeOJ+7XOIVBCbRvyMRcne90HcZnRGd/20rN0iKt0/8lkAeZ06ZmevXHrT1NZV
4rozADpx5NO3jaHa4gtdHneDuEywATsyEF9imqDyrO9nNeZn6Z1fM4womWYMk9dPrbAWV3omntkT
aV0Vd9i5iFYgccZqFKAOlA+SvrnU62USZZpW5MoyJed3D4PfMFPVVGU/jEujWrOiAsjgiy+Nxqg5
YUlOQnt0wEq4Ny2PMzXs7guRUGeXvF8ay6D+XISz9cd+huUfnzAsV4138U+hvv45Bgoj5zP8kk6B
Y/l4dEA76dRYrpZjMTc7aPRFduOG4ghcI4zxsK/vd/yP1v/KkmGbukS+Px50c4dcF1+V/YkEPGcz
f622vLxCFhwGsdQb5lc9ObNxF+WFqNxW/Gswlp+2wH/CMDuNWXrePelqvvMcDlq6iGwZpYqIgX2N
WPZ3u2f5jT9WZOZzAHxhw4gAyQyj9iF76PdI7zfi0jayE4LyH0ZD5QH0b+jA7e1w/fdW7f9ZWqz1
f8JTEJJ/ZV9ZzRDp2AVnwqWJIlsvfZr33Xs5ZV8Tt8cdFDFLY6xQqBoKK6PF0ScYXsP0ccocIcW5
jWUCNobPFHV5MHIPkUS2p8whn8CrOTNdeoi4M3NffphSNsOF8nU7zNIRcY8NebkUdwa9g1H5iRIw
MqWlrvIY8aonRQFlwfYzSK6aUj8swWvDo2zYLR3MOETFLip1N9/C+KXFZxcu99OYagVGgJHdFoOI
/wyE8zawi0ZgN9IklsaSf1egAidTO0XFF5sLDirNYArGRtMowjWWWiKI/OxzbqUz+hN3iJn9+sCk
/RIXcJXaeGOtK3upCh7fCzkWdiqvBqLDCK/JAPgOn/9YEpjLusef4O4z4la+nd3VpZPNbWwnD4wN
1D2QPG87yi7BN292LfyBzjAeY0gbxGG4BBrdb86SgUQQlSXxUXVFojbnbC2Jh2/1CDTJzas3yxMz
4BSPQqDeAfV7IOUyroiGmysMUwpziyg9aRdWJSyqGi8nN7DR8fXzDAlOaRfryr21wRjLOCnssJLT
7oP45rUCELLYMmFeGtqPR+ImWgbP8WtM+b1sk/xcp2IX7+EEY6H541J9ckttMmL4fuelFpFABW0M
Cu64HSzPPMHNuT4L/8QVCX0st86HvyNOgCP1qjCoFFkSlpOWu963G0RJsJkih1Kd7nrzVMriP6G4
j1wpTNR6rCovSopINJnU+M2eZcUXen95ATC1rWjV63wH+lDEN0AXJ5rXvQpcCFvSrEOb6Dn362K6
++HcIKLeMkZHW3xV/VAf12GinoLm9QTV0WqgXxsvuy3H9EkbVoiv+wUes9DkKMkUrf04pcly06cK
6+k72St2qmZj6BGuIatKnhb8HGWA1axOMYy0J+b/e0j3WBrEHrHKxS5Wv0FFehKeGj/6vTL6gqtB
fRayLEr900pZXMe3gopuQ6nZ3PrP4NFBBxs+N/aUmxqDZJVY/tbG8foFLmp4I3dnZ/vVKiRHTvBO
TAI0rtyZwm3t6jIqRsIcTzV56DX7vOyFSVjftlORCOtx8g8hboc9ynWymZuCXmg6QQz9xpeGrQrc
4CbL8co7bzfuhxg/YIjr8De7Ts/i/58oOzhKqzfCUOKauMLKv18v5TzERSBRuAAnQGkHh8RproB9
7ssCfgsTeShpN/7cext1FsOiD9sXqeqlXy/Nd6+TsZo2j5EQetRmg0Sa/STQLtNti123rhmysbUa
V97AY18vcqTWtphjNEMw0MsthAE/nIxyYylvB1lntk9sVyu61BvoHtRquHB3SVq/7a8KIzKC32NV
WE/+BvvrE+I9og+ye4lhh0efiGbXjcrWlw5UMN1pRLQgRTkTj++TMXzI8yl1Ypnwz2MAcgwt4tZm
l0ithBEutSK436Wv1EopHMd7/PB2M4hcJDcsHacOqo3CboldQgD7gSfNxdafnjyUHdrLf5Q8bLQ5
7Zh73Y1p+PJvKwK4SW84/6WcVZF4PMsQf4dGKJsJ7Mhf5rw0k6GP9Qx8GyfjbIQc/Oo2S3ILVxEH
YaLpPFn4frJDAvTxhfnZlPeDDvE22lnbhlbV3iP6sJx6pV9D1Kzph6OMLdq7VzrXy6vS/G7JLigI
326mOWIfnvbx+pZzWUDYvgrWethxy01m3nxZ7Aqcjg4c6YgL4oiG3KlKFnz3LGrOqVhWP2q8woXe
5X6ZDU7DJtof9NfHqlVTOBAxwENwCWZy2wBnvLIsILKCbcZhKezr9HI+H36FUJznf4ZvhrU2fwXe
kgxfeC9IvjcUPVI/O09wtPlFJ6icAjgUSWGTj1tl5AEze3F2lzFkYr9lo6TVB7k6ai4MdFJxG9F8
sVEL1b9VOdlVGU0y3arftVrJhYT4wJIb4n6U/dPbnhzPCeAzuqcDokYt1vbdN0qr8bA7bfz7r9XC
eEWQio3aua61Y0FmyFH1RNhbX2G1akoiJQudyWPB5dJT+dlxzX1Zj7stM70tWKgSO4/EDcqZ+/LQ
cW9UDLtvkz5ZF/zUBr43rQ41o5rGZrwPhrvMVIoRvxjXnrGxD1s1WiExSVP/ITCunRS3TLcLlA2u
nRk1Tv3BEbcpnkTYuoYbzLWK/Z4h6c5jRpRu6TuD2xAJSKHA8FSwL+CH6GIOS4khpsuRr+/gmSAk
SkmtKaCmuTqgTQAHe0S8e7sBlmmyyc6mP9YJFH8jF33twc8u/8jmP7NZQ+Vh0VukVOBeSsbq2GG6
rEDwoIiRVErGhjK+kQbHkSnGEt0MIMxDykwbwHtJmnekLzdIjHxqQkYk8F9WMGcg6hfMfBSRjDT7
1QkSE5g9xgbxiiUbThLTSkQTAxd31qpa5ZflmBKMWASehvUiqnM66vEuvNAcZrDLDk/OFW10ceU5
RHiqcsFjvrm+HmZACbXd5vhEgUhKnELGJTE5eJ7kmGHvWyrlq9AyJ2S5BbfnMjGSbCsiGmUJeYdM
LTzy3oUdmOLhW4XmLY4eGHdoAklYs371yNk+4glZV0fyMHPIshQyOlvovPYiYwYNeuyqp3Eq2Dn2
fMUoXvS+XKF+BziMg5QNzLy4S/zO2NeNXp3mOmCMh4r7fvomhOdEjO6fY8R5dfQfXK5nlo1ZURn7
Yx/R5wctSoZpKoV5ND562vtefo9Tq2D9c9CFPEPXqM7AXrexoBA45zA45fNzoGJrsGP6g2koZwlg
dyVEbRbnKG7Q/2tiJb0Rul5IRiOTgLMm6CX1JtJPwipcj+meKsp+dvWy5PxGnPo/dYG1X1CfVHSn
cLIIlqQQL7RfC2cRBiz775+xkUG1g/oIogYX39+6A5poJzSa0ZTCb3iAXFlqJkK7J34a1RkVp0Xf
ZTlmHYB3ALW5gMzzRF4NYTGfsY0SCTPRavjnkvdOqTiHT/S5HUUdPGm26NBBipoUGTESzH4sxhNq
n2G615dgrQwxf/Zu7fVyqep2ZYwsnfOf1YcQJQhiTtbHsIt52omvNYMRQo5JRU/5Cu6H0FveVfUf
p2Lln3yTSrlzMowDPTZEdtzVoyuWRPpFe8boOU3Tz/nWDEgXCkZinOMrq5q3pWjvaYTonPqyx4Ib
AB2ffxrut13ddsUJRI7kJ68JcgBvhjCjmGH1Y95gkKl4Xmgi1KMiQj6DqRdU34C8a4EcUDzEoDoA
wAFNPfDie6Ar8WPRoqSz7H9GHkyq6AgLcHttuH/7xcIKi3iwdcut0BgD76HrXy/bvSE4vzza/Wog
C9woBboNEA8+M0nHz+ae5FsxzvDMIJdcUAg2yQoI275h2HglQ9pWgNJJLuqkGrukH9IfJ6iAYZRX
vytSC438iYiuXOBLjK1OxlXIrUSaAljTnSzMx86EtLuTifw+Qw/BmeQjqhBzSmRSp9ruNkwcAXjk
HlFfxdvc1QoTbn4b2VUtchO9WyMnodrXHPgpZwjDGzIZds7/b6phcksLh6o4WMC1QcgF9pL2pN8K
cXkEIQslumEHpfvp7Uo6TQLP6mPuyNgo3LIT7O1YMjIYshwAb174JJfmJHS+OE/fYGKB/jmA1d8Z
RFk3eAYcLoVhU+2SpkWlusoP8CQNQ5UKzU1ATJarV2OnfcDUX1EpQW3MNxJ115mAfHIlK463VeZm
jslwDg9gWaEtn3iBwlL3Kpb+y4M5N+luM3LAiyhOMQNti+be9TghdfwcQGhbxG0ccWMn016lTtwu
rKSGPsF++MDjk4PpLHyteOmuKigqEDsVf3Akc38VbqNjMGMijp2qDVRgoIr7S6+Hrdwko3VR5Jlc
Jpk/KoR8MZPEsB+0Iw98CiIQLfmBTgZJ9DmojA6Y6pQ/DKa4ROUcVRYoOR0cnv7EPZBY0o/zUj1U
Gcz6OhHwCAHKUZu640d4gqBiUQhBZ6Tn/zkwjkwZDwdArQiGo4l8dwgl7Ik+i50WWEBWL8L4uMOu
UiK1infvraCw85Mg+zf8+LquAIpkcM+xIq8odrTE9yDTF1kqUfeJKUnUSHhV+WfBApTIzvufhNeW
yGv1ub4KlSXe7fbMjvDwyTQ4PwzM5QNbAV0SEjiYzPpjqQaDjFfvCQocwxVsO1o/RP7yt2YEbn+x
PIdah0zYWy52S4hZZaKsfUf8D9iZvB7zVez/StuoxAYwBuab40sACnKlFfaqRQIk1QXCSi9SkDIK
25nsvevGjtT19ym+63puullh3RgGzTuUA3htjAt4kdk2HA4mQagt4+MOLSkyIROg2RM8xCq6sDJh
FdbrAO53fRBSp8TMs8DJVo0oSbjifmir8FGF7iJnTPH6DfCSO/EYZApca8XJSqJQFulrdg36qF1c
ebvLygc5phImlU5XN+xes6yryU2H/s92wPbTnL+VBYR6sQ/FIvVAlit9uDWjVnqb+UUOVm7vRrxx
TJA71P2I+3jPArK9aNt1sreyHU9gZyvzBm9lAkQ6eUv5eS/gWKS6HhW7YHAHdImYA50kuSh4nkhH
ZGmvqgrzOaUvF9Y/aYdKuhcbf7sOK2uA2k1PPMs42ce3rcDjYiPBpPYhU5cmRtJhdUbtNdwwz1jl
3d3Y0za7FwHmASQAbI0TUiHpcgTcDpu9xTVNiluN6C+fhYas+roi00ZIvi3MPOrw0PG8YydsepsK
VG9Ti/8JW+PJiHGS6IJdd1oYiYJPb0nN9WdbHqPkRdU/zz2EPlROVhXMxf4+ygfVoezTB3B4VrDG
2py65vinGMA/pb2QyOQr38EwY+OtLLosL+3BLQD3sCLjm1FMHxIG8qZibtzwh7j2aGwJuxZXCEu9
IIMyl9kx8XTnqrBrSIQptivzOBC9HcJkKiJXz3cG71hLQFm++UadzIHSPyT+y9sJY1nwcVqcY/2B
CAM5XjrI+QaPOHQs2XIWHeYTC5NcX7/IbP3parIHchHwxJHciSTs4bkTTBC4w7YPSqxzeI7A/vwj
b0q3SCbas2cIIBvSHtOXcPN6itgicInuVZDeLhe50CzTfjinQkTwGrODk4JbbjYK2UBWRuqMIjQe
xlhsV9L7xcNQEgnTOZwwk0Tss5KypHZO+//AFxOrUKo6pFOy7hyMRlgHc+HwGvdY2f1Qx+hw9l9I
mBoa9fM+DfxNydNjegEQmEPuoGZLxpCLeQuORzTHLWTFRnwOz/s3LkV2z+ave5d1ljOVw7x0eQ+e
ceiy2Ic0ILpgGrbZnumI6iB+B9KafjI0D4iPxp3v8QhEWFnVVj1RxW2lzF9JWfAOOm+KQN8qgSJs
pE2WAdh7RsCf1LnFP/52S7yIgw4PAPMwpXS0rivkb59arh9kvGUXZ4fKwSf8wm3p7wbFq1jyiBay
KghazLFR+gJxoFDE2fxWeGtzrgO18NJ8XOf91niI6HsuhOv3p9asjQ61OzFD0wQ3EDDGo9SNhD1N
9XlQsvz8F6wRgkIsrCsvxxACa3haztlUGA3PNDDTcX8dykkzk7ldCb7U2SCneCtDssNZA30Mw5jV
Q22TqdEB8cg5uyTmyQgAz2WPFXMkZStLT61VXQRJh5OUGaXO3p38eJfxHAckCqoPlRTbF6uk+Du9
EGwXQegYa2qH0Q5I9YYCYHtl+EtQBDwsrz8yc2NukKkawcTPYFh3Ih4N3XF2AOMgYW5WcDYR8DhA
NNlY9pIfQ6r5X3D+9Q3DhoYmf2WgGljYa30Yk21xJ82cbwqllooVmFJwf7lbye9zZBfUj1jZbdRY
DcrGq/aFgjml3opFYtCOeQVa2kaTrGBfrcXgGrTk/D9l0vS9NSxH3SpEy/sjmW4tDxvhxcGSgqtY
8qrlo6fyATSC0ptdJBmHNHSQZS3dfe9vSQQhXEl6T8+4t1GrAoqHNCcpgbVDX6DPyKxDiO43IBX6
I9F4ttE++/fN5qUr1BClXQCDns4805IJxM/DQWkOkxbrnrg3+U7DQB/+ZkZLh90ocXhX5y8y6VRz
8lkZAAd+kMolEY/R+MX+4oi4lSeLdGQIQgbGbv4HsgWLt/oIBYCeHYinD6yDVWlluQKMT+MjhX/e
EyF59YmN2Mya4N8vUisKJJDntzJevgbfPdJydnal7NZECr8uQp5lNYeOPZ88eKue1NxhpGdLIGB5
kN1GWsGfmEMguJ6A0FMj1Hk6wKRcXFMqmOuv3nD2pXasFU2ayRtwOPFVzshK4pe+/U/9PaNek2X4
vGdf8P+XWCWJeGnVZSixUuxGjmteAHY1/v28NuDJq8xb/MJBml/jyNlAwgktRRi23m7i6OiPowGo
lvLSjnL/ckddDoJm6fH8bVicO4E1esAsBBaK/5WgfDOB6/vXntNoA0OGwYEIh7M7DQByChR7fh/y
0Drj7k42inB4ZgD6uLREqf5xJchW1oseq8lbKU/jTkXAqap4NID7XVTIxrqFu61RFxPoVBMUwV6X
XSZLNFE5pTSwCs4AD6fP2bjwiegrPClmCalm6rOneuKLZSXUR/wJr+1OZsNqgihN2zIJo4b6FFER
+JWNFwVobH5+oWvufnAi4zOkNFxtGWqDnHVpPXwrP+Y23i9Dxlw1+vpHKhTfwtenBKt9EbE843fI
Ya2l7Q59RbYw7WVTdD+ThmJk3HjUUDNJXNo6bNMg298IgAtKQQF61qgMDPYHF0qrOeX3eu9+6Tmn
WdSQugq8QYnhma2dB+bBBiCrAtBTapE6I+EcSCgQ3VnRR94kmwk7byfekVp6dPp/nVQPIfhvFnDl
xXz9wE/D6fS5xelMZB3WPp4I9c1Fi7sP5hggjGE89FBTiMm3aQC87j6nrpIm7OwwRJNQHrRp05BX
UtKQ36cTaRj3l2uGCTLgSYBr6jKMJ8jTnsfxMzpSwsIotz1p0gucYNybuDc05bq5GoerS+DSGu0H
rRr48iYqHIF7DTIQkDV77Lm3r8VpO7IchUafnciQmSwdSKRcZEnZf63PXW388R2XveYj5K2qUICJ
zlLIQKtzuVAdcxMUyQHDxtlBbuJbdof+LGAqcBJkdudR+UYcJ/dWFabe8hXQK9agBrJuVJNu4wsM
wgUCs+ova6/Abcjo+hot8AUEER5/tM+GRbAdcOLlkyJQo+8mK2pzPQT85zAoSg8Y+zAK0PTLtugR
0wvB+qfJ2aAYvLMuiM1/fju5mnnyG9/8ylt1xuQnRzVX/yXgHEKFKRQ9foG/oeaDhD5qwYg0OiNJ
XpHkiYbTluWg0/6++m92/N0WjDeab7axYfQU2rh0hNPShQC7lIDLoGSTQw7LgfYXtSkiLnzXYVyF
pv1nEKkyQOKDQFtJXqoyHlc3ew/aSIzMtYekb0zRhC8CQqIbQm4rY+Wdu0OffE02Qd1Gq3YEDiCJ
02bNJ7M/yDn6y5R8LEhe3gS3eA5BLzdL4pke6F92mNhFE7fyFlRDbGdkvdlAqJjH1uar5sgh2Eqj
s6FB5BhVuZq1UL6CGM1JtGLeDuH83CNQrUo1o9qLq4G0MEFk7wmEi/gbP2P/zl+KJS8X8wTQSBQM
yPdSNdyX50C8vZiTHLUJAj1L5C6EOfXTaz/plz2DYmhHO3K3lHJ7huufm4NmTVd576rnU86c3W0A
TqVBsr2GEw30TbdMEFmUoYKErfWn5TPEmbHNKF5xJrDTpBLd4nQmbC7aC2qwYCkOUtjdo4aqXHNG
3vwyWDhED5oh9sGo2jYClpRcRevvuTBiEbYasBLg4yhtCgXgelcNYCSWNF5G7dBvHxsQmy9S6ZQT
p3UptkyxhoHYndvfQRrvf6Q4+BYyLaMAMHhWbSl+tZqUo3w4xV7RYVmMD604NlsgYtUaEFSeltyE
1lYCT5iGYkcBvuMcqrm+/a4ToWa6GMrQAkhPwXwe2aotnZqfd5UvvT2CHeU2BUa27HU473B4NTFi
kvqemgmPynqzB1H9ZyecpzUutAv6ocyITGEnJWIIlD2deQk1fH/ZYRqghpIkbMOBVmuB3mbicXgH
t+CPCy7fa+F4M8MKO9C4Cm6nFcJZAOY3IDP07ra2qP06ANh1TMHpzmnIynhyReoXqIP6dZjjWSsp
YJ1czlHshIzIRdDLOEgNCcTtXAB3HGSigTzJL6B/FZxRDxTqhOIAC7jin/dXzE33H1ojePJMB0bt
LQJPOGP02RRPsKvt9kGlO0GSfvtCY7YydjCemxyx96yEesmAPrAEgm6IAgoGVPOMRY3dmAABag43
695v157Zfvopv4bp+W5tX62htxTeKdrERN8HUZLhz0Zc5jzyDAJEi9TJ2knXoO0+QZWa2jkrp7ib
QnOivvcFIbj2rFBtN8DTdbwkjiUzo9D2KBb4M4ADH7ixwAGtg/n5J6eTJObWuzKMxebZjDxDNTah
aZ4QiX4IweMJQwKicVmI3CzxiGcKRev594sa07Oq5ySKTWxObZab3X6LWaCB4ae6RIkBrdQmKOmr
riHMGmD7BP38NxxtiW84eIXswwhGiZiWl91gokNrdtZlsOpCM5wNKM/elwBC14YisYsAeG+NoSkh
vw4ZNZQbH0MIetHgsCCNURK51vbAJPHCfMeA+JOsFXwFfOEPJSe5FG2KG8N3Ci1FleFTECqNP2Sc
ACXzQ32qqBW4rqu3ulAGDoyQ0MdfRntyVudkqsiXrJohASiPHedgJQLGMWn4eCaUiuZ1KNOBnTDf
ihD9KMokHMhbCA6csL1JqE8G1wkixDcKCAZxiq9NUKVuUoWPFZ7HlaeO6Grn/+TcxaF5MbD18bCp
Y8nqFdc+AHEPti63T8ju+XK3+SIwvl3bj7U+b1jCF+HfDGEGmHnewDtYRjJK9onbLlJWApBzfSwT
ohQdHBbMeqyxXC7Ia6iHmLTzjupr3ZTp9pKPVlUgiYXPMiwtFPgBdMwjRUjyBh6Slvk2/NyC0zfL
nHkrEe9jCfLB4wJTJwB9y3txjcLjlIPDmOS79BI26EA+QptyvYnRwJqhCPB8TBlRqa33ofi4uq64
FdPPC9ny2gpZmaSpsRdDJFLGqqCaQDI+Dp15KzLB2nOArhMYLe0ULHsAf806aTZZ4MukXvmwTaMS
yPATP178MIZZTTt3nQUyaFQ9TcRCJDiO5O7p3ARUwLVr6jduRqm9KPCGStJkEke/Q7kAoDiDq8YQ
gl2NyysVmbtoS08aTJs6eiEfweVM2WTAVZO8GGuOfEzjN9d0l3KwvJvApI+NucI3VOv+6BoUIyEH
lFn4TvEO/vXGqnSPHj+cLrY/OlgjJn67ijqbrIg+lnO/vqgLhrCC99z54Dzxpnn3YaCZ+VqCN9Z0
8ri252/DKf4kz9Z666sUdB/ZDCkpqAm0fD0wHTKu0mf4xhWoi0/OiWOUDmRzvU5c9xpe33C3qfAB
mR+7OhfN/q/hHUwH5ZD+hr3EmbHZi1duLFKFMrO6k+YLINSFysfCcZqjVjzLXz4mfPaNkh0aMYjv
1j4I6KneFkx+FgutJESqHlup5CI9Ccyn2K2WJbB1coIDUzIWV+ykpRjyVZUC5+V7wnvh5LbUKF7P
0lnvfsfDTjjCMBG8xj+qyWZ9Te2MdinLUV3suHgwY2inBIOgNxSFJXj38GOrmCZxONVQz4veFdM9
U4LMkLCE1ztRv7Jvn9c6Lr7JtnynicpDvs/1F97wixbvB+YIFXjl9m6xc+Bvy+Eeq5Pp56qdyQbU
85gmohAE7VeQ0gUZuOxAgBJqOAg80qh1JmkM1R5Tp3Q+KinKY/m03/OVVgCMq9EI4BNRM9Y0fL66
ZW9n01OqYH9x6S5wFKorOdBziuOeVFunfeqeVZ/eZbKWe3qVWKFfQn72KVMDamvkz0E/IR3aPu0+
INw04k03/eiXcx1+9X49ymWN2BhJlHAEXly9Z7M6XwU0jy86qrs85AQweXnAD6BgbyawJzvbIm25
oQpNRHDNMCO9shrln+4G2W6R2PaECKpK3RWlzQn5MxF7tebh9epjouLxViajnvd1QZNtRlHU4zcL
wpjJh4SjhO0wXWNlSfZf/eilH+zavuipDaz7utOSKxPvRwEzk3mzXhYSW/WIYHmSXe00+Nfftgi6
gpHsUEnMKJtlAYf7CSZu5IMs8pTrHGwGaPHcLBvXZbyPVfHnD9vtpfrXBjj4Kx6j/j0iNcv/PlLw
waNeCBdHuSoQubMj2UKDqv7q+SqamP74djWNNwy4K/xiekIDj25loMkoqW00EJnTlVT5g+C9HU1e
ZxS6VHQSnQn4og7jQcB96APOcQbMd0hVI0gpxS/PZ3wYDYZZznXQukYlfb90VrWrXXOVO3A8F2AS
2i8IlVw8rRxRz3yKkB1XF5XJ2JrRn46y3nW8KG6TUF7x3xhMEePNDaZDgSnx7yDkQfJJckqFoH8b
/PEBFDMSiCQ8t5YiaHO2HIoWfZkCvzJRuyPDM5juLWITtgdHhEC2+AwvIA36/KKNvjHIVrVxwFzw
vlPvJ3Q3UtphSjzmWtcreJgSkdKBX1rjHzJ/qbiI6LgW2bu39LrFgoUaejWn5182bYF84jUG8jl0
VajqZE0nV4jSaEnllduk6dbQz7NfC9W2FhEdceQptli59FHvCCZ+Y+VZ0cjiK8UJ+//Blv2qyh3p
T32nOzv8IgQUs4ptu8h9mT0CbhsA6WrU7OkGsPAqD+ygnc1GHU7wI/gxA9JraE9ZERx/mRlCZ3/g
+XUTU2jlWYeRl9hE0ioSE8AuLIgXO6fjNMsNyS2gocKZwoJ1iaw95oaxtWenWxyDu7yfwQ6OY0Oq
K6EAV7Ki5H6O+gqZGuIf3G4RaNlfbeqRLXBKgDt9hxUocfre0u7dQJ9Y9ZsSgvF2nnpwxpN42vCy
A/zHQIfVj2SuQWs54Wkb/orwNcucLTNV+gbQEg3Ol3WKd+EiTg0JFRH+sxLjookHjw39ZAjKxNtw
z3khElEGonmXeWGDzSlPH0brkHAGRwkVWlFVXk8XoMNK+VJaT/UvfPgZ1As2jT5Z7wbLK7mTcDhy
LdrMdF0EyAmanmgnT2LA+J6irToP05xCLivVURmWmJroBqb7LRxvB8TYWmggz0QjykY39xMiHZfY
P2LgGimDHXBe3VugM9QrN5VT01gvr2aqkGx0I4IhpffLARqc9Awrn1Si3SePUbCC3udUv4ClOnns
JkXrCOcCuEZDyVh7PiGagLg2AkJJCiXKpxlU0vy0ufcI7Glr65NSKIazApdj/0eo4OIXlEDLsIbM
2h3pf2t25O33ZpQyG2hbbzvQb41jMY0kRVbo8C4CMNYaZPSux55OflNc+a+wBSc3ZgjspiNwMVNr
2Z2TdJa79YWSiamN5nklEVgwQvU9quqsKBSnneX6tm98BpmW6gB0CEMn4ZHlaImjtxpiVysTxhum
LzoyhpW/yrY2GXLKOMDJ1Z0w85JdSH+fd1ffwN1WQHHaX9bii6MW5nQm2iwbS5OX8RMeTGKVgeVd
sg0uMAd7u29hEM9MBORMx+0hhjoyjBBloIGkcbbrFSAqbQCf3MGz5r0ASiBqaXFHKEJW77XtgPEW
QIX8AUL+fT8FlE997DhSCh2k66oh5xuU+l2m+PIjyAr5tAmSPSqcCS1NkM5nmL/iU+SS/VDtHOYp
Uc4jYG3QoH0UB8saRLkLHX6+SKnFlhreCq3nAw7xGTrh++UxFS1UiHSIlKB+XBuyIMtvLcSbBl+v
qwWSSCt3+GwjKBgdqbHC5SQ6gBMGUZjsM/gfahzJ1M5VbLwYm9rVSmONcT9kOCsbPMKMRcGp4ySb
ghQcFWEbRZlyC4RpZWNCuF29lYTA+XwzN5cIa/5oRNbVn/wF6o3O+wRsFIsgDpx+jB65L40igSWm
0Dm/CrffUeuci1AWV/VIPGac1WK13KluFL1iL7MmXRmZWSMj/ZLgeoumMaawMQMb+abWggMf21IO
X78iIaCaiRpv/Uq5A5iQ3pCgY1VPs5Y8PyPgiYJeJCNq1clpPgbt9Iyy8dYaatw3dEKXJ/t4/tg5
F+xZewh9+l1JPWcLwFof1WslIkkevfe6HurkD3qoIPSBm8ljp30mE7SMTzOzLVkmpDEgk110EOFg
lRmBHRxMMQRzrgbczulrQwLkHPwBegcgMmQhayWOL3s3tFd8qCi48kcYE/+qFLUasStDe3ggBpq6
LEVbqxPOeSw21PjeeW2KA/41i/wimmurl1MffXM1GV5XpuylMAnhLGmxGWy3WO00xPjJxnbWN8ny
8mTk43aDZfjq/vNxE+GOyJXxmurYBqP4EZ/QvB0JdIc337HN7X/3enWFWvrCFDQE2BUr0A8cZTEx
GG5C0eQHzzdRcyoSCAEgKj/IsPkRpKgN3IPtU38a5qDYq9zlQiI9lN+td0LYwG/5KHUFeM7dYIuM
hFyzvI51Y6dpZWraq5ROAinQtkQqblqWi5fCC9qeHlZQIT5bph+JZMjOO58fUJSgmrRI66hx+tKh
l4Lv1gj1wxLfiiU6vMsj5l8qGCAe2IGr3L4l88UKVXnVTl1JMZVklm2YBmhHjDvB/beMe++Yk76i
kfzMH+f0N8gqyn0T4b81CrEwlbddwMKihaw4ZpomX4o/CXWDIUFrm9X8z3/wU7DSCOMeXuJYzIoN
Xm4luQ6tsS5K1hqaxBPEmZalGJJjg8GO8cVJRoXV3ifY4p8MJzdkuyD6SNEor23dLm/8/9c9339Z
FX4hWjF544rRLFffhnF8hgfMUZ+7LJa8ziHXd2wKtI4RuUjOl1vLtDGKCaY47L3/cFGk1xXc3A07
kHGa3YTT9pYJuBLNMM8w9kFTUbdBiTJaOhkc9e/O592/AfnXyumKPnm2PObOxUTltkfJggqzhWKB
xRhpbK6BNBGi+YFaSyBuI6xAaomllN0QqSKIliq684lpuinXzwK+rAu8fuBKmjJzh+QWstIVPzbh
MIcYK4UM+gBQQ9zjlYw8KBOXYuCP44sMeZgkwH1YohxN4twnezHrtfoAMDT9sv/cfosU+t8teqNp
WOqvsw+89+E6mh3wBw8U1+eVhJZzehEPIboxz/3u3+wxfY60GnR5/i4EhHla+MWIqEciQJXWE3gX
qK8b+HlgIOPMQY8j5QvZYt5fPix9TctCWc1TFlHK97fBXtTGNBNsDs1es8wODhzsYiZkRqJ7jJmE
HaUJcZzS6+/h1m6lh8Be5djskp+7DVBf/VU0bbYE5sXImHFOhV60uuJjMm4JR0F6KeWRS/q5qIso
ltE72g87wQCfDmckXiIeVbMe6Vy7yDveeR+MFlEGLjHNXAqK9bGo9LZ5H+IKfmNP6tR4Ce806tKX
t2+hRl33r+qwUYM/sUeikCPTKZ/iUejIluctVwRj/A4YcEJ6u4uKY1tpTjgJ/gAW53qI3lezrWE9
bg3dawFhUn0P4uZlB8RTe8nsRsvQEqTOHArg7xDgJ0KuyFWTh5qR+kWTRqmnkzgymkt5lTHbdWHe
BhL65Ti2kLnpl53/JmePoy4AmcLC3zrozBFW/UnsmeepYAtyDcV8fx7Bh2ipzWci2oMDDdqBrkWP
r6T/FBl1E/9FEHoqkQTLNv274081JoCvYouDpgLOinn6g2kKY/YjJ3k1vmQ7P3rTYvpENMxQAc9L
VQ/SpRsg3rv2+EHavUGEvC1+eYrMfJeVDNNsOFzZXeR6ACWBke5WbsEiwtWBS6/IWs0xLc/A9y2C
h4lX5jBssSyVZfy2thVaxCVUdbdkM7Tju8FJ5qq36v9ONvwzEsQo1dk7oPzssrE8u4+JVt6I7+OB
ASK5SqFIXnUGttZbkm2WWJ2BwuGpD/KmhQsa75tCnG0IO9ZzVis/BTayey/4r+xuV1zsm1MbiGFF
yj62nLOx69LiCoe/n15YJs5TkClYF2Cm8S+of2pSKUgskwp9TeI8N+ZpX93+bKqsxgSIGbpSTlRE
300qZwD599pUTbwnfNR/tv2mRkhg0KM3FZOBfmz6HZrd5YtV38i9I7ePZ1gXvfQ3WOLmUbWQMLQn
25YS1qpR8fBm96Q5DY6M/tKGbegNNlQYj0enPHdcU2ZmI0HlcevkKoUWhKW4NWeuhf8AdLOlaYYe
WIHmDvISH4T7XFg0ol3gTWxJVrqk6lu5JtqHHw1U5XTXCgY6ntr5QCSqlTPPJdS2Mh7B4+MnnxJT
NUrvHAuKbAYOj2QKmnDXBobh5S0QkZinM/DnmXn2Q4ObGjDZsf0J2qiQfQdmivQlc12ytMWETqhC
pPR1ZVVtjLt5PRNfJ/9h5HpxVWHwBf1xwTxl58ynIIf+13pOUMv4ONqE/c4xW4001ruvD5AJ00ON
qz5QtIIfKMhFk+MSFKkfLS3gi+NSJ0ivsHFjdEoxG1GL673ggPIMeuww1fUEu2N/QwdF8LDStug+
SPKZbKjVAtGZQVZlAJiURep/L9CQMZYtcKCOLKt3hL6aAFK0ozUxlRHTO62u7o1prSp3HAoRlsa7
/Wr6oBE/jJQQI31yVsy2gi8At7TfTf73fwFn7SNrCIHuzmliZyw9g4FJJeW9r5Y6aDOc7o/eUuLB
gprim2bNt+pbGc9KKKtr8xA+YV+GhCazlK8aNv0H0ioZ+Mn9QltEm/Or6Vyk0nOsZtD8WVK3MCDG
T+UoelWHkTsvWNzwN0PVOwdx2NQZbe/FldvxzQTm/37BLZZWViuPnZRXxapFNoM4yfvgHTbzxygi
Kl3cnBuhNT5uj//JTHwIKUTrGsq8hRFHdsOQ24xVwq6ImyZu1XVY0fRyq/j4VB50oykF/nWDy5IT
maMv1lmJOXrI6ywkjQV/PfdnIo39YYuNL5XtxPtfeVCa9R5MuV+vY70XJTOlLQglcU1FmrnJie3K
9NbJhZCv1lwUE39bfGmJbaY37LRjH8oRmSZ3CViszYhT6QwK2Xsso9R6DSPVHUlYej2+8JTWhO8a
ryslbFkhh/BC1S7S6yNHEM0znGjHmKQ6O3xTzrXA9RTSTvCi7iN9u1zivO282EcvsCZaScZSjO/S
Xw2HOxiM2w9CKWJT5xE1bqw1ESblOEAunFbENqFWyie+Ns8nT7q3KxPXy6amE0O6tV9nBKg5Yy9H
+l1R1zeqVvbJQd+hDPb5xqyC677JJR2eziaBhuYkuz9aAaY8LyTbGzCMEG2tJEhrCeIlybXTOEua
P+QQdK/BTpVaQtt6SJNntqtLIEoAF5aiYWHxtdtXcLXk7vGgDiGp399Slf5ddvi2cK4JCM563y80
oXcJ3kKzWH/W24KUxcndebVmKxuKlYqEv4yR6R7MuKkBfo7teJ1qxfSsau0862OEZg9CrXvyBhUF
XFeoKLA175/tVH27Xzb/hDh4OwIl7CP1uC6TPTsXbnIkFV85sHH/xaoaXkhis3oZIpDo9MDOJwux
NpRB+Fen7M9DfBr0SghjdP8f/wtqUv+XThPxpt0Oj/XOuN8dw1sADiE+XjUMhn+8erVjGeLXhhpC
OP+8q+n0DR9Ceyo273MgL85O/Clx/+DUcLCHJPGgLdwLhBc0oLUeOLgwdjmefqeKOykm/0uSWQRf
JzZdzJu3vhRL2rxndGLnoxLSAC80U1tduslNtCxi8YOy52cBmSaRcIaOmCnJpKgDu+J7Kze5Tnm7
7sb7rFQui0Zvud0tl7Fmiuz4cYJOGaPGu75Mmo+37gdZ7EzWHWFIZIEhoCSODuF4eEfaRqsDqQax
0GWhpUsBgJjS9zkHmqg+uvDsSOT00Vd9UwK51F1/EvFRiRAOcDR3+PUMmx5WB6fScARUaYr/bFO4
oglYOf8fOvPfLoQIZ8i1wUaQsI755c5bTYyqr1LpH4er5e1J1Icon4OoF7R5bSX9paF8WpMcOOxu
Vu9oiFxYRhsnqgoewK54lkD1nLTa2qVFJyDrW0QNpD9fbkfxQ5hEwLqyQmcsQCV7uODi0dacpGfE
q2ZmM3Xp8IIieCFzHA6tdRACCY/PXRrjQw2x6uRpzqQVsQ1qEgJmL5aftkB34LDjJ5RWRrQEsul3
fJP75jPvz6R3vdvC0+aMkdKqdvYvS43NAeZVLZXofRJS7Y5KJmGD1RahARwAu9nrx3D2MzoVyfrR
dHXu1rSlYqvt9533dJBWe1zHUq1WIC3s46r+5YUCBSfvkXIMMCdGGoqLvvOqwOfX359of71A6TYD
F8MoBldms1JQXB7EZlqsLl2tyoJDkXYlLv/TNIHNrT+BNPGPLurocD0q+xEjZjy+hZtK1L/X+j5b
K5mBFLI1JJc+uRvJm5f90iyAEoJutc/XFBiCq5bKJ1psvhs74ISy2pdiAHehULtMiLPw8Kv+2crq
Qsy3qB7QSaao9PZrUzXFOAOJKpKZ7GA9wL4Plk+omB3VfFOfhNdEje0pLoWmbpHWCQg9RTQf60WU
zyN0fSOdcU9YhbuxL4xPS89QiCCyhOxJPkc28heFYXipGo/Ct72z5cTzdU4/jljH39VyvA3WoenO
msUN41tZkZ9ScZ9kV6x3+E4uMrxUPmFUIy8nLo1mG+6EZFQzvlG8tifKMneksgGewgq7ZAu6jZsW
1vooySvBWrunxUPEcZNLrfkugWC3j2nXxmpWTwTmkQwtWT6VbCxgUddiOXK3YkHPQxfLIgaybZPe
72Y3Aj9fNkHMD34Hlm+Se8LirYCWF9te4+FqTHlaPaC8W/FPoOChps4AGIG7mTAG7xYKnuowzDy+
4M9sH8r26qCgpHP6lQlHZ+Kau9tjVyM3EZm+YYm7BBfVM8NuCmkQCPiZt3qQLdlrFDlHHnuPS8ls
8qENGALovlcHKarui0TbHOoh2ifT9YP6GGEf5hTTc8ZHMrXzdFKFENNhdejDuuzM7FyW9YyFaf5c
CN3gOA0XL5D/c2m1O+8iPqAjaC22AI1CjOOZuu8c96sZW6rFYfPqyEUq2Nedhw02Vbsl/tFe0Lss
naITHvhQ5gNHCjZ1F1H5iwU+GpZ6jewnyDmlP12uguWuex+7reFwc/4dZG/OBGLF03+9GbC/yJLh
8LraybfxpCvrQtsBjEwK1/9Iryp4GXzhLVgYyvaFYVmvo+t2orFWW+0efDgJT21KURKln1bXPYMR
6tCtWvZPFPXADAWdE5/7kQU0VtxKPlAMqb7Wo1qCBlD9vArfyfNVUO9ZeMOYwipelVbGniZc8UXX
FY02F/sY+w1zi7ejvmH5Y4rka3Gttjr2o//Pk6CJStmqu+KFTCqdKrdM203Q+Pv4GvNmrKrOFbR7
OfyQCuJaBcyUAqHINs+NIhqJft2J48/0BRYjZ6fNhguj5lbo/DfLRe2tCtYqUAL7SS46qHp85eWq
bTadUndU0hl0hI6RfSPuW1TNOLWpPWjE6t03B/RXRka5liMIqlq0Qg0q2DoipxGrn7NfL08bkJei
obPsXMQnrv2kChMr+q8pijgl+nsMYGSUfHZNB1lS9nAVFa8HOUqTyWTi5FSdIW6l1QlvNwNogZB9
xLObP3Q8t2LYhgwra84XazlceJHoRv4jzFp0omr9seS6JV5sMa3irk2O1dSrfQ9QRNX/Cfu5qvn/
mP0sMxq0RUxqMw4bNxjA4KgV30QZ8V5nTtD2UzOhPUCp3a6CQf836DGbdNyCiFRqFOa9Z47mQEEp
TAHPSEO7+QqSPkhnXu4WUhX8QDyfw7DhiXuFPpT4lsZ4wR0UxHywLKcjciwRUvZqBM4RuSA0wOmt
cjkXQx3nnJJRYMcESdX/1H0Ir3ZUuLMzerXUUvLEaoHzDN8az56R8ggg7JOv2WOyGM1vIssMsz/l
cPZOME/orpK1tHELHcRPmI7V7Ni0Q0HAGvy54DBCKQzq0QN3w4fgy0hLI1lynnraGtpGjlaUHyD8
vFamk+7oivU0YOlzTA5gxY7xfzd3iMJntoWxE6Zo3Io4JoxbC+JweJPrKFEBUNN+4FU1YXirFIEj
s1OJtcJ4v/H7B2zFuqoquTXgDJCbT/258ffUkt4Z0rOLQSa8lGDF29yMba7ehkXTvet/3cSDBwzC
5SzjRqzJjYNMkehLjR0Q3qdlOycLJFz+4TTEljXqW8Fgf/ma+FwfRtOiBfFjdbvr0p1iZqcrfgj7
emBItakEyjeg34qxPl4FFkxCt8IFHgGT7tCXX+jSBxOW/H8vOLE7w0XKEnoZYOnkqqqgJpUdNXDV
v+1NQICbak5JF0bRQMW/wUQpmvXUbs30CUY6LbxUJd8Wj55B2J2H0zYGsJ9syFILsCeL6OL357wa
uCuC/MQ+y9Mypa8/PbHvoXXW+enalq82cysFT0Yr0GlPyIt1Rt5R69AhNh6eD1ES5dxdUj4X/RlB
TJcpmcCVIIUI9FQLXuTVzRD5GiN4Uvm51jyPWVtfhAyToZENItihRZpohMrX6fPTpO+G6urtLQFo
EQJE5yk8AoxxDb0kobX+9UNRKWGjy3iprhE7qu7AVvckEG9z1eyne2djH6RwLi0FPd6PlrsVZzGM
PIp7dHeVyp2Mm6u2ZICDGi36DGGUo5HmIWnDTnCpjZG0YkdI8drMIlsyHq8rjBcScigJ1A/V3yUL
bKGo4SL81UPiE12+vFbsrhCpMxQlpyv9BlCAy84JfpUAzF1uWU4P3a3fSEchD64ODHtStiyQ34in
qBvXgtyIjPFGWLlvmCtbCtYJrBoqBHcoTAY6Wdhhpl2AERyThvZwN+dJIykOEkBVImkYcoNA95pJ
wc0VSMCfMWZbUva3u9NjubsRXM9oWlvDXWInHO3pWZ/WPFae1OMDO0BRt/iIgBCrCmaaihNbebS9
6O4kiPvD+gNpcRjuaDYdHMbwrKdUc4WbLPF0q4XtErxWYF+b1zpFrxx2DADXv4V4qUK3gCAXOdun
1xDRJD9Cdqs6OshqTNrkd50wwsduwuicwz8RWXE8YnsICcoh3nkiJJqIQfmTCdayzLFDYisNPC2C
dZtRwwXZChdaIH+6BT5Xv5uI3Ng88dDiWKKR3XBKjYd1w4yfMgdBDlyl8wz1wRsPGYTx/VazsD8H
2OzgVzd6n35xwviAaB+9GWiF8a4tlWUuq5hwAUDDXqsW0s/E8TlDd652ue/YEEEC/hgmMF+Sj4Xf
UHH1z9td/v6pe/dplG7/Fz+wSofwZ3CjBVbddztj8ji3dQN07VQIOJVn7Qn4J6XUm4YvAJy732q1
EBrHfP7GafdW6exogze152EkvrHADuBJIXaC1JhVSVK4ywFnlL/njZw2NzlBikq+G5ak4NnqF+8X
TMRsuHnJVgaCV9YqI8XLorN5yHWmOZEA8vgbEvm4KVsqYj+JvnjXoOufHiYbZHZTy+5wJ/1sty2H
AgvTPUvX5QT/PvHT8FVFY7TuesA3T5upfzpema0rEZdi/j087gii8xkfxpjNCatA9ZIu2I+JZXKe
2MCyxaQBWPqx6DmoFstDXLCjksgrD2p+QjXDaHasnm6Q879V0NlemfGIW6347S84iMeujE93SVEw
HpCysVA/2h3meGcFSHYOYIAz1dbm/2YiRfGTqk4Z9eAWEkHR5Gsl7bVBW3Kw/Pn7Lo43UskiOGYC
1cHj7enkxper7VhUiiwyV9rUb9OkaqPFnKGA55+M9dItJPIpU1uz8NNmGeRdxA+xRzFcXl+t0jY0
aXIecm4z9wU7T+MTtHb+9PYqENcfasmb0TawcqvBf83o8z0s7rQZ7g4C5+i9VbRcnnnpH0bwtlp9
hkJSH7AKWRE9MwJ/WpdkWoAdOfONucDzyWNorr4foigRt5TelB+iGkuikrDgcuI5Rqfjvjrl8rct
Jt1qr6fGYGkrrW/bJXLbUERbAnsdIe3aQ7HyLgQQr4xnkKt1zDzwpdKPHjLf3tbdq8LsA34jhPof
g26VM5AIjCrxYyfGXffN9+pHaEupBMzhHMop/9aYUb9nMqJT20i5OiJB7goZ0QqAfzvLz6XXA6Vc
4fMor0XD2TW3o8tHOMp0NRl/qsEltvlfZXw0MkytJi0n3gyKbaWCxQNLDWe43qqFZLNKzatRKzx+
Q4Bl/PTC9xYKcEe7kH6B6wTZZzmAmkrYS2Ny7qVYANjKR5FWLo5Jbg4w+RUtFaY5BxnIsJF4RK1J
C6Qa3GCY7uijD25GYZ8rNSkZ2oEditZegx34W7O8nhQfo1oEyRwy/puQXkYoVd21YJ94l9DYSZf8
pw05KqEwAzRApAxvSf1kSwz0wx2DbvrRCHPa18TUjQQ2ITOTP9sh6gEm+qg6VokH10XsKYhfnrvu
Wj+3Snw4xqii1/Dgsl9uViYO6yB2zgLLvcqWgfOTOUNJ8c59UFOND5tXNOphudWzjFHeHawOjDZV
Wy/dpah31m+iM+nUun95+9bzOIuhrm258Y9BLeZ0ua8KTpovAgD7X2oWC5xiCoCVXlEUAaPSyT/5
kHJnsEM7aPGL02QxLAcLBs1fA+SqMirOa/c6v+9d1ZtsXVD+ZlK2w8NDFfFRAM0Jo1+An2u4iK1y
eHAyf5Pm5RgQIuaxqzAnHwwSx2wrqdKL/I0dDjiYi3/+dPiXrtTiLnExhMqhd4/06uH69kF+m6oH
k/E4/Ywx84VCQuEDA1aVzq3awpVDjMDMJmgKQmGsLXwUTEznKNSOJm+AaRAFDIMMwoSesduKuQLV
aT3TvvYPNc/LSJRnREL9Uvd2CmhuI8od2PzA0bWTHdGQ62Xi0e7mB/pL27DSFbRdAxzUopJvcyVi
yu0wRNmoCJ2jVmra/Tr4V1s1WHO0+Ky1vytVqMtTVAphoYHnUde2UrkPx6F8wVZ66TcZTASrvAzr
rpJoabZ+nBIOFi8k36XZwANx4PQdyWgEB8StI+F/rXB2KlfrjwXRgOetZ/zzCLQJl24W02iZpzhV
X9ycQjT/ogaH7aRv4zVPc6aT3CwzjHJHO9utVkPWemsls6v7ObAdJb0mHtChq+pdQYheUTdz4rXD
Zy60Uz6r5jfGkAMFnroOWBNE/QAyI/l3xaXovg0qRIguxSnqTtLfR+TSChTxVBqradwchoaNcU9p
kP1dJ4gxcIXtn7qqFtXBS+sT+AL2EIvTm070IbmLZCYWRnijNSabqrpsatwmgoB/+NVmtomUyc06
VfumjtR+rJOUQyg8a5dn3DI8QbHEL9RqNnSWgsSnO0/eaDtiV5G8HHwky3TwjxT3r47hH4wtDFsA
lMk5Xx20kBOFRCZt/p4QvjjqnRWceu4utmxd3ROeVUxFi0/C9uzUKDHwYR0bvXMXsmGFn8FOMTkt
DmOwXdv/PFVaB/JkmvaS5iZaIiZYGAIY4UzyIYCciWu/lGz3UO063i29aNrbL2gtp79uQbA6l8VY
ApNsBn+rc7dBzhftuCt43JzZZ4yzu52YZtEy7wKWcyvGySWFfo7JgKOZ55F4Pl2/dQ6wPmqWA923
6R1/ZcpH6TwYxqKmcVkdNQ7Kf5CaUmoeXKFhDvoRHyrf5VTpVx+3fbN1w2FvRbsIbvkHnLBQlj5+
mLIJYV90h/XJ0E1UCIAuzs/Uz6D9uRLxdtuPTDuWy517vcUKQjJUb/7HS9mpRgup2GAUUIjGld+U
IC9ks84ku/F6+9YaoePFCA70SkY0Krgvvcc0/PmXsD6OfUKTTGHjkg2MUfpCZ27sFhfJdNB5Sk8c
TICIb92vwsd+6VG57HCTtwv5Kj4W86BGlgTK2U9cMPdaLoFXC3rmDlsxt9nF0KqGdiBf3T6G4oq6
kRtOrCGpYp7JxFxe/B9lUSIqvK9vQPwWkHQEi/h+IDWMWvIgiYvkI530QjcZszB9cDZ6SUsVR48Q
ndz9KQTQj8476KSULNLjQI+phsC3MfRfbclo1Oc8L7ApeehBkjJFEvbf/AB6AIGQNL20XXogKz7E
+Pek5m0sNlDYCEPxWPWQ2NcQrQOhkDPuJrUHrC/bUdu0akz2r47Dem9V1vaqAEYc0uT5uYwLa36R
oN/pDOzOhcH3ej9OIlX/2pd+XcUiynX1EXRsFo6aBcQsq3z+naXW0BTMW0WnTSQr0DepHYq9hGPD
NXcz3A7OqbAhIKvjX/SV7yX0WqLCCNkQ23HtQMMowLF5zPzH5exIknuI4FiJHqK8C80I6uYPpjhD
G5zBQe20oGGadxvTywPRZDMLHD3u+N6E2zv4yjmo/0yCc2OAc06V9K3HZtcYazCdDVxel7jFYhHC
S3GdvOM6RUzdSwfysnUPrlaypi7bkToWc6Nx7Z8/C83RRu8r/nR4NhyUb1taIxUjaK8MgeK9mkEH
joheVFRxkKIG4+16q9gChKa6Ba1MHFEh+BLpcESOTY9g1coZYmqphLsLaIYlFIvfqiYlza4wa1hP
idXPybhe8QxWiPCrLhYas0Pz9UUbHTHwbu6bQhquqh5lNlnnTK3zZzsQxtR75LVn/9Edyl5jidWJ
X5M+1e5Yk1C4dD6dQG89+E4JMd2XacDKqZt8f7yuVYlcW7wjwKtasSNhGMe9N+VWZOoCRg5mZle1
MG1ei2wFTM9MaGtfdK9aZEhfY4pbEIJIZmP7YNZGzqFfsImZdQbZc9h4kGMh2VQvHpDe24jY/8Iy
NJRbCpI7RdI5vsQGeOM6Yg/uVulMVhx8mIb0VOZThwF6+uQGXm72V93xToHe8hH9u6zn0mdafrMz
tgrzQB2e/UEmCgqqUDBom3/ujv5DIA3i5ec8oxlKx02+unDXo+g5V8VSMO6ChdfbO9wisG6VHsly
7pZbPRMNIiFDTtGAZ2Uj/QaM9pzRdzjOVP95LEiMAVoMvM+2xPUvAz37jAHV62uA/IN46bQDSCoE
v3gkn+Bd++UUovbNxIr61T1uWxLm4RQHkujPaQnowAMURYGmVxlrnYwrE3wiyjO6iNyBYw9yeGfP
X6MR9ydS63a7w47DQsB52+VEg2aEJRRej9j/UHRLKhPE5x1pDVz8iKYEb98knXkdyjBDSmw/BrTb
b0/Ea4jqORNLBShbuaBlMYSGYDcnzEsArseHC7ptmOokuZ3fdLXPolLZCFqv2ID2M7zL52odX3Y8
V5TmGqs9pWh6UcZY1Na67lb7rfQgIQtIUIfkTbsMhoN/Az+XREuY0R9DyqY+0e/Q8D5HTedI6rkk
vr2fnYR9SJPFQx1EjXb2C6uE8pv8HFEyCdrhXEiWGrE/gFWaeDtnXaO0+thTgIhcMTGa+gbv//qE
eXEusJhaoTVzMPBDaAwd/dg1CDZnlq7ZkKs2iO6eVIi2RUtoFdq9O30Ol+4n9FBXD6dcwYA+lq1K
BSJHE1OQFNyppvfQHPYI4wouGZpl/FO8LKkio9qO/t8Vo1TOPajLtLexuOsCXi1QLYzVQhYTAOPc
z77bJfjJ42JGcyPtNfBK0RMni2xWHXqrXwERWSgycjP61DnfBdTun1N/4AOUEd1CyJwnvjWE/ivP
sWSrB21iGpcNaOjjmdQEf9vPDbgKx82qXxQTNBtIfRm4U1m4kEUyJv3YleaWvEmUSDIhqPhqArWo
ayxmZfr+62uskzOHm/881RwTm5QCXFmrGMjsb34XK0NjVojLyoW4oRI4wzUQOKZxw/6dYhdEVzGI
A9o20LtmD/92N00BfPRPm/+7GI4ijguuysqstnssuCBPPiIXQjmME2EjV1q6MWYD9kfswaz6oMmH
G8NpuaX0RL7vTrYPuqCh30KC6R8LoEynaOn2xdz4V0fzJD2xEcYrqg+5/cxqgfundBV0uCcRojtp
z5xsxhfgPqqgavzCAmxkjc6Pj8c/M2H/jKtrOPljcfz7JyphknAyuxeRHSbAjd55KvYGdVdUVAVU
bc6z3n0y1aUnR/+2S4gKvuuZRsj9VvoZ+AeQ9YA+9o/NuUw0IF9mu5knUb5B2VjdK8KL6Bocn8rc
Er9l9sSDikklUFRLA2xNXxiZceSrYfFosyV6zfomxhpDiwNznhknvyk8GDn8BltYGEdu4TeSFi6q
oOruLYkKtrQtH7zp3BQ4yv30+lvAWBiyvrVzbDQL5LPm5rRgdTOZG/P/VmJibxuFFiRx4b2+kWOi
bP8/t6nlJDop2xtE7+mdTGapH/sF5FITd8UtXDwfSSSSV6DtBeWiXtHuv6/27nP/bvCth/3pM8oz
/UXhraUqc8BEGYB/b5UZNK8RG3KSpz9jVRDrY1zYa3AuQL1Qt6bkHLfEutDIW5Jb4fGnImyxJ9j3
OqzyTwsZPr7IfSC/I+28C3PpHTmwJiD7mm6u8k8kDNUFI3Rtb3oi0KB+RNrOaGkCvxQJo0EknNW/
7qVuX/uoUxnyqbtwLUr8hmCyj5bS1G/9NerlwKeWHcT05hX5HFgfso7tZ4zu1R4nRwskp3Z+h+hQ
yDZJhXeM1S/gihg00+N2jxUvFsBvKRpNs3748nfiwUWAlI3IPcnmvv2cT/kZ/ONAbHGCBob6H2Ui
U7WFSBG1oDQLIFT9OvSZrI5ZgCs8Er1F60j0I99wx40XEoEzoF8hjPSVdsOTS6EtjbhTxHKdNN08
uOeLnYzL5pGBG+J5lw3jghrOsQP3NnW4XvprZWjjKdlodbqwTue9phZNuEznOGUoPTnhF2OIcu+B
znOqA3pvBzVhENCELPgXPl0w47NpEx3kTmiJiFcRTZGcXowPgCKOxbTsq2IqDtnQiu0oY9wcTj93
eg30u5axemkiy4STeEs+MYLiPmkwIx5nb/OPBFHa4kfquIahaMUJbKSps37ktnDVrGrAXzoVvoRH
rjFhHWgJ1JP+aXItV5iB8Yl5IZ/y4UFfjvy+W5/4RbBzdW1pDGZCbTg7fPCOwSITHXCevxWND7eQ
h5NInJanSw1IDC6/+gwyuEwsXWPmJ7ZOwbSrjIg0EdWH3QMp+ngi6geDR9ZnAmPZSyJNQAN+JuVP
CZIWj29K/O9h4KQGs+5SPuaDTTmUL2eHKxRCX0YErXBtxCwhYDpi1nyLugCedG13LQgiwgrfIbB+
oDUiwq3Fi0ICo2FMwKZCmRsJycLAZaOZatIz7SplWWMrWG5FmXrUrYbLUAOKtOmF11rTQ29B9qjR
eYa2tIL6e010KKKVYUNjhO4pJtvwqB9HTbH0ELISHqJxEGaf+vQg48FTXNAhers7AhcApMABoeQI
embiFILNfqUXWTK3MWrbBoiQn5nC2BHI1YYCv7aFItXbSH2AlivN8STmYD6N776ZSTxOYrYycE6F
7FcbczJ7idyvIVzZ8bg3BG5dEDwheGXcOaCYCa/zcnAFfI36Zea/Ba2/3ocbsSHCcPe8bcC7djb+
5PAeruZOIZbjZt+JmqGPM68+nZws/w/hNY2IoZPUqHjQXVwxp4FyNwU6G8UkGAEmGU+0kHPYv8BC
gspiCrbcTODYSXMXcZf4bzYOUiuGIn+et+x5A5WEwvUOdpRTe682RUImu5DbrppGyPDrzS4k1u6r
hnJyQjMwDqLBtjxsyRcQGiYAZQbXitChEJ6FIby+XQVUbkeUiBYq5UNpO/P613lcYUJXuRIK8/eh
AId5b5e0sXr4w6Usrj/St4lbTehZl3wtWxmNvZQEwb+fkltGfzhN4SxZ78fbCMxFle6en+yYSrXv
TUWXztpCv2SfFuP0EnDqQ4Er8kf1rgE1DeVEaztgnqwv5tQ5BLTqo4Em7sIWXglrklvl6Jn8H+Zd
xrklmVRU5cNQ1V6bCX0Ks1Nkxkdt7inTSGBDICIfZUd+MhtxIrLwMa/oD1PE9T1teVNfv852DbiQ
rFpvvSvadWtF5XbeZ9oCNe/B/NjKThugHfht0Aqe7DYOXpIN3Zdno8QKssrb7gDI6U3HX94c/NuW
XlIhksymons0BhP/QUwIbXByCicUYpU9ChpqqlLtSXGdM1PY34LF1ARP/Ej7RUQpkGdyUKwhT8AO
D6Ls4F744RX55LyDm4awVMP7rhWyLBgA2gnZ/u0g2feNPY+Hsi6+6tCh9HjDyHan71JAWSAQ11je
xFqK7jcQom9dfRmMKN09OcmyKBhtxskcrecqzcsPzNHPF0I4S/pMnlVl47p0mKtmDtNToqqzr0Q0
TzqyXmHxB9w4f/ejNROZHjv8cz8UVNnq1/CdhHvEgbvE1CxynX+PuE6aKpwZZyb/Hd1JGzdH58cH
1AC+WrFNAL99qW4J/78c2e7g+B22hBAjduv5Xe49R5kDqpnISevsvWA0iy/3y1lxO6bRSwsJRm4P
zM3tl/3MoSICWnhYQl7iuN4XLNQ2LHGOpTKUNS8AL5OcRxpAI/8mwHH3bWUPzj2s/OqlPDQyGbhs
Z8RDK1bqns/sndCqp3dyEj6ndeeNn9Kv0VbO5rU/cb5Dz8NpKYci33qq3J47tDsVHkRsz676BgZ5
ZADs9MXwskzJjI0mSmrqtiFTMSlWrxE+2Hp7hl0hdIJxP7UkR42xFPHnVKXp2skXXOLOrLXNH9zk
HiCaEu2LKjEPNSlWWNjvTyz2vADdZj2clJhOyCt6RU67COp16YhTsN0Ktvq+cRe7zTtU9VHcGQrd
NusANY3b6qj51mTwvUTrM6Koh1O2DWk/0X4T2/oaOEIkL2IVI9adqUNYGlfn9Q89fyAYwnO+R2br
tgbXa88GOb8vVYAdXdwhUguJ8cMalIQRCQ2NOBHNHp/mDIHH+SlvSQvGBy3FUKRUreL0ihGTDDBV
cUYmwqn1qkadVStKDGvEgNhmNvob/nWOqim4tB0y9s0u6HlHzkKzbcM6kT22wV20Z1bKnixfVEJN
hmdiYjak2U36RzUTsW/4Bc09KToIsjtroZfHhf4W+/YtaEZfehh6h6XWafQdJd7ngxGVc+eEQ+BO
2YWn4EvnJWLIIFN/I1BC4MEZiNugepVx5IimH+EMjWbX8yd39Qlf9M1KLr1uCrkpZU81dvMEF0Jh
lGh3DFW7pI8V8/hER4UQ3FUOlLLWzeO/EZ9lZDW1hvOz4quseZe2W/6vfK7fvF2oTfHkdtjzIZHy
p5wxjYgrODsd62Yru8ivVLdcwhg29mkyKohZUckQctx8B2/tq29d5DzNgkGqr/f2vSEJUCwFm/ji
6+QhKJgNULUtvWED29ajZoxMiiMYf6IOx0MVeJVcpO6ucpWLv0BgbGKmslLe3kp1hf4A1DdnX0kv
eR1pgY1mSsMp41gOjEf+saFivGko4HULUaxYDPm8yF2tc11ILhVi6ldPoIw9y8zV14BIjC9NbrFV
vASY1ErWmZnjsF/L4HEG8jL+RUMdaVUXn9upyRq2sS/gAgWaCCXxvZI8IxVUK4ogVnUhhBHdRMd+
0/2OM83Mk1fq9/yzr2JEoc9yBeUgyh0IWfjZPUHm2ntM3xstYbgu/6KFZBBgDxCigZupAjQ2Pq3k
0sxPHy7d1hZ3XuEX921DEmIZXXr89D7KjPcuFCRUBocrWMksQX3MOsOOIh6VHAgJZWa0QkY/a0XJ
Y93NdDijYEphgo/kLNOQbdsH6RZTIBSFCcfPoay21IKbCJqupUvPYOtzcjb/oau5iLAg+SFmNLlH
IklOe4rKdk2h8tuRwgwWiR7vEUck1A7dpzVjubzI8Mzxk4Q/f+yA4rLCK85rjh6mfIga0VehJKzu
8zOMzDst3Kf1rmv3Bprv6oq48vuabcdBJLoDzqYrJVediNoDNzdzwwlFDW0vJAEwyGtrBDNV4+Na
hBO5sI7ATbIir0QRmp/imTfKYYmzhBbkRoRe6NHk0sUMaKeS0+C4E7DJQgGoQh6V8TqXWFqLzAI3
i30Bh/YZ3X33rXxUytxxMpgo/P7XC1FH014DXbma4QFN5XzUzzTk5XuLfuAsFe7dl6pp6iWWFXMM
KjFt3fTnmk3gGBk8dPCGBnI1xAbAqLE89u2bjYp70wMTAsAIa9WeJJRvvjXcBychjqiJlG8t0+gk
lKHDegsKH0AncHmMk21CWbNeDl5Qx9cxkGhMynh90L1X7IRrCpMgpfRYIvlySS2lBscaGj79crBn
ALYlSC1EugXfl8fXEp2Cwj+VCzRfgmjXIt9D0OuHWHkzJLf/kA7r14qN++5Ex9V084/ExEdxOkZV
TBH+IMMITGWzXoaDTk6NDdbCEwt5MvxlU0tikh2Y8kbBnCJukNSUi62EAibmDqYGv/GcSwGZX3LE
22eKWLMT/E5aCNisJFNhNo8Q2Z94RBVsOay+6p3xm1SD2ePkoMbYVCjkMWAZk/LMddPKGN/gctU9
ctyxwK2Q0pjdJpAuKxgpdJHsGXaPPxOJCXyvJO+HTINMQE56qa/yO9WY3r8eGPYeOSobCJfvmdbe
XLCYKLAMJNHY2JnvGMlBXNDikfimJUXr8ufmpWQSX/lzguxYDLESVjxKTAIbwsw0C/dkaXhqUROa
hEUGqmh8wSdl1mQ3VnX4IeFP1XNlDFR1NO1awr5sKc25/gt9nak8yJrcoQ2wsyhflCIFgpSdz4kt
716GOq5yqLfKs7AUj+37CqSg/ztLNADFVCPnP4S4su19O25MNmWqD6+9EEwmasMJck4GRo9hnFaA
HmUG0I0ueLeSp3Bf7oyqOg4VkgZaPX/dBTzoCfVGfmE6kgtTTPU9m1jnMZ4J7dD34Uj7v85BqB6Y
q3Dcond6JdpPycKp5ypwI1bfUM69VjHBP8hJIMzRQpJSbLV8n0Xvblo67FgJ3jUG6rhxZ3Fh7Ojc
9MfZd1hNBwi6ze5phmN1Zw6sOfcLvSYVwpk1bk9M+9wLMo4bqTicl98gpIyMlnzIO6BWYDoAZah6
3sYg3qtYN2SUGEdq/YFsnkl2xrAXAnFIHE+nJYC5J2fuLDcAXhl4TkAavp9C2WbiloZsgfV6UwK7
m/+3JG1GmILT012nZIMp8/wcnsJp5W/5+PHPKPiggTr+LH9b9gztoJsb2hku5KI3SS3wK4VMYQSt
Bz3UkmFtoYxdsIOFNcfM6YvcC6cDtB6PSy/HVg00leeH3WLDQD5CT7oOajuQaX8m59wZt9w8Cn4p
lFgMovxShxw3Hfekb2Iulu7efBZs9dJUk32rk7QSOUs++nsFTCl8x5axN2E7oX37IeHQ9LJNjdBQ
fFyOjVml1fyMMOhzpz58mMcmY6se2hhHIeQ2O3LEEe86K5k/XXl+ooqMtCyfmcuTZG6jYJj91K6y
wUrFpTWDra8LoL6fVXDcXU4tySpsIyk+npJYb1MiMNhV7l9BweoPw+Q19Bwq0/Vpui3CUHzvjf91
YeJKJIxZ0I9is7u2jB2oFjJXs3o24ipmmGmSbn5wFxItIURMtVchfCFBiF1MbpXGR0YfAtJ4i34D
XyBm3htv+OVBJ+RGGAtpBf7+uFyNfIg6IAPU/RNB1Zbfb342y0x1RhlkgDXmKeA5wpNNjLhHbSAn
Tr1mQcV7744OqOl9z6Z6/m0KcnkEmDO0GM3boNGDY3o1JcQWk4HQNg2LeprcBacjJT/wWB4BUNEO
Ah+TyR1MqqG2/bkqJMrQhP+fK429w2EaBbuX92+TYOTmWrguX5HY5bMgydGodYjhp565A2Y2oKxf
QKKTKb5xH9p8k7TXQ0kC205DjEcg944zp3JSY8wkyAQ38iYL8ZsaLz+dr6bUTBWQnzu3VSSZLwoK
H7WnuFMlTDICu03+kVEm7uGYnVWiCnVL2IEyiOyH4QvGJtOkA9Pc50JaJZm7ZMEjDq389qnOaFoV
uhO2blnCRd2eTJuPRNOzi9lvAa8DxNvU/ws4WLq/qNjCxok9kV5B2e3vGBXKnEdRIs9Qg/GthAKA
NNT23Mj2KKERaYEQJ4uhTLU9JHTZbRnuV7cqRhLzK97AwcEz8vC+eFTD1XeV864XwJ32jepUDOYi
g5vNP7LjU0q/MgKUJAQOMHt7vX/zchdsvf7nRmk4Wl8xBCqlhL7cyFapSgjZihYQzk0mOc32u3AD
04htYvhqjDckW+YkpReGHI4x1OzfOUTJjXgVY5cq2uMnHwfPBCodaRiCRti65tEXepEar8nIwIvc
AMJtjmCp/2f2O5g2nZo8AwAS4A7Pd7jXvXxW+825gJxgO5D15rkYgPi8R56AIbIAo2a0Gpng7OJx
cNxUcYDSp0ABK+x99viQKAwgAW4Wa6Os/IEpoafcjfRcQqcodY3uhstqAoiFj5Y2Q86q/NmKAO+k
A8fWKrgGZNjlNR12jjTW7Bz1qnAcGI/u8MDEAk1C8owffJPgGAuTMOpCm4ZtBm1MiOwysvcdknuH
xWJ/Qb8DOM02VLA6OoZPgtbz9sVTFtABNjJCeIzFWpqVfpNwzT2gavNNhB0j6yNXxuJaRzTekeeU
KcifBxG53sd0CWkQnTfyYRABQ/2fvoloQT0lPT03wtmniLzn0AkUz8FqjIU0JpcM91Mn6zTDLzOk
QsSsxvD1Pryo+0F6UbUwZ2iv2NC5iPXFkmcaBt4E9j/l/s7b5SplWOvIk6D8rF4wYEJGJNRhROoo
uu7ezEmhAl2aeGJg9sjHzQcXpm1htlVHFDIMEN+rNZoLvZ611+LVFYnfTeK1Ez98veIDH6vP+MDl
cIa1Wl2+5ytzaifxMGtpIYzFGIPX2JYvQh3HMqQYaGABBQBNDxu6poyG3p9SurwAREoFnG8Gs5Fr
1caGfef7qxLP0Ok7L47Sa7ohgJBKurvOzOTJUK+yzJB6E/23NFhWZaxlvv8G/58LeBFH0T7IbaaB
dc6RhIaIatflUhyfovkeusmkW2VXuUwADMogswKoXEQWBCh6yw0vv6UmHNjYyBKVgcr1Zb0HDwa+
j8OKGEB1fNE+iBBJjvjCHbFETHSJQvW+YPA8pyZw6xVFv4i/4+fcvwxHP7nwADIv8rGwKR3aqI1f
1auobrHsx5VFRbz5mVFAo8tMF3Y5tOl9UnyiRDhzWbnRa/61p4DqXSqOmNRUXOop1EAfCHRwdVBo
Kj0StPYOOsThLE6AqgZW2q3GGAfoHWnplowHdQdc7iOvrW3Z8w/nHMrKx9v4tbFAkY3ePJ2RgEnB
YpkJ3Bw0F0waV3cyRqJg7QhHzE2hMqgODbBeDmvNlERicosguxGcf2Qw46EOLQOODYXHr8i0RIWP
f/xXsEXBA26vScDTZERfah5sWXmbtU0GZUMAwmSXf/naq/DdRCy4EyQKYp/4/Sh+ffsYNbf5RE5p
a3P6NN77f7hQL4TPGrSYYByIVniVSMJMUqoiVZEQ/QOq3dc2zYH0mIbybs5mozslI53z/D0cl3tC
qOAS+5Hrab7U/7Br3y5TjtDaZK8UbzfPffxL9YXcvj/WGmobzL1OIDkG3aaAvpsI3W9zqiH8861A
ezntQR2P9I5EY/FpSg4Xrd61WV/DCpBSMOqVt03XVsXtLunPvq1L15cYoDNWQjTCNysq2cjwb81y
JvRaQdAvEI20Ek3YrynRFZEZ9CijQoYfagWiLLC0B8v0RQ8XzoKnqW02KexVp6NWHukJfK+cWR+W
pWK0zqr8BDhX7kieTDskkgMCeDeXZYyasfKkv+caCS0hhnrUt6v8PuujSSrrZzDhxbvgOv4mp+nZ
ZsvhnesJz9b+vFYAGWH4Gk6BuVs0zodz1xGkJFQ8H8EsidxcnnYszVJbDdugeNonvz9JQ0qxMHOQ
gPCgvfr34Kh/ydqW2MX3JjCm+PM3fcuFqIy4TKcVOsLm0VZCERXhbZyuBQu6/DYNVSlsFJ9+0Vf5
kENYR8Mmx+5cXJ9as3/C2BZkgeQAzixCC/CX76/1HthdN4yF5ldtjIzseisoKgZ5M0QBjyPdwH3+
O+zXscJtDgrbwl2ppuPFeoemBj+5em1AKsTayxyo+iRG1DA/2H2+MtdSsCFU4OsdaYMrRj/yU+Yb
8688w4Y0IrqlIhBBy7pASM0zAvbVMT4aX9EL7AtG2WDerc2vUx+6P6qWb8T+xcIOlknIm+wQhb9T
QtaEQWyavnntMykrmZ6xLyJdTGbfK02bZN8849jD578nbWsoFPW3475ACNs2MZqPTQQLkhpAKa7x
4/EFkz3m4k7OQFWicDfl3mjWSDtjtL1ThC4akf+VntKjk81o6E5I8ZgtmotuOndkPIyushCSQtGj
xlh7QCIEsSTdTbZ1/XuQG4J8dMMeJpyQeEA4oKjt6cLpRtKNMWV4QtsXD9+Gsx6j/0iSGJEAJqpu
SWQN74sCysjYIQ+atEIPHT4JjY0ijm/HwaIy+9tYSxkvvEiI41CqX+V53Z5tXUuu9Brb6cLgrqC+
/3XbauRNDWRhuQJH487T1OzxrvY9kcaNOlWgsN7mQrLMBhLWRBMdJm4/kWBGrEwbSL1leZiM9mT4
FjsM+lmr7q91XpjXRXD0HJDg+ndCJ9JDgtjAG/RL6ZVIV9Sy1mGeq5spHhN2COSv2vgWuiqyg3vm
4d9ONBQtm79o3ZAItqTExL+scZoJ+m69jO2+A9rIeYgiJjYqgPIlIInN5opJfL/A+LNYHXvAh5rA
jOBgZfTOkJteXsXpbfN3C/OemHPFeSpbbXWu5wkC/4EHEGzztyyVBsxrch3mrVsYsPCuyM+jzZhR
zXhvRo1FHnglPIJWHMDoCUKzBjEb9fmiO3KxZ9eJrNsiLVRyUt+xYjvuEYrpFntIUH0HVN9yahM+
4QVK4oFJT/FF0anfofuR2u3Uuy4+55tlsFMBIWJGQkNZ7WCpaMs52fgyHyvN8B1RxllAtKguPUCH
YTISA59aGViNDSDzgbCR1rp7jjb6FgNNL8J0kwpsYt8UGc4Ktk6nvPYMyddX8aFpHLD3LRngyCsB
YpnysWG40cL4fll5fFkjtx99DhYajgYTIn2kHg/Q2ZS+8ouXvAp1RnAOQW9uLvQVkDYHOEXPPy8c
95IdgMLDzh35iNBbydJxZspQQ/lbkMcpNMf9dqX2r5Ve7WlX9hzQ04q/5kaOazUPJ6KN/7OxNXA9
mP8BCE76eyi8jpj/sr4M5iME0/IHYyReV+lROgaHymbhvMG+0jCTBcuycV6ZUze5PEW2DMVg8QSj
x/Toi2LyB0z9jQtDy0tH+ASntM5Ss6emAgQ1N+5RQVCR8eOCiFRuFxIH1uzHhjQL1cOiGAMXRrTG
rIeEvUY3q51H9qagpgEf1W8tpcfNgnAaQQhYcUUwnbpKGR/C6n05kNa7HUFWALMP2eGjvr0o8zi3
uhuTw+nAKrAWwTxbybK7Y+vgUd+uhYRXBHo4yZBtpSp72u9CYmDTc1cRKU7/VMl2tzK55iBhwFd3
AmaAztAv3yEx2uzukLZYUGw+WYu7svM2qFzZylRdPFKxUgrP2Mt+ZtGXImRLezllOgATeQC7YeLy
bkKMfvafCQA6bsKh+xsvQTMlUUlcALvZKy0e2VlYW09aQfaH6/j7K7FWuIoCnHi2z0aE9G/7xR8C
skHvBUV48KyUm3MzfjMT3x0sFwlrcDSjwb3W4h9N06SSiUEu7m7f/5GF1PrvpwhNWhf8YCFMxWKd
HFLCcYZDQSDLRO3XPGGRFBGIBgUAw8A6p6MoF3Q7BlDJGxH/XRIqWKgJ+TfzC+yxRyl46hwncKsz
9GgpKgmk1W6Or0WNsdW5RSHnmasoG0cfqi4Zml9KKEHBia5xJXFWZc+417G5ZmyHXM/REdgCJNsq
59fTD4hh1tnCNdNV82d6vr65+yFcOIsz84pPSMMMC/ZgKJg77qPyESOpPyUsXszQ7cNAPKaxGOra
CnYKoSdJxMEF13M/S4nOMYJZx5h9tbkQl30j1+r/U2eWJr+566R64v27mQTC+Qa8nwPjocQGR0dV
El03pAoAoEYC7z8Hi/aBhcPV9fAY5OGcMW7TG5pOkukdrf9LDHZATgQxvInedDgVHnspoXpErAg0
Y+dtuSk3xgP8LWFFB6htJvMq2X40OTBb1WWq0UqeNY4gaHnZCbq7lcxnSrXcGfjrTaRgiUP6Es0Z
3fGONQC33PxMOviFS9TWE0hOcXNPg9ipxptayOHzHISr9HAGNqZV2DK26LSUulCD/cNQLnJO0CxF
BC9pnPa1yatTqCUTxPGTz/nGFRfVubhEMTDS/u4qvb6Q0+9Y42Xaf0IQQDObjxLYazBbAmh9LrOy
Ll2cLWSrdsSzNXHjiFiQ8tteKxqIlK0294pO+ewEXEuqRLVM3K0reVxtu/RUrZL/TFe4HzKGI9Mz
TG2taXwGBGR+aVYJ3o2QpeiLjtBuhU71b6BdWQchIxTBkwlMbiM3OcodHBaOVdW1sreCvKSU3Kxo
exNVJLDblRdVTvAOqvV2dQ+tV5YtB3vZwzNdIalp2SE7HDfdYIabgMN0DWT33ecR88dSlDNk4Is8
MVrBeZ3YKc5fUE4kxTw04vFdOhw3v7pTpUNE0thUB5pnXAE0JuJSiB2NmxmQnYd1Rfaa+fxUHpIG
mHz6gW6Ol1oTDa157sT69HBfrwSqCnBAstSx2C3GgkNCHjWHXQCd5UDxvyvJ8mcNaeS4SyUnumTU
nSuIpnO1JQ7HYARxq2QqjgGCSPdNCfg02AUQ5EzKQ+w2xBLS/DCM0m1jNG7Neewo3bolyYwUovnN
JRmj/pQxOBXwPCCuvfx0noTeLw7nL750RHCkSUbP8i6yGHQ+gcSuMRVQO/JomMM95YQtzBzifuTB
EIdfdtpWRDi3t8rHM+K4dv/jpoWfZyU1NR7KcsU/VgRRfb9scIkyeJ6+A1rPUJ28Zucfwz/N1GIU
yZ157aKnp06X1HFFL+qU1T4CVtf3IXVfFHDPw2ZtaoQHkfqz2V4ev0+K7N1QZRK3yTWPO071rO2U
ZR17EqMzS7CRxnCC5YShl6RQwtYYz3CavpoSW+E7pA6Qqj4Vj4veZu6HyYspYjkPRtp1EFTzW4rS
ArkcvDXfm1YbTbEKvKAni3f0OZUUYNk560TeFJl/tt3xmC3dDKeUND02CJyJ4f/M/+EjWpR1d6Ry
cUjjMuuKL2vfJXTw11JDj2ldohF+8/dSe4c8ovahUgfLSV+jNCK80a1GvpqDa51RKloLz3amtWz2
+TGUgqJ9xK87IiaC55/EKec7l/BAiPmmIvt06uh1gJjK7YHH/soUYg3v4HHhBvHizzWPW9ImvAiV
lw+S2QkCq3gUa6md3YRAmUu/aXNBaFpN2jGigl6zV9GtmC54x2L1brMfqqYSZU/MXSUfBoUl2Mz1
50+oETznM3XbY+147WGcMlR8AFIwegfs6YX686hvBHbbXIciA8fTKKD9mjG+hO8aD+9tMHnHQsdf
KG35bjTLaO5kH6eD2Yg0tmuAh+WKM8SmL3RCpZ9z6MHlL3QqKGmkioYr4r9686b5/3hEP4SSgAvL
bbdeRL+kIeuJOgs85wAe/Kr3Pv+5/XbAMS/roRYPa050Xh231bqTnl5MO31j11JgIhKA0/DWhCfE
nHIEabriXRvK8KO8dmZpSIQEPhQZjDKdSaB2fwijQc0EoC4n3pfTbynEPm9kGk3NXLTueKA081/N
jWoe+dZ/MgrEXzwFaw2vwDQ6MOUxLAZQ7B+lijpZu2Hcd4GcOnsjVbxvICkMc3U6Wdk1zNgDV5B4
C/uO86mMJq5AoIJsZOKDeVlyX+nC74G5OX2oXqAsY0QBlJxg6xSD9rOXp8mgdHuzbS3wNDVLfY91
um2imga6wgbvNZf1xLUVRgDeDSQj0qXggcOnnncPAPtL2Y4Culm4qkNxdOc2NLK/F2rxblO6TFpi
rNHjJxua0XVv9HwesV4DynFgo8m3/JC4I6xJzdwCSkeFfpfqdA5SvpqhjXiICa7LIiptzJm5Z0Fd
ugBQGUALav+xuEOgWcM4e1x8w3I9nF4NTOylW/h6p9dp+uEVArtQ8t3dq6pxYXKcv6ScYBMIgF2t
hSGmVrg5F4HQdY2TYaE3IFz43IyNlXHVfPVGyxe3ev5pwDNkYeaTp4spRWe3uJfsSA9xWH7jb2Zk
wY7qE1hSZbuQN0Evkn0P0U7/WuxgDGzeoL4X1Gg1+wwGtPQyqtp82rkpHKNsI36tH2JpGSfGAo6l
BlvZiWRxkM4t4VmGZQ1AAQNSMsnjfXiDRm8V1LjyZ1He6pKdD2e2am2KuBRl9Akw9m0RyPxGg/K1
D4dwIz5uOCFAmVpGsgMVS6TzeRTI+2f4H7OML67Y2G3UBmb0dyiWmyL7igieusfcZrQvwFeD9JK7
ZOaRhywnmU4bHlX/P5QxSnR6ZlWhonuMV8FzDI/UqKEXtt3UsUuLh7XQF83ga+iPV/Iju2TqUMyk
cSfg9D9ipTMPhq07PsMQ0dYmI2zfRwIOzDYgYqlYA369GxSsZexcqqSWU0G8+adNeYQeixnQ1w+Q
0kGxEIaB9gV++5ife/1hWMp8ZoxNILATUpBlIPIGc4vgfzsHYlY6tUcZaaE//w1i4GPTUZlKgnKv
c0ytPZ19AwSYLs+3ToKP9HqUiNUeLMi/knvHXCXAv111N5LNT49zwee+9quaQZ7ishbYEeKx11P1
aQEmOWssGurfbcFuCv+2qSr/hthw0ce4z4hP3BD8+IGvuPICUzr8BqXzOKamNmoKGgu49Fj6J82f
xAI7xJQSDr9mEnGxgygz+/WAWl+wWDmEtLgrj8xuM7wPFOKBsqhvfAd1HFaIgqJtOeyWT42DEheT
wU5XT9whsLl5IxxStpXp/Zn/msLT5YxlxbWYtVJtIzJYrfVHsWSqejEeOf7jAj0o4zub9rxPjYem
A680r4HmuPMqKEXk88+pNuEzRbl72U8C/xGVNVlDRxHxkZ5wJqLzC0eUB8gjlj5UCc2/ULjtHq4F
yukkaRrb869GjyjxZe2e1bfX/pUpJ3VjfSrd9omMilzCF5BqNNSWOx04+mQbiAPlGA5yu79VfoDD
KiyDIx9H/PaqVigx37YDfpZuvQCAMKV76spun58euBUNWwQ+sbQ+pex8hQY/BEWSOEC+geIvkHLr
KGKSgTvvOC1rdvp3sOFzbSkayBP3rkJYmzFnM+KPqBBtwWfIgkGAcHK3ZGlDuKQhjfmB1PsBM+5H
xTZqy+q0sW8fRYh0f3V/WjoQAuJ/i8uhEdxQRBRg0P52T8BcvBm/m3mFy5RetD6u39A3rg8XGMNe
PhxjRqIRLAIvr+jgCFynsVoFmhkBvynmclvbGElSXUp4/XKS4x88Hdan4L0ud8sXN+vNWi9nqPTS
FHWih51KygejFORAXh/2u8HJxuEGOIVrdthKsk9lnAWntTzIT+8+IFwrnUknm+8AAZ98t/O8AKvX
oBlwkZwOwf3BxU4c0SNu/7puHFCiQYIpISaxAIASaQMjnW5hzS4sl2y5SRrqv2DPFvSeH5ch/+1+
rrTDnvUVW5FEVT2W2TOeYAQM3kRqEyustKFRN6WL6bLL7pL8QTpY6eFXIxUXCeoteQ8DKYgiBRG5
OVO0s7hk213yBYtAIcNiULxk0TWcMQTiSXDcyVn+bxjaQ0AkxptGVWTk8oNXYmNJCASFEv/C3hvu
86skAZ5TI1IEZpB5qqsw69mHaGmvsHlDxqzeluZbwmlEwNCz3O382zkLdumU01hgBc57gnXg7QqX
GLGxI+R3AYdikHisZiRuLdY/UwfABrDr3LzhW2MAUcUiPlBxo3dYKvRaL9x6JkvmhVZWDUt+Iskv
8TyWgorv1aO0VpSoyJ1KezSKRNaiiNiCXEV3pvORzhGPvGp42l1Lr0ebybEJfRJ7Z5eFYHUhQ0oF
I9qBVhRtPQiqQYkJ1SbqZveP0H+IMVUaE+Sk/1qdQUbzXxiIGweCkYzybHKC3mas6dMGhpbdb3wg
CPpuERHoOkZROe4of/szhlwGmWeAacyC9IH7/eXF9TOgW5Y+zEDXG0Q/ar+gyL20SDvg7JQmaThm
nVJZz8tCuyuvx4ND+dKr0QyAoTWWIRUzF5mVq9HTGQq1IxLIVOnz1T+Y9d9lItvzLNLj8+dFYcrV
iBF55hGRJfa5E0X8DITdlw+aXLKznwpFEXY4PynTCGWfAmgibTD8EMSva1KhAgZ8xA5Ocqx6MlGo
WMU4VMiR45e7T2fytJY9wp0OtAQA3xEYaD3fW4tRVXg4BXd2kBLiodrd96sy6r6cPYE8rjMRhMxu
kQkuH338RNcIJDmaAt/XIyuYxIHt+Ae6vyRBdpaVohgjsICpQKkInH0OMNiauHlIr5o9zXhqXS0w
iwnikrjiUw+dRMCiRMIVZqN/B23GyYXhaaGnyS3XRnOJcThWtrYDrJoXeHJZN7h2iXnCYmfS2Kv7
nmvxzNXiYzVG+unuFxF2C/UTnAiEGY1noklEgUPDcJrssiuA85fKSRDRF/XTOX/TPcCBnFATG5VH
oDgyq0eqncmQQ58L6DYQ8DrHCwH/OvGfRR6RDav3GTmAda7x3lOavRHsIvIh18sFTBQpD4Iuo88N
ao4EZESf5FKoffp57s1xid8GbP3epz73Rer1YkUYldEJ+w9itWgbkxmb2bdGCgAzeGsY+Zv3YwAE
D6ne6XxTRyXoO6tWQsHCgDseBzBTnlNlbfUO6HLRoPwJ2RdBTqKApwv3v/zTL+VWIxjAnsLSkDWm
TLSFwkLXgIxUjC48++8BXuCBCcloHAD7fDcWAEO1rs9/7Zpq48tXeBe7yL3d2Tv74qVs3YkWDz4D
98+RnHTrDCLYASIh+1xMRJEO04SQ55R489p7ocJcfkq5sHsHU/tT72jl7YH/Jfu8jqkCOPs60sTH
VoVeiJ/6CPvIbIO+5iqpRCIfhzO9Kk6gtZphfRkKjed6S97j5Clb4OEljFH4XHHN9rfzBsho4BTH
iuU/+rQ/L9MNd7WDbIuu+V/ItVSxieR5oPcKkxitfhI7Gj8ndnjHvkQ4APg5g/SdjC2yve+/5o11
eeKbN0xZ93YYcTRzdfdM5HfhAWgrFGEsCPsRWoK/1rxUmYzUgpLpNxu49/eGxaNR3QXV6msijVlT
TnF5DsC4nV7QtU8wskiuxbpTvE+Vt4UAek/RvK81qbPNwf9fE2E1zpiOCQMEZtYWxzlAPeciDKuR
MyPyeVjbgIYGgDgUdxWxa8jHmjeVjxaiTRBCoDWUBzG7ofbaI224lQx0Vt3AJvn0yxzS/YolQDr8
RUUT4OCDhxjinzjU4fAK0rqcjYHArfpDzCHlQU9d0kpKxdOwdIzeWJ3Gl3SNb+FdpWBX9A5l9Ivb
OlftbsLCOh2yBlqRBjEMNHjyBpDNrO2VRxdRV8InWVcSTwnji/1hSKrn8DgaIz6IgTUhfmBpXsN9
YX+xRbj10otaCWBhBZzYlYlJW9C++6y+pjiPI4ZgW7zdIhjze1kfP+8lzWixBYLjNXfr3iWx3dkj
v4+Y8FLjFlp56c6FZiW56hGAg4uaCRpsztT6bN9kwl7yzQ4FAEvoQd0MUtiniiaM+uPRoxd3JNbn
9yDrFUc/pE5L1jeBpz7OTnlHrwJD7xhMQENm4iObPyRmNN5WSdUfYCibvN8WKjxDWbWx0J5n9VCu
p+qmprrHLgUXKWsRFGrpdA54PuBR9y3Y5ZwzzWW2K8P7huBXdakrGa72JUwIvoB4M18sFyRWkH17
297pwR8NdYx22Za1NbPdtELCzeSP+rOefWG2/JutJg6SjCs9lcuShWnn7iKHNQVBtkI053CxkuJq
9YxjbqDlTWrwyUoiznGUZ6g6ft4HJLgwwGv42lVsh7IA+ZbowDY38p9J5JJNJTQI408zpMfGX4hB
jP17sE6zjc4W7/RV8ud9gqq8z0lysr1jsATD/I1WaLQ/ikxNrSdIyEIvpXng6G1E8B1CwC4z+vZS
Hhd0v2GPZhw+D+ggcL4HJEsFkmymCWbsAOpbjIuLIbkmbusYLWC+2w+MGhzcOQfhbQytheYwugGs
Zm8+7iOjApMxQp/X8YYoX1ZdWvkyBj94PLRSBt5Z+oAOE4YJUQHpON9r2l8ewKIdCkPzbmf6KQLB
1V/2NIcFbJ2Ipjm043OR0SOxSuTAAf3ctQKFjpK2J8bo87XGWXtS6F7Gixay1HnlfG7xroiejdWo
mch+QUAb44i+IXXkwY+qltFfpuLbRvf9NEqGaKoY3ZoTt3WuPA/tNg/0aab/rSt/nfbSMnmZ159v
LbpS/6vVBSASUTAQSM4NPknWQLppDKvEFSHEXCT8kQsIyEP1xUTGKKhY7bRJDwLWfXiQm5RJ/8mq
h8/PsH+j+if3F9W461ulR8zwMJ/DQ900E/Qoed+vMyl/UqAhV1y03s1Ak8twvprhvEsajEqyohND
PUBX0DvIufYETYdKsyRuMsOJXDjhYviRbK+sHFl6IbMDdPqESVAaA3OoGBWAooMO36vzVKclFdeK
1Pr6sh56LTx63x2eREi/+gjgXSiwRymtsq78puSHDWC3OJ35lWetw9cprCe4jPSPn71TzYLMtV6w
FpeE9JUCom9HohqknaqMhrNoJjgXGHcOi6gm6cquKyD+FVuox0ikF6nALV7wuTncMf3HCHkjs/VR
8k1y1BDdEC7nNvN9VHeC6K/Iys3C9zu+N1re154yqC+uzYw6b+Ol7eRZh8MAoTL+x6XeEwLsDJt+
aUHxgA+9kXoRQp1ZeCo2jMe3uFs41wyff5PIB5M6raoQQDTUPI0UdKQP6NOgQQVxYFX+1hNCBXGG
LhZU3d+0I8p/8JGYRMl3l6GVROzuw1dDAZMmlbKusfaxkY92jRc9TxBrVtuVLP0kcJqnd2JfyEMI
Tl9pk6zcdjRU2N0AUdjD+M1y4nQVvX97EHdPrlFHFHPLmdIl6g+AL2DJzJ1B4QS2Pmh3bpo/QbRZ
XWju0sJJ94kyF1mCiHNP2wXTwS2pLLDGbYbUmqAiXM66+JVW8LwV/rplfq6U1RpNShdd3MTDV/TA
CXLZuX+keefZxC5t3vJe9puJ6FBJ8+dZdcks+pgxMmsz6kQjV1EVXxHu43gdlaBD8rUjmZuPuMg9
21+xGcp6nGJOzheWQQb6yIfPcF5BLWWfLvhDlukWBjsOJrLwmj/XF3fTer57KfippKr5FLeYrQqR
cr5IuB+yYef2ZgI70Aj/HIvqhi2bp1Pjx0Rl7jSbFsHIXAinz1XmsW7CFneIzGCwWmMyZVg8RRD0
J21QiXA6td5OFKvsjaTDpaHAncWX6EEP7LIBLMznXynBOpwr/A6QtI3qlYREgeBRFt1YhrNo8rXF
bFluLrE6o07PKZFfdq9U7k9PwGTSTaV4vlnTFQzlDPa947xqsu5qqp3wZwwq/C1ZedZCVRGtdmMx
VddmIcPpYiVzwxOxQYr8FUiyxO98aTG7TPI7xHwxKLIw1dlfp4tpsdg73APibkNtWP7QZBmrsK76
rh8whrHxB9ptc8GgmnXSQffVHUQii1cIFhh3fYfEgaDOVYLTkyQCAfDFxLm0tbRenOv1PiOCsQCu
IIiGpPG3vpM18+Vu5cuSM7SorLXrHmrrwRRPfN885R+W8tim7prMPaXxAPi53rcufaHQlU9nWyqv
3mF1KzuJNTQ0FqGZmAosSjtnHr8Loklny7vrp/d6zzyQFwIahkrJhtPgCoO74v/5eF9SBmT5hPds
UIdT8VmmZUhoUzMLi7h33xsMLCxWOk7qnqfzHZFCX1TSV5Zxw3ugDPYAz5g99FGyvq+xvQRrpYze
rt+Lzm5F3nafYxUMZo3px5a0BosqNwsrFGUDbJTEBUpNeN5NPvJDdI7D+4sej1bNFMwJRS9YgCkG
jshToV+IkkgncGyENxrM0AGkZp9R928Pl5uPLMA1YkVP1zEwV9EfqlsLif0IXGwu4hW76QbxzRrj
KwNxb/b5jctiVw08GKhV3wTUKalxOBxo8ZBCBVOrxRwcJ1JCg4QvUaTw7N97sZcApRYTYLvWUZfO
tznDNS915lWN1KsPu7XEEQTecvneZDMPt1wVuUd4XwxIQPzCavNizR0xedsbeZZOeubCuDu/AI8m
SdeyTmAnaR7JD3VS8oHrJxNYrv/jxWAWmFuRRXU5omiPN/La5PaJpKsscc3UWmglf9uKZG92qf6o
izCtlC/EEK/qwB3PAfcdTpBANxlW7MIBf62qA+0fAp5UOblXsxCu8GMTZiurmKJugR/ZPji3zjWD
6gaoh2w/6lJk2eyN2LMxqotP7PWav72VEMRAoLnDQuKKnOEBNujSMeRiwgM1GNi5XMpFH/wOuT2s
s2sh4Xk4aewIr0PBlQLQ3aDlsfEiQ2/sbSBFGj/xrr2z+bMkfjFk2sEYfR7HRgX96v5glxuBMsci
BneJtTGhzy/oTVZarlmG6oVA8nwc3vJZSWUJIvsU+CSEH3sje8RfUH3DiBnt9LOb++ueNBxbDaS8
VuxY94R6tFryoeIz7Dc50TiWLpVGATyKuJMDRzXCuC1joG7J60EG0o3Ww9oEA5tK7cPi+wwYx0oP
03BXXbErOwvEcvfE7OG9bdE24aBwYG6YiVpAumrCm58JYwYLBPrAQapGmSrLN5tb55b4L4fpjDno
VQOCkvIs5u+Gx2kJMJAjuTcpxVsmZ3u3MKrTjHqvDfz7Cj+PTyMmnP1kMKKTnZh6XUpOX9huIYAr
ZAentYCJpGAMbyN+1Dd+dcKWl7Oc1BKPW9hCnhhqqJhyai8J1plKIIEE6MxZOlRnt6YJ3hgPPHAy
vGnchSCWFGiKWU9Sz9J0XeqF5HrxjF5KL4aOP0f3BOw1o25gkAT0cWTQ4/Ca7yg85QKN0OO1xid9
GCHYpa7O1SrdysMBJoXMZEB25Yt1Jgmzi0aLM36lFmmnUiJwsLNPrhigoZe7t5Od8IPJewDVe8Y+
hOPHBgi1g4zzpd1WYqlqgS8NQiUPFbyFeTvoVV9+zL4YnFhYYlRd88XtPbyF9o07+ccyzoMhJ9B0
h3pQSfkkcmVf7v+eGMkhQIIgjF7YKlZ3dYTArciXwIG2/8Q/bvel3cOJ9REZWOXzxbtNs7oY4F/a
KzqlkQix9v54bXapVf3sTcDhmMoKp0vciTMjHjuUFRWz+OBqukCEIktvIbk3ltPvz+V0wRp3RkDy
QIzbs+tAifMeZivHc5+9xSSL4xqq+wAl1/enNOxvdCYAQ23bDbO8wJhWPDT3Kz+nczbJXTMaHOg4
X2bO/MjmHJmwVCax7iXdhdOHOGc8KhvKs+BbvLJ/tGpXknJ3hP4PzKqRa3Yqt5MhGhYJ+Wp2opvi
qa0eZG2Awakvqk0RFeFDQqK4xBG13DXhEqp4C03ahYOfuNgYsOe2I5v1563kmO0uQ+cLENJV+eM6
e8RMcYVbd4Gjmi6TIC8DpD2L3N/uUtdAGYsIOG71jH6Ll7/lLPtEhamvwHPhC5u2+IOQrW/ZLa3n
msRhGLEaEpd9PVd2UehSy2fyT8rzpyM+Jcp8rfFnbpyhUH/nfDzW+g2UpWSgR1J7Hp8042aWiDQu
5lVrt/ZwHOujY+E5CjdpUTQKpHa8iWKnzAR5xpHKv3DI0kzuYvUT3PTVndaZEG2AEQPV00pZr9M1
vqhq3KoELH+H7VRJlMfQJn4sZlX2aXxQKX0/HFJf6k9W/k5EIFZdN4Of9lN6HnFXarVPIeAATQyt
2lAvM3Ec8199zCxjQFUVfe8NIS08ZQYTOKyBXPOme0ojFZ5Zs0ZWKN9BDqMIgRPyAUFqtYdBbTxS
lT2m9aBrT7ZVAadF1gvOcGm0rqOTAhsHAvRZRmvueA447lgUcksFS5NAY/cS/rs1xXqL7r5iy/fK
41OIHT7Xr8Oc5YyHmVpiKzkhtDAl5ISHMMClmpfbHB/pySJCekraXRh7pVEbkxdyyGo8/DJKHwJd
4OcfDPyzRSj/54j4b4QlNMgosSuz6hQxY092OgmXW0fWa5jX+RIzfMtmWXqr6HQRge7RTU+kcJJD
z3b9iCX3ElnnnyJEOIBtA6jsEPs7k9yfxkGA+UZFHKk0gj27WHCV/jQTsd6omQWoVpYL4wAptj1r
bp1VwL/gg0xYzHCtxxbfuBlS91ZnRo3DIxnmBNuHDRt7vTz4SNtauAolU/o/TBhSC9IRJ98XY03m
tLk3In/H+/k42Wj8oCfBlFlqU+1YLcsDfcCTJZmar02hYCQXEi4A+nk3J3U4uLqfXbA8ggxsDd47
d9W7ggL+LZnQOTrlnX6HpnAgosCYcT2Ht5rNn2PQcyvYD1FDAdpB5nIjRY1nnHvbjB1TJgMYRZYO
xWJOWCdCMswOt+1hyBe+CrhrQBzq5ccnd8aInlP0cQlQ2lWget5p6A7M6giyrVNDCRKe2X3736jl
mZAzM+LD0Wq0QGLIqZ58/AfomYwq2CZvPIZ7S+Hd/dZD3WjFGfPCnDMc9NzGrHFNNT5Frplq0U+U
UiFc2xZFJNzEIkx0s+RW+BeesU61H92V1/E/EKJzQxfXjZ8NzO2Zv+C9+eRvPvA3Z/MCzW6sffOv
qvCRqGuNvScTLoPiL3HQgDPXnrJmly3cyi6DQWIcEzj60nIS30+newYD/CTKAErtTEqUnf1xqbU/
AJuKnxgBzBKTG2vq1IeIQvkWKi8uM9fboaEIy4ruD5sn6E5InuFNtDVXxzAJ5PfEH9geHjY7HIrT
uleuU0rNxMkBooDslEUInCvuJiko6GetfZA6UmulQuvDxFbHH5mBLpFrxUYtsJDq10kiBLT1XQ3K
53WZNTZBFrVW0R9+z6OIwai5aTOhShEOe65cMTs8qO/rWQLKeBOMT0+NdvK2rxgcbFi5IBs296FH
3EdqVWvt0T7PAXb5QUwzeYxbtVEaDftUaVQDGol4oHHfWH05Nh3BxLiC2ANLfoeRJpQz3cgqyCX4
raOi3aW2KIcZ7y5B76BqZjVP2fURi5MYqW8inNsZtqtcxGptEkvYLRBc5HQEP8lj2A49qMQGTxVf
9k/7IG+C8RSMdYG8E6R7svBw31VvOGZK0pS8enuY6Y9hl7cOkG89PPTdt/KPd76oh7DkLUfZ/J4A
q7RR6VbH/7V1TDHGXs5Lu1b1eIUOtCK+YbRzbdvYUdipI8KqQDqzfRwbGTh0Ub2Z00cwfSULdyXg
Sd+ntg6r4omY3kFiRQH9HoUusZXtz6eFl5DYEzKqRCYll1WIznbt72eAKCV8WEl0zmrSml0QTpnz
CWuUrnxkDFakTSf/jOVOm7HnnFG/mSdqd3HfEiKPi7xF4ijdXUTmZ8WcxB3Y0U3p8AK06DOC5Jvv
VtO+kaSXDNuu7/h2yga1mnT6pLE65phz+SVjAIhNZ2yT1X9/wGu07GjAehqrMUlvg1XpgYs5yAG2
OnN2fveCKqwEhjpDKiRA+jlTTmi0x+F5SiyopM+vkCxOiZW/VB44zj5CbBJvnAX0EKjsvHB7WYDr
O3EbMIgDSlRPrxicM5o+zD0HFu6OYGi1P/4sKGHi1kKyKh4hND2w8lX3QHmw7ZTgY3Y/EaWnnfbs
Bp7+yNpXM0LENsPrI+rVStN+iCh/pk8quxQAHPeLnJtQ8wZsZtEgLpb+cTw/73GHcY0C7QKoocR6
OqHUGK9Ed/K1kmBRwrDlrJ4JZBMkw2yBhD0iMA9UweVuBq5PX9tTXgo1fD2z1vpktwzeWo7Fr2IZ
avCQDWUDJ7aPdfmmf/bvFkuXeB1XFdQHpgN5bDcCrvJaikkGNoAZ4CmpCfiJnOVq9PCFcppT0+eV
TLVgiBUjYJerje2HbwqmHchzr/K/E9pWP4RLiEa1n9luVE7Ly4cFoFExxZPDNHZjMf1ROzbpryJi
sGjgLs9lxVz6vETwkDSkfdSJhBdqPpZPZBFEVZ4gc9c98CD2QVOv0xZgZXnexVE1LipyzlNODUKh
8joToemOrTKNOLy8RiqLo9OCqxPb9YhIS9IiJNLxAmlOIYNNFWEhFfd8R3oubsfDVsD6J81RMETE
0z7zHKWBpvD+4soExTV+CLpCjb64HW9zRuw/gjAXs02YPSdNg51RTgcRdjqAcb8g7PFyKtUHeO4H
dgWKxYfPgHWeIIcHzQQLeSpFnBUtzNVFt+zuVUkHjpZlAelu/r5+shiCrmT1p8vEJslwHXbE8azv
UqNvuSI1V/nK5mVdDsEWwaW+KSYrztgiq7No302SxRGtfLiu9UEw+vcxTmb4eiqdv17SGsPLfiQ7
1r/5XqnbNSkQeu9Go3Zj/QUJHOJxCTLWV94WaQnMeCbCOWMmqly1eadyCWKg4vc0CY2AsEdPqNU8
UEwzDqBuag6lfQrfGK/i6uqw+onPeeVjxilSqe9z7Zl2GFz9ovTt0HggBP7BkXePWv5lHw8r5UW+
RV4jXaydzSxH/Io4gNkwo0dDGmprbcn1iUhXY6XcnDVl9DneA4++Qox3e4hJPjQtvqaAruBBE6XN
OLo2i6YZJL72mm+uHL1lG/sIPiLwLQsgLFB3MJhKtQHDn2lDNVMW5Qv6cuL+2JvmxJIrOvri8+vN
jAsZG+cYZ5BHn2RyqwfL0hJdKjY0Hawil+e24URTFPOcyF5h/XuEg/7w0Chmg4iewHTQ0gRc24Tp
druNZc3XUfdse3PuiVzIyn673iB+QBUjx+t2oks0JjgYPzPJA3mEV2Av8dgl1pn7ztB2MgTe0hKr
HIXtLMfaRSPyO2E5aOXSzyAVnn/aeUUqMOYCr77MLJ+AnKt+DiZry1DKbFc/vB/c82GXblFN2wTh
WVxmDHeWZV/txyvxRAwT1s9EA4ynQvG4kJcA94Mz4yunvyKqZBd2DsWru8MLpOg9UXT0HsNOwW+n
DJb21TnfzkEChk0kMcv/hsatRkS2ccXzbTljXXlBahYfH43+lLtdQ1lUzx5I6h7W5Cz4TOx87r7/
0trDL9BhAbtDu267azkpdudjeHLZCCeOzf7uw2YSrjCsxfqmuqX3uM995w44X8wxFztIDndZkbt/
IgnKo1sl/c1uPuqXpPBTCCOrhv0DAjE/XJfgF88hTscx/CPnHfezwYbHvT9H+zHJOojYNRLSz50M
gp0lwrp4gTA/fTdFQs6FHc2HcTvriz33ISu3l4HtNzg6PnlDLnyqdYheVfvqUZ8djOYnDD3ATBcL
J/W+1wAyrgFMDXsvqIzMpmLbDg68qwgagEBW09abDk3pDwvMgWRBxzbiiSbPzWNqSwUVwWTEX+Id
A2kUAlBehnzoyapRevke438Kv32VaoTc2+gYrLncHsjVl9GyFAiNBgwX945otSpBNPR1C9f2A5tM
IhNS0gOPydQ6byiOex++uNqNe041jYeiPyUU4MePe3YDBOxZaRRWmDfvendF7MJsm3ETQwo7X3TF
DsEQz4HdrynavLaaboLiflnBOB8D/l6+5Z9VAFCJigVl5SgBh1HtUifdnJoaDxyIJY+F4Swqs/PV
LtDTyXGTzkLLuVXzmsPKEFl5vs+lDIUPWt3U/FkbL9QTg9E9ZBVSjK2D9gzU2wL4zoOl49g8+gRq
TxZw80V8jkJWsTuRIYx/nRoPTUeOI+IyXBB3LBp/a1J89CWk+fAh6EbnT0aWdYoysvtGzBbysOP8
24KSBFBn4EHvhDE3gHbf0LN0S3Y4mrh5z89vmT6Le1HPNaE3jo+V2WrvjheSBzm2DKy/Tn5KahRa
96H8D0PAKdBDZlf/I7pVu4lHFXggj5h2cYUQU1t3qwZhbfian/oR0q7Vv2QfHvBUrKwzZEZBXbvZ
1x0pIwjqyfJtJPJZDULJ9a51kPpI4Qf/pWZ4To5kdwOOAPuYtTGGpRpYFWiuT/Dc24OZfYYI2ZDR
Fy3e/WZTwjpP6JFyN+FpdP+aoth9Z6iuWbBcW3x3Q5llsHXEg38tc98QQh8ijofYGS66/K7dd+MW
uDqOXEdfhUQfrVRAfnAO7qGaS3Sw2ydv9ph3vlS9SOVpAXgnym21gR/G3evRD8/3ubdzKtGP6iDZ
Hk81RI9MEcq/ikKf7uVsVhFapoLakt2cphHX284aP1k9pTjbosc59u31thPnECiCE1z+E8EOvEkG
7w8X2uhk3utqDbP/byD/PWFnp28nAdfVoLR79TX6cnnIL9kqiyYqAMMNZavfOgcd0D89MpeMuWcL
nKddqZg8SlEO4NSqYIwtbL5hAZBC51IjvdYtlbAP2Gqqc7Ogg5zLSpKC2dPMH2Ose5/7qEegW72Z
7HeaYQ2eAq7zkbAfH8Qd9mkUdB5YVPSii9Xj5Yd/G97Zl0wskoddwj2RFuarFFmXdRfII4VXRMKm
+wJhu3LANr8EbcLlvlKOXNJErMuwSdg3gBUAlvB/6VUSB9tV0WyZ1TpMsGU+1v2oCkovr1ES3IsS
FuoKL+QBcc5ClNLmG2H8iqE9fyGfx8FPal+99n+FAC/o/SDn+fygc+uz8f12uJ8R1rKO8lQB9D/1
vEu5grDm6RmJZNW+GwsqqcAJwFSQFWmfHiQX6RH2GhDlAPfjaEVyFiZV9jROlhJkItBSFMBp7qXb
3uQ6beSnAOP0BpjH6BAB10eScuGqfqGTomtjiJ4Ul0XPYzKKKnaSnrKEJ1C5nnPw919yXFDmrIPu
f8bGx25S4enkCvnFYx5V87/z553FFc/YgySQhh928+Tv3VPHehUfviuerWwcqT24zD0kPc1qHSs/
GxSNQuvJsiA4MGk0dkda0TzcRJDCk8v2M6ckbhhTcBKoV/kIbhKM+ExsFvVm74ZSeGjankc+4QKE
HB6xUkvVwnSPd2aJzyH8u0wCBhC2uzz1cGW1ibvEisO3WV8qCz5aNVEBVpNeCnrS9W3uFoJaZ2sC
XVcjAoTiIyW3ipO2dgkejpVBJWQEsbB45P6lvw9yBo2n6uqTUm7lQBEm54afsMA+PfZdWRrokfpG
Tl56HEqoPBOHguOFVFEcr9Wfnzlw1i5+2i7Jl5F//R4NcjxMCjEu5z9yWZRarV8JvW7JgBeOZ/Ne
+g43002qcFdye9zPWBWeUTpbYZpYJajtW8qePsriEsx0vBEyjDta7vvDJJ7nKoG6UHRuxZHXQr61
fsOpHAM2GweIEOCT+apNyi3A7cQ0VTt2GE4TtXS+q2n9JIB1/Ub1iyP64bAgOpqWDQpU3yrBRE0l
JaLLWfi/YvnQigCxFt/Og3u0eeCbZYAB9EN6YfOvJAtDCzGUkObVEBNIMkz0cPhN7G5+DaKs/hTR
2De2uXxqOc4ZAdzjh6FI9NcqOtVcGHkjClFziVvT8c0gfk7vD1/9rO6IK4+hsZ1A1TYip0ANls2K
NB9UtfWfwkfbMIU+7rqxn5+fPsxkhO5kddIP03uG1n29X9Mzin9adqQ9+JYq6AAsaRALAfjV+rFX
ZuSyMF6iOXJ6agRpU87UisILDBb2nzCN+FZeRnwfwBVK1fdhucQLLy/xOD6Tdr8XlHsM/pf2J/Qt
EPngp0oTz174w3Fbmlt+4d7MhaopQuZ6hk87hvmfLNj/Z1O/Vuq7LI55cYjZhGbyUfdfrOHc+pyT
+p62Yul7T4SkM0tSGtrMLIWZI9XHxxus24WTqQvYKIUMSkV3y/DideoK8UBkSQeFGIeEiM0sKymi
LwbW8Dl+nbdPzvLl06KzAwjhV56NzV6O8913S4LJMJ+ABNrM+l+Dv5wsRtYWNIUZkjsxveset9GI
d2zg6Ht40/UyE8dJQK7FMUQF8bhkLh863Nu/3AC1cZ7Y8k4LX6y3NU55ftYVqQWPLPiavgQMou77
ta2C9N2cNk22yGg8ggkL3TVFaNqLeIrUhkhCDyMUjDVRyB2W7a2HG9gm3+0bd+Dcm2tDeJSeJCAa
Oi3uZrsMcm2poraXmqsnREU0oOM39Uxoc1fXHUBMrWUds2lAm66rwmTqSzR+unva4Y3OkFc4irpt
i19A0VYY2S3yJZJeXHg/gaXwMW9w85lSvtASK3SX+YRmvmHeYSU8/67Lk4CTHriMhWu1hBKJ206P
8OFmPBvLeEj8zie+P5HDYthi37/RCMXU3ec6JmdiODjS80d0gGWJT7t/MyqG5zj+3QdVG+GIQeev
JSJrX4/poq1JyVWs6fUR5rDeQCmlv07hRlPpY29/vfkqd86gOeRunNSDa5thLxqwU6WaBeaxAyWT
VMUsIu6GC9ZpF2u/mfrJTkhcf47PdceyBYWTLTbPgTVmeezcYQnpKk5z69ubfSnT62fMYGaDZzB6
i9TLZdqEoW/pi3Qm0UWBGETAqMBZd0O1dF7oUTaslWORcJX/fqeIp0jD+OTGiLzvn1k98OGbKkcD
p6RjAPdbO2yzq5BeJrXVPejCV5yDKCTOo9CdBkgeVaq6hnFdq9VKqo4EIO8Os+EdsdBKObCL4TSg
Y4bYeHJGqyF2Hc6/j0psDAY/0bGQyNXFfTkAaQn759MRkmWirKffpIkt97zBWIltnzW+vQVRagjz
x+zpIB6h9zViTbGjqfdop3jZQFNBmSU80syHBhNqW0cbqLFV0/ywiTnoXeZz6uXCJrMRXYO0t1kc
Lw3uMGw3N/8vTn1rU+2IbwfC6YDpUHajZonuOyXbUwhg/URVk2lKHiOYvhpNpGX+t+Iu3uvqt2qJ
6fxiNai0Al/RNJ7rQUyD20Iyv5/fpxb/zGTdRB5pi4pkD0gGszYTVdnq1B8DFSVW0JE1MfajY0tX
cxI0kB6nRjgjIABBOscwSifnrR96wieGIQ/sgoQ6WX/qIetw0WO/rCRW+mU09LU7QWBiCFyvAQng
kJA6L6+sAeq3zTqT431O3kkDX9lEFx0ECK8CXjZU7TQNGUqB5CYRPbKuDykS1/DxnIEd7yw5Mz1z
sjgY04yVpA5N1X96tJfVZRFtlt3wK6Ka4tPf0Z6+ZjciHMGJbfrwuInOmQn9YKqWHFXLeRSXrkWW
PbnI+jKemGPOpS1pjfE0z8b4DsoCX/0S+YFEbYrwkn7dFCbibXokP7V02jDdNbFApee48KUKCBDU
+K+DyhiI/ueZBtRxxGbi/aziqLpT5ZsNH9UdF9dHy1GrVKMvTnv+3OgSbBwXZN7KP0wpgRmtvwq9
D55BcT0u2Qz2hj3T1Fjpc3gIr+phAUZ12pkwyjxjB6kVS2FncIKnuWrWe/0+u+3VCk9NI1+s9QLb
faNoYVxfyOGoMB2YM4c83+EfTuWhuGs7PAf0/PAgabKA7n52l8poGTTXtpS3s2PjgRV5LJ3bKzwO
aMM8faZH7YnnmWlfZKwNEjuWagUQ0NXcwv86D2vWtNlfRBgIyRPL2NYzPiGYEvscsuGyP4nkXptW
ltWwLSb1PQfFqdIb7kOJ39ssCZsKzcokMgthDDSARhCvV3/Puk1BrnWlN7pupUkInARmFC+9rii7
AWYPWYX4/yHMTWwvPgs6q8bs6zjyk/c1YqcYYcOhdnWuwJehn8uEIXe9UpxR1pdVDzZL+q1Z5udJ
Yq8TiBwkGwFfPlUFKMhYUyGOtBXjp2Z92BG991UYlD/5Hdd0gV6NgK1/aEq9R3w4YZYX7ZPFmWxz
Jw7yCiqfuJdR14pxTP/r0TzvEt+V+T3YBMB4Fq87T0Yb4HiK5uzRpN7qxzd63W6ZgaEX+BqARX0U
yEZ+A9O4xcljd4iBVqd5XWc4dB0pTETDGMnw6dZBgFZR50SNoxmDzbwHLbs9WGSqhk0cBdeDQM7/
3qnZhURqgkS4nuV/1/awIi+iT+Bt9fLvuSOBPv0n/bVoV+LKhPjMV+aJ0hAdIl874V/rafxp5YMh
0N+ieGfaNY4ycOINouYagBNu/0wwyjkmYGlFsLMF2RSM7jJTRqeN2lNhuJ3sH6qIQ+mpwiPz1eZD
VWQmo8UhAEF35aiPoAjuPKksuWel+Q4ZXGTFzOTzszH2iwA3Yp43Vj0qvYwBAOO6Uc2ngGXG3qGH
iwZFP2npeBqz3UJdk0P2e+6Xa4n7uECNSGGXgNyc78M+eWiUXNG9WYvGyEphwZe0HNleVgi+g+0C
YO/6LI+XGlSmRRL5mNv3TTFWGcUGpBMezKOctFtH/ATKpYGJ7g1qEmkqakgSQC/e/ommY8xX7gN5
GP1ZNvt/ZIZcim5WLTPNyHyfHlZgwyraNdNn/sVmxgS40pGUPnSh+5wA6aAM18k0igDBWlcIx9Tv
fHRY9VStq6UEIF8Nwh4CmxqKcfGABb9LpEDxwTUVMRPyFLC1KZ7JCe8ZCY5hBQHtE7tqfBk169IB
yB7lkZRZ0p2WQ6TvQJjhwMhjw704ff5bLObyinlH4ZdqPCaqFTHPq/IMQAbkataDEepv7gCbnQsu
yVhJq3UxxGyB4UY6aZgx1hUn4D47me3cggZaaSupkHWxVHjWi8D0YynfR2EdtKofKewyUg5Oek+u
IZa4HG/b+Mb1ekK+2QhkXrFmT38xuDTikFXx0yxEyN+KE3EXsCS3yhynzUGNiV2TLSmkkzvOvtix
/ZMgqyTYIDMiigygPzE6ypyLy0EwdxBWcYtrztVWpIQkVvdXUQS8Ht/A5OyXr7ZYYvdYBYx9t5mp
5eoSZZuND0c+EZH1e8KuTAIclA3vYG4TdCIB6y0V8iAWSKxhLhm6oKRUbxRv6sfkjj0b4DmlCqBQ
ULltFEtzD8S7hUsq4yCql3hCLq/vhrjwohXniARNNP65LbI7iZI77iz8f4xpc+uaX+fVmb7hOnLM
ZCBbBnCVVWjcrbZx/nU4F1Bzg0ubH3GxGVKDcMCa+MhLR8NPtyexnx4QW5bzJ6z0M7ejp9AOqy/T
auGJ9RBwE7gznuTSx7nFyO1U9hvimh5I26ZCKndwTye5i/YN8F9fGuMZBNAkPcxc5D7VdpT/mKuA
D97SD38fDWi8w3gkfnDjZBJaGjrcvkYAAj/QBKGdD4D2RcKrLc60KiE+GlKZ+e2rJ8cq3lAHoWKt
Wf/CAlwUY4hm/pWGi2RigLAYi2XPL1E4lRlP4DWF4hK4QsvFAtWC6QnkMl+fR6wyMnzMFBPyCoWb
dmhWBgIekMrpQOvZ8VRGO71sLt+i+Oo4s+CpLJBIz+bsZf6b/9/md4DSvxX3j8HPbTIeeAP1mxbw
BJMLXlCpFKMZKYG8A3YKIjlC0q8HKVgyt/ey3PJxL50RZD8ESlATn44q6aNd1FyJRzYO/xIUEAC3
SDvSN4AYmzvnweM9i+u3z/uo4Rvc0kKBCVTR2PUUjQT7ZMA4CoCkcHoYfZ5yDKKUZpWKKHoaww2/
vhGy/o1YspnqN8pVRmCP/oouCYzufFtFtSrqp2qbsalhSw0keyNKOAmIZinTKgce1bsEvf8cBXHL
FoN1oqRJwjp5udJGIueUQtJIzwv9WWraojh4em8p/1gUT5qP43dTiZLk1sd6O95H+bijf6eq66pv
d1BZXKlkAyM/nU1iD+zL9tFJ2vOr0VJ3TyOCk0s0LY0gqS77Xj9mIMQBa7z0y5zRYI20yRQEWLP6
DuZksTJPfYrS3Wlb05YumGByTXhXSfS514bwmlwYXa/9uTfvBEGQ4eWzdkkvrLhsgfEzFA0rJRBx
mbkGyWZeK0bvX9Mf+PPjiG8Rb+yi9M/tToU6M0Rm7G0aZeO578vS9UYUo9fShk3oMNAtK1xm6eET
X5q1eKBtAr1wj2fzj1y4ZRa5xyodan1JpxMfvG4pJfCPYRSHRhFLscvfJEo+4SD9CBpOUOdTQsMn
nLHozDfh/jBKJPx/pbZPh0FF1PMpuvi6PLgnPIy5F+AfvUgg1i9pQrT0/5eTuYdNbwOZPdheVpWX
/n2hKTmTg6uIyfFhUU4McuHwthyT2XwI5oe3w3GTv4AKsdAW/PbGD9wWtTGBCha8lH9t13slffCh
IvNMJzNswzK8kG+tcaaAXNLXMaECTnRuT1FgCUIW9xtAEC5cmGbjRSUOIkivspkJcLmXfM7Wk/4r
ehm8q3HmD9iETabtEquTwEse9ylz1tCBmONFyuNGWZ/c7V0U5OABFtqdxyIY1stL1GpttPfInz5k
1mvhT/3BUZoSerxkR3uqCudSH/9tdkhcvz0bxtKLWGP8BEHLmYtDh4oJDvj+XoDwVld/MTeYnUnL
KRJMetNgmfckLQYQvkG8lPJwvbVItiuwXqoTPMu3APrJWboJNsCKX61L22OBBoNA85bHqJp6yeoZ
7iqFhMaXs6MOtw3fyj3Rbz1omkoMfwOwa5YdVjTtXhxekt6PGgPtd6L8QAcc8YXX5N6YbdOU6YcD
jfWRyA3ToCi7sy8m4tu6fSkysxhhMEwh8BDFWWVmRrpiz05hOlwHnm0Y4/pDppezHwKZVOTiCAV4
kpc3kPCqt6DZYlswa+qCF6QPcDuWpnsVvU9kUwepm1zHihy15nxnseU4ScRy/Yrdq45Vhupin/o+
2UPWCDdJRb4Tb5e18rKSCpvlPqeeo4BfZeBLmOKLNDF1qpC52ghcLLwsoNpmwRvbxM0Zv+28G1QN
EbkM8enn2uCwK9L2rikC9+5JEc9NtJ+QFAOw7LuXGy1AlN5PY+Yc6N3WAyXnFz5vbaBU96P2zjf3
WaKHi084MhnntEvJGTclO70NgHXXglpKNWbWpDzuzuL4tMwXJFlcFK2KoJ+PTKDiyBM+6pWxC2dJ
9WSeEFnGv9ovxdNN1dgyVzJEoMEKlRTWQFwmaYOzNrBOywo+Nd+zXlrN6fZHPo+Fr5jwS80TnxVP
pRXiZsaEUxLxIhQDk6Q+z5vrNlNgAOR5l7HFNW3IqMlVAz6CUpeUf1XnzHS1CDQiNirVlBfZt466
vTC3+9zajb2AaV524p09WtioNNqcrdkNd9Ifk1SF7q0Vvo3NwJCjM0Ocuek4SQWNvJCJ9YAkKeu1
NdRzBm/QttNZXkU7KMhE0DBqqvlXcWr3OPtmV1HUW7EuuF302nqTDcvyq3Y386iN94G9J/8ktqyS
KUDk/nx5Y/ulflMyY/H1WtvGVUedoGr14Ci5CGufcr+SlRvGa/1YE5SHZOWHPZ4fQaoQGoKeQSyn
MQWWTKhQRLLcDlPOjEjgsZLqsD1NPVsiJsLLpeX3oZTQ9jqLkClAjgekL0gSCKW95SbhBxFTLfUI
yPd409iT38rX/RIP6+F6wra0xlJbC7UuU+tKOVAJijRmsRaO0vm942giQE0A7YT93CpnLWiSp1Z/
/ztDG5aXgj8vSULT5/Jckvu4IDG8ibItBQvjSj1KEUbgzSA4r2hDT3fwrbM8m4wJZ1ryrXvpyoL9
KDrg9FpeWXZWFd7EeiAikashwAbtfMtb/LoIUZGhfX64pu0Y0STE+GIwU7iGC7EYJpiGXJAeOG88
qaRQJxxbJnV04QPtsP5WOZlXsLZIKJZptFXgUjcbVor2SftTLCWj521LZT+fR7zONJLtzteukzbt
VWC6zGDtDgMGVr4qPZbL71ANbpE9MBd5NllaEgmEzKJBSbuYDZdf2/beGnEXDJWeyXSy7QQc6l5V
9bRkZAg4dfxarVITojol7FZLbTRzt9dvgTUsLz4BnZ5UT3xbgna54KtySg8CSQaJoSMfcuQekm/P
j/EM1bhQd/tJlOilJgpIvYHjbcDZjUZRI7JfQQBwd2xuVaiR1fELj1mC3MFBzYWGFvu+nnoH3eKT
bUsc8OoRZF3xZ0PMLValzVFZycPXXlmGY2Y7dLoZNFXd3ks/7e1p5TYWn6dI/8cD3fFESqLp0ORt
r9BKgf1RqAtz8AGCAoBkyZO9apoIDtU2D0bCL2z4ce5LIPS8eoq9PWFWG5IHv38LBILjeo3LohgA
CJZhO8slYa//ccIAEilcwDoMGzBkGZV6MzOn+8NY1tSCEUSVrFbxfnhiaWnqAiVYXxWSsqkL54SP
8RrHrkOZDGvwOgBrSi9Lvur5iuNIlcXvVa+o62Hd+uVlAOCNpJh9lLAm7/9u+eNPwqP/Ci3NvXbg
5lRaYj8dhbapiGbVgthXs64W5hkwvD/qPe6cxp7Rw14dYAQ3oj0/lsSb226P+5LhveYdkKP5P97f
sapwmf5wgbZxerb6kH18wIKL5u8ge7aeTfwNckaBxmfB7aJSZxGJXaEfAYeytKlKtdTQ86FGuOGv
xvgsaEZnPk75xT4DXEu5u/gmBSRT9hXO38i0Y5UFLY3wCv4T2AihN4cYEtVctwdxsJauN24T/spr
M7D0/d83rn3imUpgMZ6/ABA/xfGpqyevuhD/qvAeSzYyQKOct5gyiqi/a3PsailcFdMhiVFIXbEs
l2hbFg6LaHz0TkpheG1fdvSAzg7jjO1YV7Ln46Hks55uWRShJb0UOnBkad1ZjRxZUL2wgav2LDiw
bOGCfGeGxC0+U1IDXxJT5B40fSvXmk+I1LPd076+l0IEWhn582Sck6ogtQxUHktoHHzQRA/fs+wB
Q3M71tuUgnpO15fd9eonvVj+PEXaNhM9t7Bexc9j1oF8TRkR9T9XYuJ+dkMXmXj3BCvgyDLb6WQ+
qUM+E4hhV09YuEZ43ypfq5pPLuKduSQNXGNvzxed58VwWUSE5b6d7gaWAEsUaWvQRdL9dAfTuQ5a
R21gLST6kRkd9mt14faRN7AXMgjeA+veqQFdeWlhB4tKRR+oT3jLqjU9UOFCpXkgVO8jOdsukn45
B91E6j07znOqr8CjY6ORwcnA0SZqPpNnSbCNTpn6gCmPPwnkkSHhObo7Ec0t4bqMGtYDa+OWiibz
86uJq7/IAEyAMXe7koGqTxOg9rvwu4hAE/P03dkDgVfU0RbOPH6JcNjBrk1jxa6snTFn6Iq5R9LL
PPgx3tsQUcwcbn/8AU7rnL9EMgFuXba6UYu4gx3K0UckVONOAjqaOrMf3LT8IyOZITU4v52dQ33+
SlcC3tfYRVu0LI+E2EPPz+zW567ADy31Fxq6vkseFFSzvc8xe/yaCJB2p3nC84xcNwLwfGSbnT1+
0JbnzaDg09u3HeZLCr2Iso0Z1Tgx+IJQHPgMe96wWyQMnQQ34uAaniXwXsSgnM5qgw+wjULhqaOL
0IgN8ZWQeCAbtEqY8JurN1CiftfJJP4IAqwYBUtV3xJRfAnENMhSuBMev275CSQy+HPrixKAICQx
MUV3RVc4xRBKHC/86sfmiIFyRLzllDnT1TAY7zJuQoU779+aAkLjBGvWEXySY09zHnCk4JfQNeyE
opEmRFEODUKyqkTcXfudaEodQlcc0Ql2cXzqyKNU7BmJ4qImjiEg+GVsgS0j0yrg9WFanudIRwIy
RpxYkRTJCf067M3CbPxFX6SFztx6xxVQR5OKyQlO2wSmlC7dJFCjqwjkavSWwf7SCNaA9ou3Rfdq
gGIvt86Vq+t7xym8BxDEd+U4G0T7FEO9z50okjWZj8P18oTMzzbP7FmVBj9JugIUBdvzu8DRxxbt
yIZA9YPTUEb1gWRf8Pnqa/JQeLmA5CxUI+t4ggWoKM4UaxjRigRlLOiT/B22iQfzevqCy3x3igKN
09zLvp5mRLVWAucJmIlmZ9ChiKPebhEXaluLmpTC7bCak1IILoLgZTqEGcOnPlb3P5E0VPVaqvHH
a4t5KlQsiVdJr3s/oiJPmgxHdUlZ1j0XGsQsy0zlIFT4ETAGGwUI8TUvVwQOqzBnig/HQURNcG7W
hFrvI4VJlZoSpIIDAai+DkSWFZDLjzpMhJAq9w7Jt6C7VvyyvXyLOQyxDyrAvM/a4qCOER9zeeAo
b/29Al6e/cepZ/uIUQ63E12jaZxlIlUubmugwhmyH003Upe1VMalGIWsIT4yjCGCnXx2a9ButKsn
MTxP9s5YuYMoApZDP+yM8hbwy0yUNgOMEmxZO2szfrvlvO1vf22LzigVHE46jC/2mCZqDlh9sIdI
jRn2IMJQCoZqURIzZafKtBfY9dJJD6ZTGb1Dux/3mTLT37JqmPw1JqFzN4KpaqmOVsZ888jjqWnd
gPc05lBbLDHvdIpa8aFxwvb0zNxXlb0MtS4kXr9mmjZBkvYxmNgdUfffogDa/BVV7jMG/YgbUy9N
IE7OFGGs6GLGgWiNMGcpHkfgRloYTNABPh478xXNoxuu/9LEhcjCDHViYcvTdYMyBmTcDqt3hN4Y
QPUq/EBpvkFcEOjOOy5Ixj2J8SjBy2BkG0KTIqavhnS2mPqRL9z2dFPhquG4Rc0HuJKfIT9rizae
8t50hZnM3qW1Th0IE3BwalKTm4+uOnQbBsUStYBP9ILt05wh9VrJx0gkzzIwhDFOW4Ey3EKucKRs
DobgxIUZauFVCoFRQCwyY77AIjUj1CJqVsmrChacagkiJAg2cu4nlgOfLu7DB5p77gdOqiIvLJTa
OBiQCgOhTz3RfEy31pHN0py18aeSsguoj1pJn0wSiLIRRL6OlJKrYcJlUTzPzx198SPXltBAEM6X
lC5+qVta9mmPwbicT4EbyMcwxrC+WlxyusbTQJsO3S3XAXX1BRqKNq2FbnrcfrVv1mkyU6kSZ3A3
1JpGv4qoVRjIrrfb8nMiqMoS4h4Fxj9aX7lXI6o7FJg/Lh/fTnxn+ACZQEnJVRzPJ3gSN5FLDHSJ
NnBQjkKFsgYiW5XY+lzTzVHhAsiflCMdCsi0E5zLymyOHoC96VhhJfGenWWT+yZeWlL1yDjucWwP
4BJ8BQoAAK0Vd4KdPg4Zcb8376eK/Fp0PIf33KGrLM5JkA28gI5jAvxBfMcY83Z1LeG1mLDjXSyy
muU55hMJsDjoaViDRG+bVM+zBa9wj5mFNXa8ozCauI8IEx24rOBknhVlFX5/2rVk3k6y5sNyYZqs
W5Dkkg0IZsVwJHs4BHQgVO9nIB9b2dwXBJdcU9x+Cb07Z2bddD7kMX5wFdCcGtjwSsioW2Sdif3n
Dngig7eNJKZjysv0qOT8onav92rcOACkuZgoPm3F5PKntxrEL61QYtbZVqqdx5HpNJ1R84hZ00aJ
3Qq5O/f6lleWXhcbGV9upvbc5sSeho5ksnxpg+HUxDy37Eh6bBkr8tSkah9RrWZ0K3Egg+jNe1E2
TGS36VZvLk1dCv7IVO2MM8uf/pCTWNBZ7uu/byPdwhmvX7rasexzAmHnj7l0yZg9TLt3QtlH+8+N
7WAdDzFGPprMhAoe8cYxLsbcF53GljDCnxDXTLJxKWplSwF/WP8ETI22Oenfvv1YJUvjf+8WcANM
oCQUUdj2v9rx/WtBdLHaQnbwJ+EqooNK2xZEGYrIoWen9DqYWmd5iACJbaB/Wf6MNPMTtvoGGhoG
dBxr83AwMbHGDBhnogGbNXlgihwO6nQ8GZ2d16zPxMQoscsYn4U2goWsiImnzfqM2xHcWBDZPzRi
KY7bplmoVvd5Z7jVA6NRY/QvnrAkpKbj4HW2lJ2O8SCl6xMCP6Zo3xsJgUcRbcnd42nJI9oGni8Q
4DXqPvZ6JcWbYZev8X/SnIq6cyfyO+9/T+IOZHRbNXuNYmX7VUmTb3CXm31jON3BHEU4kMn81TFs
3BFFU7JlnUgWHJ69zDI3lnhoEAfGgKu5LawREzz4aZVqdMfPnlYn8ljc7s//IVfarWOUJmDM5w6j
mSrp3/AjCRcLRqmjTVfqzQrJPT/Xc3Z6kSi/TYMjTwdVFAYiu9Pa1LytVJvzjBdiAs0o1agagJuu
5YVbCM2wf4MQl496zT4UTD9GrP2iSQRq/GxD+wpvoLSxxuoynyOBXsszVuZwxsHMvJdprZpZS8rE
VsuMCUpg+YPRV+WzbSMqHqO++ACuJGjL0LHaafnUIyQUXdTuf9MupgWOyTjOiYh0AsiYIk+Cg4OP
WCC298dfeSPCLADIOLPHTfnFpTQsPlw5w8p97sdFOiPTGNobVmG9PabN8OZ0ef43EI8QQ1Fafu0U
IQcBUvg91OSw1KvBZ8PMPolGA9sdCVzRTAdp0zA9ewECfBgHUBxggtBfMvGzLRH9wdxdMETmc5o7
ihTnxQo4f5FRs0I5CN0YZisQvGSsBNVg/EpIbkYMtlActdwxN/p5CqQfMwKYCVWBLSgtTP46B4WV
nm73Q09joBi9CqWZtg4NcjKaSUOlev2dxKIQnRrfjDBjlGg7VQ/ETjsK7LTw445hYzgapvL+WJ4g
2kQaIOyxrJsYEDOJUE9iNHzmbhPJsC+1S2woL7BU3fA2tqnYgNnlBU/J0q2fxHGZVyarmrhPfyPu
mYAEsnRQzdnqarpBmlxAOneVJys4a2jcrvA5dVYoii3I9CpaQp4gMlYs5OdjSeiFvG9KCKDEZ1Jk
1S4Ew7Yb4FMFQWqumFs7pNP8kqAP1qpdCDxjYCT5J3P3FvNLaEkBm+FQr6WOTatygUkRJOsDILMT
QEaf00c13RtmNXyVwMUFAaYklr+Ul8cQC0Vi+HA3LrELpcOJxwR6kpJ9nRs6jrKDBPx0MECsk3ED
ViG70bgUkKVpQLvFpDSnMcn8Dws3fQTjOfErkKg6CZqv2kT6vgtXxXuld8Hio8cg5s/UyqH3Xjv4
u8yrQvANvEb6xhYsrdKdo/rJhX38cxVjsjmzNDDhI2+IoS4r/eXG+f+bnG/PfTM5QVyNza2Pxqln
sZCVAYlESFv6i66J0MuA5Nlx3MTK9SpajF9R69xMH4o6akZVqEewXDxevrvCt8tI5NRCWHRkcjkl
VCldRzLuzADvt6k4IIzeSabnejF040L4ff0yzH1lHiiqbX9aRHj9R202+KIawalZLCZEBjrBDSRy
CNbwY/RXM9A4nSsLcCwWsDtjrbuRXjBkh9e8kL9t5XXeCQu1Apm6XGJUPBN8OTih+i309EUz4Cf2
ivFf/jEd4O3WyhymGcfQCbzP/PfJ4BNXADBZ4mF2PEdhyuiNBdgoR8LQC7X5OI4FxTkU0Lrrjn1/
tG2iJEw8tD+TUu1XpXLJTLx8/0C0odUImgDos8wR/zOYzj0uvqu4BkJLRxqwkA4Dj5t/Jq2NXOXb
Pmzo40isPzLmSitpxleQxzlobj6+U4zL72YY9d1XNbXlsdkgzbiT2iAxOF0ez3cJQAgZycG3guQd
CUax38yIfVVGBufrk1RZhO3MGOdN2r0zncccR3yY8gZxcyq6mIeD3J8S+jJMRxUDQU1vJbdW4a5a
opMi7Wd4wupKAikkux1FKseH03LNceSCn6T8WLnlqchlaw6kWUzfQDXeQ5DYCuKmvT/DE1YbqeVY
TgxwXihvGG4aSGdvC3D/vjGluCaeqi9oD3JV7baxw3kBYfthLg5SA24eYp4JCRgifhewj39S3+oh
SYeRH+jsKWns+1rmGZCOToiawhES5idrYUFsj7SV36Ocp5NFXdt51qJxtlYF8B5j0+gCbjhH2RCA
OnDq/2aqNujVvhEJzAkNZSERAp2Lgpc4H6nvsB+Llw+2pvKVcUPJVUk4hFb6CXxKB8xefLybD0a8
Qiy1j7vEO72OQTsF82s2cxIIMO3n+JNL2zJwWEvgbIJi2CzknkQOY9XVVBpDZbC4DmCPGNc2CED+
bYCE/xVSyB/ZJMo/PTEnV82HiIk1Gu2kSBnXRP1K+fHVVYs5zGfo+UGQcu6cXjMlK2Me+qjl3Xhj
Cvqi4dzZkEqMflFhKQLhzMKS4qxHmUXaAwTGbxB00A1sAqPpPRx0EbW0GLmGMnjqg/+rwNdRAbtb
nBDbmdmNG27ZxmgGZeKvLFITrc2kUcelXowSmoq1T6UClIrntOc14fyx1C5Wl0rpfuUY2MASmQvb
ajGNDkEBhFmNAiqRsvcqPfuj5JbJBuEdp1KX3cCWSyEToJFzaBfgNW9cwO7lGga10VJAE3xLSxO6
CUz9UG+mzU8s8uFMRKms7z4vI7QRgn4mdnp+HkIXHT+Yao3NG59azf1G3KNbLqWTfPg0IzGrS0mh
mYH+fefBtGyEvzi79AymfZ0iFB2qQrtrbojbM1g3mc3BbRt/4F9ivanSq7jzhM7/G5Ma/AiN3XfN
ddIhBmD4eNT1S67+CFInvGRxO2s7+hQRPJUcdA4h3lDOo1Tjuk+q3gzLttylbHwp9XE7NfFXR0ds
Iza9qmSWiqZfShWfV4ihoUPLqgpjjW1HiQiw0KP5nLwYECKnvhsingStlBvNHR69z/5YY8qaY2Cc
vZKoFX9zxmfaoxxeTpEwck2HiedG607aStRmQUFV1nW/Hy80e/UWNy6PH31NCyAo+ZjGG4nupsaA
+ebamOle/wKyK7VsxI9gxk8NuJlx5I/0X/Ph2Drb5Anr2CDf7+HCwhv14dBHoMPKh46bkeeOJXIz
p/Z+11FPB7eT3+Di4MNPeajwVrRrEUyJGC8pQyJhBMX3g3ZwEwJpRZ90NIoizt5QPLBk7O6OC36g
85Q/vu/H1ss3+C/Eq9cOv2Lcc02B7d1pSd1tzqAvWWLH38aZv8sgytIm6ZmXxcziciOBrYC3iHKK
eoOOBATo7bjI2M0N9EzjEXoYEF0eeizi7w7pW5B/5tzaoNk53ED65dwvRuJLfqiHoVTwwVssl2US
LEN76X1eRdChXPHlWsHOIJf8XJdK63dD5eGsvAp3ZIK8+Xtx5tnZRBhaU+gGT/pI5zrlqJET0tBe
wnLcwIEnA+Vg6g2ywDux6y8SEs6YOfzORreKXugW1G+axl/rsUzs2zXQHddTJ1rCrrOavJ4wdYF5
fgsFjMPjcji6voIemYnikNH7I+IIhUIHl0yx/5BA7sgdxKRUrMTma5kTTvEoMlRMNkrEoZGte9tZ
uIzaYsGtPYB3Q8bNwQL3I2h8JLLSwFYhoCeU/tGgSlIR4eUgBbOHjiv//f889RMCg2S85Zh55fC2
5V/V06R0ckvFKajSLGu7JRZ3T6XNCXZnN0to95btYZ55DjnLgMCbXYeCC+CP4PzXRP9s2Pr+s249
h7J90cnzphojUaZ+Ll9xwaB0ArWU8C+0EJMiMarJhaBpvI4TZkFNeYNNyBMJAk8JUl8FctIhCC5t
nrTvgv+QXm6tEu5Pqzda+p+8TOXtdzZNB7pXBugz/OyOCX0EaGOvuQj7oX4JVY4Hc/LIUxreP68a
Wq7bbU35sOON9UOwO/4tZ7JGO9h0DkUsq2Wef9HfyUtF9cNii0EnKp01ER3h/NaOkDpFoWluK7dh
RYkGoTRjfwBPwgBeZwGjHRHxw9E3B6kyntX8gdDB1gXfL1yvwNM3fJ6XKBmEViZQVxZSQ4knnzP6
YmOweLebqyUnzhsKl90hNVY35rvBDroHVQ/f0u1YcSaQnQnup85AWG/7KxxTiriVM2J8UAJRCegJ
EsxdIHwi2rlowU6asVzLlvI1eESNk2XANCT2Aq7QynJi1+oCRjqqRVTDLEY+uHzfM/SEqlKuy8+N
lcKf1T9AGFm8CeG+LZtFY8fID6E2g4NqT6SNoQvBgbUA29doVpJ9b3ecWJB11RzYTQZRtROaAXCr
h0aM7cuGtL7X6FiC9VIZE+rx4rIDjj3OM3hquNoxu/F6U2R1yTp/POa1ZkH5PbvPU3Rb0Z8NviDy
jd2bo6vDggnEAS9Vinb6jBxFLQ2jyV/BsjFxqepzJqAbvgsdbRe8t3y22ghAAhP4wlWFsYCw3McQ
SwqN/3iTuLnCniuDP3oCfefbBFn7WtbXeFdDN3AzR7O5aT3YiertdWg/WiXZDgqhUVk/fNebOAZz
2qVlMIdcPpepSDznpXjU/D2yEAkEfjebxxkC6sD2jmffz7z8wYMbuSwJ3EvdB4gJQivYFPzOP0b2
I9iZTRI8Gy9gdbBjCSnJRpw/d3tV8jrqx/89ZAHY1+PU4dZuitM1RvmoA3Z1W4QwU22eBB3s2VdX
4aemJCvu08FjrdZlqAJvWZdehpL/lt6zyno7fkO0GPsTm/oX1LIRZQGhM2PMrCl3kGCLXHvI4J7Z
HQyXkOrtuzYR8KPy73FF4cmACbyYHDfApyjpYDR8S5aX1nzx2w+fVxroZr7eK0sTsLAe9bE7XTpm
hrKCuY9aAcc4RRcSvJG2LMTpNHWq573IOKp0O47QBdLP7FE298rFFq44tEwu/L5pDFZ4T+XyjylL
D46ytqwcShcNZP/nNyF6Cmgy0kU3XvxMRJlK+rrgh8PtOM6arb3DQwILL0uUm462YLEROhzY+X76
oUlaJ1CfA0J+6Y6LtUhUvXBqTqt9paB8vD7ERyh27nY55cJ2s2QpcGXQsV/tIpgSnpV0wJlmdU6W
ETpnGb7y3NkM1Zr/908srTaWzWZRQdXGWkTV6jyUvGa6zER4P48/REHjZ8RThzXoGR7XEynnMVGs
guqpO1mxXvpwIc1tQtmLjyVYotPvbOa03NBM//Ixub3BaysS6BeHSWJnjs6F9QcUrkbDxfPpvzHt
ObaS0v4rlDHlQzUeQWcNMj/+C/3sJ6X99ekaHWhV47ec8cEzRpVlBrdYJ+iFIw3Hne2K3VyoLLxo
7S/B6dSEFZXZ/yBgN7epCL/Vj35AkSgHN6TidtvUhkd0FU9cdRCVmTDf7ahntoL0JfqkayqJzeIE
YNLhi7zRwVEBjL2TPy4Kx7p4PswDXMBP1OBSeh0lzksAV0mB3J177vP6iYt5GI4qak6EigGJrAJ5
3Pw05Zk6NTs+grDxN4lMatoWNTC4xy8R4eGUzMfBgosWPuxomE1kMWjW9ARliLO7hW/4o14JTSEv
opn36SjQLz2cgld8xXC3z1BXIdSb5vWn9gbBz/dg51hJRuC5ewpt1JWWJXrN+aGKdqB/2dKdfKHJ
TgDd7gwDVqAb7rvssThbLGqMyr7FgHBb9Mj3xXJLLQ+LNwb42r5Az3h46+lv13x/roOI1UtpTBjl
Rzpq39MTaZ9BWIYnKItkyza7dKIiQ03CsQ+3aEwMq2dyeo75koNw0vxufAGTUul2MIOQojRv9Qc7
KRKfcMhHP1yJuamzK2iBYrVfXrpwggVmEsqyjnRSWhks7WJy5nzRnMZwUGvZqdDsi1poCR5ZSJGp
3IDTvAM9XTY/geK85z/MJQ3yPIBwO00uNElojp7OuR4G9KHCX0w0DZDU7ZEeuw+IwVhB4h5ymrgE
kruQkfBf+thZ1E7dkw9/PMjT0zy+vN30XXLHkNIhEeN7Blckq8PL0rYWYja/j5r+2dT57iMKL5Ye
QfqsMkJ6m69oWva4qo6MTR8u3A4smTy25DUH9BrmLMT2Vip8ioFfLJJb2QfGXkfms4NisqfswLkv
EJ0tNUEnXiQ3O/sf76F6kG7BX4LagVnQ1f9OQ5x6Ote10iv6xvrjgzPgcqsNz8P0R/hXPAOINFYp
WWB0dRC+WDPxjQzsRh2MvxXtWt0p6qrbzX3PjcchwxtVfnRbMkCAu2zXIWqiCFVHxBCU67wRUnlt
LCfpO/xHYXHqSBVamKUAoayKr3uFWxdAR2+x5qOSCPQ5eU0Rhmarr8o6c6KPUWJyu4UWlRGycTPS
SkkvUkwV1DUQ7Y93Pt/BxWA4XSMmlg1Y9LBU5Oh1okcbP+zpUNAxIMd1CrndqltKWT5lrtPUW1Mz
AquNpcpCrervd9cKoURBr1vVToiYqUG71kABJ6juVM3YFvBkjlXUNxwXPkcqifGYsKoAfK+Fn3eD
YHZwaPzwtA8914mUXduoLuPYgVn4rVH8FBSQxJ7n7WTy2DzbGNER6vaRWz5BANukDw78UluUZlN/
3RHz4GZxFOzn+B67ijM8KwKc0YpuIootHqdVbsc7h6CsdiWnfb2xMg4hAvTfdhg6gtpjI2XTtErG
OR1epCO2dzN2SXWyp3XrB/tKzaGCSJk/J6xu4N8lJh0YosBt02GBRNrRJDmzN+rFjqIuU3UU1+hM
F8Sfv4rgf/3RjRnzyfjKj+pDkTNrdmRAIvlMSJVkYjTmRVdXuaC0y15J9mbSUqOp/0jK1h40lizc
fv27tP3w0yHLI59aZ0ONNBJfVK+X15B4Rd1NhnTyIcMoVcDz9FaPm6iEU1UveiR85BOsinfTHAbz
KQVLNIhZ0M4XZ3ikvtFe492e1HgrINsGuY47FBz5nrRgNxVWVNhbra+QP6jWVRuX27QLRG/+JWXI
DeBR+wxrbvBEI5nyXP2xND5SQqTDGYq7fWUpcSzHXEr5VUzB6qoyQFh9KdVEy/KJLH5zBKu1plTe
Z9dqecGGwA5b8BH5C5ISDbtrSstMFYxBumWvioiVri9bgrfKTLt6KMtW5WuDYoRKGeOdPHTJrFY+
8pTiBWaFqMHW9dpJDieJ/rQgQqaob9qU6Xlg+zVUBIVRQNQkZJ3ykXJTr6EefkOd2KZhZXvlXEYN
RzSFOTJcNwfQw6BHb5Ry17+/3YMDi+3ANsqtMYuWIiOl/yf969nHUB4aJEy+jKOA0LX6vlOv4iWV
50T9bAgtxR1Ona3faFN7XRUvKB2d0lX9hj8cKs/gRA238odFzl2oWvE8XKX9MRBrn1M2pkZ4Q7h/
3PnGGjsPPG5I9F83WolXzSnTp5g0pf0WfXdkamaBtino63r0ewcmxH+AXxPtLLmOEDphEd3aMqXY
6zHxhD5kXg+49PUGJaDqcqj7gAgqkkE2CHiNdGQCPVitVOycuT0KHtEHen44w9lDNhXv/UtiW0xp
WsWBUyF3UwG+RT7e0BeUznnQMVUHGlh+ppOlWh3EwoTxYJ8wahSKuaHZEr2EQI3nlKBvKg5Zp61j
wb92uYSWVTmzReoXA4KFMWl5vaPR5FKLFtes4FAHjbG1TCRpHEguZ/3I7a8gHExF9mTEvFYqW7ly
xDIWW67kudjCuvcBjp+SpDONO74il0A8aBv+AgRjG3gL81S8RgE3bB0ZPbg0HzLw7NjS8FD/rM4w
OEliiGe4FwcAl9ORI+EvXRefHSY8wOgxOXNvrUIJAwtC7nK54NUtdx66fVU7T7367UFKwe2Hu6d6
iAXRx1pJlKVOfkUc5Ge7cNMjGLaC/cEgyKoJGSa6Dhfu4pThCC2QuDd8ARYkcJzli4SNTMCxrvF5
aGi32m71ERVAvJixfDxpfXMNSpxzDgVooxSnbe/lrWyuABrlopqQj0ZObg8IsZTkOeTTFYl2Ssxo
VABHMl6relxF7B3WdLHVbUK+l0kyHnNCkaX35j9OOK47X4WK+8V+enpcZIjKEx52rITQzERML42p
BcszcJI+/qUzJgFsZV6OU/3Motwy472zDYimfZ7dG6jhUc+ZSH/vbk15rqwaciM7mg9tQ0104csx
7oOP+4PBg8/r6kzkq/ZOqVQdg2acVN0Qw9hkZR9NP51jbsvvu6iXfJyJ9yDxKNSnYEWsTx062WNF
00On9hdK42no2HJOHLCC8ARo+mZXzerqYDV5t2Kn/Bkoo+jxc1gh24guDuhTJB2w7DC3qI/TUyGA
QG5PSu/nX0fmWZ2x+GlX0v+k1niQ6ggoeM6xDDKMS0oYjmJUlVNuEE9o9hwCg+35kgcWciem9eMl
VfNNmSa2rwHADW/9L5eO5GqWeR56NrcfOOJSlZK3mmpCoKyjp4awAWrBBL0kpI02rZghIZ7Il0N5
B6aNuDMzCqLxpOCS4grv+nzK56MGDUKThChuRu69erQDJ+E4faL6BacvL0byPH1bSnUi8ELyTUFS
WWKqLGLzEmlHeXBCDmLcV6BYbUKbqR993FDbP/iKdrPl2Vl4ya1hs5QuIkelIRgp2xzA26LFNAeJ
chrzRRw091+qPTdo7V//q4OIQ47PF10b/QAHrd9HQmNnRFu+hpltRm1dLVptduM6AE57+aP7v9jC
ZF9qcteEraj5MW6Odjiwrlo3Ge8QDFTqmYrUSDHYlqIDX9ZdxPVnhOqnHnhQ7MvD915if0t1zHDu
1Q1lbAmaA1WlXTHO+oWHWymv9u6XRcH7sA9USg895K3k4uulwofh3pCP+I2GLdE27avI/Ab0kdBG
MBsqrN3H+eLv0GxheYsDY73cqExRqbTHLOtHi09K6OukILupm1ZVKgRFzhdCdx8EqEyBdrHdKZud
ExX7EL/iizHbm9WfUmQLpAZd715UOR8aNSRJGGrXzja0jf6mbxcWAPSztzd32b8rZsiDKlrBdk+7
zph0bq5FHH6gK8gI+nIyrMoX+ZLEZDGgFBeIks56O+Ew8hDGN6nvxE48Y948/eYFe8cNBpm3ZWRT
dzR0DZaIdX18BCL4aA4RE94BQ5VSvJ20SScMWlHx5MPkHIZ2mdV6svNxJW9KzsbHe/cuIqTfXUR2
xDW4MZUhKqAJozZ66gwfJZuHq1og6roUrxp4ODp1ToNSeXpPv9vg3HpUUscSJPOg4/dCEQUZ5TDu
N7TKnwLsleUgkWbGa3i4exfgI3JWZF17Wzw4FYYO8BXcbJsn+5yEbypBEmn8ATTKdjyQ80H3LEIU
a+QOXWnBNehpIf5Vac2H9SeOaXyoeR/sevgty3RKhtuhuxD6UvkdgWYtK3HfEOl9z9ozZM6w21K+
3qtKWtK7rHL43I0WV96yv4M9Z1Paey8nhvqzU303SKsbjMLvTmur82QOCq0sQyrayKPPfXgGnVHO
7F1ADUXhF5WXphpfW4SwxFUFPlIOFBRpTLXy9TkICPWSW6qTysv5DS9dzFTU6wgR14+hxoJbaLsp
JWSd+jtpHilryuxQZM6F+3iZOszu6awLXLno6HnAkV1vynPjoZVI173KMH1Z9geLGEnoJf8fcauI
3GQXp8rVy+QImCSbVPWRj5knQtUH3oRCj+OstyRU8o0zOiibxjaqBhw+t0UbAse68TF09YHnMwi3
k+0Bvn2Tx9g7FbPt5UU3mnmwJbUk9yndbosVxbGWTqipqb6gU1kmyqXzl9+l5QLP8NuaWuHbflDC
qw2RhdZv2gIyXewnN70m6eYoOJyq9Vx9PB1N59dPME93KdoPf4vvY+dBo8VVBZVlCKM7ZNDK8Kj2
Xk/2smQ6vSO69Mj2hNUH2OdblMRXOVDslRUvIUJcO7mZcGW/1I69xkHKBQIjPhZw3yCTNBnA4tyQ
EsBEhhgseXMbGh6GO3mdSY46Ng1eHD4FKS08w+KznnPkNDUCPCmBWyUMGgop5pjTX9ztTTn7FMoZ
8ojEwUaxBQhJHHobh6SQxMrLwSd49qcwLkzGlYBn0PPDM1d28nsJhTuP1/T52YAZPW4APTdRkwGO
r/7yXoiGbOrfx5NBwXj2VjLahD3YWbOm6S3p56EiXUzbOLd1lTH9Txh1lMnhO8hSOi5eDO9Ke4D9
9/hUAx4JjMiUNjL/xjVNMehiIqZCPxZ9lOftPDXaiWIDaQR55cX904tPVpWA0rN3rD72mTwZsM10
HF3AquZMbjRVDcNjoqO/QgeidA5bTutxzAl+B1VWid9i2PQheqks2nNDP5z5vHZieC2gcDlnLP32
CdsfRS20nndnU1VDywsdHbkczwQlavX/yyURgwbCD036h3hMhnd/k3KGKMGeSz9ARx3Hyki5QLy3
68f/frKT4w/QQBcGiYs9j4T9MoTK9GG3QKpbl/oZTSdn5QUlDU9lmH/ZpMAkQkDuwAZ9SDpdFztQ
huY8nc0MSpCZLEpGprYood7nsYO7MJXtlnJxxAVOSSmzjqbP5cUTgj8ZeyQZRmE6ZQ8lGfJnxIAE
46cojof53youvMFA0n9TG4vVbI5Va7n9mendPyGyJ21Z0basaCpAk/R9Wl+fNAoW+IAYN0PZnSje
GnQwMJNttojxIY4KedYNw785i4yUKXE69eNjn7M8NPP0Do25xXQemaOnBSd0DnhsXFODfC5Q7qnJ
F3noZP1oOhB0m0OwmXvfnGqT5kKksjvZVq2qsfvUkO8nsOOhz35WkBazn5IIgK2P/Ba1ouea6dSh
g0xIOiEKD3YYylOjB1IC3MqpHFzqS/ijZpJbCQJxVkDWre4keP6x10utnaBBgLn/PsNjule4aA9O
TZHBfmRIELQKHcOAd4+FwlIZ5yfWaBr4CBuo7gEWyG+mSVaDvcSG4VzOmIuDHYywAxzJIfdQCoqD
e6cKbj3rxxqCavpy0NQD6uhhlckWTaWNt6MVi+2gK8Pch6+ETrDx6iRmWDUrYzqgyLv+RjsZdkZg
eVeXfDvbheYHqw40uGtUVkmwkqWqEjpWN5T5EQ71txD3eeG3wTvkY8OEcKJ3+urtnWeHHmkrt0qx
tiJuyEC6HgRDTPNZ7xulRFHwl+QU6PH1ewNhbbRkS5Dx3zTFNp9IAeOP2WU4KwaJHtoeMZjL6HZS
7+O6ZE2y0b78R5YVZnZkbby4KZICchfCeaDJVD+1LF8B/vE1r3wM+R3m1jJlj556d3I94MOX9iw5
+sSS2ZGsQB9TLLzV0deGb/d6n+rhpOZvK8gUm/dVsFNsswnO+2DqjHg3I9Q1fQ+WNSgmcmhnX5Bz
ZC4mck81Sc4uKWF9uiiwkfKtyH3jl6Oos3nPnm2TFi7W/AxlcXNgxlxzzGnvF1WvTD7/pejdh6et
7WeGnH6uLheTmkMvf20a4FmSJ26Ss8Zw78hndoNMdPf+EUFH9J/P2EVIgE6S3YgkIs38bCw/wUtI
22nWHqVPcva0kERZGxAhHa2I0pqz3HOzasdDuGy+z+Aj1ucuqz8TrkduWFi1aip+0Huwpoj83teg
iyVt3XjtL0vkHgn1L+S0kAM70A9vQErfo2rkNEG/1voFoc+rkal3k6OnkjMMKfzvbi6Dxs4+BQya
t5/mZk7DaxWTWN7CQpbR8yQj/n+EgN7w3UKX3rfX37F4d+pf3qrspTza44qEzC272yocjOWs/lDB
1mBF0pZj9QxKlOaiL8HC59E5ivJKfzxkK3844Gi9/9TfNMP7+iYSw3ZNz9kMQa+r4vSGPqUO+hzi
MyA1M5d2GZyuRZDxeZke1y6VRDTudiP+26dUJhsJW2PKSmRCWU4s2Uy6zfZRf+R8UgE4WdNoDer4
cmFwOxGtC4dpChNc59rcqdG9gBq0sZvB5FQXzgpohdlV1HplmPCGxXJsAOW6aauvLE1jdE25V8I8
dhS5eQNi5bmYNdhxamyfGMhtlPuLaZTKgZrrBZx0WqYsvPqMkPyAos+x4/GzreNKT8FctNYOYJ4s
Q6KH9vbf/1rEV1N3zgA6rJkifn9aHqpKEba3ejy5O2X2+RNFv7urMvegQY+/az++LhkI1K3lR6xk
4pDcp2dF9q4xxQ5Q8xQm8cmFLFsed3Jn3AYY/R+9zo/5a75w9P7nAvhL1Grn//3gATt8YhnSPIHG
NLYmdmLPjutUWWqeFG8OuH5EDFM8CcffuYtv2fZNebf5IUKwGGEA6k0SHv/3jGeuU/j64Fl7X/iA
C2Rous3oNWrn2vow72Tb1yqNUqYM3hd8Qy/gaFSQHCp4u094lTt79LlQYapaUev/KL85cCvTuudm
ULiq7i93sxL1yiJB729YEJ18ob7eZtSdUDWUBcdVOEhNF172GjfxcckOSXA07R+LGYvrksWhhKBa
UEwFjl4pWxTuzL09DGiA2tQs48110Eem05EtOadysm7V8pdUQbusaxLxcGhBs58GzHO/Q/XZX+HE
pmhNiA9pWVAeCYi0CN+6craTiZP4B7a7/oTySQWJ9D5Zccevam2vIQcuLiO7sLPDSLtAisX3M4a0
QTDJ/TDn63G9D88IbSrY193ovyN+2wdV15lylw37n0OBsPkeWZVescT+kWMPAlAWDCVDmVcb8tcw
dIX045o676xo0nK6z++56pLehsg8k4vYzgsVjjDCmvyRPPsZhWsOfoboKEhvp3xgOStiGeyRBpkk
pYgES1+MrQRvHQZzNpKNvBXvSqgokMHK8Lr2vvSA82fcstO/16FUauRcsOyYWIjD0n10BUwcncfO
dkTsR7DT0G8Ukrif2HxJWG2ifsH0zEMvEngXhfs7VCG6b+NLd8wDB+cRsibqrCAmVwRa03lqW8KI
dCVQ9WYwFH47XOJUC6fufzKcbepwpozvQ7Zx1gT7toS+qT2Ff9x/npnBp3xbOWFUorSo0sDa6SCk
ftKibR52Gr0Am6vxsrr2HgWEyGuXyfkPQGDhhT/lvZiB3j7ZpPNCSBLercaKf3v/3ApBY+MNdgKw
2ONHE/D4a2v/Hex9wVeya51Q8AkrTKmHxAz0tQCCExnX/WlyaF9GVr/YuQp1zfHoeMs6QZMluSWI
lkLak7OfIgLQzvgeXHJQXQmoYsoOYCQVoq8kqqSgAHtSVIwp8u+A+Os7xBL9TIO7OWZ49ZMahipH
8y3pMZ8/h/XeEusefwr9TOswf3VJrU9u21ilK+ujyBqv+DjzvytzjRe6ryPczTX+M2DKMpCWLiEY
iIkj20WWXWZ02KghlWc/MogkdKsnXez/CxoxoVvezOvdkgRKUhO20nJ52nkHyoTy14PSrPAmpSbt
oPITY7MUWK7NpGnapHtOM8QzjzgmOFYX7VCouRXrz7FTb3xqUUaPymJWwLViEErBoW6F0j0lpdKi
6pQ9oYf4aAJ5xtBCJg/JC/EMc/MqKJ/NL2i6ELGHVp7qvSaihi15w+geXDtpTGoUb8fSPEBpTLNi
7oti6B6+rs1ZuiJfjmXc19iIMOBw/qswuqs1Va+h/1cO4vosxIdv/QlL/LmNFUwxosnL0mR7nqOA
RmevYsYMuQ7DxzZnrWtwBwTmyqITH8dTI9bvy7DVJm++1AbboXw4kPVaOM+CAOZTtChzAPpIbEAr
5/K6GA6nIwlmCY1uHSHmKR1Vt/9lhBD9NbAxIE5d3UVKoCd+dbpRrojZ+m+3F8v79KTm14cdgVOD
0tSz3Xbbs99PB99HbkizyocuKbSI9hWQIsn5iTEuek/Ig1/vk0bMwOFAI1xdjxoAxfAuhzFrze5U
vaxCskV6dAqbvFrPQqCaT1IMuM53Sm/XAWaKz9pyUTcNmeMJ6mEM2EH4g56705/RcreJmYdsan2a
dfYAQMRMijNs/jAx1I/wW/RkhYkyxtSi9/vLzM8BPMul3lLC8KQUlU62pNlkiKN4tHJDwQVI3il2
wK9OziCvW3YqIiKJLZosGkoTpzLo0WHexURetrcTZKGj322uUOIi6pgmhbGgICCstXdrDrI8EtYg
4gje+m1iqpzruQdYCDE0Ivwiqdt7gbKTxScTliJtXIWrLz+hvgNphV4J3Jw3VImm9VN9TBXMYbK6
CJxE2hwb+5LKTEop5FKQQBTlP/NegEZfda//cn0DaTRPH08fp5ViQ6FTH4CjGRHnabNegRDQABg/
WLZH4ebDNMOPSIIvVPC85xkquTREAwbMPXTq/ajOijMYQz5kGJycMlHcj07QB73FHI6mHKlgg23B
R/92xt8AiOBX/+T10PYAuNPrPgT8xH4a1BbaPSb5A+U32LIqUYSI8ipATycvvMpQzkevmHakOnWH
VkeMTDCmOqC2Vfuw0aXTDhZ2xxJfwt530AGZgAmC+NJ2DKWOhfmLWXMJIUze0eKFNcwm66RAISC0
Xnh5N2dCWdWZu0MEKnp+X73jeyRcgh8yrOZJ6RbvJRtW/pGxzq20UAcYJp53kKw3rTGYo8HY8DSj
buCcbuwQry2tGzm/xYsGBGYoQzvCMpk+y+taEV2MwkK9CyvOoidE2iYsZP0RR+luPhH+/uwUN82w
V1wY4bd60giBqbHr2q7KCXhV5lHCfXDjdIEg+GxiYqBu2nbOxD5JQf5Ab2zvglkJaZVxQbxGCvXW
hQPbnGnFRSwLlqrV545NH5e8IrQBAQyJ7vy7xxNKLzsBNjK8r6WqzXKpKAFWknUgouFQ+ZQLgDLz
oen/V56QoIpvTd5zCg4Qz3eQdWQRy1zCljXdauSYynsyxoSn/evsCtfWPCNNuHdOgTSs62UD3Bhd
86iXIb1zGkYWU1nL8cplIhLZSW2ClH/le2zZQr97ROpgEfFOV6BBc0K8oYGSDeDfMByl1/D++B9J
IQRbK3RY45BNQd4wmCHBrGXSNTPfJJoFs73AJokFGNAOYK95w8u6HfdSsOZpxEun2Cq8szw9fuDU
d9VySTjVYCzo40mzZfFAqF5whC8FYuZpaDi/gE6HzyuaYQW1etXTQJWEXMO5ZKNSBd1VfTF53qag
K5fbNrR95y91FUt64n2EHe6TkGDBT/ZlLiL3yaEElb8K04L5ussvgi2KQatmZveZOkhtcxQ2FwZd
+XBQSMYSmI9pWTnJj9m0Dhrmb8kPVeftkbsp2Z7jRQga+krWHUuz7vF8wbxK+LY+/XMKj3NHjoNR
4xwlBhgiGsZHLpdnusocwFOG32zl4NzcOKk5XLi6QjDHb8IKxSoYaLv8nCHjKZB1e97q8EdfUDxb
45FsjQnQnlZLvjy5Kpm0bgorv6b4MOwFcCCclHyIAVLdipbNLjn40UkfQiTE6g0WroZIGVNcBVct
/AE9lCWqNcubMWSU46ql8KcMxW7EGuwJLN471hWkvIJ8wjjfmbN3qwk9kE/0yvSf3b0Gaj+pCmW+
DL+97CzVt1IwtbyovD3hvyKbqt6QpHZbyQkKw5JMBY97ASL/yBGZ9xldMc1ynQMvFUiudRbSAMIO
K8XUy9rYjJOqtDSCsoRmNxMHf6AQiqRaLingBsjT4ibYq1Yh/kvlUsjEXLlMS481x2eWDCDOrMqx
/LgSTwSfctwnPfo5e/oGi1KBsRT3tk7gv6WFNkHL4yqNX/mzXX/hKpVHM80MjjxDJXjDtq/KbyOg
xp31QtFZY9YYPn7lqjMfmudJn8vc/1qvQtXtCuOgeYkvuoHxwsxwYOlsWi6DK3CUPYFBULcpo853
Wnv7AdrI8vvE7LH2UioUUd5XDnGGHHspLa3n6zUcgCX+69CbntlYqvsHiACGkRxlUsbM1Sw8/94m
sn/7UJDqi7+OtFT+hoGXlTMaDVAP+WQ2kBApK6EMDx16wV303M5XpkyKE+ZTJaRGcfAT1BOMAAhA
VXkRFtRJ1aHB/qHh8S9sjBRYM6RfBQfhR7/BuXDrILOrDDbymSKqAzM0OH/LOKEdhMDavIttyktW
4XcwUYhc7e3lXprrJdi9+4QOticp5WBnKW3UbtTx88W6i1OOLotQhMjePWXw4MHTOPO/DhJ5qgyG
UKWcTT8yJqYy2Yd/WygU7at137FlXZlrd/qeMokm1z91V5u6fybzFrI99PDRMHpJP0/40b1as7Cx
tzf8ohTtYp8G6PzS4uteXtkkEGAwrVojtaImYFvic7TtqAkyYLm6ubdW5q8tdOhkjYvrqS860CE3
Q8hm29Y1FOv07B/aFI4pT7FVu0Q/fHu72YN9tTMYgDFXYSKglLFOZYV10MhxbJycKgMgJ35u+3/w
AA35qsg2rhz1CmsDmfpFnk23VQFgNxT8kIgztLXe/fdTfONTuUajF9/Sm2lo+x9eJLm4d0MC8qY8
btKvS1ebOWDHz0it24OC26BIwUD+/4WmBKfGu5lw7F5QOHAud1jDidHV8NuNfl5UFcP93VoutkjM
ytLLz1yMSAkEeFbpnkOhtqWRrBoAyhZcfEjCEdyy+EWJBHnb+dxGBsS9O/UnCA+BSUcJCrxcO0yW
Eqw38tTorEvuzePaPs9blQWU8p9X1q0wdSTAUQi/24OXWqT0Jb5NZNHpRcOoYDWGaHR/wZZPjpUm
+3QhfCAiCAqMgIdNoUsGtXbVyp8imHOMDQZNqeYPX3Am5yH1J5MD2pDMqTF3D5PttLqMYBPyrnxA
sggkgSvkJVCiLgsbhv3INhX/I9xxbV/Ua2El9BAfmqTI0kdZ5i/AFjT3hb3zECpWAn9nlj3CiIXB
hauiBa+4JOHPzvYx3xF2Fs/HKaXBy5ExtEoLqGSKbilbQMEOxsIdfN6/GR2MM9d6H/67CfbRb1Tw
kmzbwafwyjhiDa577/YhoobufDFt86NtysCzmM3jbdiTzPP6745LZPkFGAP9Mx2FwNqCc2isP8Ny
9RxpxzldkeUOw5G9/r6v2b7nnKJEdgzDLMH27FVFf7vBUbrudRsYN3xB/qFtfW5WCWdn/wPU6Ss4
612uuOzdu0ICSfAdL/5F+t8ynmrRzUDQ5K1hee0AyoFbH9kVqanGvKtE+2t6hiQU/g65Gai1u1c6
0ALFY44swl9snZZN/vtjId3vufe7fq1OymOga9ZtycuAh+hdDUdd7i9WwxVgTqKYUtHk/aVygbRa
aEQ7X3gCt/YrlM/JDRt678Uw+EfR2yhDn1XjT7vnN9OeMRpN68+yHMJDx0B7SO+qyn8s9AxSPFTm
Atooo2+GVs3S3wOxDc7PU9vLS6PNnvCCe32t3/eHGToalHvyOwlZC8AXpk/AJ5cTUUocBeSuHCU4
09pEHk3GcYZjft2dGDhtfNYkeH7Agbvihk/49FKLwAsLllCUJpSykWJnzA1pexkh75/4Gmp9f8b+
o6vY1aYS31NJze/GpZsAkbRlY4TrvHBdNTbvwlDYOMXaOdwDqy0RDrf9vSZpmOwwBV+spKM1suAO
N6et3B5DPnekAGv7gjfpvNtH1cY4i+LJY+V7tWYwV0BapfF50vd/7yJGOPN4fofYzZmn/ii26ac2
TyxPmVPuMXvVU9tM6zxcvbKnEPMRJwXBgWnccnUuoP2de4P1SKPlVEjNNlO9TF56Q0KVN7CxweGT
RMi8YygyByIax78yTiTxJd7K6W1KGR+En+4mb8UHPMiJ3p/p4IpVyQkwJoyS+b7yul3ZCMxfRj7L
slOpvwI4qRts5AS5VumsNk94+M35rr/mhxri2Fmvp+MrLGK4vPP6LI6PZDcHhMIG6PpUVB28bw+i
dVGazcCN6E18tjWwFxBC4KOz+tWWw8Lo/d2LB70AH/w0bzTYf+kxFqZXbnfwmddZvVnYKLNBZrcm
+uMDusDNo/Uyl8LagRR2IHTqD0JOGjg3g7u0wFlQAL0sEjWVNVc7tixG+35ZTtQ2ARLM/YbiMLTT
xsXZx2bcpY68TELVvHrnSTJkdLHJQ72VbqatfCw/DIoYdPfZp/uC6LQ7xULMjXN7TOOSocSY3ejT
bLeQVqmQJaLUBAuoPIb0XFoHx98qEUMtaswQSKW96SmN420PGTyiUafVa8QBeGm9c2q0nEJFy0J2
vAHemSQ5pV/YaLM07VgSZY6+xlMRBc9L78QA5pTnI+hrbvCn8n+uhMyDyYcODwwm2iBupqZESbDp
m2tr+mHxhy33VavRFI5Q1tD7FZ88KCdPoZXF8mrRETYnFC/UTRvZgNobhHM/9GRuMf13hOYAuld0
qrmYMoTRumyId0mXeN/vEuOqMR4DnM9dtWofLEcPKXZiwXsPI2CY96RNTfhkj8b6/y3jJIqRsX4Y
iaoCUuRfrG2oKvuD/bEE1w4KF3bxsrQFrfiJIW/Z6QiGKz9vZ42CzMSeaTa34QNPzs1a8cwExQOc
xkrdQxtJwip+5Y3t8C9wEDmsV++QusgWCU9hB1W0qFauKPMUtzrgMFWPRPmXtotBbyqSQdiT6Um3
APS5N29mXUmhniZsrPW09VS4BVO+WEfez5Ge+A06UNSyUx74QhGGuKnRi9U1qFO/PCIWm73s0Dh1
FYO/UMx6e8nKR8A1zutxhW6MMA9TzrwgsDP+fXjDhoaPlZkr++qtB8Av7p9eOzdL7mel5M7bOA90
7OwhWvS+ZVYzzcHERJGGY2n1WeRwdbuKwe8+wfcnNWe6NV46vNytRIEuU8u0/evN8bpWm68H5wme
2aYjV11xXSwlszpHqNq2uX/RCzX+xzjJLMccQ/3TQ+uv1uHqeclkd+VQp/0Z2uJi58VaRUpx72VL
9iO/VHQTDd9I2jukYSALWu8lRpqW62icJP7rlvAXtnkHsA8l2Rk0Cj+NtumqWmUtT8pNQFaf/p4A
RqHBzNHVOTNk+JcevTxNGuvZVmAVrkLZ+lK51IYHxg4KvTafwWCn53BD99XzPm36hU76fek+Lfu2
kqZkg28r6dQy1FDJpSQWRFsTTn3Fkb8aZo94IexfbsYujHCr9hmzzuVPlZYfMg8Lus65vLOC2AsQ
T6pIYhLJ+DQ/UK5DptZ+8qZLL0fDwbGf4riDDn9ID6wFQLCCGEC+7b+IcN7gE1571Lw+PPDNMnPS
G8xMxL0YUSfu1XzM2Vru+dQH4At3riVVjfXelpkM0O3fei7QUatrc1+9za6SQOcnZDKjY6ayPTt9
NlzTAZgqqrZW0zECjETkRw/bMQr60LQB4YwvQCK3ba7BZHBdc+rm2C7MCszBRwZEB33gY/g1gHBv
HGrvObGuqht8mtBIZAsjb/dv4ck9S1lpgXvNHWEFG9Cr+XvGGF64km2yb6FAUOMePrnaiC+m1vTT
QmuueMuLOibdU3g/sPvm1vDDISztjlIx+CIJYYsUaO08lOVTMDJD3MOTW/NDEPuPnEYkglO/Q3Ib
ab/M8kFs0g04tq1Nk4PMjWZm66kTr7ZeWG/HpEABSXUzYtYYed4w302hOgddz44QbPQIFON080Po
L8kX/2ELlGUNvxSVlHR0cOo9vlOTdSJcgqqPlmZ5CZ6+ZVtn+PyVpfwbZMF+Tyko12nDl2UDvanx
Awvf20jWVH+oZpDwixZdg8pNNCsy4WldoapTKFDjqvqY3gGCHRXfgN6mZbQgtO0fb/ULSYHC7j5H
+mu85U85llYI13L3cHLi1hGR2cAXah4B9gtOyuCM/CXjIJwAir6KZvbj0zCPV5zJEPyStc3QRlyF
STWgUk5tc5BiJUsc+DT461UjDNzvuCV4etFlCiW1PZNV82qiVyOB/pzSznrIqcpRWnKnSNQDq6Jx
BWYiD3avhXirGqFEUZ56EutaJdVBT26zj9g2k1LSSsgBXs0YF3W1NYQx6i1P6M/g268FqpQJHFei
jsIP/PIGlnB+hHoFPBrCMa/1B0Avc+fmgRLZLg2BWxtokJoKMLRKwow00fmzXsqRDY+8q9EHUyv9
vb/ea9D9MgFVmSVAKxabcyYBI+qmzFg6ohjbiHK87EAz5kG0JWZ9iczW8KsPLni0d9VZ3XwngWhg
vRyp0aIZxC0Zq1uTL4KVq307RPNDXHYEUAb6Z0SWVYE9iqD8QYVyLFTTS3rJgDxS9YcP4GlIuME7
zMSkBkpR1ogAVOpYVZe3OTHJNVUTsaCV64rO6bVIzDxdBK4BovyMb02UxBhmT4//JifUpoStlzez
J6GDtm4YmxuE3ot4puhcFn3Q1NyFXerCx3rflMccThs+Z1A45s7pCH6U/0LGcZVFYucePPGYuqJw
lbsNrLldbsTJ/N57enbUqKL1wkHeW7RGmU5UXroT0IIc/e17Ll6OBv9dWWt8fu9ApOa5H8I/BeQ1
ynCGufIFf+3rr5iTHmMA8n5cxokWnNcbrRZnQaBu1OG177GkAFCdCjdseaSXsh7EJiYsnLltcgiU
mM5ENSH0iSKcpL8VqNq/YyfqG69XwQbihnuFsNSq4xbkBqg0F1NDg6k4iZlOMF65+Q3ybQG7qvCm
YHIGLYYCgnAPxV8d6h4nVDGV8OGSMWbfuYdnpaRQUvDtQc5KaGgYjPDkD4/kDwyN8aMrN3K2DOKB
+uSkCnWA3qsKhzAG9f5b2Bi6lxmKBH4YAEwXkpsjE5T0D8ZZe0TjM6p/6sJWnkmdOT4/yHA5zp/g
z8MIzVYhUWuGuFxSdqcoA8gFDcnM9ZA5MPusYP+88NSo+NVYZVGcaYC2hG4w295NebJfVXadKAVg
OK1lCTPuBsN2MTg/2V1NybodDIZR6n9NhSaLYX5bXLVyHWkgFJ6o/WV4n1ZYFaL6BLvywwMte8cN
kb3ZD5SYy6ld8vzraESMMqcRTC+23uoyXl3BVfooxGiaJa1363elIvmf4rqoEv5ipHY0MpmbLHLq
GWNHg5hnZGqUG/zQrGFJ2t32Lxn3g5YOl3O3D+KGYAKh7AlNG3FEAbjfJ0HT6QGliuJZU40y1iXi
gMAAX8xQHSO6Ib/4tUxGKH0XYLtYBQJJfZN+iQGg3uhWiltoleN14kKWNhpYO+tj1pocUmF399Yl
33nyJvoL6CgxXjGv5zPq7SoYsEsLVYG1/nWOYa2IciPUV0uFHmMe/NZYhMSaNrZ4QWFQp3jOOV9d
ZjUaxhj5ZBZyxUa3GXA0k/BmumI7SpMvSjlfiMrPAg7BWsIsmEkfmaizuF9TKemXMVPGk2WOIeCn
dkWVgGJQZN5KgRgWxzxu/larf82njs/G9WReab+nH8YSQmE3PsLzNKeBz5r2aNhfvkQr8Q4v81XV
dWqw7VWUB2nVYq82cZh9lmXhpH+DWy/ogNRD5Kw9l2P7bzAi5gFqxZty8el677gtw+HJTk972zMI
pFajjuxUvClap4qm+DxnBbRY0ops1SrLN6Jf7bBu8EeZtu9IOP1eagt2P5CpYOYM8g1WOp1BRJyn
iFxnTYafLr+F+u0520nijhPRQBCZOr1vcEK4z7xTxTOWBoxNV1zR2u4I8JZwRw9uAuBiGH8LVk9C
lyipmHRF467AOb8hRugf/iNyLKdlRG5c2IbPRaRq/57yD/+6zUqLTvz2dq4CqU0ylre9dnaIxPK8
S1WHS7mnAuBw38U8KcfCFn73SyyKaSekDeu5Ac0K23W4xLReRe0MsMh6nVjJZ0fYbZUH2XkHmF3R
u4Tk+yWPuKJW4aUB2xudn0CyVLGA8fjLqJ8u2ttOxAm9wF3dUSAQsUGl7MMoxBAY4wgV2CW4Hl4K
/n98h8kW8iyOGVzt6ZFsrNrlBfjBSm13MQoHuiOOVGT9qW7YCeShNL5qpr2WMr9EDAVJARSZtWm9
qPDY6zQPRk3eLNcS2zLbyjdJIbjrqGxFWnS6MUj5TxQK95yLHWAfjSCxi2bNGrvB/Pq/hv8uDPEV
lmTemC2TCXpyIaCrRfEsBELnUgwF+X9HWUSgHXRZlrz3B3hmAEsixXoEvysYvNYrNphSo0ES1A7/
mBL44F7P0h7irwQ2duUO6kkOg0alAArLuETfMmHuCw3tKT3awGQgfWjmcCUu5d4D48tXphoV5dqe
XLfFYkCz7r6rVqkDqRTvd5bQVPZIUHPXv60bmakMkeZ9OcwwLRCcKvU3LXB7irlRDXqq89TuoYJn
cHwruil7QzVjEzniZehmP5WgPxVUsWh3osNdB0xBTDl/unIaSrIh8p8MiIB/hTJBSwnqY3DVGgIX
XUHcwxtycPGpcRfCZabFenAqzjH4NkbLQKTG/3/hjuMUZfVhgqYRHol3PQyLMBqbAEiSVPeQXwCB
fU5OrT5/zpNhh3yKThku990v6HRfpe4B5fq9000OJb1sRwWMgW2fOUF2KqIMcIuHe+mG34aZYuzV
VtvNRFziPknulv6txXPUSNncyjN7qjjTfBBUxPJEb1UvaijCL+182804a52zoTyB68HT/HB6znKJ
qrlG8eH7YMMiX1rPSnJfY1kdxaz9Cl8zSTb0synmEp1/u7y6zo4b34lH+HTU3NTgWUvWLnUaXbyh
6wCKlS3V5fcXQljfixwupWd74H9/DqwCy8UrvWGNFDUJNcY3TDniz+s0DBfg6jQSzFPwk3W3hp+y
xKtKYk9W96pQl/AqC9od9o869mL9eqJStaoe0lZnN87cL+5BbIk49iPslLpekoJdhLOip95dPmK+
i4qmaIRqTq/WHDWtfxbuRnB8hTdtzWfImw56VOsqi/upCLxnhyVQeubgqOhISmAJXSNOYYELckDE
WOBGMahwhpPQlsZNnwehyOpiFnWaX0+mAP4emPLVd39gWcBhMQU2/5Zjkix74kGzcmyOPQXUE5J2
agPdwiUlb6RGyq5To/ma8hQRAjSwHKtpbN9MqmEY+yTKCoUXaF0VNvLZmvuiFUzUSr7XYi55AjV+
Kz3IeWa0609I27+5jTVAbzkGP/htDeNoq0Bpw8/Br73QzwzxlOQI4LLXGTYTWTn991maSvoqlRs0
NozX3owH9KV8LR/Cv2lo8aISG3ccTITmTk7NXouF6GVhLJdjKZyh+uj3uJi9vZU2TIOBR9mHlNv1
bgePIQBJ0wJ9V8vwHM/29nXoqmgSdxlh0EZ+JmzqW5N+LLZCgVIEUhoe+J0vG63EYg1hZbsAbX6i
fD85e6eUu3GYoqyH7ZvNvIPjMUEwm/Lpsdcgf7ewQnxO+iFoJtTEDYbozpF99zn6GHKqkPN1iG/L
jxDJyxarJEjfeVTu/tx7WwKI0G8EDEqL9ZcF6iYV0sTf+IVm0fdCTMfJWrZJWl2Y1U7jqOuNI1zy
Kcui3fbyq/y1yKbEi2tmIfSjCF3GYgBp45URKNlJ9ypboBS4+7XQUP66NMHQ71YHkhr8/X1wKxf2
Ap3bmvvDMwA+oIBcBwO8sPcpUp3yRG0weF+40zL20Wnu71uOBvKjVKP6J/vUvl3UKQx12MJgZMTk
zQh9JNEJVmvyGfazEhpChSd30IeygT60ahl6m6CoOOVZSrXPPsuQJzY+8EKADz9F7Q4qdGk7NVZz
yHEMNFilf9OhVfTmNcUZgeFwPk6MI4CHJOFXUoLTWG2V77KPQMljUx73h0VDWrAw/2Stmt8h/Asq
MIyRWVK2M5XpB9WL0RbjsZU7mT+TOhxfyZTXoO9GRWvDKJYV4EuuxaRKmpem0xKdXPCIkCZv/TGp
jw950J5JMuiAbuydi8CgtE2yGsPHGatsDbf6H99N3LQOrJU2+ydDQ83WWJT2pnU4CRftCotAyc3D
6rlP0gJAZX/MvQYsBRgUrz/UnIJaJ/zX3YjN6tmKJeKUh+VliQvbf3yUJj9daRGn1/PqetRQqZTW
OG7/mVRIlzLOUTJ52cfiHvvUUDpH/o4ErGCry8DJneKJ7NtPhxEagZ4SFGF5zaUuIGvhvi6i9Bmw
w2+OlZ7hd3e5FtLYs80IDgpSuXAsn6P5nlWV8QPCiC5CxyHqayBWCtqGNVJIzOmuDwWTf91PJlt8
XLbQBpzXcUHpHM3/oeceQ6c5yhWV0ktUx8dUjNYWPBGLw8EYz6sROJud34bpax3rVM9UYMDs8LHg
TSzQ3DENXPfg4oBckCZ0yWWAWHaE/HnAGH+sXLQdsBfMSMcj8Xf0qxMkFzfqdGfbOivjO+5LYm0H
00NDwHR/tzTuRLGB523ZJm6wz7ghQXA1ZNW0s8gR5/evJ/0djpQ31nIoGv75Nk/dTWbuKXaHZCoQ
AG++074MSjN0OHYH+Ed+Qrrsh9/hi8oZaJ/UyBEMI+PxCp0l4tvp0noE457dkGhOnMTYcvcfY4wy
yVu76oiPpcRkutWmuAGIZD0Wbo4WFW9/HGORYRBHfHmttyjzILOaMlcoRdXUKmdW5pvSpclLQ2j1
qnB4CjKWQ5Dj3xQuSEMbz3cpaTaXCVL7CQA3fGI156yeWX38yrCBk1WvqEJ/zFGneZa0HUE3RrO4
ZcK9nxe4oIoLRCguwjtb4/uN7xUVzC3xTd4bmM/DI5A/Kw7V51kY1bGf31EAt5o/JV1Hi0t1WMvT
bqsFgh2+vKDPZsfmD6dV4DMu4JAixaqUOGuhRW8ogb9J7+n+OlfTXVan97EIb4NXVdkBZ7n4BO7c
HSxhcE2CY+9C+TmW26VSXw4zWNdKJko3zZ7G6xxPS3zanQW2seM1Z/la37OYuvS9Aj424zpjajgj
zLkXgExAs9xDiLdaEy1mQi0aHoqeIsxdGxleg6wvLtD2BUh6xSlQRoSAsGCS5M8L0CfZwYkzM98K
LT3BUprXvLlBSjnIwMU03t3qC0Z30bPatW4w2bz8Nfh4qzWuVXWLd9V4ZHhGmUFpaknSIbOR8xxy
JmWaH2KGTtcBjUBeybFrQy6lzs2EBP7pixN5Tmt/NECfUHx5AaNwcknXCpbZ3AsIhBP38775FbPy
LXp63G0EZOSdg8HJSjTWw4KXk/qWD7Ek6kpJbT/Qbb276U+5wPRQu8gdWv/8f8ok4tGAtULZ0cu1
ZaKIsj3KyMn6AxudY4lDqIYkliTfaP8BwgNPq4UHuZ1RfoYq6ZGYE1qP8LkXy90wucSPnolYCviH
cShH5PH+k3ChS0jQPK82tJ3Q6U3Zj/IH9kSbjnPsY7Pu/PxAgPWnfGS4W8cxFGJoqhfhxz4NgVYr
oj5DUGRxcAPyobupWFRpwmgplicK90bFNO+e5om6Dq/tluKBKICC55w4TwxhlyYyRsbidIHY+k+r
sPdNi5iUAOpJuP7ZhrYQnNX3oXN2uhV/bQi3vPI5wqKRaAWHxvMlaLi0fHU+az6kvreWWTwSrR6j
IQnRVKlZQDIVG3AKG1ZxaraXovUDUiao2n6jBK4sw8OUclquXuBFXSLU6rRHEVyV/KmaDJW3hN7f
JQYSfV1mCc2YC5n72TbpRxFh4ewi9xitVYm3/iH0DWiPuA6oR+iuhD+/NOzMWDfnOZJQphOOYnls
mYJaFdNwGmSGkgedXB44+WVUXR4dh7iwDina50be6t9qs6ECWkc/eDlhwEXoBXP90IBpyzaS4dj5
NpX6YhEq+hF9sAtyHHpMZxx4o0MBGvtmBJuyRH834rl2dMErbdh1gKzwajOEKJMXPQKDWUuMVmun
sgMOplW7XvrZhbGiIANbJz7AVb+Ba2Rsit3QpxEf/LiTQoiBdB7FmmjmJul07z51L9HGBLOuGpbI
bGiJv3UfAlpWpGokImmPXOZ49iZwYqKZjoxEO3g1wVSij2ti/u64a1goBXLQ4mzq1YryqB4CnUxF
tdxUyvI9KJVNPxu+sm1OgFqVosu4NNK0hbKd6MIqaFWJM1ERz3dRe0YseGbMWy4O95OMNg2ly/Gd
uGdGia8+7GlUbfG+DWj8iGK8Qik6H7GdMUsKDLhRucJWHFWhpxXsQ8dgoMW/Jt2qggUmkphANOi3
WsM6mrUmZqGLpBi+HB7fjo1be9lMKvWQ/VMJpZV53OmxDkTYV7U6vyCOnmiN/meB2aXrjZXod/M1
INlso4tSEfLNSmwO/j+9kPEvJcRI1vLhF9DNQch7V20CovUIVxdzv+e9SouVjWcQcewPzfDVj3a6
P0ipY3yR6RGQvqTxrWClGzQa9dgIohO/wOUhDAOTq0THv5zt+jVol1TWpAoT6RtA84JDgT57hU3X
bWE6a6GBf8hrXM/73733un4X45C5TdtPSzS5ScffhWKdDWBzAHPugebPdYYjc4vEzKrHpkexk4Ra
ZIfVrzT+RS4fKSbZxFK4YzAJhjt8EQcMw5fiq2M/mZ/D2uJms5DmeOlXHzIKHE3w95HefYeFMBq6
wCTWGkrbCDEL4VHRlTPo+/W0vfCuu6qh+96oO2h823LZ/ltNnibcUKdaBw+7SikxHPo6GQEpBEN7
hB2+9fUrZ4qxGTBcgHCJ/IVQ3iAIK3NbhNHI8rrRDUtjKKYAjo1CHhj7ziC+nCVteOLEe3en4PBa
7X7kULeK20U1f5NS3mjexCUk/JoCubAcIXRsL4INN0LJfVFgvDxfHqTv8zm0MhpwceGDBe0yKFPb
7lyYNP14odYZ5QG/wPJS70GDfpt9Sid3icftx/gY7JLBMtw0vRYSe7reHCUFSd0msDUbzxsP+wo3
+5y7QTWGLLO5q+GCZ8Skje2ntH64/HSdgOCsjEHlH4fuUkhJrejlxGd1i74Q8k8lbLPTiVNLjZCG
qKT0iHUYiyP8ekwNE1RRqJgVDYcyj3G4C1tTvrewT3JDZMdjl7QntIOSkOJ/epiCRGqQnMczS0IM
7jGb/2m7vt3BZbfziU0uIXm/3wNyp1dU05KP1LWw7p0L3OT2Hpszm7hoGUf9vF9cw7pKu6uxb1sE
ca0o2kTFsFuqwizosk/3hKAYPfl5bH5Rl/l2OWXkjCUxND5AC2kHTVRm+DTArwRC+su8n+AOZyy7
3q66NtGbSD53b9+E+N4gongHTPX78IbP9STGw3VIYU9nyPNQ5VVL60tibNDQ9i9sLa3spULvsytW
rZUpwe0Qdls/0Y+KZTmeR0SF6y2CRRZM+NlWmorMD7hvPzYv9m84HrgPF1Ud1oyXY4/F8BEa3DwH
prbFsFjiMsuhn5CCMS0mVk7VnLk+aLIjYtfTcGM4tqlMw56ySZQ9tmtmV1Gruo94yPvVWlweQfHX
QuAx4t6DLudleQBEKtqiGIQFKdmqhXGX8MVlMJKdEE6QOP1waNk+30JDIjys0fQFD6eyTTr79oFu
FcUr9kr8UpiKP9+kUbokKmA2MOiM2TMquFdEN5iCu8W0JtZl/uOEsiTUS8q1NIrxElVJ+JL8xBG6
2TWVK3TBRP7ewnsk2HJEVlBUpBOGkg0H33sOFEPSKTzBJ8XwplbAR63Yqrci5RcSnZrLB+MLVvAR
sTuAbLhWlF4nab096Ye0SmI04ncF/Ek2HiwhQlW8o1HGNI6w6N3csn6eTV+0jgd43PX+ekPl8jMO
8u4bdp+tJOQ/RP0z30enMlK58qTtD8qz+2MxPxiYXIxHxXQfC5vKgMzdWT4dDTH80f7IxW1zoYko
cnhUGCBiipR2x3IQPkIXyToWeYrGsOJmYOCkm2cQugkG9i0sd4O8lGn1XXCQaylhpCbhUirU8i24
snVpt1XrIKHy3AcPyuQx0sLJCpmZPCcDay/hcpJlCuxL0HuI4QxwKXeD+SYysNr5BanYb1nt4pIK
AOM4TqK4warR0DuikmZrZSyPE6djQ3gSX95D5Ax0KljB82MK/s67umSyoa+kUemCXyFogpNt5DNy
MjpxLESE4uR9IAhC14yWFISgHaPkZkqf4tLVjeWvuQJZTl0JNEzsVXBuj86RDlgR8uebeCQBpt45
yt00KCCwBcVUpqPM2lWRJg0wozyOzw57zZKQlpXXHSMkBurcHRWHy3/5aURbvIaluS83RLNLs37K
lOcmnzyB1m8OeZXhm3DfNhenldWNgbpd6zdtkDeDFIzoRPWNJhU2Kh3pELFEtxc4wxVNZD6HmDV4
6Zxa+sBREitqnJms2hqQIlUz5F+nIgJVwHkrqT+sMG7GKr7xeEU++V7JMoloj/Q/Ezp6JZ7QjdfV
q9ptcxUmEtdCbTsumVbnjI0TXqJtUPiagxbv2TY39SaUEpktsp2yVZl0/4DoJz75jW8HFmrt0X79
YvxaG9BumtRRqMBJHTbBbeuT2LX0UOURyTcB9TruvoVh2CdffbRFT8/WmG5zQjouBnveMOvqMw1X
C87H0tSPh1oZXpEu7yuRPgdCOUJUQbeEn3BCqRaGImeexFT03MbW+aLbW/ORYtUJ4fuErjnKSeap
J+Jn1kyzv+8ozmjzBuWn10KI6JFTiHKO7N8cruAfHcGi90zWCw1NgWuRFNACr8axmi8g5JC/fYiO
PcwuxmohgfAA+cY0VbIrAeQKTBaALa9oYqbIJG3HbVj7mPI5RQX/yYWbiasQeNLgj0/Kt1hAIbxw
GFIh0hG4+DgNmZgpHQmkZXxeIDFHR18m7Dw4HV2tCclRoSaGKI4tFjn1BVWiTk85FYcecutoqNLJ
0Pkeplf1nDpP1hEU7vuULbjGxa6DoprA3BwLyA6tv53V68+pPJ2r9egHev/4gqa1yqD5zSxJXO4G
RjSrxp21Ae9aUOdJYwWXlkvMfrVUHGy9y6sM4D/3Yh8GXYyMQEkPrxfT1Dmo4y17w1uEoOauN1WN
tZ0X6Q3j9m6Ul+M8CKjg1O1skgdf17lmVx92XaurmPHy9xwRHseT4TgJx1UvYVq57InFGvSDkXjR
1fmZggddZm0SrzHXxkM9KZp5oKJS3jq8v9SUyDe+k35/HYbue1cbNZRH/lnuelwlhAAJkDllAdcw
qn31PwPFgT8971Vu7dBRhlmcmDoxOC4MbrmYYpWCotj31hk1oXVuNto9McfxacKwheWBrMqUcpuy
U6qm5zt7c67Ze9kwotZnUn9zHxEae6t63Z+pLsY9Jz++9kCngcG6cdBD+/XS3CmD1U/eStwrwXZG
87NZABKgt0iy7pIYDMaB6VNk908sTCUTHUDr5fvXKVae4mkZsOuVJA1hWg3FCs3LxkNqccV2juos
1FanGsgvOx8fpJCzW/K82XIhwxGPonQ2nEkURZ0nty3M9JAzuD6o4ai/ycongKD+DmmFEb7ol4AK
MCOIsj7bv20fOSxbX0RWLmwt4XZeiMjNT7K8YBYV3EjT38J5ShBlzmKLLuOi0zCnMrtdIggjlDKI
/vwLusfNlP1eg3pKUyGt8uik2YttyNsGXdVqukpIKjDGoCIecuZy4e/MVoHeBvN54c6EvpQ+fL58
fks0AajNC0XRzcNsW2cO7gmmrI1KH/W0jPLfSPL/dr4MgvXlClajnNytBm1QpjshHYrD7sUGjbpi
obUONEdS/h7n03d8MvwYhBoUmEoqEfE2LOCPcPhVGMYJU0eKUl1o3QP9U0MKzviiu4qVtvDIr7Ty
V1uZwuxKc8cGxIZwzcj26DhhIh8jzHk8N1TVDY0hzMZJf0m/8EpSjgAncJlbp9rPCCzdADiQgjJx
THwqNieneBeQAiKBRIllBMVziihUqXM1Cihrg9f77j9h7BozjVRDAauGLaEsKrUrMtxdz4Sjqo71
i6dZ/B/ikcmrq8af7aF4zqWFJAFn5sd3Xi05rXzE/uQsfnkYp0uZCc7NyNrpYVrSE2EhuaPTLo/w
kt5Zf0xIrHWCIQF0JFi4uWE7EBMw3fRV8tcRSehvU7KJOJdPCmCEIAvyXP3MLHyuqC92Hw+2Tb/F
hqXKCYpe2qqw/fUxdXDhLiBOXDP4Lj8oyCfTdvQr30mwqfcuk3k7sJLEO5npJvSpyemnUeF/Dxf1
jTLnJY7K1TERi8hWEyRHB5EDmKwR7RGvNV1l4eg7Em2RrzI+XSsrzuDVzAucWh8/mcz1VH6sc8aU
SVLaxmnekNBTNuwglpO7iimpHGc8LT/nIEC7JhBzLu55VQve8KOByq2YTEgtzo2juX15NIayXyMW
+rHOgKj1qjexFtKyA5N9ONEVNLLMPqMrBm+1cHOC5Ta4z4kOtyRqJ6H32Vadb9ukmHAgPSZZfn9j
Nyq6N8YW5A+cCDGwjcetzNfJRxEU363jnAOepmDDtH9DrzrcDqm3Ao6q0JHPZ6uJltBQ468K8krk
Y+xMwqxOixfAvdF6/vrUeU8LCDGo+Ba2MHa0d7l2gbep7Vh+8Qv0FOEJcrtbhYpkNe7x76vAq30/
OdgXyXez5GBlEptw3mIJgcWLK7YWQPixcZwdIH0Li6xN9z7bUr7DC/nsBbHqa+W0sOTi95ky8wDD
3ogXAKPvWjmZO2g+ruVRikZzhQpgSrOnZR11FmolSpZRKMpkedeeICqaRtweN9Z0D4fuqrMcttaP
u8M/F93PtLRLQZDs5nBArw24XeneLLY5Wa2tvNQ5YDpAGYCvSIPauohaMQDUrtiNMd3h7iXxR4UA
1Y1+RQWWKggr7HZPVIWyg69Jeg84kF0j/gTgdk6bpfFc5TBrJq1/jyz+jjfkGmil8gFUGBWEA13W
ZlNMda/O4lWVUS0kk9ukj3GOIN3OUkpFBcbE54s7TS4CEkpxoY7y3LXMq+/vNQUdcTlhAZGt9XBb
tifoDlrXWxUXrAdZe0U5fQBKQKBuNJ1NpBuFqz/T60p+wJ99UjOzR8yYBhQQ3cF286ZETGa197Bt
jWXcDJmwj+W2wZn5jQzLi+OzFMKzZO1Efgb0468/CZMo2ahKWHfujnThJTKVPQ+ksO0M6KuZChN0
o+OaJNmqiWBE58gchbsbLa6EtrjzZByzFj731rX0Jy30Z81l/7FIAI1ECh9CzxY1fXuyO9aou685
3jFS1FR3SBlnkTtp+hy8pU7MVBXlc0CVYUWzxpbMDR2FzfDdvnf1vZeIXFu+XXmirz6a24waLzmy
3rZ8qV3MTWjHBX/PUGBMZzCM9CQHD5ytlYNR7Py/yVOeFi9nECrVRQmrBkRDF8ET4ZOE9UCB3nZL
dFI1Een3X/nuqGIcUDhNTBEQ/gT7d5m/M4AMHtWyP8ntbwTykh8QTuU4PJWXEnFNkOnbYO2GB3u3
YuRKVD6DT4YAMzg2x1BSim3OWYNLh6lIsfNBMmbITwUXjHj1mE+24oOYdGMkJZLtCAfRDzPlTLlo
Rzc02m0uQd01BCrE256jhPO+qaU2hQRAoueD4XCatNPp/+jc56JAtWggUNmxF4rj0nnO1tOuQ2ZA
MVj3y2fHtNqP2VnpBTEJ84Tl7MkauNBeuXLMnaqVUiHLRua7EaFkj7nPWIFFX5jMUz+f/+3ECilY
+ltgFM4VBafsMQW3uaCtX/o8LD1LumsHkjASUUqrRWx4hInrOWmWdfrZfNFAkZlhYG7mJYcgl2aL
aG20aw+hfRAiC4gQPU0pr8Qcxv7f2KHF3LM1x6ZVhD1aJFyfTtwVnww77oRyTJcnl/ElSL/mCWEO
VfT7wYrupeFVKxVG/oRePTFMgsTrBC0K2CjJWOu7KA9p23MIcEE2YOJIQkIuViqBuFgKd+mdxfAe
KnDzVLHN5eT/eS2zOg1eNETiqMzu7YYy/dYe+uaEZOGwm+IQoyNu9CxlmcqlbUsNGNV2VYTjoCrg
Ixu1HAGfbQHtM/E4yUglHKbutxWmhWXAsrk9JvNw1D9FdoL4pcou16VvR62iwIWp+7RbTe5IbTTO
7Lbith3FWE62WErzVmSGsYlRxhLrHuDhtyoG2a/cjOmMMfrhf49tQyqlbRr/AuE5OFCaiIOWuPdR
RVh0E3an+cnSMCagzf0lx/QmM+em/KYwcdRqsQDSCuAXld0goBAN4wj3J0GH36PxtstmfwXKPHYj
y+u+F1VsoJErr2vmYcGjgg9EyOdW0XQjudY6TDvxfKGsfHgI1lBOEDHSAAKoV1W2S8IVDiuLqIxU
L6fNxghDUVTorJxxXNPP4MnlS81V7tGgFMNhFICqH+X8uaOvGNGU+xPlzU9KlwDziz+5SnOqC9aU
3vznedTnV1NRfvIvUiRzxAORIPZL8kjcUqHv0kQAqlxGNjTQVVsjEQ+8pD+wqK42Urhx+8lAzGZa
3+pAHZP+RyuIvKCaESQ4UtQfOLsgcbPXPVuDMvXg2D3oCJZLXZTZGqm0FT2aPMDGNT2fDelYSHdK
/5PQ9B8P2DjPQ/cOhPK8OdjwnN8tWcKQlh8yikHVTlm+GHrgndpa/llZuEzbr8VDa7UiWshEDzTV
gQCBYNkis4GF/oMSoHsaCsGybIHO+7QEmvZoB6D/ept6Nml0Y+YYmUyKTlhfXeQUTEpYbnigUGe6
4iGwqQoFthsMf9X5AfHSGo+izyt5oTlkXXy2P2K8d9W6MogxcZwu9yZCmwHauRXgyfR6IPjbcxyd
1Ttik7gjbkekzOMzljgP6SqM+RvR+uSQVDpcyn630ayzgzPyJ8jxstG9JduTgOmNuNkmWpCzu2VP
nl6d9MVIb/4Sibh9BKtvrQ+ei9k8vKENCwYOz4oKxBveXNgSlqPeDuYxT4Q15hrqkqZASBT8NkPV
Lj3+mGICGxqY9Ce9PpJH/sm5nctxxSDJ78J7h8IRjcnQzQ+kl3AYCepYLb56sHpliTNrYrvf5KiV
OGiCXf9OrgbpL6RuKOIrHpQRDuEI8iOKt8ZjEcJlRNPzLlcBOQ4+9hjAcTAxuuarFt3IZhn3aszb
eI+c7TsM9KRgunv1TCArfUzHebdhI5xwoDB1KZ9cvo5mMrsp2HD8cwJOMO75s80jzku1H2FycJ18
LjzDSKaKB3VlSteoF1KN7JQsiPsicrFB+Q6hzaRldNu+OmI6VU4wmfhLJj8Lbfrd3/XudfW7Ghmt
e8argpcxfd01qGSDBk4RL8z7Q3bn3jawZ5JJF8nwVgcppbddA0Vek5gVqcK+6YEPu3RJoYyAv7io
7VGifZtwNWVHqPdCiDAeSb6qMVGQumP72IeDH2CbdHza7iN7WbBpxtEGVzbC0LhTwTZIDvtCt87e
a0k1dmfsSAE+SpdpjM2ec0/Kx1G9WFwMRU/LqBO5KFDnTzlHk1brkmjqVtw8CD/KTseFhFITvJqn
Earl6pPuKQLe/N8splelqorsjvIiJUT0QGSKiUx0DjyiJseE8l39GxVwF1bWKizV+EB83nbzPWDe
9JWZ5W4T86EYDYRwHuRBb71d3FFnb+vGbt61vTUlz77YDLPm85+7iyDMJiHutqXZPrQ2RPn35VIz
EHYDciZFNvihrhAuE7bgLV7DL3XJQ7NxPgQbPqArH8gWFUb+22fX/ABdJUAs3BMpDviqQIdcIIqy
tTbQ/qOuXt0bT/qQzaKmxUCLchLbF3rgQ0oIW7lND9w/zui2xWk+DSZgt9YwjHo5ZxT+oSXo0iRC
J5+E00wBdyQkIWyCUEhvpzP2wCr7SzFNSRMnH9bGVpL6vDg4U5psGXEc9xB8Y1wo+J9mlGfZBfpf
vlSmrxxkZJwfcuNenG1hbnEBnvhjuc404LrUCxBgXVVq26GBZeuWUlV87Y6KGg4CIGtt2SUlDHa5
I0Q/G6n6hRCej0kGCX7cjXadv+2T9yba70EuGzDemC6TMq33+jZCmtTxWrQj5WtP7uNeIp6jvPwP
f5kd9vzcR49ui7OioSnL6bYs3VcZaxP/2WkJLHZct+6GrjWZcklG9GKkGllAYr7Z62ORhCDZfEqp
1eVKfC/l62M/6ULkdGVEXb9yTzWPj0lWYnPf3ogH7ul3zdvCsrYE9QrQ0vcTw8Tv6nnn0k8sTVe6
wXZfviShEC2yqNrvOdRcPu4tTQ4/GHXLKYsCOYkP2cc96L4ZijcLI6wkdGma96zand/uHbb0dxqL
q2cOewMEy1q4VptVbUmu+IKO2YmquSTDdJAEmsHx5cQWcjdL9rTwt/2NKyMw/17YLPz0jKZXeglW
NT4j0eRrKWwGIPSciyJSzR5sSs77jfYuqvVyk1N33NOF3FCgDFs/VQXAHOIQN3goy4kFO/udE2SY
VYVlHG1O15ktkeWx+fuLjQhdE8UjOJZgulTdOqM0KnL1rVqs13OClb96wuM4sz1prjkzlvuaY/Cv
5AYhZDV9IKcPdprtmXWqpXQlWyqdWEL9Dbv7D70ApObRv4ajHgZTlSfxRr1G5dulBAzJkgLHKaZC
lNhAZlxfbs9svdda6OMBq7LzXurRrG19cwL0aSzsPRD21cOMTGz+C6LUo19wHoYGIjtMWGp3kxyz
LL4dvC+sYRE9IEDNdAEiIWVc35kWZHw9DSxrxsgZIp08nAzl4kzrvHB/rL30GdFobW/Njp5u+wR3
5OPcMiiBLQzkFDYGQ/N3FVS1bT0KlmPcue2DBXbUGDl+b2HlH1fQJQ53TIgizE/j+ZZgzKzSNrol
9qHFPx/JygZ1oAWRtDModzXX0RdkJS6pFvlh5NcKgDLQBd7Q0Pcc1YMvlTWuS+V0dmWKtiWxrty0
kOJKHiB4IA3AoFErpwSqhCgR0GjfUItx+I8m2s32ot6o9fL2grJm0hQdgQ7vcwaNylu11940KqWT
wt8LwQ0vXz5/6YT/ve0hISNa1wApcXdOtohofWOugdlvXOzoGJW0JyNidWYBpfdJOQsIGhu3e0SW
JED5AcPqYQgIZRWmMKvb9sngaqAnsSkWxB67JS+lj13SwSMxBn+YbHfYNg7b7TKgljF/y0kVlqWc
cwAoCGE2ylnBgJOLUBLLHxwlugEDzAxJn1cB9M47+2riwluwKr07d/sqQqednsukqBHJ0W/96xyY
KZtLpGW/9HglyUUJRPl9s0inQUT5O8754c5VXzObg/eg+Lbhdby9RYZpT/BrZymzkKX/g19x69ox
VmGrkHG+lRIK0f6Q8LBiRkNyjwEV3hzGk2w7Fvi9z+BKRMXwtHCX/6TgswwXJ7xQWpUohc1tOIM1
N10t+78eePvqBTLzwpZmvqQcBO9VEXpKUR1PESZxj0UxDy/NMkYh+Y1acMQB/SRNCPS85r4Zjs96
F35GxLH3OqE6rWmCJvYRJ0QRxHEy9qdqQV5QejqqadKBrDSj/CCktgCT4fRDDG44AWgTglO5PR7G
faOYeq+/OPunbLAkh5AOV5cSghTTYRPlxRDBvPJ/YbT8BZ6oHjJZSrJSEG84WRRJ1oxccpyb5OXU
1/8GyUq/QJ+xwrAAnvu4ksv4rSZ36RHCApBxXrZekiCIO0m5nRU6jVqle/3gTB4Q/svHf35fttWE
mV0nPTjc3ImZtK+GyCl8NntOmv8QHBVBih24AC5pTqgXfTUx3ST5za9Cv3HlVap6lgR1DDVte4Cd
1jGn0mBK+UsV+IVPHpuxgZe1DAeh9BjZEOL7sW4DKSq3Ufw7RNDOkpEn/l+kQ3cPQIehSscvV3zc
RPWtxH58GEYpGogSLGgLe9SkIkMvOG+KKigEmsnmbCqwtwGUioNNgN9nzxSf0djQRrh6dOEN97ky
k/AB6joWtLM8wzWXgd8SKAj7EnY9TlpibZdgSdPdO9JkUnQU4EZAZRLZ+d0CiA5vWBzsKRz95UjV
m8WtoWNUNiLDnRSK417qHoNjNhhidX2QdQ3HRXDuoGlo9YxRhv2t7i7O4sJejdBiheuXEJ/InB/y
7UfpHWHv7NVDLrwzmUJOnNdlnR4pCOCEWm/Fnf/gDW4WH9LEBPZMjqJQZk5RDf5TFGzWV9j2OVr+
Pqjx7yTjfGMjwZQjbh6fTNs8RTPDQvVjZOeCgP4h2ETFdP06PdZHlblz98rcU1R7RtGwqo6QPmU3
KdZBpUA4Qe2wp5gK4gNNNtzJhevPRmHIw3QOPSRUQDjdEDAwjuIVC+xwBcN1TrOY6oot1K7D1+ml
eWoszDZn5YLlnt5U4Wa9jZTFbafqfCY4iwOtf+qc2FyA4HtB7vncW/g7JO2SFRLEEHnash2w1ylx
UJjDm5J7kew65u3JRarPcHanSV1wcll1Z4/Tn6n4FGfF/FutiTVVCZVYf3cRog9igQaOhG9ghz0F
HA8P86BhN5CzFNh6+Ym/eJsnPhaAmzedSeXwUIgGcnN8i7P6WqbIcHPktNSf2OjVfCsb+YOoGREm
FbOAcmS/v0jCyOh5t23YwWlLuFLEsQXDv4l05QnOpVxSKbC2JPPnpijamjz6cJn5gecFYxPX9aPf
fvNslxkRepaNkHCX0qAy2VKeZZ3uHLB3jXRC+E6QZDqyhMzZjDDZeWmnthDqWDJNHc5omJIrguIr
JZ4hbe4wFcTpNpEJ2o/iLIrNRFD76Q33P/WhJyc+IpkdnLqb9b1+mQs4u7usHEcQj12EIBDN0HNH
YotJ2sVFM0oyf5HuB9MR2uuiIPGtp+seyohJbMxpGNOsEmgLnhnXll0+nRg1dleCw4UEcCd89nzY
d0M7lTVHpPWgXzkergqFx0BYyAAdrx4c2OiCfs0cAT85WQQqBfKQiYLG647uxGQRNEYZVPj07ZNk
wlqmbQ693gByLNAFiLJK5v0lYKd4SWixnhh0f9OaTBGGpyx7E/T9Z8q2sAA/EYJNgCjiiaXNgJCd
qRSRHiH0w3TX4XAxI9snI7oFG5QtSTPJoSfLdBodAo55lXrgUrB8KGAsl/f+4IwWLzrTNyobmD0P
tMSCz4P5yrjMi3MgZoNSvhs7+Kjn2eYZU1W+5rlwMp1T7PEwn7+3YCjy1aLxgPI6kF6e2IjLf5zo
W/eWY1zB7ZzpoDf8SNoewTQ/3Wi3h+nDxJd4VUB7Yno65npAYDRpvkj6No29vsmoRRBfnRUJLSs+
0/rL1ag9uJtn0BV39B2WUrBVDfItyoWAtr5x5GwRaNkXjRWCx/h2MwWuL+/bWcxC5R+jkwi5TtEq
5zxHgP8yPz4IuJLaXBrj99rXciiN9OwQgL9CAEsCfTKOH62e3Ewu5HaCtHP93AfOB/YptPqwkgss
gd3LevxpWE7mDro80CONNgM5G21m/UXIqasI3YZCaEcSA7+iJRuFn5PRPJoJ+oeeCmkbNmW4QtRb
+Fj72Fh5g3+BO2IGsdeUXIAeMuLd7FOfkxXWPQolBFp3VhojjAZj/uiPeHRMgPyf7cojqPqQWaYd
5QxLqJ2XjbP/cNUYgJi+Jbo3lHHPdULztJrOY8yeLQRN3RtdpsxhXXK0eIY+WsuFxaqyiuYnBkEs
ilYYCfw/289fM4JpCw9xNikm2KOC0lwcLzgmoj3jPgW674KL0/IEE7T3wdiemUeVVbLwUUHURTY3
zCkBYO74fBYh2erUHyzKrglTtyJnO7F0yfzWcdodHu3iFiTcbJMIUgiKT9r7uzlF4J7HpuLXH0r5
lHrbHYUKdjvtu/VBmYojue8G2HmuedyujdF205nHELHy+rzviC9RInGzyxp9cIE3jFdYxsupPF9r
yYxSB2VvQom+iMheFElrrG0NQTl/xx07KWu04Z8HYaxgLeNqn3aT1blYDv1GDrEBqWN8Fw7B/mkJ
+4z/53gSMZprQJEb7teFGvxvAUGt188FoljKKQqnCWH69ZI9JV4TLku2gJiENV5rpSY++slLbjhQ
vYrRsxSFkczdhz1zX2qv3sFHjn4QQ3PcZr7MWIpM5Buv37e56ori4Tr0EYbzgsCMPpVcr8BngjBw
ZkUjdx+qGbDR/Bgo1jAnRAquNzjG0G7Nh9qfLwnQ9CgwgMqiXsinrrI2/8FDwW27zlTyCgAKNA2f
eIuOpdewN7WdpPHYEo+76W1gXraEDYFWK1Bd4ERZdAU9YS69NkoPd8mc//z2JAtah69piBEt7FUy
s+gSXc+TLtwmyp7utH5D4uIBB26gLWzgO+SU3nVOly0qvqSLXMQf7u7uiJM15DU5RmnkwJuDfqoo
zRsDfZnjxlom6fDlLPtsWLRZwYJFvnHJYlIoeRPvOJkwNrcyxzRciwgQfflyY5cLYzkVES2Tlx5W
srMej4htYaPFVuQ3ho5JgjLPkxOwpFNHJM3n/HuOqVkrW1TYV3jG1W0AIYtFPMTmoe3CKYkv7x6x
whJfLXcLU/2svC9+Z3qXzwPD3dwyOcV9vTeKAYEeqGEcfl1d0AMh8PKKKeskHyJnLpL8o1Eioc2u
N777pBFVRz6MwQUZhI+JFhwf6HEK1OqwCo0BzU6KaTXVrLDi4KUlYVlpvQ3m8DGsX9+pXogJ5nSK
+s/5AIMZV7RXrprQ4h1wHbCFHrAgazV4/MsQXnWzXOY/x7crOe8kZymQoAs/AcR3P7BufMqW6b+t
Bz5X1N6nlp0TL7ujbHGi89IAt36BMaUo0ISCd3sH17viqAC9oMCO/GJ9PxYbJH7/kw1/m1IZ0EXW
CQRk5K1q/m7k9RFdZOdOSDdLqxCPwU0DKI4SI2SU8eeQGYT0TVLiyMzdPygyjSOaLPUHm2+1Hsmg
3kBX6vYfoUFI1gzDGcrJ/d24QSWJ5exMTfIOngAeo8s1ua6godxvl6oHG46schR2B1ctFhrhBUuC
yn2010LX0NqVRXSiBpsssOhYsCAuXBinJ49rJne+LECMUUR6HqqcGJP2gIbbi4Sdipn66tH638Kk
sc+tMbbj/LFVkKZCVmyOflMdjxDk+WNQD+v6JxVAGwu+fxfSmVI2xhEKnajzd0nODKgKf5mU7Vwg
ZH0VzdycKSb/WVI/i6yLGMrckuJfNl9Rd8cvtMeVsEsfHMTmreKf70qkCHFwWO62NqfglSyPWLEE
4I1SUnYvrPYj5dMiyRdJMlaiNXIoly7XGHTCT2lHrRqVy5JQK8BjO/s/dpK77+GO+9gB7rXX1bfN
am86tZePlkfbIt4ncOXJfnAagHG/i0boRLmIY2vl5GFzA3Nsn9KADmQOwjrR/1fE9xmuq9liUVDd
qVCwQGIqNa0NOjC2JCcRyF5ue2Qvb0yE25ClNIdG+lI1xdLMFpTg3kKveQhuHpS3O+hjfdZusWVN
d44SH1x97THJyGfHZQGFA/y6A0doXRiNJ1Kk9X8zaUEpT6EOIHdmdgAG9rhFJuBZdvBWyKjbYeYf
diDaFEIoYluthAzzkFqzOCtf89qUkrbYqGLOS0nlOEGhxQNbak/EqV1r3ftYOkZiqf4eGBVKGULK
ljLrypqBYyji3JsS5FvAxsH20QnL4isGO5y7Pb8muNuFSMQ9lrcJOixQ1Na3oT/3kvPp73rP9MaM
zwjYZucfL0r1ov4uS65EkA336rjuw0moiGxwPhCiR0i3hforykknaQDld6EVSaVlUlujhzlvJP+Y
M+Mpp32k4LgcalPgU7IbMmRVqWeiZS2mklID06Q8tzjxOMzk3o1r8YqX3gmAWi+6oxqODxKaPU9S
OQTb7DTsCuGjTsI8nzFWra2kMONqGcwYH/DnHk1QRkLOBg0BUXZa+7qiPc6m+WClKFJg0oKmAgo3
S91u9l4PqkDvrGz8TG76W7rJUQLtMVO5B+fcpe+8MhE72eVDqAsME0f7X2DDUtFAlDg2Ukp7BvWd
HBCBw21M0jlKUKdUU7vapHAqJ6YzUnFQaQm2g0bkiqaQMGrlRp/60AUwcrT/Ifyr9asa9pCje0ZF
yPQYyuPuPpgk0q7EzyVKvQz8hdCBb26KeSv3QbpD07xU2/pF+F+go1qwqKy7zat3EMzjh/X8asNe
3weZXHdHCyjRKKClHYCtimkJEKXfSSa6MHlczvPrz868oYsSrg3lc1I9dH8GCYBhqXQhi8ItxM0R
0mSDWXkFBqWj/uNG+XINJsmlVt6AByaB1lroFY8gIpv/FQsXDJ8g2DHQSRopEkBnDmClgScuSuNx
3qQb7iJXEe2YUjAM5QwbxsFqi74d9Fhy7EnOv3QreBXjRzSgHCdKT9MgpJq7FFxaCtAp4mOn4v5R
J3Ani9n0+45+sF/wtpQH3UzCPmbT7CcFSpaT8toVtTI/B+GLlIQ0DMTvP0pKw6cpeO5wWMAZvbsK
uj8RhdD1KkNn33kZkBp442mSXdrysz8RNWydaVtLy2VuoInfDW9XK+dHwoWZpNqxRGB48mtyrgIQ
setkudILXunim2a/DEp5N4+ZchKMQjInDMr7nyQDIbT/s+67BwTSmxrxl7hLgdKpzUE0DI7UTNHu
blG4wwY7xhsiHhc2auLZK2wCvqWFsg+1//slQKz5sYFRxfZgZSLSOg34Fxf/7GND0ObWsa3KnzEe
qR3Ef3wDtHIPJaEFjkjMjZuNDhtbdEPfLohYmwMbH/a5gLVfn+1lniUTEYHXLzGfu7zsExguwwXz
i+/ML4Ftu3otumnVxbr1BYQF+DDGO74e43reC+obKYuuaIG7BSe+swja89b/LSlIfV/ul8ZREIr5
3mpNehWvBNNM8soILrfgJdI2bIez5hTfE+bMy8XEABLWbKn2gjyOWZF59FHyk0h0njKm0D9brImX
+ot0TGwzhNhg41DwiLU4/9kmaMa2IEAC1i0/TTP3UBj7PLrVBCnhrKkR1WaJLWd+6O7jhC5pUNTv
w03uiNTXDMLipLtr/tV0kNXVFDLWbkkTmqGsGtIbrKkRwYVMGZ/T1MR2ja3G53OoRim6oP9ywDSv
81CgS35rmIaqB3vJ7sNzC29dDRUOBQgv2knyyy4D1iOSZa54OX6WjduGQRQMH4F0nta3hWWz8R4j
oVlj0yyI8oPFVfQdTId1PCDPZ4vUxY6cziTQAhcmLEJnQeDho9d34NFd3TsYPuqH4ZfhJhuv/wpn
gbCauA3OsC5nTbVj9HMUg5UB5k0oEPBsYFO9XsUPz3RZHXIvzqfjDLZqNNRngxbhs+dvzTlGXRht
/ti9cAYdCGc9HeHl6JQyP0AWiBguEpzPFsWTX7T9IN1ESSRhxB/+Xitm2XEKUkMjC9tny0qLmTUJ
npirZ2zMkMmVsEV11hSnfjPMlk6qZbwjmtD1UZDF5OMi8lSkDDFDgwE2+ApL594vGcRtQiz6jWha
w47Y7BAWNdCe1/ogR7uvLYR949MaUoCqiXlzH7pJ26HnBN1BiRk3Y5h/Y2ET0o9ruVpLi6DRWqxt
7C0z7kCol4olC+3D3Hg60DRIx1ctOR2jkDtEAWk2fN5J4GkK+ijOU8nHnhH4n9h1bwxZAF7BHkU1
gCxX2/kJSkxR3TRCBtpS7LcnKdx+wMtXrY9GEMFffTG7yrFmWHQKG1pNUaURv5A2gP6CbQEyUCEP
HEy2cnSyp3W2xo6aL2VSLJ0FJXLycXfTY5hsknLMQ+03zl0th6GMxI3+Fg5ZSl8+F+yhDEV7M9GU
3+gInYS/qlzHQUqdbdyN/gcuyt+ekysDWIuieo2/wtoQHy9+xTocDcxBvwS7PITDFR8+MZTM2vOn
J41LF1bRRyLF20GoC1PREMKFGs10mW3wioHvjXyC2jhcCxAqHAiHGA/6XqcdJI48JwgBIS6qfLiK
yyGWh0YI/z3/K/oDff+B2TePFAtyNPBCa9eef+BVidLmPclGGm4SXYVO4CqGPxV4EwLeB58Fdey+
WE3nVccK7Oc3XXKFpi0z03nsYfAiHBuz5TqJRxEL0+yDKk5aJynd/EGdgCJgBj2dXw9ea2bEYVip
auO2C7XAkmjCaMsVU2kkU7y6wpezqktZMMt8dJ+g944PwaDnRQ5qMbo1qEgDI+qnikYuLCJVX+vW
f864Wv5O30j8KrwfmOSCr0TQSGH9pjnV8lf04lw3MXwISVLur/rN+ZojkGYpS8MuNyYV/ozB6di4
GpyDvziph8JQZl7V9O4LYb7IZ37W9j8siqjbN0KP6dzHr3RbZYu6VyS2Qkk9kXUQvVY87N/D9Eki
W3W444n5JhGRA59qRRInAGlV6n4lgYsiExd6OAmfErjvs92cwpWWA4bjg4sJY7Agv3fdo3yLtl89
Yyj6eKf1pu5pIAWRmR/Jk5o0xOBNJheOFSYsSTYC6vnG8KSoIsE2M96YRxNdGR8giGr9LJJeTHgz
ZMP62/41b5ur9rTltz19CHo5vhsGj9QLhVGTrMykmrhdJIscT/Bx+xXbrqajV27uHB1ojxReZv0R
UEjffBZ+W3gOrKw1bS1nfxOynxtAAD3qEH4fHpiqzENJ/KUrCO2jetNw4TkspFbYqretvhUk8kBV
CWwzRX2OHt2e9yq1fCk9KqskYQVGNNZ+nkmq37fzpl7vQ1g9UzArtbPP9na8Qrj9/M+w+16blCKK
xm6vDsCvub2fT9lO9UdY0MsW5HEq/TUka5dedZJw0dGUmR4WoPZYTs/MeWxqIfX7iZYR8+wBivyY
++tmXjlEXGsWy2OxyBYI3y1UvTxXukLIDqr+uBXnIF7WyD2NlIrXzQ5kbuxj2BbfjNLe857tRb94
MFNlzUDllVl8vsRXd5JsidM7USJlaz4GbqZVI0Ddh84z3KSkBjWyTwG6OUvhrUhT3lMSrrs8aKS7
gDT1XFrws5YYJxMcsyM7EQqRA36thUuicXpWfqS3iUUf8MEVTnCXc0ZKXPVBjEfTK1l6EQAv9pw5
2my4A/NE+GT+1nMnPhUmVRizxuTLDv6klW7hAe9rN1QClPddwVNlbWDESYQkLt01bVqB/14SBK4+
6Jte9UkB1DJ/olZp2uvzo0wUZYUL6pMCIhcajh2WysW8joSw5bR8TTd5TnToEtgNVB3KFibasm3D
vAkiZY4lbP8Fzbev58/e8SxS2Ajh2b9Wmh6OoZ3W10GbyW2D6tE1cBvkjM4hstAE2seq2TO1/LGC
2S9NGx1HNrO3Dp8x2aoD1Cex6qSai85xUE85uJTffV8z/4B4m02ZuPc9+kb+t7j63TXVakra+/UM
y8Ww+/HKOKvBN//KC8DgHvp/e21rRUSjUyei15ZoRZahRjwRGJR0F6q/CO4opKW+kLAPpKt83GfW
5KikLyidxLW/4csHEABZVjrDZrEUaq5q5UhUVgdaiifIEZZ3GcWSx1oAjvnE0kr1MbPNqC+yljkB
ySGOWk2VuKsE7s0JqVoGSAzCjj6H077rdY6rHSi26l057DGCqkixd27DqmWaJ/+tXXCLMvOFppfL
oOOKfj0Dr2HseE6DsvTf9mhMyzsAjHUYBquMF4S2Y9YRPH4I19CErwPBcO+TRxCiIzZFv7e0szSf
WTGxp8Q+wuEbUXnpLAMefi60W4dWhvDpub8DvMVKBigqNBk7Or1Cl8/2fAYsnMjWY+dI42DiKDgB
CWH016Dg5tOlI3Kg4Cb0vxMBMcnjouuyJg9jGsxz2u2YLbIEqeZ8e0ptkBJztK02YnpSZnPf6INI
5WH2VW+xv6qTTgvJqmqV0rQq+l9XA1ysOiwB81xbku4i75TMBy58EvazEos4P9o+RACOmXjUyS7f
m7mQNTM4fxrWzBh+bo3gq9ywZpDth7hf+7ZyqMkDS3BDTok7kbEkt9yaHLhDu569ZCrxR14mLivD
sHyszJnXcgojdeApygIHKqwVobO/DTQs6+Mt4IMYkaOVVYBjoHFQ+pKxMg0RIKcmcyolntG4hGDH
VUL5ELqS/GCrYs4RMG0gBtzYD4to+qNqXEtDuF6mSkym3oHsz6yXWyac6/ykPXHayRbE0a+a7PZA
PnCi614H5V0HPRNr2ORMo+AXt218leMV13oFcYIfL/PVvue8EBu5DJEBVDPaazmSYFZFmZXF9taX
+7pLVR5xOtIrWN9wOw68n4Oc8Osw8VqhR74lSVmQFxl54ya0JL7deHLsxfecmXygvgB1j/PGQzT+
RfwO6B48wp4/m7Lr+/kxONRrip+tHKTi1ma9bOgq3F93fq67REZm421GgrSI+X9PtI42TU3+6CSv
QHgsrxM7ys08DgyGXHPkapYsavY8+hl/zY+iLGXQCxOd1ohnqxPiLWbjCzU4sCdPuyLgYUOQzsFS
hKPR43rpyfrTJNwD3AV590xOmkX78TylVFhxu9EnNAT9m22iKXqPA5nTn5Dx4zaa4J1prlw7pNBC
muAu2tSuQN7Aw/Xea+SbBZQg7XP/YHz2Hrsm4tFbHQeRUXOixX37xi9AVhUrt04EENR+Ufu4eAsY
lbUqHMvvqV5dAC58rY2I0zhbwx4/R4QJxNczn8s2CfCXFKmbp6tRMHcbOHq+HjwTwKZp3MgWuK+p
j5X6K+QFPoVCuYFE3o474Egcpp3k7arXOm1syUluN90pNQcYwAGQZBfWINB5JJcoaYgyUHtUq6YB
ahrjp3iECMYJ2Ts65N+lk/4S0u4k/vlHCQGoOBLTMRJnCO37i6e52N1Vz9inBm2pjVvRLHnxDnbC
jOzR04LFh4RU1cBo9F+nq3zeDGoIlVlQS2rG+dIrBZe8xJTmzKMFXrAhd8csZOG4IuesCrmxrzqM
58bqzD4jqgg9QpwNE1eJBodU28syisIHdISMCcMoH7QQLo5wQl6eNJC2fbh6v9kPHJhKmImB6152
9fKuhLm3+gO/kABXf0MgMLJ+3nnIJYrk2pH9Ql4JN8hI+eE+rvrfFk7FuLnKhhxqStWE4xZoqBqb
e7CgpjALKtZmJjSwYeiuxzINLTYuuGrz7DLdeaAOjOmmEY1EKhI3FBywTW00xyfd98FCrLukoN+9
ObK5KID7/RHajx8TzC2AKAui4w/OdCLM1J/piYdSK2DXVMEdzAJnKBZvPxKRrb64HWrbeEwMCBgX
SdES8ZlGFiU1MZGS17+vnBEc7Hou0bOvUJ+2UlWD+EDTP75rt/erXBmt1BNaZqXjoU//hjXNwxIS
Bv2sJ7rrwcw7vcunQ4xHVwyzJgvpvK0FHPuFDv2CfVHg4JL92mN9rHbfrWTt8o6zb1XQACPsRxnG
iigbIu2u+4rzCMYV4eOIXnuGmo7UoJ3tUSAKS8Rot/IwnRCKZohNvEYCW4/wL9rZkvM+s2LssalO
9WDhExbAmsgIfPTqF2+gOuFf3H5yKuNYhj8Geq0WJVBflm4nB989gu0FH+xlHSEy6SpC7YL9QeZ4
LwyX7aP+F0DdmaRZvI0k/pxAb6sPuRNu8lnDTDMOYTEVM+N1Mf5qinlCZNfbO1k+aZQkAuFgTZLW
2l6xWl2uD0ZG59+IUZJaioftUTNYhRunmUcqhTup2hjlTclo78F65BCmxzmL46/0PCAkfAhW2Dmf
aOsqk76wKFE0/xoZZohjHdZy4dD6dECgbKLr9s9FgHaB+lZbjXxtYybpx01BqyxkRX/Xo0XKOUwe
EYT6nUZ7UyVusg4D+CqCT7zCIdsqqLebONDX7XXkVSNe+kEYom8hHFt1xbf5keVVugx2wkRgnymR
oGICr6YIelTrXEzlZsKQNozt/umZqo1BaIWyd+wQfPb37GAruFyTfyVq4kmfEVLyUPNpmw0c/Gr5
Xgk8pnNzvE2gL1PuHbinUEYjWgCF2d9Uo+vsRHk9P4JEG2tw1npGnKsnM9HAXwioDEb0CwFNNH7f
57ujcaSp6sCp3nYXrBm7I844Hc3FSpuq8X2xeEAioZJe0gssE0RSEfPhhcdy0ReXhYlfiCUK0pcy
yWLRjiDuqo9DgVl8B549fsygIYYwlKROCegOE/laDBeS55E6S3Np3lGzOf9XSm2ZQq5qY+SKrFx0
k5/5qIC/0Qg+3RVrww7aP6QHSxly7rH+fLFVxC5T1T9Txh7+BVpgW9jNv+4V8DGXEO2OhIrwa2Ge
DwaOLjsYLwYfF/h/spNP8mWBA8zRZFEt8Z3aRicmWrSm+w0cbopkUJVbXf9y8y/2PTC031fPPw04
ABQvyW/A0/7Qf4psBV5+9q2JQvkeLZFGl2WN7X3C3X54rf6bTp9NT2FPd3w64hHCutSqOy7Lrb0u
H5e/vdxW4s2kwDibZOrMWJkIUhmnkpcJnB/YAA7Zpa0G/6pEo1mcuXV8Y0S01+AWsPx1FBejeggR
c3ttmt6cr+x6hnGMer1qrNci9MWjI4vTH/tcDLFph7Hopnw0arDrEtEw/5lPjKlxep25x8klmDus
3zmGQz2sLywqbtpRKa9AeLQo41LSkv/++nCxXiCmeEva6Z4qvpUATe4eUs+ShbBerIcHxqqp9J4P
nqeRzYEJhtxaChnrd0EKJqnuuj/EhZqAxsKdGFnE6EZL9WhrwVDcZx6TZXhEI4/Cy9DfaV58/i9J
XdmcWd/6WhTQl9KGS3Qm5kgs4WblNEqdBJl/cj46GRMFpZ0qId654HU04Zxiv9ji/p7riDuJ2Z9l
rSaOV7o+XoYy4Cg3tpgA2J75NjXuA2UQPkP1W919r02ejH2Y7IINLDgO/rTFkq2gcjupilQtEyJb
/o3PRvAl+JbkUKTA8uG5uhtgqqrb+YRxMj/87ehjrW5e5Um/Qjt72ISd87sSwGcWKUXZEzc89+ij
ONl6VBhKA7B7L++207sz0UTv5TUA05eu8fMrbz+6fhkqaEBpi2dqeZ4cx/wIgf19YEcGLEQ9kiRD
MJBmW1woBkpQmr1Jtob1Y0sC+kUvbSXDyQUotFwabpPxaTSsb4znsnBGd2YfM8cnGY+NF2a7YPGS
z7afdpm/e3ysCk3mA5hfF/0vvxJMA3A2X/toJEBIAE6K1+s7bEsBeRP2Mpz8//HrZEFR1ErcDF4u
LSQ4yKcUwuCGE0SfcwvcUDF0nn2ut0koTsvwnPwAjvVWDMug5PlZTqi0sVFiGLE06jb71nDgQQyT
Agpt9+m1aTJyoDge/JUfK64aspxpmxTkYiq23/TdXQScNddV/61pL9WM1HgAx1dEY5iHAW/frP8X
xhfblwwKbJ3eT8dMysPkhIBNopd9kMwu0Odl1AAtu0ZoWQCoAFDmMVMOqKsvhronEPp7gtpss6Bq
v6mMbNdL752wRL8YtaI4u5k+Ij5au4Butcwhw9CqLlzQrCQjPXpOKRTOBL/fnNtCWSvTzryk00dH
snq4oPI8erAlBH0FqIR+bSNeLP3WUz+6nGqqJkhTZKtNSZLhaeLBSCj60H5u1+0HxhUZcyCJK6ES
UuaiHXLYHqLWEgJgjFaTr5HbA29/1bB8B65FrPxEbdju5Q2F3EBGURS5IIojudP1QIWqxB+r4uiW
fur2vpI5DEoz9H7ek99df0kmFEu+eCsVZiByrmVy3PfRyzNFK/p0z5oVipqgFkzJcIFzrzDq2zMd
YxvAIe5n9p00jauqkL3x/MlEDcFnYDC37ucyt/TiPJQiwP67reBDKeHCrjmPSPftjzfTER8E0O5K
/L5sKuC2jTGcATuK8i4Px+cL0ifLguYK/3bTMM+7fdNHE6zp0TthsvOhCPmSeW04VVQewkmOvZC0
D83zexgoWSE4p7vkdfI0lquWWXo3ov8kvEwOkvye7h5q6aMUwr6KM2+8aKD7XymL2bArejPaDZqj
x/vH/BSFg9eS+0++1mnMOgKwa69lYLVvcYHaqPcmaxIkxmvsn6/t500EPSONdQ+toiX272CZLMkg
OvUQmWUptRTxRR0WDIhjhVx5SYsd13E2TlWPkNmHifvjwXrTVrM5gcxKj4PUpTsvevnSczHQ8YVu
p20lmGod03nWq2StOKQvmFER1vTkQB1RAmcoKlq1BKdaJA066lualOP8Rxibf6NYS/VQj2XQ3Lcr
dvUtDcNj8YajTDBGFbBHWw9UHugj3tO7QOhPpwDt4zPxaaMnerb9psqeHn148/uSgH3QbrdPV60q
CI4X7ymDcKcnvpEYOAr4NH+rbZHKfVlMiJ9hVyomUgbur4qYpLDGElGn0r6txVocEi77mg3+GROg
GOIbkBYH5Ap+aUGrdn7tzZ5ah1RskaN+ujlx+kGfiFkRssCeRoElA+zui4A1G3ATw6TCPDgxt6Fn
pCzJoMrb2lHWWJqifIRkpXPnP2iLLaIA66hmN3Lxjd7jeGU45JmGprZWK4Ke/yGnMSbVHUv2Ad6V
U1LaCk6zAH0nQJV8ORvJW0mUaO5tHCQpCq7WznGx5SRNK9OOdJMQEzZBYFJo6wjKmadOLlsdhE8B
B1QdjUo261ANNQXGpZV/h61M6pASk1t4PwXF29xwYfa9qZCnEEQGwNx15KsPafacTvnHT81n48MI
948uNNs8kfTqwC+/+CNDIAVhRRoLFqwcQm1hAa4PMRDgRQw3UdxYV1TOobpfvONbdM04tDF0jQQu
eXIzFuaBuGuM1WD76dPSVt+t04gHG+ZCVz45paoNO1dFQCQZofw2Qyz0cWFuvhI6ZW8l74YlQABF
aQxS0iBDLVdeVDZEecOu2OyZAz52eg4MySbIWT6/kLertoL8moRFVsW0OKCjNA6EGR3nJG8aTGor
RVeiOYafOPROH3zfbvGC5s7HQEgUYO8/cPkmGQVQcMMpUYDTk0pUmV4CM8cdFXZdqZQbXye6zQGe
peeu0c7+w81nq+sXmzYgSmXroJyOlugW6s70gMNoQgETm9ZzU4g6bDQrF3zpGwjxyVeEFbccW1yk
5an3AlPO6pk4UZiRzh8IV8IO9vaJitA7D3LZgn1N/35Yla9obzSXvmI7XRPYSTQq2VHOlR6RusRz
tkoj58J22ZNg9in/UarEc6rjpKIeUW2UbjnJ48DW5OHwiEOCWzXs5oWvXZ2AbKs/MENPTuDeWvga
R+LELTXKgD+5JtjF6oX69xQsLewYBsMEn3BZGc6qHvtU3MwwUotLCC2NMYENQ0aXE8tGnmeDmHKG
VCjN3PW/W9DhWnMHHXNXMmWJC6QNROPoKTqTSg+I4awN6SCqDGC931lrzL7KStp5J6GamiF2MarK
LBcbegTdbp9h/lAz6135mQVgNpFkfKwM26+jbK7glZL9wWCABVFAO3NREdR9jU2pWOoJsi0cPSa0
O8bnMKVepMF+Wcgn+YJoNqYK5dgw+NuBOnCN90sp/yZaLm2v7pjc/ueIp53j/3U6fab6ZyTGhC52
v1LGcXcuRMKMs9symFq+j9K3VDwCMt47Cr9ioB8zbrVVNJ0yzkSOie4PINt+pKBKUr69WXWT4APb
Pfoga3iO35wUmcUx1fTOHTIDy1yeZwGmrbkdqmBQsyf4hrqVDvw2usvi1yhUbH306tACKPrSTB1e
3EiwPV3OeXuxO2Cuua3Fr8m1mzBYLP0xq45F5JangStTpU1yZfkIusivuT6m1FAx/EP5RgF/qPPr
Evxt3/OdDUyUxkaVvQU/B205ZuvYyOg1V2LET0k9IKN/ENtMalVyD7lBjoYsQediQzdfBMAfp3A/
12bkckTYwzE9wew1/cm4u9xIBgK5IoIHjw02nzJPCKVzRFdXtEiVOqJUL/SbLZqn1CsXEQCPLCr0
m08/0r6r4FJo/iczu1R6sSQ5RU28rIiOWXifwXkakcMGXuLpLr9WdYV3Fc2fKT4cXSZFRKzriFu3
6tqHrb1Yme0NKhIO6WsMEcByGWHdKyQPcVPPZXulE9noxMNpe3NxSD7vAkR+SHBP8mXH971x3sNE
08y38C8gzV/svO6YPp7jeg5D1jucJFOS5M++tPBADgtwPGTHFGvpsa7Ji7JccoZWedwLjez5LAFo
LyF/UdSRDRCIDpgDy+YtvAi5KUCCMjZhTvyI/C0zvSE0lUGHa5ixWSIvapLU36jOnHha33MqdaNV
B4CPesMvzqUnG6OPuV8MIZxeS/2QhepwkvZ6dzcMNf5c9x59OYcD/4Wl5vpcvLjiF1xc1yuTdoP8
kBWufDrQSAddaAVoeAAKfmXGVMHmPXPsEXctIhJPaQD4WyZYgD+/NqeO0U9ZMTMZNxRwc3sPxPWe
Eii2lxdv3TlcpZr2neAaZoHzPYjfAlHRiVx3J7f7y7TO52ubP1bOCN7+aoFURZH56VC5qMd1pY3L
cDKh2YNvEHMLpaiuCMPAMOSiImrppIhEbh/bsXEp1PkmQgj4LZ5BmKbDYxvUmenTb4/5qiwVXgJR
xs7P01+ALf1g9EsesNUvFey66ftqQ1Z++vbAYpKmGpUzFI80Mw2rKWb8t7SjgQkaWxDDBFwM1xjL
j63hM8+E6oWwH37oobvRHWxHI21Q+Xlmwwz1hqKfUEtYF3vR/78MMR19pr85ojp90Ja8NHRFAVLt
qnCd7ZrAp9RNo/tX/TJEnU9XC2zJz1ZnMWbx9+a1sbnyuyuFEKdsoVFr5WBG0oODj053qbNBzOUv
lpGDCrB+LmJB2xqoCAG260Kz+IPeprau6+p8Lb6oOFFs5o4QB/F2gIiaqt1ElzOFSXZ872K0krVT
o2XijBWI+Q7kl4dLxQZrgzUh5zQ+sw4CKur9ZBB+5dAXXqiSVfIr2DYD+U0WEMb6SZu6NYpujMGr
tutq41qG7oPGVZ17ICWROS1acwGB8ynMZsbjZUNtOe8bqrQ8x9Ebr28iDfWo7A1qVsHmNnCcBtwl
aVQ03Hkbfx/4qZTnRgduYssSIwWScjO5MoElgzZBw1P6ArZ34Ed8QCPIas0wrZY5IH7OO9Vh41oU
TF0R7h9krDhge6dKHsbxIXQELxxdZeQNmqsyv4D5p5n7Uzc9196T0XW96uF2QR4CQvb5bXQ/IUwG
MVDuT4ca3zIc6dfVkn4SpV9u3mZj3xRxWEK9h6gZB4zKonAJYB6Y5gJUcfiXIdIzOpZQ4LMsJuf1
oHwjblMyVV2VOzMwQMhoq5cVmE7YT8IiY/eO32ReoV3iTP3mQ2DoaURIujvdWi1ERcq7hvv5ulGm
11takm55pDhmw8lpCQnqR3qPP631p+vZWZViVsCe+NIPpVQg3P8PwneQJWzsrSGhTBRPg72/c9HO
fUsxwdEbsvX+KoaQfUi05UMlyClMook/g9ROWrtjMac9XXodURLtz++2SxOS4ZAMlUZvEGcydU+7
eclSXnMFVUwuh52i5gxHFnxb8G/GQPaeeajEsQ7SmG+2Pih2CWg3EsCKlYpptbWQxowNMAyXMFMQ
5qsOoVqQ4IFU57wzlqzldqI/m9pSru3/VScrm1pC2Qb+ZIPppLSy9RiFwUB+HTruPvY4p77iq1K4
umJwus3ci8r983FPSQfpSsaTLICWuw+5z916PdZ89ufsDCmvRrlxEME8RTohiBBql5ahwZcdaqTh
PaX7TRlKfTbJA2mepBK1PUdkNlaXI5RjEl6y/UcK7l5DPXlESG97Tf5E/m6N7hAR18Vo+QeHmGdl
iavs7jNbj1s6s7xFT71mLvAwtZcKxz8A0YgzvgTpf6WL7PEY8dEKBC+X8/FqFCwxt5HOcUlfprd4
mn91rHELjn5TLOuw0jqnT9lymTHSoxEjX01c7Myt7oZFeZfPf2uAwpmOYtWfxEzwBPcDax0dFA/b
CyewgEJA9oSyuyln8dJrDC6eX6VL6JEhwtlC5an0D1cg9pWhEyVaQBsXHn7Y247KBDcMPxXVWjwQ
0ZS5J3jnaUVpC5vCmECMiIhmIUP6cDymacxTwMndgyr5ZEC3YtTXLe9BcMDm1hxhrJA1NJC7e4xD
PZlj+RYfRu7k+6Gd4PytSJ7Z+0LQD4P3JIfZX1tgypLyEh725uIbxLBuhV7Xw6kImIJqS1smHU3e
usJ6SuEf8RG2CnkbeHzxFSx0ZBfm1iTbkACpbY7oKkCCQNvzFHdD+Hk24okh8bkbAlUp3X/wun6W
f+uqPa237ginOk61H4XD2dXxI9fMiAqmufBrksbP5vVGpAJgzWGymWivDhdNPKFjXjO90HOA1Dvw
en15gI6FhW7yiWLvt92hx6PBACnbu++yr4HAoGcO15LyJEYblvl3lP71oi6NrPAk7xkavZiHgJU1
JpuViOqpK12leC7JcReiFqDSSCQMPvXxqn16uzi/5/LMuSYEKsv9Obya7uYUIgZm+4nquZv1rnaW
XLXoUIlU6YRGQS6+ex+ndVkfXiiOnpqLF6pV2ECNH3oa7FR1OEUJGwr0oYqS/+lLYM1+WXzD/+uU
X1M8/mghSlYSWGFzMXUJnEhRgCl0RheXkt79oDvGo+smrwMEz9S6rZEhJsi9usgi7R2FajtT5Sdb
yErLVfw05/5MztA0j5vsHVzh9QdNNMeZ0Obrmy8xIY4d/wSUG2O3as9CuQmdbxjVj2cfu4CQ/evv
bjZuIsEbbqNF/dtm/tZ9F4xGBXzUaLfgMHpIBBny5T/mHrLLa4O2orI8IxGhbbhes/fOgX3zUbpC
XEVk4djObLwL8t4xxIRGRL+tczytrM3Ysb3aCFj1JaiHeT/doQMDDX5apCPuxW/xFd1jYp0hRxzy
drxzLkmVv1RNZw0UIqzXJvIhjldmVAs4ajIelfzDVVOLwNDkZl5WGYDSANGjxYGNTgFRPKCs7Pag
FpX4FbrqeBRHYTKx33Nko9uP9mStrVpDTj6kxlf82uPCwT2N+uay8ABJ7W6WlmBwQzcd2X/NanHK
DgM79dKZ/fwByF9AnqaptW1AN2TS+K+1l80v2ZDvvfUL5guGgwA4kO57fdWocCp3cUVGXoiKInA0
u1G1Oe7YvCP2L5kovXB+3F//IbEWhBAgqt/xHVVJn4qeK3HYeauWg/KAPTDEtMFNHqLS2G96ozbq
BLMIEhOZMwOa9DtHMICHIOTo4ZJ6YrmdtzDG+o8vZVC5xB254wYe+0EABpEQ+0qW5D/cFfcN1sUt
OzRZSz/iw9u5BAiAi6e+Cn/pNsZ9UU2RQl35qdnuESTP4eXOnJCNX9s2h0E7HMjKDjemC9efEFyI
jk7tGZ1rmWo4S4H6poXJyVMp+95IBVdrFk21kCy484UEIFOTwQq06cOxYkztq1WxuosS+/g+eE0H
BFIqa9nuymVgLDHl+XMfbJrrfog73LEC9aIf3qibbSB7LNne0UHDlxjVPMz/G4xEug1psLr59UVB
oYb5JCDjH08EW/HCoglVnHiljgYkJ3OdRt6Mc7X9s1e3RgIOj41TCoHk3oH/Qnabzt8+ZIEP4LuT
O0vJkrXmTBQx8h3fPtwBKjGqLwJRPyG2vsfRWHWdm/0Z/pCSahosSaki4iHe0NoNYuBCc5T+xOFc
TZqHUhH3Tj5WBY8Hpg3JUPg9g5xNUnidOikCdByuVzp0PszYUuWBWZ4CV2iElM7MyKgIqgjA/anJ
9b8hBG1bC5K/8qnFpwiBqqEGh9iR/xwFQ9D8bGiEKW0/8UA+w0cMicqAQ2PBKFsHiilSiLGOXyN/
ZHcHfSwRF8SQlXx1Rj1RhT2U4Y3CVUTN3SCNApqtoquC7kDfmu65EzTkTl1y7f+sME7DLtWRxz13
/YMJCJi3sMr2a2guKbzrhGtxXxQcScl8FLLK6zxeDUD5ZSj+FRzEiXIL1ZjfwPhlQW1K/aJIkwO6
HSpn1w6QG4sUnup0ZoNxuq0YtLqTsNyTrMmlzu2Fr5GUO3urZsOaQeMVEPYo0bUMzm1PkitPH0S6
majcPfyl2VQkcUZ1Eyw6T1iX+qTmVoPdBIIg1qJC/oFhAPdTT4GFggOuSL8s7NDym+jIdjcvmNtV
48IwI4VPdxujsjzbdellMeh4VAb+Y9i7w/qbsrdhfdBZVJuGYhzdiVN9ENLAcwoJoGVCKHBBRREG
PzfKVwrnsdyXIXOyNxlHDooTTRoiRJ8K/hBRll8XyFuBBmXYNqq516+Kqk0DZi43mGS5KL1ilQbf
8lxDWSdm1Vr/RtlO/ykdgLRQMo2UVseqC5P/hCvqG/aPb8xkFCBU44N/3+EjRnHpB/maRmjTO0mL
KqyVb7Uc2VGu46cU7FzJ2/+lSeNT2imZWd/nOE4luiMTtE6HtBfGK5j3nmeVNco/AeKFCnnAyisU
k5Z2Duhw9Bm/odM778U83N9OT28TFVu5l2SXfgxA+zgTKUcSo03WEMW8T4hwvGbOHoT3xMAFsTdr
+vB5d6eSvuXObGRgoSnHmDLp0eoKiTQepSd+ArFv5D791CT9Un/Qj2D/aDaZ88e8aXJDjyDFIUJm
qZs/bROcKUP7xiW/J77Da7NpwCOXYk26dDJT0ZbfoDe/kUBKbrCRY1c9URfwEZ8XchXSYLeqrAGQ
ClYB+Do6PqIuJj2rK7zDCHvgxCbx7eGchhLoiGWN6k1a/0e+qG+GPaY15yQHXq1y90Y/ZxAki+uU
DcQFUsoC2wda9u6k2LME9V9S79vmL8qkwiODzi9nFzfxzEbUip3w2wJe8vL25eVTvTkSFTpNhdJ4
3rp/yUDiX+UzFXGQukqhrJUBBVCGE9rIdiiD9PIlOLpC3P34pwPZkPNL1jM2ZaUpc1GhHK2/agKp
ujFC82X7dlV7dD2u7Fymx/RiP8W8nvxUliqhuZ3LGTLjDGEMqrJl9Mse5yiP59TGJ3UV1oVMXivN
Y8sFd6uLkGaq2DFcXIaajW/p64Vy5zjP7QsqClbjpSCF4ciTtAzIRdV/6KLMnu9ovNl30R1YPR9e
NQh0050IAGtnvjzUkU97RpGRBVqOEX49ijowmj0Hzg4+blycQ9aLqIqzOv4YN9et6f78sJlgdnxz
zeVrVOWH8Lr9OtG/9USLDQ7M7cqHWIH0DmpJeVNfj8Vbn3DRi5iMXSgiV73mOnBiWw/PgDe2Lb6g
3xNNvQOLNjMcwinwZxNXtnjz++nUEHS42LxYV+69Kc/05NmRsYxe2WoevjodP6fSQy6kcZ48A+/j
hTPKE0BFdQMc/+4ekfWkzZgRNgURGkF/UHXVkZKKsqHfQheo2h8UvBGZJ05caYCfpbr9vCS6isg4
OnETalTYaRq4pwSaCl5ozme4tmC03ygQ4l2QBVrkxYCS22A1xse8LExCbDmN39Rb3iWBqyIqOKmm
XOsZH6c6afpkW0yd0pI0D10O65gY5hFczmHfuiVBSrMeL1VSE5cX8eWQVXMIC9Iu7J8AW5SWA1GL
EeSrF/JnYrmzqZpejvi3qIXXkHBWbkFdf7EKlp1fH7mmsY27DaQSRjAKo3aOOTc76M93q7opxwNs
RLtJcab71CAW0rcbyGvzvrTzeUq3LPO0urnZGRcywmfZr85Iukq8vgdaxb6NGQnN1YLIQKvXdLKf
IHAET1cM/9Wwsa3zzDJZvCQptUV2tay+4y52D0aWEU4XLJUQOXV2B7/s3U4pdMX//WNzg5GiiEfq
dgoCL93krFu3iGBzU55WJ9zjgjGfWsWAkUNxstgatTS5s3cPzWqUCsco3d2KJexkGYV3Y2M0rma1
NuqYD/Sf5K2kSDqvba/WEmQFp2rIpo4EFTdrfKOQONsR86CfSQ8gt9YZIsNhRjSkNPGF6Xhmqoyz
AA2+m1J2LNtWNv5t5oIFrl5IcsfKk2oQ2Brljg1uP6mxVYQhgJS4jUz6IAiplg/Gasw+EV+93U2t
PwH4DIYXS5znA6li1ggdfM5O7YZTBDWeRhIYuoh2sugHtngZmTc6kHTd1xRfYIBmDJJ4SMOkQW2R
OpAbL7Jf0fLKDKv9NeR1aK8jnh9rwRpmkZ7NFRpS563e14vBcl/1SABbRwX3AjReQrJuXLFp8I6H
iofRDHp310xXgjtphAl4ovtw2CDDW3Z2cs3LqpCf7SEhuQMu5sQAGrA/1bVcebIf7yy4stRZkcV2
uCAE+W/pXgCN/+NIXHD3Bco1Ztr2YECYpopdo/NnxRurXBXkLXAdoFSFRGgwMcJKVjOiKfIulAmT
nGZ28UXbR+7MXEuyiLZGZMLCVUco4JQNm6FSMgqaxvrUF9PlczbxbBrL/vuWNQi+pe6PDeAAL2Up
t+5wwWwvXBADwUlJppQgUbGp415eVq8yyqk2uKAA2MOF2lO6A5Jw9DCV4HRvWuoOLLlMa9BITNxW
zcAgHQw7Tqf7yEA6KLi4INtvBdlkjadCFJv56cxVvdp9JXQHJnrmZzIVEzlvoIdxiz2vbPTB5oDH
/nwTbkZmRzTu6YHdyJ1DFLkiM3HnZemjMgVkdabkxSu3wwN3XR4UVqF7dWvmTylY6mnPjO/b2GQ0
Wtqmyz8mtAclANDOgCj+p7wsCdOE/5OL9vWhtMqlf0cXzSkMlp/npjfyVvEol2sKfUTa83isnSlh
JcsETjI5nYsG5pPqnm08Boy3L3lAfBSdS5NxxwL0GHa36+Zc7quRPkXCf1QJOiq0KJgYUZAni4K8
R+eCgeuWlKO5jXagqReNiNWwZT9iU0faGY3N7QdGSsK0Ke9OfWsmL0o5GJpT2Xok/hotHz2TNWcT
x5B61a4bEiqvW/ZJfG0Mdy9hEcuJkuccsUKqwDgMpSebq0T/Fg2azqQyvQUVcX0xOgNidQHNanwO
RGCJ39p2V3zwFW/ggI9+9rV7XPo200XYuCHl60CQ1M3jBbPDUbwnL7ihWZZVJnCsomsOA5HAcN6l
oj5KjWMnRjtAoN1MeV9vFKkkb1F2f33czctpc8a72LqJh9T/VflmTM8TPLUbYeJsvTKT0cnPWXiE
4DhGezQcM6j9Ud3Xw9w9qwhs1mPa9xt4OES661oP1mvxD1MptMEF1HnlmDZ7+pJVlYyBdyCP/oPw
Wyv73Co0zw/yuwrrcYu4vF2M5k1GwLwjupTTBHUw/ii2svvJD/D34gK/PkSSjkUAvSqahw+/AycJ
zDBFCDisItzLZassbcc/eQF4Lz8pSuSQyoGG4Jd3pBEkQAZ+bneZot9qjB6JOsNsicuNu4SyIdoX
yRJRmvOa/KSG5e0SvbikC48ujCPVNTrk2UtkJiECq3fNMb17OVss78vIejf7Z+w0CXqrgpltpHLD
U2I9/jEuV6yTyPmx3YodCEEbSj7M9Cw0MeVV7xowKD4R+U7HnQAqQgSZSb3ttHCJlmngvBEFt3v/
PO/JGffjY/FwkEG0MEQEapHjoaBDJfX8Zvyn0ePFfkkYVBHpLytzr6jDiQ9xc8QPauafOf07WV8l
giz7pnL02FXbumo9jzkosfaRPjXzB1D4cmMxWYA/I5nYVQqJ3kbjr8lj9ghnDOJQZLIVejkkJ3w+
kT6t7+/XhI/sjdbOdLxDvoUlBm4x0zH4+4hgVAOcL0+mhPKsr439PqQHbOpc6mUh45WbxZMXG9+Y
3erZCMbDnNujuePWYhrtsf3LoL43E6lbdPHxdtXss9vGqq7rXxEyA5/B6kq+I+8N07zdQwr84yPK
aAkCgva3/Tp1evkFMOayk0aCY+8zko278Se3ZJD5NYY7+rwjVpC8D/1pexqkcC2acw86hG0c16Lx
lshqiG9/OOLrzdLtT4suICDIMwYysVSqDhWvU/L9X2gi+Pi7fvlE0UkVitSIKSfaM6tmHUfmpKQ4
njsAhCR8XZqQBi9t6Tdr5pysNkzZx3tkndXG28L0DQbijyj6hpg6xCo9PzR/sx3Dzp07z3eC8Zvr
qzk2BHcoWVXVK9GrJbJUBE8PQxgiyc5bq8tKw+dUL2hTw34b+xRk2+piYuIoVS103qA8NIJeRuN4
FpxmnLcrUQ8LOF1gaZTTZ1GJAJOnftXGDUEe23DNlzTA8ByvXOcNMKXvYgFlx2mtcyjBeIa4q+gj
hk4nG2aDtnui71iKHcZqQJoF+0dDD7d0nuxc/CpNhrFgTCiubHVuhu8GXrOfR85f95N46S9WVoi6
qN95X4BA7CJZEgRKb/YpL2W4umiHGo7cL7xm5HpajXeAHuZyHSpHh5RHsM7NHIucPMnMvgxmOtU9
mNJWfBNaxvte5nK8yuiSREhs4mSU1SGh2/ec3sDN/V30LnU1A3oL++vW4EGrt/rc9GC3qpy9VW//
/v2V4keZzQsrNKqc3h0b+xUNFrrc6IXUQe2ECflxwZlgBvHngx+67bK4H8RscHpoBSBuC6VMR0B1
84q7Vg5xc+/RteHaJaQlJSbiVStawfzX+lOJ1vFqVy4wxNHuzdg8aihcySs2W7xV8Q6L1ek093lh
LtWZijPlnIlSA5Jb+3bw+7TciseTm2UJS09T7YpImeZI2m6CuVmU79qFnyjRNctIydgm34AHhBim
TIW6Ec7CAuUHpIcuMwVqtkVWipbg9V1Exchat5rGcHiiCWWlvQUdP2E2G5lRSkgjctAJbl5sWUTN
maIWdX1VEz8jBDEEjZAD+A+MlykmZjvbaY2jI8susSAvYWJN/ym9iFDUfSdPsVJUd2ZufCaoMN2h
N5YKIxGI5FggDMtHOAni/juDMHsN8LJ9dKwNxir7KITKBL47VcFmTMM9dRdsyDciTAnQRE5yJQfp
V8q91JjYi4PWhVcAFIOp8fwQwlr9KrJlM2QF/IxH47hTjwwGOIo7TcHEk7RvoKbM/46kdVrEC/Eo
NdNLy7kJcFGUbreJLLKIwWnVlrnB6a7y6cE0NEkUu0SDUMewL4iqLOGTuuXpVx2h+AOh4cZG9QWA
14tgmhmaBcaClL2cgf7bbGoyX9Yw87NmK4SaytNp9dykag+ffA14zMGIfX4GqRPvibpWzrPWd101
ytxlkMsjm7hZnMeXVddHvJmfStS/UPlOOADSXs6c2pMfjE85zQ3+4qM++G2vYjM9sdQTWdmrtRAJ
Zrw1ozSSLOc/3LkEnLVH0Obj0cCTOQRD21uBZQcGFj1JZpWTIlQV2TZhhcgK5gAngxfY7TONqzxg
Nenn780nYmsBUZh0FN2+a5edFV3gSAGQXBlW+sOIiLRC9qC11wmztmIpM4JJVNOUqCbKw0dkuWBP
ZyXVhD5NVDKSzDWPYXHkKWiz6Lgas8VEesUw2HsKLyhbOd8uGXz3JaqR+sZMWyyvh5iUl28NTQo6
i+FvL0PWx2ibgPLcf4R6AsXh0Fthv8KjmoVAVyuhtdm0g6MRItoDyyy0L8fXVsNQegwomWevSBvt
G1x7yJA3l6mk7RT4a1rdfbBQoGdyKWHwz4Kb5Ijkr5+Uholqp6ZR9sx9G64jeqc5YyefiByJ+V08
049xVjLX3GGOLp4ixfxTts8/0rlySNvIo7D9th6Lqafza8WY/hOx8ul6egXCZ4gAVpW8I75Q1xoe
Oee9GYCqCmLtcYhZfRW0TusspZr/A9x4zgrop0X+BkONpl4gJRBs5JFE8xJMkVDUIEOzEc4JsQaL
oOZhd2auaArDV+E/52FLasY5PAqP6/hnepDmwOCEspth3Zi8xWmMcspkROqdPvv26ZSmR7ugO9mi
b4FrWOuBo+O3AOBSNkFWB1Bcxw6Z1fP9A8WNpNXy9P+dkBVwpEnBrfQNdB9UbD2neLrP9MDM9NJh
Kv5tPeSj6wo9Z7ChXuef7uEgbTKXwP1pXH6XJvyKCqe0jzZVIcl6hfwd0RT2q/SsAgcU1RLJCbBV
kpjNc5JKHMYigcK9ZXp2wulhZsfgUdMg/+p7PTaMszXUQfcO4Aj4lt2So8Bn2WNS+K8XHdc0rU61
Qvp3/h/Stlp8N1JhC2DkQncD0NbcuH1dQzl/CinwRshC4gQmrN8j39BtgGgpCPkRyL8i/D5FpY3b
y+0ruiy3CaB2lgwHRf6yZXBeMWZ2boGBgYiH1FsXuUIP7CM5gXfdZNpz57uQhgZq90WBTIs0r+cK
Na9wUVdPN6iCovHB8ykqoeFs4hodz9tQd1p3+f4xZnc5AI1cq+NiZuDtwwqVCZ1TQs7exvAnM6rC
mz2ilEeHVUnjqGI/eJ0afS+MC0xOrGamqXg/N52ZME3RgIFMO46p21U05jlfz/HyTtZW1GHI/eEs
3y7FdN3HPChaARjfZTqQkYfbkoSPjgzHAktluTx23dPhc+ne6/vzPOkmgZlRTTzDPTBTKcVPWxLK
3V4kNscW1gx+jTADIYWrwTzHkbR2JtF731eChfiDw/pf58I0ctirOXtQ1ag+YDI/LcUHOnBqVUpl
o2mJtHIRbbtb1vpdqcCcwaQpEganbbz7b6NnJXgvNByo09J68RF5l8tsGY5pGnzxJV3MF8AQL+IN
GzVm0c2vRGQ82S7dJhGxkwBiWbbfCl9wQsyOVRQ9uiDJDPe0TLkksLXlQtBhHfW/vgviwklYOg5A
fbRtZ+adzLeSa2Vz+jB6wNY0QJohn4OAdbB5/u/6SuF9SUK8vANxtIvCSLtGHHz/VkJhhEyyWO+X
Ujcr2XtzSD6BIGDrmqPOMBwKQCrAVp0tAmLmmAyWsKipYEkakp4jKopQ+ly5LoaECu9mkLfahAyV
Nfr9a7BSjp2qzJkTN0S506H7TiGaNL5mTTCzDxWdefvpS6ihd2KMgxyke9zwiv2XqZBdoNNDVt6O
se52rCvuVF5NhicTXhT9hPk255AzMsbqoALxSGR7kTPwc8vjDA1FXLuxsESROwnH5usR5yLGmGNH
rxwlPsjelZ9uhOrfC1AAdzaQ/0CmQoFiERCKXBsdSsYIWqUNJPNYdmKhc2n2mhbwwvoLD3LCDV4P
CWQ7BTQhdAWL3CyCde4lkyhxaEcBDVeru9XAxt62fvMOQl1PB0VEBJlZ6Ph+iHHq5J2+EnCkMWMB
mBgvTjz0clAjucDjMag3JkmJ5DDIUQ/NYVwOb8qf8+94L+f0RN8uhIuoGwQwTDLjKZqkr1mBwmi+
+AGaBS3YyiDH40FZfW4/QSbszeHAvuHQg/1VFP2k3p/G9gBizo0Sl+qyzrHg/2jwIjdZAzD51Lvd
5ugH8Xu93zCldDYjZkErRsdrSAvyK71k/wk5b09Oiai3qKlh5ud16ISb7FWPwKOFmIQT3WbLsoHS
ZQUCPe6HTK40kFu8Xw+ZeVmogLwzFcb1cQ7LYQxvdIZkzddMP+t6+vh2a2Ii1u8VQEG/DyAVuNEQ
QoSOTK5hjOgcc2QvHq5CDmDN+4k7NfSpRuvDGsDFrlS5ImjGaqL/GkW271ynC2YFOmvypvKL75j0
BfJt5avc5nEED3+pQU1QOum3+V2Yg2imJ907PPBS1REnNYIXRIwzQjRnk0WNRjZnZCXmJIpCcsmr
h8evgTZMeQJoLR2qTil6t2oavOd2FwwqNdtSilSmQURpYYA2OLSAOlrebfA4RO/DxTn09Zxtvquu
8Aj+MMIQcBfQgLCi1F5koT8VXLVrh0ZAWmnqLp4qiVldK58HE1LMg//lgqJuz13epRgYNzS/QE06
DRH7iHQpAZK7Vl5hpqP6G/P0KOdWtgaf3ww2k+E/WtTA8rjHa08YSgQLsDqccj0D0GqaLYgDkg/Q
kYg+/PO95fXz4XMiRtcm93X/mwpxaZtv/LVJ2Grh/HT0Dj5T/GrQ2fFjHULp6aD8GxWqY/3fyvqa
+MaMB1ryVT14dPA+CuW2gT5O3oGxMGUGTIOprL3Du4aTA0iqpNVCrAiJ+AwNzWkNWEZlBE/mQAvG
pXpX//dlj+nDY8KlYHqm8Ho8AszqzOLXAKbyqU+l6/SHAGqgvx1+zN7X/3Rju/bqoZ0mcEhAH61B
TNqt+ut4IqbZ1ZVcIUQw3U79WydFVC/jfOY3CtAnpOZBqqAUSDwbEyoUdZEIPKDOh54OgSP8bMRh
4yRkmJ7R6Em6k0vXbj3bc/9J3/W4qTJDmZ5S2L1xTIf87p+39kHJbYvBAXGf5pPqclpX3RJr1gAm
XhrA6ZaYQw282npsO4U1WasRvpHU9jInfeBsrHmLw0bvF9vXNEHm1BbAp6NxZ6X6A094XVsgpx+X
7trBdSzqeRUE76QtD2Qdqw/MVO/wq1mWO+uQmVsMl5QT1m1F4HbImOuRcCSFI3DwxfbD3JAnocEa
0U/7mBt9eUJG10f9Usi8vPyI8FzrmLSF4zcHC8cYJPvYcC1NsTWW+WvlkNqd2ZGW1Tah46K65bfw
/e5f3qyU6qKQl1AOtWP+L7HpNtvhsUJghsFDQmAttrH5Vrxot2x97jftZ6hO28LJiKSAgCANbyJv
LbQvi6sBsxrzEkkPv5qNH5GBbz3i5LDCOxm48HhYAERI2ERB9ZsKp3FwoUjVT7qSWWNiExxgTHFi
DcLBssSrETY5CLnhsIDilY9FzWRIgznQWFD5vyJndVWo2op+22kDtfCbRPwvvvuN6yFW6OfNqiim
8PwKKeBfVeHM5UId0OkWbSW42WOC2nrOlh6KClvNavkoLz+vD1WqSGTCNsK0oe1R5gxjwC8LYDWT
Gy7FN21NoxozgNN54f+m/NkwvMumMeX4fW6Q4MtcQrmOLdgIhdkmVnVfYgjL4o2K0mHX3/tHFbjc
32pLN/dsd8TKBm391Pv2cg7slhZxg0Z/dE4XfdOe/UEib6OFLuJJHSQruU8Sh9gTXTJd78fKAJLI
MmS4gETqtKfblRdAPylhrCrk1RrPCzxt/fedEFYTt9Ie9p3o2XethYuyEjS+zurkT2NgA3Blmyah
qnImikJEZKz7MJQUGQGThAlp+/kJXslwYBeH2a40pnWIuYNv2Q8elx+KEA1YRCCJStHue/Jeed/h
kRcsTxUSMR0kuXjVWB+tH+Q21KjfGWqudH1LeEwDX532Xn3N8uj45VVvzyxu6jD8lnIveFSGjDBv
jjSoHnnf4091hQF49czk5GwZmdsLgSC9eoF+wpjvNhssOgo+G+A0MgIQA8vL+sVuNcg9Divcp5KY
TXmY3/fx5zLE+gpVNvl7vIPvHoT04067kuClYwWs0Kb/Vu1ygzeScObPoP1G5hMTwzVu+jiN6/xc
zYC6VgYFZCPGV+9LoV9dAixg/nEhPBDntIlieFz7Wsz5EruuRFfCEbG/OqoU/PnA5LziM1Nkm7Rn
eAYt6X1y+E7w+57EHKAVyfKTkUBqFoVcSfqpNw3IFA5J8TeO+EptALwfXOkoK1C+4Gb1LvxMgd1P
M8XgHaK2LCGn24DPvPcqQL4nbzKhuqxJYnXtdax6+02cMO6Ogh61B3T3M6KyB7Nij5k1w1ftYoh8
znNkA9r8lCF4dIk9q1IJu5yFl95j0e9RF1mHzRw4gZpPuKvVtnVa2bWbLTRBCg6aKj+UkBVCePyK
FKyCnqbntcazXbcQgZkQOfrKxiWle2t7svQAsHCmo6XseSXmA0mUOGXF3Y67YarJPdwvOTzJv5Lr
oFq3pMOxx0VueuhCOSDUfRyftXWHJof29A23atsfFA0S+JZsxZqgABOf+Dlon7V2EQ8skQqF7zkj
Gri2aJ+7pBhlHXUdJmxaCmj+6wwj7H0MIJ201EktsqnBB1DfzLxFAuLYPL2CvV4KzcnQzfEdj3jh
AF1eGEOt8OQbrvDKvYkkP1mBXjVpt6AdqvNFQEnyhfap77ODmXvIe26NIFGKWwWybZQfucrKKH2n
S67cWdkIqgRxOytTPLv5vhIMLEeCL8Nydx11vXowyBHm8tTCVoAGx0iehm1fMRGV9+yMvZvBBIbt
KI+OziVSDXzOoKe+Kpjy0tHVqdAUxXsNlUQPa6km4j50oqS/KTzLAN6S8fSPPy3YEgsmpk/Q0bRI
BOGpf654nmfChlelO4eNk8P46zuRZBXaevDWMFS6tR+tHLt0ZnuAU3BBpppdAR/eKVdGtGnNF40E
4fV9cJAKTGVKpwncJqbj7NadQfaAbDEWNpfMKeZzN4dHXbBj3pWLo4cWPqg3Fchus/fqKCdnrEvL
j6zkIQfB6KY7DBv88c/BTwRnS3wnIt6DWce7r24UxqCa65Euyx5l/lG0yvyEEKYXiZoPT8KLQrqC
vW2cHcT0njv+9ZzjtMnty+EUbwlUVHaZMvHA8hkjeW2k7j5e2ofXJtRFRDToqwqNB4rFcfiSyP6E
ns5uK93GcWcrhCY5aA4teAa8+Td6SvGU4OjM8a+G/DjDb0iYVlfhD+xT5Ji+/2sjOZpgb9oQq10N
9m0cfQWzWLnzTPZeU3D4PsomXbDfBHUNCwv2hF3OmujPANcMPpMqU7c/Gb2If5Go+woArs7WTV2j
cd0xylAVzG5eWc396CN88Z6rUZV76JjQpQmdvMyMkaCsZUYGDpKP20jj9BGjs/swUxQOn+726AaK
ORYlkSiQqVBd0BPRKeJt78qtrDtC/kA85b2xRwuA9eOF6VVG+aNjjEPPPCcSDsAz9j4Oo/2UaVXk
ATJLXD+LrmeBUh0GYxRdVEH63b16nlcJ3yWclcM05/ecxGqaq/+dk5xcqZSghzUPLU39q6/8SzYC
/UIlqx07j4CmhHudHHpzRTEKfFB9L4tlr5j3vR7/8biulTgit6roGxxUwbDDiWaBJi/sm/AsrVZN
MrsFLwzpPyv843ch3xBXvXQwqRBtlFQdumQrFrvFYrmYcMYFbEGJOVAVVW/xvdb31v+huP8o0DfC
qzgXEaFSGmK2fdG9mCetjAxVwc71vKyLarSvati11qg3t9wZ7oKTy1LACNyYg3oW2vvxTe/rbYxS
6b9Olicw980Jno0nlHuVigtHPr/l7NvQ8qGBy1DMbqHktUoqmyj2X5+cTJeVb/JVFVWgVZaEkob5
Adgf4zjzDR8XsZSVZjeor61LVZ8lf2QD9PgFVOpBBoK1tj0aHlgePZqalqlKOLjCqRb4qpSp0Gcl
07q8aZT+1kGzGMnn1BoJ30x8o8EtSzODAgo0L4/ZaZS0uCNgE+jz0umgj2G9muWK2KlqMRLArIIR
QE6FWXDfC3NT1sChlHjC/uPJsJ8vZcNYg8dABV8Swx7sdq0aJ2lyP477qC1oTWnx1oqy5Ohe3UEh
NmBIWRI57BWWvoIyNOurjODenNmPEcqSadKH0/VfCqbawJVeQkvF3LVc33lud5rSEefEF2j55Zrf
1MLVL1gCDBUrFpSW/YwDPdi6OwjbQL8Nw2HNhoP39Vyp2U04rga7fVAfG2EWwhDQ1T66+ezg1Wrg
0B5c/IQKAdicIs9AwUNnxB5Nz9CvNdh4JEnNi3tFnCacG43XCtDgVTgEhZkFMnIDLNggtKX9cA9/
R3ZopZm86aC8f/PeWbQFXx+71E1u5jf0Xt2lSH6AW07lnLGMS9Bsw2xqqWlrdQupt2fofB5T9sND
rZ+XOwu/WbyLgiFnSPbEgyMZCdQm9XA98XAmhwk54tzpIMTnkxyvn8zArcTsc6pNfNuX75ZHd6v1
eNDm+kxIpwkPhgQQU415nKaYydzMo3RJTiyRqDy0Yi2lMnBXF86FO16CUc5Lv1K3I5ROxs47OUWz
8tTIFqv7Nr4jV1eztKhqxa99W+ydRzkhIHa8fwDh+4RDnUOTbfiR7tkQA8fKLsC+0hwB+hPiP0EJ
7baRfuSDfqp5xNX0oFksn/r2QkyZf1zWYOsYMkT6r7l9xv91iBShRv75M8ISS+QcKbC3HmjDWd60
z35kbsp7Zb05CWZZ/136VrrsptvexlMMxuZyg6lxbQk1ZkqYY9F/N2bOiQWQIT1AAFSrj/PCxPx8
1BfZUtkK18/sY33odwUswS2G8o+NlBeuS1wOhUaXAxFJexiEM3rjUju3RixlSL9qwoCdAOAzlkcp
LhzIH3q0Q1JMRonN8wkm5v0vG4gp9vJImObyVxJ7BuylXLgcfoWhg5vLQOKMAr01ypb5rWN2Alie
ao+XgorcmgFyCHiCzokHWXg1Zlh7Eju/hwnHZS7GwjbK7ZKvjkFm/+T6iZLtmvWlu5ugjYC55b4Q
2h3eLdvDQeKAAhnrW8Zy+7b/oqhYw+ZU1ogRRoCc32ueEG3VLKIDvCfiR65ksGKpqF/V6UnSWyGT
9KyNisKq+QQ9IAOe16o1q4tDaKVjaMd9cJYs+GRxFlpgOpa1NWsj6b3hhu+HfypKms/jNWc9OpHT
FxnDWatbIH6qrIhqW9dlnrzj2P1xqnPvxRid8sKY2Fm/sam7rEv3emwZ1E02XWhcaOg2AZrjjuOt
AnMGi2Md+x8iUWmT2eQKpmv0tVjuWI8TPKBx0Q8l+yS+r1rLiPBSSmi2NIpkY7oHt704JLqMZzUI
HKV3zs57Ubh0rFTEgAiJSe9CnCnkXXaCoiIp9pGmgsDUjTCjRA/l/GF7Uetisw6WcPVsI8wNns4S
rXFE0NJ47KJYXWD+t9HEjzxIdfvvLBU33mnGPdt98wUhP2Z7lyhxtppeMXQWwkynU0R2tHKbQdAb
xuZiLAFQNewt7wzXiE0yJAlOFSSYlyTSo8R3bwIbA0ZJPXfqIAg2ojJUZsVjROdfx+2WXL+waGrL
Pdrrp9IGsvEu/lDD/Dcjr2ZHv4hnQwQ/JWqcVThGl8fdWhXJAEiPZafi0bR5HVBTaO4getE59ugj
K/rdrQuvacU8v0KGGS/cjUC//G1URgzNIKBtf/h4xUy94wmKCTVUUZz0tnq+y6o4XEMX2vr6qxVq
B4j/JO0qGs5F78eMLJP3OeWgNp3neQMeOXT+4zdWdcAYYP8dIrOMN+QMJSYueanXesupVfBt3GSM
HptoGjgQVzpPGiGz18C3KtBb/pMGxWkCA5kPMoc2dGGQGhyZhNuz69aVWqW6xzA/jd7d4a88F6qi
P6RWekGuLM76/Qa267vV7RsyMmIQU0WRJswMJ6TFbfNFhgeGKJhsuv+0/IIC0e3BsAXKs5aUanKC
UFjt0ij5Z2mQCrHZwRkpGoTHNOQqpsKwZQdwZgQIYa6qYrsYRmFwBdMRROLYNCSfijmOtDQlYeo8
MkpF+w3Fjw3An+F64ZYtLqCuZupID2IxzaJ6nPh6RDpIaAI7pNnOmyrxXFi5I8OJckkUwSAAn0XN
J0Vn7Xp5Iqp/HznAEDBZSmWppp2mQv5NQTrw8kaKKa4mzki+qZ8BzzsHnpo7558v4nMYvBU8DRuL
zZFll6G3HyJzVObXSvByOXkZBmcGlQO7KeE1UaJv2tY1V9Bpl1tbrZWnqtPxQkIpJNJxd+ew+dVa
zpsHidpkbkiRG1Kvjmmo7t68V0WNeKA37JDi3Y1SOyiOgAfNvUMDlDhcflA0zpJVbfi352nwl7u7
ynea+gJQIYe2KH7EYec/7v7VpJ95nm9czvlavbmkQIdobVR4XW5VAKHFmFSeKXPkVMaA7bq88ayJ
obwV4YAYtpjoyO8HNdJjWV7/VG8ni+nfPLeRlYqU3wd8OulpZlA9qCsBFEtoMFlXeOcr4DoxN1e+
MKCaJrczElN3L//jzj662FNNSxrTFzhxCbP+vsNX9CyqP8DD9QpdNj5D32vkdGHeDglOecTGGGZ4
RE02sQzbizyiOBthpaBsPEU/17G1pm0xZ7h5dy698DPNuLLFvJo+k9hs2yis2Dp/nNoskaCQUcZD
G0/I3OUYGRYeuDw4C739DqEkNjZXY0AxtHkzLZw3/LC5PyCMy6HYbkW5I8KTMIA4Dp1lmkJ8vtR7
9qTM97WDD6HZUeal64iDgst1XFdNXansQ9QmnFRGZhl7Erdth/ujsftdUFAPnqits4GCJMu/g0/K
PihS4j1sOPgE/ILOYvkhT3vSQ6u2AnTXwJg8eUq/wS2xRGmIiDy0Tmyq8zgatfJEdbu/wdWGVX7o
h5RmuZ4VNsCclC5h8FYWTjr1XWlJwxEha3BU5k8Qno4RCpakDIRU1copMQzV1ww4lFMah2+EvVYQ
MfWREzS/3iRL00Ffifa4LjGU26wxNI3G/RScw2ajA2j/0cxEZ+CP8d4xZ/s4q3wa3WuZvEFA13i0
cgAHC2Rwbkyh3Qm8xKqBjUx+bQGuXgJlbBjYXGsTIvoBQSMKnErM9dSlk7++/FoI0mPsMb8HLata
xFmwLW8xBbn10j9svoUqlhwmRv6DYMSNk73Rpoz7fD5FYIUjIwr78y7p9kYu3qVEB3z6K7zThzb1
5aPNQVfA3heatoW3zKwExrfyxx++wxd3uddno3kguR87ef3nTZn0ChBAHYxH5I4Fsq9E485j4QV6
eHPmLNiZ9BJubdIRjtnod7dzm1cx4CQi0nndy4IHHgwXYgwdNUWMtd3gcXYoVDLG43t0/htsjXru
b8mKmC+2uGTw9p513G+0kaPlLqpRKzebvmFAk6lR6aqVKfxnyzdl/iaoGb9eqBAKxEmje6X5wYZi
ifWIQ9QfqrTVJvrhK+MmBKt91bCRR97VUFO8EIgM3X9sjM13CPJpd9ZsuSF1zIdUuX9R2fF3yGIY
Dsbf7rQ1nCVV02bvrMr34jZesZXI6zLC+S5+8D3AF/Opt2DzY8YX/8sB3RtnNN1tZmZBYbV2aINh
XCwwCgQMfb6hdI0DVJe4eKd/0aUTmJR6BMh2Gy/TEX/w4nHDxua49su2RVxO9v8mB+ojpDua+sRj
lsvjw2yKNAwzMBtTcH8xxM5ndvULKjjJtOLjjULZjy2uyp1XsAZROVeUbWW+1MlRBuyzRqdJSWEZ
VpMsaTYa1IZhE/Q7/wRUR0pBIplcNlfqh2e+lZx/b35Oj9fca6jJahc7ydN9gD7eZPlHTlli2ESK
CL5/Z9WAHuOqLJYLjoeaN/DFXa3Z10dk74oyxgayCDfMJ4vPgDQYxEqjO+m19cWOyCGNhek/x0CQ
sTq4JmVfF4/bDbgCPg7h94jCmmsfC+GSw/M38NpmikxF+1/rAJlddQpdxEnlWMAdR7TA8JZnBL96
JzRF18ntExNpIUflOhnl87bEYDwEMNM/e8avvpTYOFnSYRv4KWX1hXE4Cxmbj9j9ldNIh+kA0TXL
7LcKR2ilM7EnXldp8KWJMRfW6wJoHnaHLnUu9LEeJaDEfiCmRtR5mmSdIeOu8/IBEA46XCp4km9L
mR6VpYeQ/n2hrWdZPi8fdhWdsMYuwn+UbJkKV/rIRn1G1RTIQx26UY0mZzjIhWlblVFCPGCfWU55
tOVL48IL2P8yipt0E8hk9rvoIbiDL9ic8Vlt9+1iDRS2iuFwlbrLsBKHT9UdH5PD5WvTL3sX5lbt
H2eqQ+cA5X9W73cHnNp6izQtoQajc6ifB6csF+7GFtcbVak+haFG6M28Dpuo+Eic/Xqei0FftV0R
lkLhL0tg82MVitS9b4LZ27iUwcmOdGmIjXLrHeS6LNd4tOyL0tlWtFE/lFFqlra/O09OYLbiiXos
Tu0Mj3LTlxmGvPWnwfCdeEbgQ8XdIaPHv6aECObPru+vWrbWahUUEbyjJ6KkD3WuJUveOBp2EOsI
lXKt8XlSIrY6K9NyQXTuZOpGR9UHyDLqyqRRV5RSp7aLhC3szrzotMkII07uqeC1CdOrCjHfNz0C
CwmlYWmb9NFUQhhmHm2I9cJXXp18J41Jt5hy/8dK2pSFHo7rZppVxHEUiG2+qp1WpBeZoEpjg8oG
u+SB955zkHUJTmC8/a4Eu3fiMdoDUAoNppxTVJfhtx7d6IzqZaTEfl4qzHp1T04mbyXhKosc3jap
6UCAwOTvZ56R/7+HL68vaAhugQCSRY+EFFXtiQfQSMm3bwfvfLYvI6a9usSw0hrh+Wq+5r1VT/SZ
076JUtTPbD4GjRuRxrKUMHN88Nu2vRy5+cOGs6FxnvnpGsrZRTA0mIvJvBQVB5BKsuVoMnCnuqd7
yuiL4UMV2F5O+Df+3BhxDkssrA09JqSfmOVLW+q+xUtvqsW1lesvFw1p6/iF56VSnKrLw7c9zv/E
l6UjpcgYIn7mPkqshB6wJfkyo94255kvYoRh4XWyRdy6FTs45a6uMLw7gBrl4zgADW8CadXpTl0c
7oiv5jqWjOgRf3cFLJM06Q1YW/R5vDRbcgpVmNFavIuPGHnMG6YAPKKkCez2pUMuOPPSU/CuLue4
1h8DqSGll5YOnY24zvPCIsB+vW2E9ZrrhVe7xF/OAsp1PYccVexoskV6b72S8E74zI/hS3RVpHx8
HJPRB0aaGuyNOhEta3b86oSZD8rcJyzlDcXJIhiakBow6Z0Grm14I0AsmPuPvVCoVeJL7exk+rqQ
8pzyksyPqn+bPzCgmrv3gzU8hEZzq8QgUPBKgUJRwzlYFSG/ijvuS+gLy0u0iTrJ+TgT01ZmJ36P
+mAEEtS6mY2Y4tzQ0JeQbfGuVDbAkrt9sh+pxWvUdWDY/ZyTgr+Lgb70C6f888vZ4JB3aspZXsJi
oqWUKT9mV17EBG9nDu8Wls+mnRsCrGbUQt2LqhnQNOsXHKc20/DLlnXbJqqFb/KpuH4cydVVny4h
7S8ip/xv7dVV6iKv/d/EArXmJVZtPa8j2f//5MOg4taaOqQXifrHBQN41kwqE4mOUrAp9kTbnnSV
GXftl7yah+8gd2mZbAQZVGlKQO5z+Ma+o/OzweKmLouck4MgqKm5Tr9spxSZv/MCpGq5Zy4AgCIW
k9XFVo0ME1E4h6EXIltXU4I2kT3DbKQYCoIPIMEpSuMUOPo+2n6yRWFLyz2SWt1LqqFVJghjgi8w
bYiAZb4vQDa0JgHoGYIc+pHr0o8zwPtwN1aWGztdTka27Byk1HlnY4EKX4L7u5n0Fgh09xYGZd6O
wkFyUtHwrk561vZrvaqr/VMyuZjD/R3cIacX7039xKnAEoxdVmybh6r23glmMhGmrB8KQliwihGv
ckCxUcupXFDWp5KYO1oaPs4MtfJ1LuODIHV+4B7U7VymJF0x2DMYtSW4bLSDVzHwFs2wXeXaTWnd
QNr8kU0oZI/Mg2mxv9NgBc1vAHTQZMK44mlU8LkP8WPd+lujKQZtiL/FF2XGzFv0P+3nOWpMi3B9
e/d++CeLDgb1DJEW/uSoRwOm7XdCfAd9IhXQ9ZTPBYlMksOEXUyEaDo7XtrXkI/bhPRKUsmtCaMy
E1hcdkWXwXEmJfLfXCHpgedEhdynWPY0ND1jVgC9ejScjqa8Ovqo5N7TY3Va4BGJucJNIrXaVU42
bbMrOX1zPxfgh8uk1F2JhTeO2zdXxIANIv1MRl6cuxRfE5dt343/mOpatw34MaUuW59+WDJLTitp
6D2UcNU9rVEsz/EmnplUofepighNxy4YD0gq4ZQUfPMOcXGdbowBbBB/JosOuTmuwifygcPLE51G
lxsLySLUlYWhNixygsN2m1m1hZ1jLHWvt7h9LLBEqlaeJipPOdRBXViLYHqNO1g6hihAPUu+nR0T
uXfiyT8ci4PYeHfnFLfd+Cq75pULlqKBLn8VyF3Sq649ah755HhyHPdURT1zo5r0pDPTPCXm+33Y
O/Hi1jOpD+zgva5wAar1Nz/Ezi0xdRZUnsb/ctbXrK/pq5KXmdOJi+iRhDvfKCv93ASg6xar3+O/
/tzguIlQFDYf5ZfTHrNVUw2WXracSS9ZiQ06QV5RzZlxp98Jk/ad5Uqpy1oOdgTNgRVszhaSuj8x
1i6UGH9kM9GqhjSXq5YaBqoklZj1JlbwKz2BPSyMWkCA5M1rP3YptTBi63oVJqNm7Lfs2IlyJV+o
2QnTJHQoTFaQwd6xDj/qK/GDTQsf8q2UIajAxD3Cuh5JCveAT4oZ5F24cpcHKNwkLr8WOWhYg1C5
XR4gla9eBh4Q5eMoK5uZ7Pce3WzXztyoReXnfxCc5gaqqBTv5e/I1+AYa3r495X17MyifHe7chiR
nLFqg10GxEUFQiaMzy5eIgP+x05azIcFxnHEve1WKgyhD8tKPkYRJ82q8UQ9JxElCs++iGkRMO7b
YrZOVfRASD+CcATxE2t7nelPAZBr/DG9CS3x1jLrsTp94Yoc1Pbqjpls2ozl3FEohpR1FD5YvXDw
/GlbrTBuYvJHDN9C6Q3niwHwHQyH0QhavzJtg+ObDERbtNiJOZ1ZNg83J78bAlNDNlh7ybRfCY1M
CmSZRcFaofi0dNNPO2WVibu3Ej5bNGUD/upQBdqFoYEcWT+BSRdCV9wZVktgg7pXqTUH4jMsZ8kb
vw4PvwY2VBU4yWiAh/1xiBFhDLNPvmRMmgOEFgs5UR3PtzW9WcPxWInpbm91gqWwK6Ur8LGcQ5Ha
EsdSxu0IHRMMqPypjUJj/hOOaZ0EBydE0QCD8RRhY5R1L2W5F8uxchRPCvsPeY1ZKbEZqEcZygPG
MTpb7i9Jj+FZ68vWMqw9AsUdevoVqY0v18yoJFLxpNqbPRXvlRVp5/dQxEoya5Rc5ey8rXwHC9fG
zY6cBlr8Dr6OwJsfgys1YTvY/iZtWQCgl6zSXQl21N2CARlxoq5vGCtYpYJTeSW8XgwxerMPUkRT
U++p1xEcrHnd2qtcznW+aclzPLrtNq4uG+yYyHv5l1x704uDIB5Yvb1Knwmq3M6idNt/E9hZ/bzz
nI2qIDzidZjtBk4GECo478iCOak36eykF08TVN1a8q6o8RaJt5jAoJXnd5mxigwPOcoPqmzTx0Z4
nuIXvx7e1mBWyUrXr5YT3VAGtDIHPo3T+66P13ku94ECHUlarCN85UF97QAm0MikrfZb6wX2Tbnk
fvBB8ea6lEUcWd+5oylmCiKa6kvLSoEf2Uxjlm9MsPnlEqS5XCQA2e/yhr1mlrMBH4/z9jHaMBiK
AXfKf8m8bHC9Ecsu/KcWMtvUKnwGW8nm0mzatUrF808Zmy4u01G6Zw9lmEakJxlz8bDYNH8ydBIp
hPH4QDYs/J6uVLMBKP4uZg5AQkuzVIZPfDmZ+7F6GcHABSAaYxQns8BvbItEK6QAN0WE4+pzBRYk
Iuybw/KBRkvs/8YnmYMnlaZl2KfJUP2PhFZP4gRSqR8YVpsMrbNGuD33wgM+Vr2+D4RtTgEmAUgo
jdeY3Juwm7AmqaiVJIVm7KPk5/D4OAaUZ346JwEnsA3KAL9UmHIyGu8+sWTmRYaq9bHW3R4qCUhi
y084TSSkYQiPCBMrnm9b6vHeTe8n40hMavsGbiK/xEfpY8eRIBjuAuWGRVEUn+tLacmzLCNJRZu8
XVQ4JeOpHePD16Gh7OQXDZTxEMLiqI3KtD5y+oKTfi/MSjTYlbOJqBq47UK9mslSkypjjXgiumtf
6HcJTrgz8duxsTd7LxhkweKUrI3nT1lu8jvw91kToKkltK4ePl8eIsZYdXls6QFEp3FeWWuMZba1
HgtU5AgcDIKApBfIolcrW4uF8Y3RkEbfEnZ0eG7ZG8xwvtj1ID+yZP2fwO5iwq/9y49wuoi8AbYM
/So2F3lBTJmkbuZ0VOOyYZnTS3xCzqy0XqULFjNIsLTeHzmwK/jw06poS442xmo7kByFo6nJRXr6
ALnfC8IYLaRH92v0umSuHyuQwvq/cG+yyR3EEPFvAf12lkofSLpkqoh3OPNDh3ht38pf0piqvi5J
GEgAJ4cqcQpjhCIw4dznDgJqiyyRQwBtG9P+mPDP8sOlYJ5XTjBUBjrh0rAbWnH0FPzGjZRWzAvd
yiRMcYFuVyAta4VZz7Qs/vnbkgK2PpSonzaiKD7nH9KRuqK5iMITPtVPMaPkqadJnbcFCB0chAWu
rpDrBxskyYLBaDNE06KhO9gKpNmNC447fnqNypaY7n6waLihcVSTabfLfTDauCG6+AdozPldn/Zt
fgqrK6/AbiPV5CSOWr4Ha2jForRlfoFMv9aJDn3eW1ATDBxnFhmsDs8Ah+z8wvhkthniVd/VomGL
SLo7Ct8kfImZRfcd9AKreedbO1tnBOoY6ly9ynHN/n+IPppHMuG4JPj+tZUgsHAf6EyJxdFHO6d2
hd9SbqIfoo/WA686W7ZrNJaOXW9tVY4brcU/ta1ZpmlN1p0MBwVFicVKA24HWrSY3qHhNd+VALJr
0PZCWPnvKNo68Np2LKdYI62LIMdcj2K9h33yC0pOE3ORh124z+ieUMqmd8qgJr+BcyXu7a04h965
TOsTh+hjOaxSxuSCN8cavp3h+xs8QD2O7wjsH3Jc0f/7TTkAS+Rbe1w3ukRZ+eVcaz6EvR257yup
aR3DAtWm1+5Kb2O8Sp966RPgT/q6PM9RL5t7J+wG6uFeRzgVkEoqL3sAEVZLhYS8imNrA57a8Aet
CDsVoGWAxefuCzzlhU32i7HsEIE/2QnzgDW0hL5/YeE5UuyUSxuN9Dvd44G56xAyp1c/pcIMTSe7
o0l8/U8JrVR/8uTdMjxc+YI6nyIFYCEp0/0npbsBandnwZ6ZpCsFSJYdas49v3dh9s9TGXjQsCnz
cDhrxJA0dAhNrroh5+MwkZvjFuYt2bd2K7EMD8iadDlA+SfHYaTErSEl/mwyZe4tfWCMRhz61kKj
NSJeFUUhH4gwGZJPHgKvEoBB+WPVSlSAtuaebfBZwbUjEhv7yXboYhWrClua/0AE+ZZveW1TVqm+
bry+wiU/jz4kyxsc/AcfhKoObhmGcsRiF+s3HGwkIaV7LjmbosGMnfSjQpfGddGAW9QhXkmG0awx
5Qq3l2UaNrIK1mIXvkhxBPaRYlBppZ/W/6ZDYuxwYL/fzwO8xieVDPMeM4R3FiWioakDZnspi+52
+gTTMoGcS15ZFZhSHL/UFeHHtjfpOlAJ4givXiKl02s9nExf4nXgodhqE37PbKF+DlodOPe2/BEr
yPtVyvzzlxnnwQJRngumzJgghYGWrroBmz9DhHe9Op1qZjmVJWUbD+LoCIv+OwqfLKHD6qIKzvpB
SqOri7T0KigoZjyde01Zak5EP9G+xdPvbnOTd22alr6y6iqk+og4yBq2vFIfPS7VRo/u8JPRb2Ip
EEQtnoI0RDTK1zYcF1rhtD3T7osJp7PVlD6fE+wqBG9VnVQEUvlCINtH5dKhkv2M5aV7LMFeMHTw
RHEyRY9K2TnyDJ+QdT1Wtop4RyXfKeLOS+3d4MT6I/j7ZKViEu2nDA3etcFNUgf1GFDnMYiF4e6E
2bWKxNmSrgH9j1jFjvHqS8Vy15ezquRMLiucYI++6Z1GZtPV/+ZCroit4/i7uiqMGdtRLg06tnzO
orPhmXD4uUg0LyWZ83sIfwravX3+cjoIXIsRJcb6WVhKcqrpm2Scpn/xCxCSmENMIGlwZ4xxeCWV
VaZralEOWO18H47PkQ4R9K7V3yETx4me1bbfxYW/wZpJqRi56XeJa7TVuK0rN8Z/vc+bCx2NOYjD
/nImMDc98+1BI1qQYAGFIztUWoiC3FDneW0sGv6BQ/TdyVKylb9vbK1Ha4sQBLv7YkTtvWeI+bCr
BrIowT6DWxxyS0y6TPRrx+44fZPHzBoYruaciXv3r/MYzKo+9kfGAnsKA0NNxCR/Fyj2+ENwTVKm
nCuyKP/hBNyTWIpWFWFaZ2FXXoI1JE4gSM83kSTiP6iKBZENO/0WLCUnvNG+y2KIYm4B4X/mvP1b
TD3xe866tOwXMEFmVvI4PKS6vxmIkzaGSVycK1wQ1DEpTgROl/ZDur9KPfZY2R83yD4n7QR2+lhG
gf2VtfJSLqNT4Ro3r5oeHgX5epIax1N3iUmssJdj2D2Shiyy6jE39h2VIxLVk/URW1AzQwWZuCQz
n0quQk7LzcZ6zv1vCrI677iZhy0aTaD2F0JqhvnTUrqAfsv/sTIf5JIeqnwIPU8bhvG5X9kx0VWL
QQOKl1oxHa26kgS5VWeHe4vpwqvvOJUKCH/Fuku7LbLNk2IoblfJhZWOi3aC66UJKy5wFRhJn3XG
ra9btzue/IgSVGdRDiWSxotvZjX7bwt7IrdbuAa3XcL5W2yqD9B8x8Wu5Ij6VtWmX8LGoBnSiY5z
R6dYnMu0k8An2Bng1ecHG5TM6jcDEFpzdz8b9S62PLH5hg3wyLRfzlHR6gkj/FkmblNmiuqE0eE8
JXzoZp8FuQflsG6mqt83x2T6398R61vCsW3HHZPr/XYJsaQFS3zhCJsDfj07TpF2+YvyP0U+PYu0
EBGYg30gpxR6LJTwkQK89GSSiDkUYNl1BulT48Utorxtu48wvlaOvKrt1tCQRRmFjFidEEnueL4U
15ePr7IXlpRIYbloaHGfb9yysdfVZGg9HhySDzWpZxnMjuD+YOqmGpiAWsISqkiV+0gkd/pUFq8+
JJ4Tz45JP/tXBa7+cNEZVnNpmIbBTay55R9OsCZOpab9z/2kSg1bXalaykam6+hosfjh1iZfI7tk
ABE+P3a3YebAZJ8O0ZpXHVlGWsxSEzrSsKsjwr7hXhXcM8QzYmRMQ3whNaQ0LKkEK6NbNgNNwRcr
asNhMwbJmhUSvUboxPZFcz3JKMMLyRb1dyjrR+kse/Zhk1Fr0Tvj2fA27neal7sqdit+78ipO+Yo
F4jTsCS/yIKUfabkzN3mdBj6iHb7eU7h4qCaYOYOacvRISA/xqO889u5MzSX0fVxwcV9KLKg4SU+
3B2gXxwZLbPoWS78GngB1GUEvwvBYZQZDfW/HK/wReQxUqklls1usf75fPvAO50GRLJLupdgljBX
GlUZFBBxsQ/7co+k7OhvPVs4K/LSyymjohfoju5GaN/2Kc97bdSLVah+Kh48km4snlZn7ZiRrp6+
M5bhXA0x8bA0mhn/KHUKHauLmUEuDGMxkqdgYSysOatJLMjtkZq1kuBioA2pUzoQUSWsOiHwBQ0W
1J0K0/Gc+UaLUjLlLF8AvLyw7KZ6+Ak7Z8GUw3tyL3DaeZYsyzmKv1QEXcHL5vKZD0RN2LcQ1iHo
TugcZ8bx+A/Jg7rBzV4dG63XWvBKcSA6x5zuXuE/gO4b1nod7riti5Ykts9Xvl379yjofVFb0i8V
0uKz9Bhtz90gk+89dsN71DOx1M7iSqKnj77G5IJz2oUf6w7NLtUHK3FWRB7V//yPWriRLVGuU1cI
ajTg/ory7Ua+kTfD06h+nt2kig0GkX2ka3PzeVi6Ee/vg6IN1h+deqwouoCXG2CJc/N79o/Yrf0b
Fv3zNyfEQ6jhNeg18QDQYB1o4C9Pc3GHSWAG5KdL7ATtNtu/nUSS/lK8yL5so6mX7yLa92449t5r
aOZVX/rVVC6FP+WRueJ95mUy98xjog0NhJq78KN5qIVtPgK8YwcJmkNi1GJPF1pfFH+wpq17uVf4
zrkwvgE+GujrCR1zi9Sm/6Ac69mMowPj/qb9ZNJjril/VRqUe8IT7DlxA1D2r81UETh6KjeI6Yx/
lUg+iqu+ay1w5p62KBi51x5q12rU299p+JlFdnTx8Alnz41N/WlIgQMKZ0vV4EdaVu3sAyjPkuFe
3E8o1pJh9EcyFTUMsXNcGbyXZ+2NpqhrXFU21orRW60p4O6MVicyezG10bY4h2WVrum8J4DyfwCJ
pgB2GH0Cg3j7pAnUjlUuOguhLyiAr7FCjH+ck/rxSjYuZDJIl88mXyIOx42scSvC5gPD87vYQTHL
Rpil2w3+fZ1MuYLE9KrLBUOBvPFsEakSygUHeHSIPtX0mjcGTIP/fwn/431C4dDZpEXxfmt1oFtH
Pn9TPqEmyhCAIyWo5CzTCx6qkYgzueZzWRdjBYPxonSHb1jid1rmDL84Mha6aZq6wUh0W/u0/7tV
CNaTXufXDYVK07ZobZ7VP0bJ/N1VsZoXNRseUk6WAOAW9rOStXfcp2wtiovnn1pbi+A31V+QXJZ/
O7YL5+DsJ0GuBDgWwPMR8kVo4m7Iavna/8cnDIsql6/iybffsULYTfssiaDQECCP/OPEMbWzgmK7
ACyK1QxzjrNfQzqj21IKwqVuaYK3qQc/kS34KLL0X3UQ0rQeJ/NYiQYjRVYDsp+Qx2MzdrQQbvsY
PP6YfHy53X5K69PfVGb2Xml7LHkLus5Pm/E2PMDxld0G0a/t0MKHmvYi+LHRhiJkhGLRNlri9iK6
P0NKrhgXWRKXdVftb0l42t+EAjc3eI9KcvRN1LhdXJ++G60W43v36R0ybXDOobkOIsvX6XW9d4y/
1iykmdqgSrj5NsGVxCMd69pewpiibHh4ayID7FATifssyxzYnYnfmOv1VXUfiNtOLSX8Ky0yv3rV
sX+9fGE8f7EL+bMZVloIgFVCFmmNKj6+kd6o37ZmlprmdRGYArGLGdlhhY6j/torA46kRvjxQCi1
s8wum6xbMMXmp0xcsRs1hg4jH8711E7c07rca8MGasYV4DWURymlkce0nSmmvhcPB6cGcxm45a6H
76MEk+bfGnWRU3aBc65bnlFCxHZdzqqrB1bImP2ZkMLaBfxVbdZAJXNah/pe5KNDUQ0Q2hqneAZY
g3yx/JkAxQ9AU356gz/RPZ7XEWVM4NI7fe3sHnnDe663U2gjtpkACl/67xDsjw2cqF31u6zUdUiy
SbOg1374lTH+NzOMEBG9bD2h2uVcbyHlS+hzmmnydHeoBLCqrSQtOQnidt066qRpboFQ5x2zCOy9
pimLA9HESS8f019cUz+HcK4XWZyCKxBJTKHsOi8gd6lQq5mHq25cRXYWIUPMUitxJVCb3JrrPlQT
8jbQxeD2VUevQ4gqKORYOBrxTEleNEahGlA1bhH+O75SS6l+Q9mUP1YSqL/oTfU+yDjaT7pfEpPq
OY0FlU7NPagqaGOlwFwgp8E1cXcDDLSCAa/OkjOvEdMvY50wZ1INapGZiMgEFXSqpaeBjFOJ45Cx
AFDZRVgLI671T8+VXRcVZloZZcZ5Zhb7qFqaPXacn0DLyRMy+/1Mrn8OeZxZmqxyZnqjtdjcTLeI
UJ53jTiIVoYGp7Ydmosw9UH0A7hVZ9mVVhAVa1KqNUoPlAhEYpAlQ2KxsdS4ghqd/SJ2I3tunUsY
f9QMB+GVIyVItpLWzfQsu91sIBgTZnd2P4P3+EYy6ZvNhQIEHQmQn7w24jl3G2bcq3q8m+HhL6r4
c2DvSg4sRXrgfJi4/EYM0P9xOzTu2AWi0Ap0BUbKHdr4UN/QlvgmA8AxayDa596CuVvZ0UKkkFFY
hTA//mE8WZJbNvaXfmW5Vzb2oKR1WCMffL3B00pSWciqrEv/cbtQikB5QnSd8O+NPk8LlS28JHFt
VgMgnHkNVamkEWYq0ryuHxiE61JHPDwnYJg2WCDFpFFxmfcpgAxFwknYRe/fCUAPyH/lKy0+pZhY
fOFxWf1I96U75+xhDmP3s2GN0Db/galXlqF6V/YDMz3a9YHomAeHZSQ1Yl7D9rZb/9NWc17jsTtC
y/b9pWdO9urOXtgd8j5ZDxiDZy3NdmlZ/K1sq8YDfgBgyZ0FOs71cSxKzq4y7WnwxWA+25faAcpY
56aYDBdDj7DugSYcQW4+I7wQ6sKGWaOxUXzix8dJBxG8fUYE8b9d2EBp0/7qGTH5BtZD/ompITtb
a9UtQ0Ea74YneNrRJ7gcE/GcHff3qZ/re0ZDU4h230MNImhoQRRxc97GJz7pbzMICCrCeOPURER2
2eiFkAXcpXrIVODCA8poLMNuZUgYx23jUiU7QyJro0v5sVqYBhsHGXKiBh365YK5mwr6Ui1/jQOk
XpprdpCd07NLM+c3CilBPA/Rp/emnvP9QWYDEK5dUzixAK0qdvr61nwYxdSF1DuQJPG6TOcG6wRo
9+j6nlZf9dACUTG/HDnqGUpMEfQVFY5FRcrXgx93j1qMFMEkTGHaR5xs0eLkvsxy9b6CRQ3tH9+v
K5RsyLpc3WUtjYm3XqOv8iZYMg3ELUfg2w8iDQsWJc7/YAN2ZunwlHqSmmq+7/Znua27s4fwjOsf
uKe+BAlIDuu/jhdZURZRxIKZYwrk22ZVKwF7oXFUYVw6SvcmkgS4FtVMrDmMVbI6n+KP2XaJzkqe
MrN0fK63aqm+qOIfVEwOWmeg1C86m147xHogkeZk+HNGKf2LiRP0BsG9VosgrnMKCNtq2qEL74tI
cftVxrZaV4pPuMef/5B8c/vYZwnOd94jm+Q6jJF7/gHt72yzJPFZpTlGWSks+K6mcYHEi8x2AEty
7RzUxlTMsEwln2LicT1l2HBWE9wiIk6CKJCh7C8rCfQU+w+p+eYAlyFTLCY9iEv30KerUg8IrHD2
XmCyi0Vii4HFc5PBebOUd3BrKYjFYfyOIisY8jaLRuMgU0tjhDZxTrwQHH/+/VJAOxofmuRbwC6h
jqSmeZaBcJQE3sK4E7zxR4j/GwjgN3fPf4fzw+b0N5xtRAtEU5gVFAUE3nCML4OC0d+P7zjjGpOy
rHGGPCMuXVlSWbkJF75NyWZcXVPgcGiAS5KNB6ODOPgVJXQFQs81SQSFP6AbzoUx5QKt8FHaoWCL
gftGCtXt2Ki0g28FLBd6vKywOw4GsNhGUQt6scpDWSalfajlNZUts5YPAAwfhe1BY94/jdCZ6wKe
zkFnYAdphjbDaYDFd5dji1xZ2CmF1korRlktUhrZtrazbXYFiLonl94oOIS0e9kVBHRSuwkBWaUe
0AB9MJpIZ32eDo6Ozqpg1Q40LeJwpYP/MXQCTpga+r5sXF+QdqThyIlY9wSurhvRe7wjoiRoti8p
n4JsbNv9m0FV6qpciKMa+uvABO7HloqlzNM7KGjDTcodb2dbZJuMfozi5oL6jQmhpVKog8HfL77Z
FwubNT6ZVMPQqMduH6knawpDV94DmuTnlEke+W9K3MvKHj8xErea+uc+4d7H0LDw+xzqGHbp7tm1
vZp2xsIXoWqwWYoOa4U6ioj3bkhY9zdPUms0XkGPO4AL9cXWJlwtyX6Kb+f3VJ+MXXorpmmTGDk8
HNWjkYcLHGNGabo+QJ/O/+8VIlJH2iyV+fHbLV0v4i4Vf21r64s+iw6N4/4EcFvTmKrtwNsKGIpA
0TJVc6eu3pU6ndeWn0edafPUcG8Kf9sT6zJpuZ/Nd3HZ/HpUchM1w6jA/ZKmLmhNWtRuQy28EkyI
SyDVWZMcWj1bwC7FPm1YeYw9dviZgxklhZPCQyIPbvxpQuh0c2WuXj5T9H8jjtwsrrK5ZG3pcGuI
to7taEE0g9MaJkzCJEjs816Gn6I3e3xLf3222XFCi69i4pZxBKpC7HFu1vKK5f5D3v85HAKe5ziY
kOJrCzE6iD8IZP+v+Ty5n6knNjD71+n7aN2E+k96823VpxcViRxnpIybrgXcn7Yahtm26LSfQMlm
eI5H9ZWN/DtYSa6mKPMjpKWHe/veC81B3E9HjWIA+9T1b2FfK/61l9PKOvHgshF4AtP20hc3CvMb
OqbdapWc0hvyOGB6jFcg5dsvCp6OZUVw7MgCyiLsAkZ9sOwXMu6OjHjNcZrkdiCAPpvMYxLE/fx3
+9xPoInobOsWppWXvK8UzzfxY+FdrNQRE+Wt3Z5gFrVy4jbEZK1zIB9oLA2PUMcx8DNRzEYCPgVP
OdEDLve57yA2FK1BBeWkQkN989d54sCzmEyAN0TLeD9sBUCt22WUkPO3m7HzmEQFDK8ja14NW1Fu
oQpExA3zWk4zqw0TxXtW22f28c8+qvDrVbEraxlPDB1aprrB2P8iJdVj0/jYLeetGHooiyHrki37
0OHjqaGuVA5zr9R7W+t0W26E7ux7j2kaWA0cLwSJJjJXCWmXjTek/vQXh53J5oD4swOm1oY7fvbf
O51yMfei5DPionpKA+Qr0hwHxXiIn4WdDcEXef2zMS5dZ8KbIVJJlHueQoy8yG2nS05x22eKoCe7
AW5Pg9QAMN3fHu7qsTCtXtHOtwJxTtDBWZiQd8mBzjE6qLxdwg1B5QehvNonIS8PlFuKclRZ9Nuw
DtxqIcV+fzCtmPuHAOWUeRms0DtzeAjPrqtunq3TF3N4WbDUENeXBlQu5sE3FdYwQV7hxvQpaiwr
6Lzxq77EBApjfSxbX/4q6sROMQEv57OlAmKBmId711VyyVPddcrEOKngzXC2uT+/m1eL5vMARbqm
pWi5dONLwwUmCebU9dfnyaY1zyzMzNAyJTsq4AvNRlv7nWdcu0a3xoM5hnIsSPelwQ4wLzOlr1B1
DIBZg8yf+CEpyJGdHqBqCa+rpQizHmMNLRGFy1T0ZzDoq80BZi5Pd1g1r6351spfnfXBZg1Imnfx
IzCDCGdDn9tZ8oVUTPUljSvWa4oCZcUwZWPLRX3WgnAP1Sasigg9XTYuxTLZI9QqhEDRMv9Qq4mp
jsWu87hYkzkXp6gWD1hx4TfnjD9GggpqamjXfpSeaDSWcTQEAAuRM8rLujdO3FOJ85VQK8mIdsFk
OI4t3ihwz9cg3VaAHbLpeCgtw+V1QGmR3XR5V6VX+I8gKi4p3jehKCsJAFQMmDNrb1e3zoPLhSrU
m8YmKSAgKrjZ5lwkumOkSGUOTkAEZSFe20Atf9FCS/GYC0wgtEGvcrxRdhC1ejClXrlipqgzdzr/
L1bzBuxNfHcgwlHb0JdfHixpwQnhpczqeJC660qlAt+2D257PqbN///yzwyhDdLCtu7FUWt3EAyW
RWTy/E67Xj9BVFsyRAkSF1CNSsjpMlGixEkrR10v7UHdI3+cE7U4yMSM4G4NCx7PBpa96CbhOTDl
1VRSLut58vLP+4Jp2ePGRzg+x9NJalAuMxbJK7gdq/9Iybu/Pn6z/m3MIsrTjDUe7jD8xVwXnQdM
Z50MgbcIYDfublS5jEi2fR3k7KsoGr7Ssi9M/gVm2lVTpCg6JmZNpnO8hk+VMIiZBh5MSk0pyvH9
mfhdkpjLkF0utBfDyxOW7Fysc5HtEWcyKTMvRlipA7NC+lq99l9JhtksJw0xShViVUQc1Eh/3HyC
WMZTJ0wI9TLizRcDjCJaEEKh347PXtMjQRzuRhVm6IluJDqDyOzt9OTXMYIpdNwYNtkk7zYDjD8d
9G4MJUA0LVwaCOhV3ziBMh5hD+t4WG9vn4yr6z/F8qnNrghnEFUFSdTdGqnR9GrBbOiCosW1SqMe
8mw4Pc24N834A4aeTSdVRqFmQADcQx7X9tZW2HdCHudQfa1qUTRjuNCk7mRdbB1SHF1AtTfYrVcC
TlxstFIIrabxhR4Hz9MTQM1HPOG9GHIL//n20wnaWvTtWzckzz2kc+1LFCNy3tBnZGCsHWobwEjk
A/Ivt0VWqD47PVvkjLO3HJPDQqjOtP/tLlRIR1XUjriOqLRcZMwfW1iRxO9ZexPM5N+oXomSKN5G
v8ZKwYOWgT3VNSPvc+ARK2FsiXKJJrd/2OvRCF7xw3BYnv7lKZqgGC5eL2XomhmaO/4XbORm0P0V
d0qbbtEDM4hi5jxCMk+6r02WHlHS++1L5anjIMckuuTbV+W2uYFfZO9irz6DqXJgdk/+o2GGU50G
8W7xoFQ5ObpMD2Qk4qt9I3l6BOvSxtI31fx0KqFEb4kMRW4t41LeeGKggdP9KG3afueMDH01mbS4
D4ZFjCCp+reI0jW5IOCWBCQoK30lvR80ZwmWkokah8Jpajp/MwWNUEvauymv/3oShLKA+vXPfYa2
yfjSu8AYuP6UJQ+1w37/jHcVgfnFxPhk+yzly9h/xtJcgZl/QObpSzi5Xiytc11kPpiDD/1VgJ/I
usl6378k9lqmSoi4B+IpWnDRKWigGquuPYk7ADyDFjy/92ainiaDIKT2RRK0f1AQuDx21fh+MQBh
mP2VbiTneAk4Xx55wGI0eBF8kQhxjWt0PEWXqmkqLZ7ZyfyvYPjGStDbJkBEWnJ/xW0NFg3qxGm1
PG/T/fE5L7/phG7IIqZrDY3Bf54Gy2C3Bi3iGIBK4Dl+9TaFglS+1Oe8z0Sv7NRpsnxYKFJIHQVd
VMaFMJtXeCswpJNuoWnI7Ojv3FbM3KDV6kLjPkMX0wMu6r34RUD8BZ+tXkGnDC6HqzxRJdc2JmfS
axS/VIYMOKYMVwfjFRIaXoEIgVIuTuzYYAPv3vNkfDkIhQliQp/uuiWdMnp26AezqpHzg+JJoMvg
NeGfQbDga/OwUPtvau361Hn6L2FqzaC8Ne3UemxbT1Z4usuU5mUMV+7eCqkY6JRJU7Im5cmAt4v8
dvVpKRawmJwGY723tyuv04wf+dr+wPF+Qe3+qclF1b98F97hwFowxcCMIGcndh6kK5Wten27g9vC
wR9FmpYGsSOW+VaaqHXNrTuxdLBbclYr6rB1zI5rnVM9BrpWUpjOY4CeYLkxyoXyJTK4xBjgXbMR
FwFX5vcViLFD3r4La0RHKmCauvgbfn1bt2UA3L/IhMDycc8KHQkiH1WnmwfvzLpfckITTuxB9vWo
6WhipG1mSyVUJyR9xwYZhQafYnOmOGaqdEtzm9AtbZc7yCoPgg1K35OHd6N0pyVY5teMjKXGltos
hmbIKFynWRq2l7EKFq1wk0LNbvK/6Q91gXPljSTCtl9JU7npa9HaGQfPXJu5bb1XmUnPo2awF8XW
JxRaHufCD6SCMTTCPIzfCqIZAEhXd7O8JtuKkP+IRWdBebgQl3u/h30eZJvkKiJ9oByQsIskH9cQ
2xahMaBnY9x7LEBVJYE8Q25HwcYM48sBuUvmZHdouN7mYUfJcK/LdLw8CDQXq9aK2/IycFJhL9ZX
79mCdpUkCO6zV8o/+OChui/8371TN9CAjaQmC5hx6A9oRbvdRNZDO9Iv+n2YLQuL6t4cvgs/67LY
VTHaPOARwhBqEcxI7MHdeMWWaIRweionLuardhFtap/9rNie42q6vzN6P2e4dTyMRoNpeCv5UAqu
j9mXa3umC2EwYmYLG0ESzjf3b4jvYfDujaqo5PThCSoJwtbsAca3/n1cMS/ciEbTuWXOnCbaYHx7
q62rXf/aUfv/3tifvyXlSTp/5LI1pTLhrxxG+yjcE8s7awncny2/pRuko3F2qQEDVapHbv2r9Viv
h8WxYNN7qglI3lgFlt6/TzsJA/HxKJubsQ2Ioed0uc8FkQae1HZJuF75cw+gvehQUMj/pG7/SjW9
O4CN9H2JmynBxTptfqB3A/fEvuEUOrSblQk63rufaDDQOJATbl37Axd+mxHhvo3+UXYxhsJNBole
oYZ42gNjz0p97Ak6WcWLjiy6d+CONbk71SAzeLn2AWw5n8pSUXzsnvFzJCnCEAhwtcWwVa+HlHTH
kyzJTpwDWt82HR21v7cOIbud3bbKTxumDYrY1sTIH0t248+eAgVCsYgq/StlcxG+Szbdwj4KWXaw
evv8QqmOf+66cNMcDzNfyyOr7VJJTqeNHQR6QzfPIHSr8JyOsXSzagwS8q/aSb/ZM7xZvuGv4twL
2SwyNjhGaBoxqac8Siiy0KREYF7/01YRT1e2vrFs8JDSCXS6OR32zs0oABk5SXgKntDIHOu+E2HI
ZUzDp/QC/+svabS9IT2BHYR32tWJQqcWN9kJ1EIm53eZAHCsCvWs3PAwwAVmSiKh6fOmjsXFzzqj
3vzCaLlMR+abjSxnVGu6Gcpf+5R+D0hP6+iq4+nOsTMNMldG8XeK4UVrtVftMcIjiIx+RGmwZzFw
nsFC3qbR3r4M7L+QO6VIFApUrUy4cCe8c4ezMcrIVvgt5S7Mx9PUf1zZzROLu4GIk6ngBGLDmmpZ
zmebBCUgFrcG06Z2OrNooRBZzNQ/cF0NN9p0J+00m5pdt1OV9LMXMopA/0+zxat4mK6uMeuEp8mD
Wg8AH/0E7L2srHA1J52HdSsssPAoHwrvPTVQo6wfNNQDV3aO0olEPuT0VmSd4WzXPpmqvyPnMTSo
t6BFghXLAuL6iYRnN1Q73E3KCxCdVc+EXZ8b+u5Ni9Xqzi6kCxHPNGNq58XuBdCvzR31s9/Wjls2
OxYna39buHUGHOM1T3U5FBPWQ/cn4o1dPilpdkbcaNVTcb69xr/XVN4vxV5GImI7t1qYxipGpXA/
25QVQssEw2azV76qCQ8Al6RpYDaU98cHhkA02HXD/gmOufLTRSaf+o0yf+fTDhxQc7jN9xhEcZN7
sJhrxx6nX2ZBeVBdYq51GJZ7r311k3Pzgk7Mx5fqvZG2tA7ZL4mX16RB3/gE/H3sPfMfNdF5oIOO
cim2x03pYsgscGJLAngaDFeCu4SqUyGK5NXDxzFdLoyb5vrzbodmdgUp18G22KhiYL0Y20MaXT23
F3VVrdtJ7VrvY0P+ehvv1IAwsYJ+esEHz1GoEer/OIeYZyNpB5Ki0crbEdgZtnm2OQWOdtl96tku
hDA3tlb/qHuP/GCItcJQ1HaVNe5aY4b8w4Qqbeht1+0SjNlQmlrHQ4++T9iLi73+8RwapLKxPDTr
GmC0/2XXy5OVtCNWWQqnsdF+o3aN+bD6iu3IoPGk9flNW0dePj72olVZA52kq7AXrGq30BLQOKjt
Ja7gUH5QELmIMMdVO+mGsiKeqsxgIu/nmqvK3Ui/xLkbusyt8bgM3kqTCtGCy5RVs2irt7iERnA2
32bOqBGEa2on4pts8NwCo0KOLsEw5IyZQD6evUn2u0tX1BJupwGfmLZInJJvFuyQt1047gVxHHxR
0WSa7q5LhXTQtoLWBPosu6SKMo+2hIX3z0VaeGq7G1tYQSNJgRJD9M5SUKVNTv47Q7qjhyBtDTwt
E/RX34ljRmnUpOjx6mafthz1tVTc5CH7R0GS5VmawzcO/LrRb/Q6FN1rZy+EK8Ycl5D1fAOq7edH
mmEQGhpBTuxmHdayX/r3er63m1qU46gv4jEJ2sE0y3HJNibEvt8Eu9nYL1qjRLQk5D8kA9mpXrvA
qs4Nh4k5vLTM08TKXNV8MoZ2zVdxxFoDWLA6aiZuuZ2zJmHPi54cENEYV6Yv/NvpXKCEW5nv2gcI
HrAZo/287vyAxPPsbPnqX6RZ37WJI/GkVdrcRhh3ufKap0rkzWRaYtid4/NUB1T71fj0rDODznnt
fD2Ba1sjFpCV+xIuwYroa9XudAW2ea5LHXPi/D/jt92ZvvzBgP7r31TCmnbmbE+tZI50ijr8tcZD
bBnCnkjabt+hV3GEbUA8O4rF6RKjZqIDMQlOTyIXmZvTsLaajkoMSDLsrw57J6LJkQasRaSa6kmb
DLMPo0vdcfV4Zq+ruxjIUwx5uqiGlaicfC2enDve1VQTJfnAS9QYsBe2Oous95fyX7/snSt5k5az
v0bYeJBdl+VfWtMeMc3Wu0nJpJXdQMitG3c/OT44/cZr2/TCDVH/fyjc8/2FHbri1gIfx/FiUjdv
oGdWwgesP6a5Lhe+RYscmMX7NyNVOzwDhHZqCHNBWA4MfWP+sC8UyprXlZRn0KYJ6ZGAB4MRSyWM
JiBsaCvaLzPv7sTSvz23/8ybQPcnq4+8bOH92AxA86CeVSSheIoOkWAS1lN2phq/qUuerAYWH4Gc
7qNmg0zD8dZMZP4AwM4T8QhOE57XCJXEIQ4jGCI/vZwIQMB7BuVqbgemCc1mcRjXjff2bdpOy6Ns
7Y7ROPhDtC0cW+gS3py+VtcLBRDQsS+tbgxPMIRuFRjXwtlgf8XEXJ0zakj2KIyUf9t70KPEhg2B
TnPHSmFqogLJub83QIdqbOPx2Qnl5Y+t2b0UjKJ+foLlvNhe/qBhojy6R0W/13VGB/0A9XGhhddx
X4CWXfIBgn84QrKiq8h7BbfsbHaOCDMevq+F3+HbYG8DFL8y1HyBkuVY5urAhADfiFy9CmVWfMhp
2LLmPt3Wz2LOIWqbUmha8KQlgNH1keJNF19TmFE3wbaUQQpBzqxQB8QdM94sUfM+veLnRqcNWHFe
k1KF9FXVoP0/Z2Bit3Kmg2ArTbzp1yIzr+O+lhw92YBP2vzIsu03jc17d1TDTOMqzsmVEQg2ftp8
9WhS8UcRwzQzNvTuSqAx1pvY7fdvbYzaqhktQ/o7OyJzPAsJYz5akKHNL6eYbcJS6RzASaxH/Elb
UpJre6egB3jCzd5QFFwCro2/ZYmQsh3WslXR0xSIxa1+lKMd0gKE8J8QicUcHzWiEGjTIxJexs62
k8rLxV1ryIpR2PmNQ5i3HJdy9j1RHLKqyop74FT/Y/PR9TCqdNy60R8CU3MmkONcwOe6bfu2sENw
hKwAPeu9aUN7aodmE1+kU0Jvk3MtM4KbmWSjMUyNsX+cvVGXl/buhIdU1h4817bJzdq4/1ftqa9P
cYF2aT9IX2fEA6DwGBfelHjbP0qOLfoltm6sbxV2slXurCXxm/Ta9u9uesFPyFhcGokV2KkJ2LuS
0ODgoLkdqzcSpgGvcjmb5qwOKtV5BXHGMpiOaGDQztCf5IWCfpO0iSrkKfngYYrhgmMZn02kZXOB
NPU960vaCL651egAIWLMacNO73/eExb4M/JDHjKRwobWmcmF13ctPecKWS16UVv8rf5AaUrEqMGp
bGn4wboRTTng5fjcmH+RblrGphvFg5iti6glF9upYNXEnL5wiXOLS1kLDBfCQ2RAJJvNFevJNUvh
boYTscf/gA1HiyDNVI+UviG1+gcS4YuLmZ+86AODwaEzwJy7yh+qDznu5VZmVLjkQRMY56u4B3+5
USwZl5ZEfeZqXr4c9z07a7L4vr29IxHneCsrE51a6lIbBg0hUIBUWbaTiqFS14iT0Q/xIMq2qJQu
3owxH9NOejJMgJ77PZPc/rzITV2RCiD1umpXZ+yNrgrk8IeZNuj0+7ff2ukBA/J2T5WF163v1FIi
lc2kh+nD9uxoMMdEUqIx08FrwAkQzccF1f2aUvAV8r1r4Ge/9WEWoBMUZpy7dQGWTEJAmOoSvyif
Z28ciYA1DLAyY4ICHrkvEsEXmALPrvdnCHf3aNoLb0kKdc8PNIBhPQxKzIU0a5jthPYKDA3d4JLw
mKQRZ5k36OFr2TUYYaU1NRYFl4J0qg5Ai2INqF1PysU2LDQt+e+3AE/j4joucl72KxYVCbMz76pi
X2T87EwDH+DKQSbHWn9TLYNGXDb3Pk/8JpzXIa2r/xg8rycVlQiLH160eYEwCadvAhGQ8CIEjy22
xIR/YsOgOjpNwv9zlyB9KREuKViFmGwYRpzCqny9D9knO74aNg4bEbl5dQaooppIiZj+9dgR3UWf
AGj1OpbYD6YfOPW2OvAKmmlwvsMd3wXXeECalA2YakxURVIaUP9X1wUojnAh1BDsrd3PoeoAVNm4
Uj58uUQhNCM8qRpFEXXkRKqc1WocYKYMApNx5P4pdDuJBx3dGaLqN9suY3lFgZiHVKIw/2kEMuEE
59ZoNPAntc1Zj4OjhwzLGkPmZKRwirL4n0NGj8jQoouFYpVbEmba0Kh+FJtkVEe2AdfPLoLyjeUh
u2HUY0tBZzlAGSHryLzx3jWTFIVl+gV7+uM6spVfwDkMb86ZZfycEv8HtVOM5o3pJdOZtP7kt/t9
uhLS3mcq2+2AbhdhifWRxxOfKIRwNVa1HhbcH7vbE/2FOBcAbM97cOvehTiuLZ6sD2pmt533kxiC
PYkflIvKU7+ZRvvozrQ4tOFsIoV4lyEga+UdjzZ8vflYVXKgehcP+0FX8gIkAUQeB671I8AOzGnr
7LM1zJaqgLJV3lHusB/FbgYiN5EItOvU8Pc0C/FzDAS5Ti32k9y9F4t6QWxnjVH2IEx8dsJ8y3uH
T8QeeKr/Ws6ai8jTPeirg26uHev/NcfztaqdWZgGxlbezVpakNxdF/unUwTR/jgHoa73zycIK7Ag
RA2GtI/TvylVT5QvfumDMR0TNks7PK8qUh4hQzdpl+D37APnh5YP6Tcf6Pyd+cHZb/5IJAQdFYJ8
VPhkBWDuM7G5RubusKMIN6yJkTXZObwmjHQBrQJNw6VJvMCAZW7aZJ0qDZLvYF6chBNPj+ztdPWk
Wd7JLmmo970YeWVFb5Cez240NnKDc5Q+/qc/ZsKPSBVSYTRo8g26rHniWnvzWQIFbRZGnfRiF7Vk
DD366fXUDtg3dxw2tTeC+6/zrBnTWAG/Z7NV9rmfp9CIDj/jdkwhMJVIo4uojrBgOeDf+0OgiBwK
i6VkxNw5vVXTybDxCjrf29zuF/hF0rhMT6LEv0VwRInV/JDNsjXlwM4qRNgxPJlO0ZqZqi/7bzYH
revWjFORDOZ0zSE5mGhkR1uDX96b/vl7ZUhNrCQ9yuDh45lFhqz4XH/CcZVg4AzD5v9+AEwS40gH
pDx8Qy4r7/Otf1VxwpAJaBL1mqfn0lX2hpulPe0JK9icreoVrUI96kH8PpbvixEgPOPBjj+YbzR3
32ESv4FGY9NbUFc+BF0rZqD7YYGEOT9Drt21mQLWeiMckgCqFcJlpu6JMrRGgZEwiwZx0isGY0Vr
n4s/VjhXlfB549tW82Rbq+5g5GLoc7y1oTaIr6/J2JvOl1Q7TPUGUpNWn8DeKHCiO+DH6QWm0qDM
P3qC1geh/rFnEv3EVCpvoi8svdom+9amPPL28x3rhXcpUZjXFpzN77GRutd1D0eG7wZQ7IYkWMDa
GCEaisPrOnCsBHs3dt3nrKe5j+scPjTwfchOyFF+pInIyWBLHkdd4Hu1E6unrjBFKmfOakYt/kDi
yvxG6Yq7UINN4O69SLeOSQv0fd5TeT5GtcEzKWv8uK3h9eXUdT7mSUJYT/Rwfwdke/KSlQwGniN4
+cMrWBiBKijbc5gdEkCboSJyCg2u37hSx4SbpIoPlwFo0oaYQs9e+mpGRIK/V2R01ZMSxh8z3qcY
V6MYX3rqmZj4Ka/LPItevk3e3SytuxCCIEIZ3AgjVlQdz2TvVB75Ir4ElzMa00LkMqYBaYLLmNJG
JpIdEa7rOLo01Gt+rEGOcR35/PJO87IWSukdhgiVeACeMVbVh++vgdRa28LJs2lB/0yTZzLXNeXG
KI5py1cbWxcAff5zVrAy8AxsdJ78r+zoR8j2Xgr0PtNBu5crKarnsGnDWbIbYcMIwvSGDbfhrcRv
AQz1HeJtoZDU8HTDA8ccc7FaT1SzmRwbuoKd31TFmscklfmoVBqjNr/00UjjWolmp9kfLCumhZT4
pBbyDj4CVgHMC4aIeUZmNVRi/zoPLLug+SzZubLic96JQiJwk9T2FfCUVbzq8mpQwGoZsVjD9T3y
alIag7PoXX8DPoGvqacyD6NgQ82b00ai7VpSf3WxgOdcPGQrxwF2ee3gLrLhEegvjyGsX5iWL72i
+BU4pkz5ORHAPwKlrXF/pQuAG0XB5D8mAghlZfCzEh7PGrqNWoTfAJ3BWQLu+NF+GMN0RojPNLnb
zlIgH+5pDKhMa+9jRVYurP7ZDYKYKWEMHxeLEDJanfKGv4INtXYjKZTzVyoEa2MKaJszrSTjCFyD
66bPix4vprTsUqbNlpbuf1HikE+UwluOJ8ncea/0qsPjzv4wqQFr3Y8yO6imCC58MBAh/WaOeGFo
HLntwfsvOxRz+3Z31dVxor3+28ZmjFq8o7aBur7F+dUMrdjOEl+2uqTn2viZ44KVY9LGsMvlpa1L
3/3CJWyR9ra+SbveOMIVrbRbvjq72/HyOkembH6i7tAhNgnA6NMF7qGuk5baYDNPG+YoRAEv5phX
e7GF4otZ7WDAo2Jaq5JpBzUp4/WvrxAfgezWARQwWG8jZ7t+obAa0fyXVYKkmZ3P2SHmOlktqCpq
SEj5GodYRyrOXlMDaRaIFE24w/xRVGj1kXPC9pYZeW6qROZAPiADcZfklYo3xoVLXpYo/RWfeM0V
stQvG9OUUdThKnYaHDtqRUG5CQxvt+2NmrFhaYciQc6iEvwY4nriZ1kBCl7M+t6osuI1OdN15RH8
UZ4SoSdchAYTSJ5BEIGz/L+B7lunDR22xkBVS/yzBKyK9xYIqyN4xEycYlozRVMaiEmv1m/SDo48
q0A2C4FvePIG+8YlzrnGe0iwZIYjzjpKEWeCuktsv9Ha/q5j793qUFYEuB1xPSvqXpr2XsGTtYoo
2Q+dN03j68x1bGJSCJeKkrAmdxliA8QOQ6KaRtKySkDSrx9UuzksDLBAef7kV7XU61varSXFdYYu
gdIXNzA7a1nrFsCvvf1loaCB0vsmVq3jIyOHCIejGvETRzuyRdMGrR/hRwmMpt9DJHG7T3mPRYh9
FIjwNHpoe4sm5dsT6JhrLP9TlJvm59NqRxJGesPQtyffIMPr1FV1cRTjnjtlIlQt7lk4zMmwzTRS
EayGZn7vNsg/+f/sGMtU0oystj0hnWIufELn12DoivFJEzSfZgEunNJbbjRFiXtmzX61X8ruBbVM
6JsomOHIA/xCoDuE/3bv0gP53HV1sFaUvRex/sbNt03mM+gkeXIprCo898oUJOw1xOSblM8ACpwX
hS+mDmUF+cNLqPZ7AhBIi+3zwYSNa2xr5U0MlHA3GoQCgJAQLuBQOdTLtzgd+NZYT5EGQyq0Yvzs
7eEb9g52o0xhZRoKBCdVP0qt0ZRZXqjVZxeNeZHTdBPQABdz7Fjgdrx1E4sI3PFwRtVmt6nPwIhu
ktNdB7tBDBKfd4V35q8aFIlSeh8bsTW6mdPlhD3Ezc0V4CvP1SxcTNfHurlZMR9e4Px/Fl7Dtpky
1tBdzLR0SOPBWBxFS8aN3Yqv44AhMMtH0vGulckxO8VjBroUyTyDzOlzb0f3fZsiOnIStx0R2u07
ebs+EtqLufLXuPWrGE90Mz0nRvbHeQjXGKONEueTujpT1AneewMkDi6sllQKyeXcIKEZBKO3gpnE
Gnse677beJvym3NfgrNpX+bAU4k4f5ay8uslhxCP693eH0Q7uFDx/1i+4yP7vTHrjA3CywrqqO0q
mgfA1/zpzZDk2b9BSbFrq0ovr+mkH3wQUnsUUYV/vD5iu4x51p6di2e5SX1Pp8u1P4Sts7HSvAo9
rgTAxcDiagGtS9baGLM0G0TOLGDim9BGeQh9MUlHpCTbjY3dfIGiCW0gVPJHvQ7r51Ycco7rTecw
keU8eebky1RR9v33q857OTrKW2dqd+w1sMX0XMcr+iNyWQXXbU0kZRvDNORQ6D+ryx2O5NMIyogI
cCBLJwV+X0R2YQcaeXTmlsyD6ckpiMH5LfXHd+Dwx7IrJySslS7iNWiOaplA9DtNw3EBk06OEpuF
raotoVCFXZ96YCzy3tDKNdLcwL4P5LDRlT6UpZIRLrFfMrAsQJvYGU/Dsp+mPlkbsHmbCZx5HNWn
S+aLP5z4HGOTkc7t4iXpphoGVbA4ukjbs10KZE9PTaWdwC32/DQKqQwsuSV3qODwLqVdsXtL+qc7
64PeCUx1cmYQRDTuYr4uPoI/UUDmnn/rfdP9O5O2tWztvDOAtehlQpNYuUIbLBbNv6WwX8kHF0DK
BPad/Ve+3FyVMhiGyE6JgMuijAzIkHv9h8/yZHFg/i5+yXOYHp+Dy32hmCvyRAHMtQmj5F8NInnQ
wfoUdLLDniNWnNvNa8enqDkTSS6c3qPX8cJpf8qFwhAsGP9dKplE9bTBtng35R/t2EAvab8m7DLg
/+GxC9nv1avR7/h4kkhWHK5LZtzzlTcmr6AHKgyhs59jdwfUxiCeDRRPUjvI1erGuZXMO23SLGWf
vfhkk1saaNaJtoHUrJiOGqs5r6tfPpm2UDryCZwPPK9Qy7TvpfNDAQ/MIVjrAJvehyT6uXrR3rBk
JCCEobhR7hRTDb/16cX6Wyp+sAc+ehSNA4IWcq+YUIBmNUVLhkHCsYT7jNDaZeDjntVFv/ZL2486
4nvsQH0WHqchcHMUQpQQXdX1Qq7aLxQsf+9n3PN5ZQYIuz9yjdvbnrB4nzckOpUB7rEy/knC0vd2
BQh/MWINi0SxpXrQ/11t2Ozn9o0YFX+7T6/5n7kMNJBTQC4uMJJ/J422gg23QRoFFvUDnKoglDxS
5UbwPQZdil2rG4d8qGMFyJcV3lySZOWBtkAe1l9WdXDs9COhjYHdTHwJl+9DK3bOcTpD1tWMjvZY
j160g1GKG4sDuh99bZVN50Iwq1e+QdXHgSj3Vtzi685nVonp370i1ZFo7oMiSkIwy37zhOypRSBS
3Allp8Q/yhbLCs/VgnTkyABEBy7VOHObXLw9xHIxAHgC+6ZkapbkAiY+YYljlUy8kcaQt2/pbvE4
MOBCtWAOPgXA4BR9t/HjzL6w2o1owQx1Olt8kR8x9OeszNQaJLRfXEypq8ng986G/hXxq8rPkG6p
KUEW8irxOREkTFnLw3vF4sJ4lixZqWgJikQ9BppxmZcJSsBgPrJRNca/gPsXXDg5ahzju0CCWy/m
fVJ2Nu8bt3kpXgjwT7I03Umph2W/xc4SsdMq0SSYAGxxX6nqBnXGVE826naFIVTdpHmTfNMbjqE5
9qoaOzOXfzEZCNbEnJT5nqtAHj3Fw+DX5bS3u8Bi3rcyXOdPtGq83NdT9fOFeNVZAZ4xALgJV1TD
xMRIJkANpMvAYcgzrwLUYRaBYpPph29lIoKh/bLMLS9UJjjaoFT1o0AjRuaR6uLyumTmcYAf49El
ot12R0ZnfCpiwnlG6zuFl4wtjRmWHbKgAXDYvISzLD5ij4bNGpsDqBh56E+kezRO6QCvXcnvcph2
Gtb70nCPtxNv9Nhn2oQbBCZst6wdtm0gmgL8cDaz0xsOhr1hs+2km/e+yprs4hPJ12KexF3HG9NH
u+yJRfe2AOqyu9tyZak7vmM9xedgQ/zUYic4aaQhGSxR2v8zT1jLPPrr2TYSYneCpMKym4+1vgac
+SInr2Eu47tO2ucc1lSkUsbCtZL48PcIKDcPKaNlg8pkBYlTLJEf74u0lvUW7h311IyhxJz83G0E
iY4WRMg+03EEauPX3v92D7zo+yt3YnMF8bNQeaOq/pwEmuOPqRuwMf4oTdnzXVhk86oPCkIMcngo
m2VNQc/M9kQke/vzqLPcMn4auYVI2ulyKjwL+R5aARrqrL1r5IXuMrg9UXenHPqazhl7dYKQs29q
Onwbdm/LTbZeXOYUocgp5Wlmt7dWgwuc2gULrWRw9WXa1GbNAsvB2p9z0heyeGWRnxtjd2Un4TZO
110uyeBQHEqHgqu1135gBSGtwGVfNzRFQuujhJWd/jB9ZOg81Il3lMeCd3DaTB38WkBCx+sI6SQw
r0QBPxgMZC2AqjuLGTOLqq3JH1ZCrDDZudhGGP9a9Mdt8oK+K4qxPyaDyFfcW/XCymnXN2Awz2NZ
DFpKE4ZB9LwLtGGQsCB9dTiR+VuXv5BddXKKOyPnLlbKOzGzvtFAwZI6j6rCaFCkfRNMyspxil86
p1pzj2Pcuc26ZhygnY7CSzRbKQLOGrfw7AIT2RVVGDLk8owJtZwfLqIeZiPjvUVoTZDtvXxyhmdk
j26JOY3MY3gtJw4Dnsa8imtv6ZrRqvd4hnKL0xQYYQ/4meEKWxe89lMA3wY4cERRBmQbVbci753N
Lr9Q5wjM7tNwOpwHrEhJcexTd7qrxFDs9JjXyuMJhteRv9axTPBOh/vcpDpTwbMhbtvLWYwy/GA5
/Gyzlf8nAPhWKswSWmskfkP6GdQ6Z+YcS1xZyiiApdLcqwkxpe00/9HfPO+Kod8+mVB3+ijkjm3/
uxHBx5yB1WG7RHTMzW4nnBfRAly+elt6kie3nn0umVt1U6Qe6A5VfeVPWbMVZqXlaFtQj/mxGltm
Gf2StiARP/FQTeb1yranQWA7VB2b7pkW6AMdrZ2H15jNNMlq9AfmYf6vVWOTS2KJtpKAsdXBHQPo
HG1NN9ZlZjK8QkIFeAxQkshePiMk+8Jv5KVPBi/TAsloz67N8umZ7miYrurrjG74GleglsCcHGU/
E5+Wsib6F5na3DeUzk1jLiJE1AoOI5KUqVN6UokVIN0RLviKA1SHejW2gBB3Mw+226tKc1TLxTec
a7NAVtYQbluCWL/sfra8R3DCVZk47c18tloIyhS6C6W6yTvEw/lCjWPEo8mqV5JDwmZiw3DLkHed
b5WaKqYVcaDB0Oe1V+4QyfLGwO72ik+bXOIdgrgMEk9iqOoDetmhYfm3abWLdkHCKy7xtcdxTuYL
aO7tQUyF5dFIwJb2Fmn3HrSYKVV0WMUZwu25Gt8lZS3hPE8tE3LnvYL/hKum8lNCVbtl4YveBav7
YLk6BFr0jC0wZ0zz/eSHugXcdDSSWevYslkf+0u26aJJO15TAqQRQCyJjdxIxFZJUCaLoWo4DNWa
NkEJWNTlgJTzsGOVX/5ih6sNIivLyRv6MK6KPNjB2dVKdbVejtXvEHt98zLUScDWdis/pXNUCmj/
Nm0XtEwapRdfhC5jUpVAyt5DkI9ZqTvOy7RkIYNn2JUcT9t8sJPhnCZI/GXTOLUVBC3T3+j/3FQH
cjscnY6iZQ4xmxzhImyiyq2iUNOW3dbiAR61TuggGAAcGkH0mOfL0kc7I+6/IfmnboWpNBlIN5XO
rx0ZUTaTWyiOCMXoFiYlZhkt80xkH/yeU4XJ/3zgQIvYzVD8aEcH8SNZ10N5QIVnGfoVHWTkWyVs
5WOo81cUSqh7pgSTSTavS9O2a4yi5f/Zj74flVtbTS2kluQxaSRAT39nzKDA2QcjliXZTwR3OvFW
R1xBUa0yIts7mVm4caFZqtT6tZBtg4S6sEMTVgu1y6jUJdWE57Mf3T/HEJzSxKMpRO4XCRwEmPHR
dOnDNzTNTJ/yBqKOduTl682bJ6zxEmZlYNEjh2tprSMhfs5TIrQNOEaLmexW7sYtAKebxgMlsKDk
QWmnwLJpYgvg8iJ7Ovxz5RcmAT4UQ9r86KA59mIJeattDSwyQcIjHeoHiT9mmy3FSggiy6NcfXFg
UD8RfXkLFK71/skjJi9evuIaD8SrbWbh/cTd8SK8BE4KB4pwqlKeKjVDyjS+FB6C9nVyoSl3EgcF
0XMSwPFl78ctrbQ10tKSMxB6gjqMKsHSGo+hNttxDlhcIesS+u5tfE/OVS35OmLdPlql5ig1XZWz
+nx/h2MmLGW2RKRvnKOJjZgcvRq7VHjRiIZSWnzEQRGT3kKBmcwGCFomZy5LReWx2+ZY0DwvbLws
Sxpn2xyQiB4GVNlji6xhuQ3DSol2JAIwHKYVP9veBd3GtIyUgDCaPWWyUSmlDteKfNnQUVNyUR2n
AYVGb/BcAhDnJkYB9LGB1yPYrk18jYbihv5GBB2IvgkJ1earEHGRLSXp9owwhrP048bXGp4X99kQ
mePTRpQQ4qzohoswjaNXUkUclBm9KasNkA+2qqVInK9FNSYFca2/Ex1OPCVESMx21INQpkLiiqZs
Jm5F8p8tWgMm5xQQljP6+scBLfkh8XLIxz0VsEZQPGFUZrdn67mU+ufHV8TVWAQnJOBqJCTZ6ntR
B8pBiWdSb2T/Zv8ml0V1s688jdcDhEmc4NVQhapiRXn+/q/2KAYUSpS8KPme3D+lxk4WLRZDqbGk
cISxLObL4H+zEO8q8Ocv0+dXBfewyTCPVqtsTKUIKCUeu6Y87jKXO1xpflLf2gV1U7G9+XMacqOK
br6SHa0R1pHZiUSmY96VYGMwNFnhQKTpse9HFda9PbmC3uXJV7NfFOUfU8XpaVADXK7LV4J62gty
2FwdqJ3xZ5HriDOoMsV09lmU9OvCNIsWioNKWd9JjSXmC/DNjIAEkL2sd69H6jCyGsmv/T7zufY9
d1YowgLZ8FbphgI1rwKLaRUPZ70RzEMQJhGjmyYNOXWRiQaYb+dg9atlFZlpHOYc2YQPJqtw6cja
zZgVacqmL5M0chOvZ68Tq+wNMp5pQWDiEx3LNDTpkfW/SddcpImt8DR+gYdCi7QtIS30cs7KWhp2
zSYnMLj3PFIvP9dbRxoeuXdufQiJsGyyYNLhKn5LQjK3zY+HrFulhOVuw3ejQK/JEn8xVaEaW3ba
WmOCcHxcTmYLorVI/8zrmvdn5JlofUiQ5iXhEXjVi82UxfVXC3AXQr36rGyxvTgu54CPXdWmUPV7
leo6jpVbvQgLJ6tdi+/iz6mMNMDKO90u00gmbDnWSUEIL2YhX2epnX10m7Q1ORHoO83P1DNUEWRp
hgXB0m8A08Y7GHB59RrQsY7fqPlWvUOPqvov35rO3peYlhRTQIypVZ6Bf/hDm3oR5gf5BZ9iW/Nm
TUnHcTevsHFbNhUnovQklp4NodDdtJ9Yl66f2k07s/cdoVISSzwY/m5HPf4gZBTPk3wv7sb6VWYR
MTJLS9/8KNx9X05+3Srt2CYw9j3HaMmAQPoxtSVoln+tVB6ZpODqzPBPQgSOiggGOjiwbRDDJ4uV
1OhqQbfqlCNE4zjbBcGNEKKDdq+ge/O2nD4U52elp+RCGo0V8QdK7rLmi4WMYUyGPccFfhvjoiaO
Nr1vIqwBzz3dfj8SnsH3IVhHiw986AavDMOI9jfSlaOL6jVaZZAsj6RuBLp4kN39+4l9Lzy6vPLr
acJpAEob8TnNVMaxeJS9R4ze3hAlGPFgVNHCO7zBmkXLxMi9zkw8ulZZ03zSChneLWkbXjEAaxT9
G7i8JpMDx3WIZmvIeVS+MN1fwvAxHguCsLE76m+LzaMIStkyFcPIlXYV0kxJ6SyOad/q+XIcEC5D
T1TqRwwSuqMI/pkv8dREbyQ2KmlKNTkZ2qlbh8XhDSkkvtaDerwnkJRrIT5bhDWtGUI9dnWE+uGo
cybzDG0HfFA0A/2ZHSaTClf38YS3ATu4asm/zRfzkiXJA5Os8j+HN+gIq2DdFRRr1ImrLc4tPwoR
wYj9B54V/S6CWdKTzBGrcj6lzwTo0kdyqcvkuK93tmbKOrMEzo7KbHGG1EtNaNkd31tkhWxCNn9X
2hXL2gJ7XaGkaUtrgzdqVwyYD8jViZzcehxE2mvkB0Tk3BKHavUe8b+i1tVHil8ugHxAUpsZF51Y
WGxtwwf9CDV+/sXzFu03AblNsLY6xfyLslw2jBuO+ZWpvj5mjKa9TzvvHQq4hc6xyx9CqgoCh9aA
sMHiU/yeVK2aqcT2nX/RJKWlkdHknmihMPYwpJIT/0es9vc681YiSlip+kllSl7R0vo4nN76J2rm
ZpjeVmaN6XxMKbeshDpDT4rioN9ywj6yM1wEvHCNvFr/hynvWwrpcLd/JShHTf5V5UGRF4+ABAK1
jH76OnfvDrPdy39igtIKh7peBGRToPOYDWGfWzUnBzWUjUeM69DIzxUlBWH/io+w+R3EuwWGLMw1
mKsxgglG8OSYAnWaDx89Gbifoc97ZSK5bO3wDlODphKVlyJYJMnsmTp2U+gtljMxlU2PlfdkhARr
WgctaxgTZuG1tzGId03HtGSJJnHxBUUeuHDlJoiDlMY3/1E5YzaC6wUfrfjZlfDNE4Hw7jaKeEbg
h0ApVWp/rBbiBX7ih9XYePwAL2gHS3iD2WgjXiE5vc2bjjRwLhtvR0xGl9RHEV4iubnqm40x29lR
qZPg2rpygGm9XKgzoV6dYdd2wjp2F9OEn0oC4KiCxKry4TvaU3+TK3mwEFmtlaUXxbYEfEL5OO0G
sYQWBW4Bj5QqmYlLk37PYislOVj3H7KzykFkhKzXWjgkwF0glYxM0eRPcgg9GajkfQKM4Tsnmb9B
zObspNQAF/8J0B8Zp4tMXJxTA/uWS4R1pvClQhDmzUnV/1t4zH2D+ZkBPHEqwKYI3XZs1JmmzZ7+
EZYitPNAoYAL357ZNDh1srLMzVHvQ5EEFbqe/Fm9HbqQl+PrbwEUAwtestZHWrh7chn/UhBhguL2
d2Kb+/aXC0Ss1jFQYpeRcdGhMtjgScEebqbPtIe1/CBYPitvvhbL+FkFUGoGs+IMlZImD6wX9sza
MxEScUhTbvkIrXbc+PHZtTr7vY2o++/H2XFbu5FNybmE+OjHPIsLha9y0QpgenYEWH0cxEpIOJEI
CCxKou33AppLzYJpfTBqvlpo3jK0Nev/KRWJVv+kXO1ZeyHAUsOTS2lA1tmYQfU7IluZXEf3uSEH
YQ9bAAh/vJ0fivq83xf2zgjpPGb11YmaQ0m+2yo4ZwMP3imdnQ5eR2rmXQBzaCD5XTexpEtllurS
6jmLYarXDvwJoaIFxJgdpnJNiUswze0ksVwobCuyNokqmjDFreLU53u8clS/tmJHXcE5gXEnveEK
3uLWiJUICc2dP2922uKm8NSJA6hls+JarHXo2nvQbimEq7fXaGip5goUOgrdBp7tkjR33lN1Q6Q0
PdH7+npt6aF4tLh+MgkAc7ltU382OLPBksiYDMc6haz9gS1adP2BgSHNXYE/E0pICG9r2zJY7/8v
rVS5JpMbx8eOnr1mFGE1yKpfeZKRnksbjm4YUgbYickHcpv+/fZPaMeFpmPZYLvHOiW4UVompJ0b
ttdbE4Ize4K0sffiqNg2MZu507gh779JYAcBipZQq++/ro91HUGDrvVycca+DdG1M00+rpU10nRd
tyXURobdp340/VmeCedZv6fPHoZJP4x4fdERokaK3ilpBQAx2tObHaBp73ABxiEpkYOKTXcSH5/L
x/mabEXFHud0OJkD8yGP5Y7DPli8F0V9NKlgRnpUycBRwpUBobiO1ejWcU5S5oDm4I2Tsm5x1kLk
Kn0rg4N/4skh6LjNrmGNDMVhPsqyr0lQQ0taJ241+i/hw5kd3NPPCC8Tr0/q4sip2Fo4Pyux1CVd
B/ghIsVKC9h3bIEY/U4QlrAaqzikOUYBv5jiChUeZgIDdRTgk15mMVn57fiJwxRNITAVdwgCOM1d
XwH6ozzTfOIEM4RKrQ72U7JEURCBbGXhUUn74q3Tj88GJ/cAXadNOfmNsbDDQxItYpX0YxuxCeQ4
qTXIIf7Xes7ZYQg7KbMeELOAfUf25Pi7UGCgEcX1ddPKTkMPZgGHypQZVth/Kn3wiIlJdjxkGt+A
gCfRgXD5gf166rTmHvfRh9yc1zPTVlnCvL2+/R/tW46UBn4aWox2QFh8YSoMA9WCgi4zQPaCvpHK
w1y3xl40uQyw5ME18eHhKy7FFclO/lLHB8Ro8GJeBAacl2GgHGb3/p1wkbkx00iYI88vHumX+nA/
z3PvD/VQZB8kevJexrLNC1CtEINNs74SkvSXjaHXmZ1b4Sz5BgFCOlwk5WD75ei9sSvLUzHbi9eo
PTEo6NKMxQT8LdwX+2wVYEHP8h9Gf+Kb7yfz+6Hg6Jn8ubi7m0/Wfj2ptzC1tIQz61jSRSFe3E/N
FRX8XJS5ykc4vLyzRMWHLvGn3x0Ah2Nmv6W+ICW7aYBprBWbZWrUFTiHFXkJ87lU/9V21yAO7JH3
Bti+sa70lVQIRQOhvdsUmi8oR+21K+3iormaeXwohgJXoTj90JZXUqhZQxc4+aaqjUSPJNPys2iX
+6/D9rhh3+2HD4FlsmFeN2MbIrKGbrxsWrdlS1X3GYY1MbyFd0R7Z8ZTXeqohKLtmtQOXbwybr3K
sAOqZ4hz+IvlHI91KGspxFjgKpFb49wlwAQzmKxaKWcXFxshUpHCqBqbYQsYwSfXgFNHjCUpUOYL
/jYfo7ViJ7QrLnx6dFpA2AsMzY/JiGYdsZPcs78withgD8onixa4u/gNqDZBMkOx+bnZ8q2MW2HH
Nhr1dRiOpawljMAdt66rQc09CnRrLuqb4rbbE5LrsBZQpDlmOtyVrQ/BQ4lnW5L43Hm79wlDxu1r
x44wBgAr2bchJeky3Hk0gx2K/vBvLa1FV3mloPa/6iq/eKXA/OfeRtsSI6LzpDMbUGHiSq2y9ZAR
0Cx4wiIpKSzFqcsmrOGBRpfpbyFhoOnqcV883ZYqqQ5gxEJBBsRZb/2kob8AykP8tg00RbBHu1WD
loQDlLJ8g41XrYV85XrXDabJxtiNidPReE0hf9S/qdzyswdclyVq48bXq2mNjCWEw+xNirzVvjKt
06wTOgIyuPu6DHBN3m2OsQc9p26vdXqO/Ks/XOxgBi/cyJ4VWYfhGTxqAZA71Nsm41v5r9FhhA54
y5iGGSFjMK0FB329dsq918EMDnywARIaFjCKzkFVyT21AYAFjI1c41xiAYi1WnVaxeJ6rPn7MkhB
ynr3lOljpUfKcFd4JXvIrkp5H502eSWDsZCYT3O4liuaEBR5wtClTkJ7sNgBvNOhAyFImG5T/nRp
zkrBM6TL5eOoeP6OCBak+Qz8+De8SyYtpjpI8SZAVqPl1YGy+d+ynzEoNC9daoRpP/cGKDseLVdW
wyGYj2BsNVj5ZE5/bYRdaXjezj97VyuqcyUwfIjuG+kHetN0lG9jq2nQpSfzzjmee6O/753OMVtg
aG0a/gNw51XEjDbz03n0pqtQK3zt9vn6ArdX9OdtnKF53o8vE6YXre63p6OEQVNqYKx7I+Mj5s/8
Cs8rnFwdusDF8DnczpzHeup/9jlfYgBBICThuPKMJdVfY/lxNNMf3vo7peycJrmmDZsXjBPf028O
Owti3uHG2RVeWlfbvsv9udbLw3BMmOBNQk0atSNvE/xmEtmFfL90LIpUim87M53BB6vDM6D4qx+B
mBYFZVeilSlhXr0/ELSza1BRiKBgRTrCHrKa1RCfBoRzKdLc1fLYhYs6wfq7th4TWjI43a3/3CSK
35BqGVEDXIz7JYXQTkq9xKvT+IVh6o9lJmZDL1aHhVHMFQ/Deq2vnnULk7n6KUtMLKNSzef8tEPM
c5uxV2UMQ4bKccqGYyo1DmmW9pz2OURJgEfdSMUkpOZ901xC+gpvOsPIjD5JFx5y/0XEy8od0z8g
N7u0FTWYE+YjVNN68kvZg1NbY3yud8TD6QMg3zwhUtrIXH/fdm/VKqWtSbt+rbFVqbfmfyWfL9I7
gOxMZDiheE3XsmP4LvG1+PKkzoA+gxYmei8vEQ3Hyj72/SEJOS9/qCDuWeTvhp1b3lCjZtoSYRiX
XwRreL9OguZQVUDHBIEfsMxLxufyZ7Flrhv7TtQHTWv0qYfx2TKHqiMRfH3sirpQTz2rpIDua/iF
SRoWK/Ec/+LkCeHUtGojPpTtmWfZW0MoYh5Z1vxxoIcdM6RxhgehH/8Z8N98YZJkJGGu03tjfkf+
cDrK5UbBm9zwelmROHOYdcTvS2r5jYQjH/vdYU1sM4vyy/OTQovaNiUSTSuHJGn5Pq/qYyhP9Mum
kwwU9YQj7N8wlRfrQq9SklKBHaEaqjcLoUypglsEaest4KQFYgNceeP6RyHhlN8EQG+XeiPW8VSD
5zEtxbDFllYZlN2vX1uE/qyByHrwlFtekkm0OaWkv88BreG4AN/rYHul7FB9oQQPwPRK+PeV9ewA
lW52nXoyD1F35xvsFesP6bK4MUoZTFqyklM30ftLve4htGVdu/F1upSMsy+gSfa7yQT+ee65DpR9
dt3VKlECpxgqPh+GxtyuelxFbhbwF5tdXhmX8/u9dmLW2rZKDgWkTZYa3dMVBB3WdMXADBjpbFB1
g1Oxdibxjwzkf8FfhPEI7SzNwOHfZqGqjb/iMWUZTCpy/KX7+fmreI5ugms1tYQHrHUovS3vBeN0
08pU0BxB6r1YLeLT2A36aTXN2Bsr39VEkSG5xxHkxCzV2EOgQCXt290NqddLmAKBRuIGpIKaluKm
dtB3H5SAGXIC8JkGdq3dJ4XJmteMQCNlF9Zr9p8DZp1zLXgC5ZXMbRb9Kp7wgqZnCZ7SIh4xlJQp
kGtZmnkH8zY+KJ8+j4PEKQfHUdxH94jwPl5FAXR8QEGQ4Jeh/FclFXMSqKr7WOa/+hTCrFp1bl9H
63Ek56Y8ihyBXjOIvzTdTlmYQEqWWwg5IeI9GasKyR0Qh7gXA57Gmp5aJ3YL/OCU6dJSrXX2K0iX
ArDPGNYWmMyTYlDlgiHK3wnLPNw0x5Ixca/moxAWKAI7JLDnV078elLBV+jfzpmp4XjHO45KMXjw
GVav59g6AF/vZxy0NPlmV+YNxS9Fcv56I7OOwuTt8IzFQ+70UjoNkmdTK2bbKB6ol4s/MfcQ4sQ6
Fe3JH6TDID8aEGglqoqurRi/SBsSuBNHm90NDvmhBkgIKGpfheRXI1rHPG546pSuyoSB3ioLGNwZ
V8NOk6TJGZTf3Zji+DUFx+yYXAHDezQwBD9NlnA/wr1EShG0nWWvqO8ia4Q1qt3jkHjCTgpew0iC
NMpMtPeVkqx8JN2lVe5qJstqN2ba/NdC3lb2EIDty+BTQdrgzm51a3jVjNdFrNl85PyactuSmBJa
tmMRjeoBYJ9rBpIkqRvRnz9j9ZxDHiiQjBftK0y8yfz/78kez/c4G+H7KbMcY6CVPzJVy8SYB5xl
aTehq+PzT4ZaCYq58wQAX8uMeKrkbp4+SNG9Q8AdIVIycU3m53ikn/7icqFSrmFGA2eSUc3/HsQj
tM28Bo11gHfOUZ135uv4IJuO2QryoC85a/1PN37tXl2zSY7crRg5O3eXZ7kUl/i5lgdGBa9dcvm/
tuDgx2Jh/z0kMMK48PmW8hPbcgn+6uvVy1aWnv2h98fhcHkoJnkd1X0uGWryYrrfRxI8rw05ScoI
x3PVId6ckskv+03gmPSpTHHAx0FwysNfn7zbXYBaTlfvmNvWmf3hzqjII52Wz2POzEW3NjANANwe
pjouHsy+JhGcbhfZqdbDIUi6eFzjJOvzrBJyROMMjvbPnnzrxkcKn8bNKTttrdcuUxpWBDJv0eaj
T00Pmsa8L6eU8AVWOKcrUJzWdglNmPDQF6AHgFQOKrKreZQM+eLuXTvznNi7ik4HOg2Ls/LS/Cgy
sr2ZdpsOaZ7/gMfRVwDt0niEzjHzVnBOqj85O/2KPpneKfmXpLqkyYGrPOssng+IkJZncJwGyNqt
tprcm99fWmpcjfHAzkP2KuHmqZ3z0eB9gkhEltsMK1AQ78EC8uwvBpGQOz9BkMrRVFcvmYhO+0ih
7onmQUVqWNU/+Flbt0ien+i8tylevGkDjPuGTosW/inf2HEzgAKDDXQ2rYDrPcE8k/ZsqH8VMmz1
4v8mYLgWIGurq+6VpOnjFA7m/GLuCfEltUtXJag9xZWdasP1CK9vMpsBbzXOuIM/B2lFJYLcKa1E
DPTVPjFs4W8oOSTdcREMrOuwIYOIC6fMBIV2rv/CZfZvY5j0+Yceuj7+MVRuL30RoTFOY7km0hvn
KHCyvXQ7yIXDdJlfx2FreGz0aWMfJaXM1dvwNULUuS1yMq/755/kekwLzvZU9Oewe8jKR14ZMEfh
9B6J2HC1YcHJaLgexXJmbOyV68dkqX0aaIzKRRaUIB/Q1+pxsFjvoV14+IhrWC6siAZiId5kwXbf
bAdnjsauTo6r2mzW4ku+iKMSldUT9y9m9hsitjw/hyrQOcRoMGI27gJNmC1bVjVETCgI/o+K2o9G
DM9b5bcntRyvEWDSa4IDV+GPypVdN5i3mKwEHZXZKWcfzJO+drIiO+m5gm29/q+hSGycgeZP+ZER
4ErfB9QtCThUyWW1x1XrS8/hWoi7RqPtTdGsyrP04dgawofh9lsXSTvN0MQZEaog9JjPeStEMhvq
itDLCNEQPyB4+sjNoTFoYgFKz5pSU9/87v0cJSdlHPo8wn7bfFKrIysi3eGK8O47kFnwaR6Oqs+b
IYmy45xuY/v7oEyTaFbG1GC7GZrcR0O776lj4Ubp/oItAi7MMRCoChVr+rRlmaSxf6np3yYxx/jP
NdohHrOtqbAIUURB86gzevJlz/3Vnr7dUnslXKMjZxwWdf56ONJt7F/HhORWFeoihLXHHzoAdyHq
4ndsg7Um13bINczZ9oAadHqRXbb4dlzv3Sq6yxBDQDRk9/Q7dM1F/B9LVBGcbUcKBqDFeBi35urN
vmvzOt+IahLsAliecwLF4DhCznMar2QBKARYCscB2crSA8xufpVmhFlZkgEPvmOmsqHTGzjVaMCk
i3nhwKGyyqGto4ka6rSnt30hmpo8NFWrzym5MeH81kOukjxqCNWEhSthmpYUEjcFSLl1ovli+oC7
7Bncu0ZVqqQk+EqgrxJKOi7r/8I4AcKcBs1T5dL97/I7ahO7AU5H+uftcTZ5yI4bltliDJWXeHbx
XseRjoHs2AWroscmvytTSjQBr6qkcbVtIlTofU0eVN+XQIsOca22g7vQxXiVKj396SM+L+ueSjcP
Xuci+NR8RqQLLTDS/x2Mj4i2+Mvz6K1gIdLV/G/pNYgLR0qRTSrBYIiAAe88unVW+YgWhCV1e5SQ
U1auGzJa7Z9Si7sSG7E0ievWI7y4DkT6U6t8GHERjUx0emt3K4E8EK1PGCq0Mc3A+EMmZq0fCQdF
tkeTmjSn4X5FWTrB1yqbyn7VrBcMqGdcq+RwPzSxT8vvw08Aa4fCb8HKCahgjErrKlbv9bq2g+p4
B0jXwQ6GCu70eB4rHGtB2yNPCTzMXs5fRFTrmtumOSal9VQtMGlX1YGZqbn+F26ZjZ+syJWN5cPq
PtHSfSgGywIkXKzam1XhHR0N8Dp3kUSJ9QGLuXjrwMgWAgUNEkjJsc8HTfiJUn/yxHcOpNhnmLty
4dzVNE/QUOZuOrYSuE0zE3Oe/EnyiFEk3sZZwD8g7TsPiBm16wSpFKbaXK8qc/HpvR3uWL5N8/zT
GHuM7mCWf5cRpb8HlxHI/HiHMprXuee49bd/Ot04R9iiMsPykW5V3lGy1UPsEmEmz6Xsziu8y7fM
kvukWarzMv2X0hTXhboV5ELw08LVTE9C1PoVk5yseyQ4oQOc4gT4VkK09QyBdCVgwqCLSFwfYXz/
3cscvOpSlFVc9kkRCX/Toc2Wv3sxAaLlPNgDQhIuaUvh+MfxBtOTmuJkpdRNPYmPVAWYnRVvjbyw
K11zsMJm9UFUNevOiQ9l4Ps1ll8OSIODsbCqmclMVKiWMhCmfSl2+zL3l5lbT8dJxAdrY4blyXj4
SemaM1LY+IBLjo0nDnxG8T+bX4BFi5LDT42wa6p7OGiIDAeKxLWHnM7Gi6o1dqAYDzbk6WVfIRgH
nyvDfJJL65/Br7WDy65UtAhlxZ6dQogQXwa+tQkZFs+YbylHL2TbmxAD3k8fHeTBphPFOxAmLWsM
plrxz2G30vc4E/W74xwZTId1HCMbcepGYo9Vlpn3MbSMfVJLdx+AnnQizfoI6ewnOm4dcJ9sPdz6
JbNhkxGm/bntCgigCARDkndFgtbjFPscpK/MAEAdodCkuoZtbrv9LriITFWjqJza/iaVr6zt0MJR
y3WmMfy1OZHRAEu0hLZaTGxQaywGkdxWa+7RSbQjT+Z9esU0iYPFM4+0+YyifZyI0No+8XTNGULv
to7+4Ja3CAweghmnH96gWevb0Exksh/KeuPh5J3icb9T2vVAluXhnj4C0uAw2uzQr5bxDr+EQgtQ
ErTcUMo35aLkt9HlLoufj98envKs96MX6DXuidZ/bQD0vGIIzx9lxaLf7hJ2Rh+VzxYnBt8Bngrr
M2P8wlFr9isJrj8uDZqVbWsyvZMDrGWKwEgTgnw0myxS6mLto6Qnsk/W1Wqi+La6wd+No+7DTuz5
Jbs93cWCV10PpZiJT92oTisc8fUz+WyPS/hmdZ8x4LUF6T4OpDfd0yud4dVfNT+EAc4LPx3rgp0X
pJHTvpUVT4FzlZUXATOPenYg2DamBh/YBytdVgc4thHw0pBNy8bLVZE/asNMuHmdk+PoW/zAwsdZ
qfNhAfopClsYjjKkojCEjlEyjtLL8CMcCOGSscWqgIYRtKNl5sRjYQw8u1dL58UGnMNRICxqCwqu
uCJD1IGJpAYtEgIducUbuIALcfVI+REAK6nOd2bz545U30YVip4KMf1PGx7vM9ansrFoTJnZlpEg
na5VWYn1zMkYtvMb62w938NARfsV9ZywROgGXCA1MJSLVa1n0sO6dyhv8wCOln8X+BliQXjRVnAd
C/nboCrmf6XfyN+iUlYeTEAwiAZ+la3JpMD3mZJ5+zvQrgMtRzdFJpWAR1UNgsokYl2HLB9j4ENZ
c052WGdohhSFb5Bao/4XVK4X8u7AVqVxLe7FPxNX0ASBRMZTiSHF2pEV9V0f47tA9LxGUerTITuC
uzTL1LouMPT1xGcmNYxaTgkD9HDe8pQ93YGdZh/yIycJiDv3VHT5uSff2vqWDGoQgZl0ztI+4LrB
NwjNwXax1k8pm+/6LcytvWF5888rqYSalOl2bfKn2vC+baScLDUPeu31CD8l3XjBgChm/fnSzThk
iRFS81zCrPcQ7obdxAmYsjBo1EPpC5gGZUhOvdQaJXOL+oT64VnsYPmnqA14+wltfbdG0V/vgdiB
n4fZw8ZnLzmAtJFnnJE0rTZ5jAZ2qLXNfU/R5J4sZySpmAJpaPzeETFva18i1o3aUBQCKmyL38Ap
Kxymw2AH29Sw+mgpKSCzb2tNoQuFUtUX+sv9uxcmKfRDdc2uvsXmHj+YVP450pHH7ImgdkyzZ9WG
0GJtx1cImcKlOCBLl8JpmbKIRtcamDxWHSeLcfo3epORrfcfShcJTBbe5gKRNCr1zPIAJIhc60Qj
Q9zI/FxSxHagSh2hcG95HWI8ubd5kuAqccCMRDw33Cs0x0cMd8xeKgBPuclOD/oFj10MhGuJUdUL
RdCZBYpBjXqMzkP4E7AsjW5OS67pKjN+EViwOGk5eRAKAgt5Ep9n8RNXfrZlkbiC7E6j6rAwpiqz
ScBOnFdgXU2o2++X6E+heKVobZd+R7UNTI6fLx/X77NPiY4CmLtSmGB/TE7wRaaltDf3xfbqWDow
hq1ggUPY93avv/J9JLrvBgYPiv1QgeUetrI3dEOPj295vaWnwOvSdqjGFP5sOh55Wk8uLLeAPm/j
+Q3qGoIvt+kO5XA+NmKjVPHOaw3xZdbdNKulma2zItPppElXuKqJxzdCDK8QL4jjO7sdmD9OLUaZ
D8AjMjmBJCDKHkGZMkHBK722zTjRGaaYAfwPTnbcgxcyihcGw+CLmL38FupJY7U3OLE4lmhheQUO
aYDVXnWuNPdMpAEJkKa2GzKrH0zI+USjuPvEYlUEoX6w/jmWAwO3TS+hr94a9N3ZiXebtRsS3OHa
FqI4J5nVKeRrBydfXtgjePeYwTIc51t0rJhaxBPrn8HnXuRDjqF6nVMeM/GFzXymxBDbaHSQxhqu
PEmWWSt+7sPKmUZEcLSgCiclCq5GR5lEOmrXUcSpSOOpY826O+kDLkbbHFcyxIgcr0meXfc6eXaF
uLwEXl9c0730axNt5abGDtoB+52++mBUV1om0J+bDzMF/d1L/iJ0EJehsDQhzQcLUDHTI3W6gR/F
CM6nownOQx9ZoCCXUp7g28/2KaOSI0rq2rqvRrvUzLZzRoSwuUdVqU2AxI96LfktnueqeKxN/hOe
dY5fXg7upfboLYvB8lYmPK9SeTfm7cZ5/mRyOUZNhUOe/OMLDS59X5DJQrklt4UvIWrPlz266UIC
N5DFek9mWNDRQ+Pkd1E0+1PKg7o29i6gWxjwHn6L9RpsrVDuTDmp+euKyiOh1RDmv9oWpdh/FaE/
degOI6g2VE4MQebWcfR9vmSLJanpQKv5Zivbq0yk8+ZefzPrjlvqiJiwuls4cK6p5ALp7iUMrOtQ
qWtt8rj+9j4O0lI2YNtGjSFMJrGnUww0FWqlnNBQHO7oxB7gsgc+0rc8HJNuN4fd2xd60Gu44xHI
J8ygCae+UHYvTN0HiTK03SEfAx9VWLH1ZZAJ9TiSdKjYUrbIWgfDamv3GFWo9VlJkZX+CHNjs9ir
sG58gqui6w3B+IxccWdH0Q+00X2/9JYdYsPfB5KY+OVIislmf32Rq0tMNV9UrjUJtYg1Fpq55F2B
PCD0O1Bfr8ZfJEN4eCQMQ+jTVM6jOi+PTvCQ+tWKBah/H3HE45fDEHVU4MAc1E5ICYRz41FCw2y7
BBEl8aGhUA2PB0hED2fEJPk7lEkCRYOv5h682R2W+gPaV+YYVUuzBCGXlA2eIIgR6baSNkRQj0TK
SHS8JYizUBN887BUPEaE4FOTfkng6l2QbsR5gc7fFkF6VjmNRPovwj2XofNpIrdJsxTOlkyaH0l3
tJb51HxgB2WUgPujIx0CwGjcUUG3QsXgzu5tgPpFuTYajpGEZDJiqMsqoTb+D8Ih1kBdH1L2Zm5q
xtANLtT++dN57ZXsqOQvxgmVJqwrxbvz49nO74jHLphNBB9D1FDJ+MG2J7ztLMr7RAUij6NCy8vA
jog9KHogp7DzXzwmKOyOc5NXUNFPlHPhSIk003WlWv6xcBxZ04Io03I6PQB4TWpX92/H6dp1EK/1
dJQ0zfGYbfqOmde1TmBhd1pmX0DWnUjqrG+JHNoyifSlyelFg3hFeRVTQrjIM9rPlWGPB6M55kkm
XMBZYu3gd8RVea3SPQTFuwBA06MF49qp9bYUOjr2lwoS5Vgva9fZK2VKjGPwqOrZiQjqKraadfiB
lhlpgWKPsaC7S1tuJA0vWmtTYsri0/pRJ9n6h45NSTPUyAYP/FLhsd613udW4oz+T+dVhUoTY2bk
IN1bbUcTA+BSKO3GpPcD5K36VjLfnMdUKfoRPNbyQ8BvJcrSO9Z5ntlw1cbA5S9mn9J2pP2wHSYF
TAzY6zQDPM5zQeKrIjouGOaekCvCIxFg1WQUaz1UdyDgQB2iUwkk/OFzCmTsAzebQ5/AZbuH6srH
dIhr/PUe41Kar0qnP9VWLPh547XDdjGCuiIMgIi70FnKw+PUIDOrPKQNNdiM6wGz3GcMegQoKkFb
oVWjQC8JLGocCpf6RdbCbrKxchubVdGPU/YexYW8ZKjc5Vqj0Bgqh1K41AwVv5rW3SphcrpLDzU6
GXQuMSf5+GiVaemvZSMb04aN16ZyIRSQ316tkG4h1yn4e1so1f3DPpJJjJpnshoAoSxFMq8bxJa4
2tYzToAgWs7zST2gwzuUUC+N+dFZcsyDoxlKrT1745xzPAfHXaMv1BK+6nhn2RNY2gvi99sorQs3
yHDr4cq0WGM7IccJB3SjUT2bo/AvORA8X2lc9t5xOrhawIPcFQLVrYMuNnammTc9XJpLn4twLLCv
vasqmwgQeQKIQkxILiALu/YR3+bHBZZgxWh6atUEN1WQkUGypL95tghN2//vNOaJ+049BJdcvuvW
/BTGyfy4Y0/AcLZqEamzpDNxva0KLOO+CnJ3GHevs2RlfDjLm9IABKSZz1sARJ1tyCDylMQI0ucY
hTWssFmEbh0/25jMGUIhTS55Gx1Jx3hJqCbp/sgD2PL81O2EcTt2HHkcWCgDnUZmW6/yW4Yz+gS8
FiAH2EabTi1E3E5cn00QB/XT13Rs7DXRMhyfQU+gzy9v8CpUSpsuAGuNa+tyAGEMJ/Z9BvbKSfg8
4EVbkWrUNkwwOpBXZp2tEAI6dxNi8m2dd0qEhcnZpLfDqMahV4vgwGyUBPPiYYKD9cDZOAbxsaLI
Br3MgWCfbq9ILQpKHIWjH16vae/okuawf1bvnpbdyeYecF+HD7ssdkVLdB87iF4PET880MTtiU1l
AUhmtydfwLsF/NzVW4arxjNbETckkcYjesaXw/Nj2aVkZvG/NzAbMYBVLojwZKFH2nAxNg0stvmW
d/lBD+G9VV1AW+gc3tXq8JBMmc+z0pab7jUFw+PLam3srPPyE/sC2rymsZ99Kfz88oOvTC/UqJ20
yYyvdUHf6+6VxOIR5LqpQKFzuLE/rnSQuivGz9KKydks/16BL+bGIcmQ1/QllkulogfdtV6464q4
Xx+NXgD92VTotgb3OYl5Dk83XZ51+QI9uD397VDZTjefWdGqaaLLpwNjWc/BvEBFQGelwnocObnJ
Z6snEcEURUobsZEzo2FHqRs3lfCa8XyExTvY5Mvfi9OTrGQIIB7wSvPrC5vMt3U9pIgZPCEfWw0P
EFheR3FyC2SDo7stnzKkYFa0tO97IPOJz0EPVO/SJF5Jk8nykfAJSvdp9DeoOzy3BOqrIpH1jewj
H8lugQgn0HzOdkfRkK5UbozDAojUiOCcmYWFji+0dY6W+U0Ht+vfLa9EtbZ/gdGCkE5+gjIQGZfG
beSpdnA/CsQIICtZuqlvoxuXv28UMmU0YLuldyUn4wnJpUOM6AkoftN2bd1TSpT9eF1f02VTvEqM
SZauVMbVWb3833mD6KeqFwE1HY9JemDzR5W2EqZx3PiC6AhueCk+HBX4UfeG/mBLoEmTHOtBUCrT
Vn4GF9TRtlfELuZeq8IjY6bzETbLYWvSe6+rVDyiMYlL0ZSe+5u1PFMrcUJw0yPmoMJLopcDDkWu
b5poK+2pahW3ebMr9/iJynwo7vlCABjxsEtlMlbjeP3/6mjZe7rjbctnloOu0ZL6QemyYeH8enI1
j7ffLpWIv9YDIJDW08mD1HFz1R3au+XmN5rbOWQKvb8Lt/8/vCcjul0Kx4YA7o8+1hN1HSVSvjjD
Ka5h14ACw8avemP2/1Iwfe82aKwMtVKhb1RkjgDgExoGDD4gj/6OkIrzJEra143aJ49DRocU7GMx
p3mB2Fd/H77ncOfL8xmwJnlkArGaUj2L4e+foGwlIhkxXfLJjtE3YogJLZ8esD4smLaVwSvDmSOz
tsMZOpKAuT69XyEQ6En8HEo6tyJU+Iptj4wKG+0D4Uk6TOEj8eEEuH+2rccLVUAMsgW58wttIQke
rtivH/CZzRCweRseBqHqaq8P6dOgjJ0uBe86gCWu1e1nveceSbJreal7BbgQxMgS+GuEjnI/cGeA
CpxRO60iaTuIBpCql1nCH6WxZWLd+GNl8YpLiBDxjumJ3sYbt73RpvE/QduO+CSs+4nOdghBdZ2o
a4YoSf8X5e9oiyviPVMmemZNaQ56JsdfBFnNp2em0mz/RoLErcPzhGdpLmYMXsYpT3TM77EZacSO
b7QkxtzaCDbEvWyVi3m1JI6I48Z4g0HIvjwTkf2sLQ/QpDnRD9pz9Lq8Beoo4HHTlDGp4/iAVurM
jimRThuMPIYnE3uEOXZSvlV8DDKYHelLqMjddccxnTrAjbTJwhIj4JYoulTlzKvjCkVPxDyatV7x
4Gf9efuxq6bWfrUg2bfMfkicNdvgmXhWjbjAnkppRMYFPvDc3bNtglihdUu1ARmiqv0IX8C56n1p
7VQImh/KC4kGscsxehZ7ipKiNIHxIfAkw9oGK/4XUSGmWea7o77DTG11t4ArsrJ76vj9LOxElp4s
MDZ/LWmjk6U5mLTf/v2zLA2ILM9Sib5HDHkiWn+WBNcGfDK1IqegazmhcU0n8ip85TXnptBYYIit
CHh3x9ezkWx7PUokLEU4msfWdKRpR199lBBufHwPrQrNvbMRaZDfMChlR+BqjRfj1JjRCo2ABJaC
slQeAUlxibXeZ9idX8p6a24wTxmIgYYkf6UUTKZB422rk2XlAqMmxkv5HlWXQEbWrU0Huw2qaAVg
3r0g0q3JFTIlbB36CzsR285V0cleSNpAOLhK5XjcIP/ftyh7zr3te3+L0thSm46lOUSd9MnTu5JU
DQREGL5dlHY38vfTzcQHCwcKoikbCLE/O1hCk4btJn432NcHiTsaYo+wpzF9NuYdTLS4GK+49vJ0
DdSstoNwmhUHD7l9xJ8gPELvRik5cv4p33WYdGC5APWrl4Ki5e0QW4rXFnt/hq3Qu9C9qzw5/e4B
2VkkvKJLTL6a/IKyVifdr/1KX5HWZg4ZG2/Hy2ShArL3i7pu+9ONdAW+6fU2jpLxdx4EaycruKX4
TZBg6/LPaWFgq4hwuefjr6rmcF1JtrzsNHPdXfUT0c44HSsuY2GlLRmYPclPNzxZ0vpwGXCA6k0b
RmFHRuj5xOIRHsApm4LTUh+ysgfEuEnSc1kgbfGYr1qjrqaN2eYaLyi0PCaGutY0fgNTHDcU3czP
AkkY9V569G2EH4MMGT4cK8WzbrB/Pke8NBt/k1m76+QeWW2pKU33BfRnREumKZ4ayXt6uq4xyS8F
9NsrAmK5Hj1d908bQlvqthygkYdh0il4Pa5oEjed4rVLUXoCQkcGcYoVDXjOJKGjMsOfOLBiRhf1
NSEXjZv1D8itOrIFBUdUzl2d3g5CZ+OSMd2yIdr1ZRfupfpyGcAtmtotlDUFWFqHZnRfzAQh3ErQ
I1UPRJQjerVqsRZIck/OOI90orkII53xkSLL7Hy1kaNFGFkEQLXaqTbtVWu1TKRAUm64fmfPybHU
aI5+LsZWbF7mj5XpEJOqsL6JIYPBmgT11zyRR3nKkOFUjd6R53h7qcWpgGVUZrIfjeW2jHaTNrdV
JSMri8aLVUR/Xaoe1aLLXo3j7x1w+FFBCAEUrqN5FBBJRzznaYd3q5J6LyvUju9leHvpHE5VSK/c
kxMuQV5iL5xIAyUNZ55rqe2wPE55I7usisjQrDzphJjBtoz14vzt9S1KfOd+9lDExwN7StM0pezm
HxqbppGYyc9ohzIbrP4bAjxPKXTm+ZxaX3fjuPIuLYFeVCKZohev9JtqFBL5cEaLlI6i20PsSsLJ
MMQZf3AxmSdZIy34CLv6zu6shuUHcSkxnEaT+2CRF5xG9NqHnZEnrnpfKvfK0jd1MYPGt1yd9uL1
c/ehGcsMUQ4oDLVvG2sKfEvuq69RlHMnNw8zj2AZY33zFP57Flzztw1lI2/Zgbt3PQxR43pr7aFT
GeL6a81dyP9RVaEdL2mWonNypyfQbNJx/gc5dCHxVShzj4yT5S59hr5N/iLUO80BZI+RNIJediNQ
muiyHuap5GBAz2CvdEHU6aHpvgeab+Nwz+1DPUHDh2JptOfGZsWh8drmcAI5h4jfyhYcrxTsnE5Y
4Z9Zi68FP0rIc37/qJWU/KE+cs+O5p1Dp/MT4r/NXcTW7qNpJ3HtQGkyyZwK0XLOazjivgt0A31o
cmhCkU1tkNUEkp9P8y1GAzuyQMk5a1Mspn72o1SbMjsaY8bFYFZ+W/aH0uO3i+EU8xIlkTwkTaIp
pplCoobixrt2Z8QHs9Gkg54sDpudWyd3b5wasUxvS8S8Ll33RG/oITZoISYv2ahiIkPD4HwLDTWJ
3WdYExqhoSCgG6Kx8/lbT3RuGw+J/nO+Y08NFosZXQsTOAbtICLePKrlpZUEe3e7fpDctx3O064Y
fT/FjruVzXMKkPqohYatIpZEUhcCnXuuUHh0J/qPkJe36m1uDCE10l9y6FMpS7AorrMKOIln9gQm
DBjJCfLf3sdL/laEAP/F16/UX49LYw/CJJlqA2odv1U5H87OMkj4QfcBi71DRYfDFQNPR0QkGq+w
Xq3QFZ9YjCFTPWm08UHTNzbYJVIhXYMEZcPe6Q26JedSA02jnjAkvNqfUyEKSuMUuuVwxG5W+B+g
NG+L4rBbmp5mYwyNFywqRrdMY59qupT3IcMqThsfvRut95sElxj9zUBrbxBhcLq87Lqa5qHIJ5u5
V0lak8Cnpt0qbGhRrJ+K37iRr1DpEyyBm2VtkVVRFZYjMZAxGYKfAh+RIzQmb4cGx36332BVAHEm
OqzqE5fVDZjD5TvzsMOqAl60o6OmoBj7j0uzxB5gDq2rlEGMM5D/d7Z4ku4hzQhodkJDIMxX5vf6
ClH5G7yshbyDci5eDjCJ8alT6qMeUcycsHMWzlkTfARWtXv9Mn8Z+4wLTZ2RLVlsUtzg/h4YidRJ
vdx3Q451RdXz3Wn7Jilx91/F/IfQflTjIJsCBeOHLwupqBcW5bkN8fglM3EWmqv/PRZTgneQxjIE
KXQ/B5zBqdYMDn4jrX1Gp4yUJaAxL9oP8ItqZkTBn9NTSc9BQaIcPydUfG29Iz9ermmmgZKT4LTy
Wae1NfEB2r2XlXQYW2n4U4aMVFIJaz2zMnR9Wd1/0oWEM8Igr7uVxO85pH7nY9LD54TQCqT/vdFW
nU8Iob/3zWP6GpNm5dxiziwYEZmDVpYk+fXVn8C5S2E2Y6nmXQg938GjtEJchH5gsSfol9Qsr0/T
HTjYA+l/+baXRzkbxtQ08RAbgrxzJ4pzNKLVirkfH3u2zqyp8wrg/plcd9KXpbFUD/IhVUrOTqu7
kmeqP96Xbv7iz5iKkiLseDf0e5CzSBpXoeUUYk64eRvK6NBlAy6vv4VP11DzL3w60iBm3OZCSizq
thoPGigdqucY/tjIgXOGpfh2PoE0VQ1vVgNFkpa1NI307XzaXxkElFnOsx+kl+NdJOS1Qjl+U7YW
cVUFoE2LB8QD2+MzRUO5icaSspS7RM0NRh+fAcs7vGLt0Sd5ClNbAtXDjKD8NNqvCvl8XPG/gpb6
PW1yWf9GJAEYV60/e1niIe3DCarx5QdPRGlJY0TDWfAmksQw6zBD1VZL/5fckG6UuNab1wsJMRjP
YTRni0Y/Zk1TmemNK28NhYGPq+OuDsaTr/SOrFe+HNTLYaRDQvRA3lqWR/+lw29VPQ/E55hSKp8S
TtsHANS+vNr4LlotWwenQ3xbZ1B4OC2ivpxecVMfFi8D5LlSYE1UYsUZI27B62D20UT4jFuy29hd
efYkI4H4aCYPrY/zc1MPpnFTXGhpL71xGgOd/J2sb6tSZPopk+citP2hE1pQE6GZi5o1fcBVvu9o
edxHNUfh0UG49/5m7ALFm/o91cRYGgZBXNBBhPTlNYoxQQ2jamnx80ZA3sRA4E8DhX2YCRrfBQu2
bP0UA/lJjAan2s4E9qs1e4NMvfSLyFgGVYa3y//8YVheLuxGABf6IiC85B+J2NJj0m2EdiF303WL
fG2BaeJVYrT5s8eA9s+VHS7saUI4f9MKz15X63pRFysFRbIu5sD/GmSuyWhHgF1uYkFMVdcM54rL
x9lFYQH/YtAlswcL6DVvmUKTlhNRF8g0U1wUhfEIvN8Rhp5bxJL3nCX7mRlIQNhuja5HSjZCJmjg
NA20/LAfZkvOkywBMQKzGzk3pWz8ae2A0WVbb1ibd0UzWHSUGJMlEJQ+mCHXQal/lHwc2fG97ser
tXnxw8zzh6BWBYEasX064sZ1JzewoQMndPrLBxqhtmfPqliSGMP/TZnQ2B1aVurElTfF/mCreWzH
VTW/ww+nRIHHEKWYNYIm3A/cXwzE7Gou7LzY2v+qXzjUf+IpbYzeLh12p5ZLQSn4P+zxTXLfsZVn
DtrtHXhTfaDTGOnuaNkBXZxHpMO1Q72cNnzO8ClkDShZ4RP7K4ZKfa/hsYz0l0w+6XgHHc+YZ36K
QlxLjkZugriv9jD2NbbWmgMGytpyFAfugWouu22A1iE0O+3F0hNJ8brufr6X+F249xZsfCoBi65u
SyQ+v6rhIqKmzFBO03mmfnsRQZEWRQrTtu28/3+tzLKB+Dp5Gv44q1jHEmo3ls6u1xtrtkjCGzuW
1p212cL6aUkAlfiUxORJ4Gy/8eoQbC3+aBcIWwhm0hPWE2hQJoJoqmjaQiwTWlevG201Cm3sROZK
y4DkqpadjVxJr6Ko3dxR0GVD9opMs7bGABesrSmsLTEZnTK06L/jPipEYVSuJ9zTXckknfIUA3z6
u0aeDULo9ao9zz4dbv+Et7rv1YVA0mtctVRtgoW4N0hlN8pvSN1UMXMevuhbfWm+nRetDhU/WXfm
+7Jds1b9tSymqvMgLCKyzA0lsUXxVmCJKFfM4e/2JoT4l/eCdSlHHAZpnpRBReKLk7rbxvre9at3
I0MvVMfIF8AakKwtF313kgWn0pNfrwZVPr1nGiYkk7TR8bSJNQ4p0wuD/W3sHco6r6fJMyDHrkVl
Dzk9XB6z/bPWi2j0IFJ1ciQi+B0OpvMbuTV+02yn+Edj340Zo/x4bI20wSnP/E2PFTczhWsiycRX
jjkLzBVMo7SJtRk6pyFhvofKFSWzuCqvID+e5MaFZCxmSkH3NFJuw2lvnn8wPXneivpdBg+QGMNH
4+ZJF88wllx3U7tx16ErdcluqOisSyBRL0ZexSFp87shdRoB++pfv4pcTPS995TH6Gw1n2BhZ+Y+
ceM0G+70p6Jxa7Tnd6SmdTTMj4J+XcQNundSsMCyzGVUAHEHb4ifL113bD71LrBkPCgHdA5yQxVw
veKltdhUFAkxT7NBKqmzCmtCqFb/+93RnaRhY1JJcNpFa3Vkfie66NxaLsiz0rCFnAxpEW9B+JGp
JB6yXpUI65us4pkSko0zNeD+PzKSnnJ9852t7YnJAko7Pa7XqxGu8Ws8UYaE40rk45nLehNcJjK7
Qxz3rLqcfYoGkkxsRjCbFOa1izZEnH+xv6BrLlWIO3/sNDItiq2JzFbnxHfdF+YlowYhhbDH3E8R
+7o36D4K/bXMcPYV+4EnfPnIyJ5NzewEa2yHCRJALuCwx7pLour7osfR3vRdbnv3SbL3jM/kFAfx
/3LHZ6RS/645v+Xw78YfmPiZkM4FefT0Iq9XgpSPfTNDP6v0aa/iiAhyMYR7+WEkYmZCLGTvhjGx
NbmEaFBmlDekSwPRmVb+XqPYrM+Tr5E3tUTCOPmC0dA9JHqhEZ7cPoOGjAwA7WDj8s1XauW81Fez
7QvC/zcLb/dvG89dSriFIOK7jXmbCuBnlJEi1qozp4JzOobTQyMJTX+zVhLnYnmeuO0yIeEwZdw8
ooDysvXN66zoYUy1Yu/q00a6z8P/XKG28YUIiGZEpevam412NtBd1kpzepzNc+FsYwh1sOU1eCSq
erFVk9rxMsQ5ezWBQbCnRB/SldTjm2GaQ/R9/VVQ81cX5iwDebSZUDV6Zh5HsvGensdf532hSBNh
lEP5idqF1+taq4hLLGkGrp4CTbiHSLcpn7yMUJKaOSIY+Qw68Lztl9V7D1JPwaOuncBI28bzuZ4I
Vded0amTH3LD1kwgoVipTRp6pH4YVOpmZq9FysZVlHz9SIZeztQFfinjFDdVoTCm+EyUnwqIZBQ+
JFHISWEUDkwoSnIhbWjk0ce4HskM99FexsWFBXYYb/ScTvOiPjzuSxeMPcmDkKi1+BZyCcdt8p11
4RuuBEAyGVszTb+rdQ0Pf5p5wNM9+HMn4rlS60IT6Vz1yTvvnuOBmjV4+SsY/J8/mfP9CNkE9ulc
DLsZasV99KCgkhDJg9geFcs1j7g2lIPijPhCZ52x9K1hbDQL6gBdrOQVTt4mQVpluvpKPkGIml/k
fClhVG/xQTo0PP2H/tgmCuSX6Tzqsq3xNj3gstnYNuPCfu9ZERbJt87RtuLSomj6RZ3/09cuNZ1C
P04xMxaxbTXD5yLHE5QUYgkvz6D5UxNMszaY61veu14FSJ5m0C0+lMnUIm2hIisvG8GQzCK6HHGl
xjJIU5I5CsOB7P0ygtjeI2aIvdwyysLdjkQosvxskimX4kcl650wBqCfxCLKuwUYMmDchdyqxMwH
DYvOmJtwNVKjgFK41+L680+wH4XmEo0Rprd8zXRBYo1/dsTl0A9UTta9ZLCcGo5rYP2F+lI5DiQU
SBeAIsFiIPxFNhj+9RWCZ+nQUoKQDvo0QD/KmpH1ar/qNnnXnH0CMRTLYTfP32irYcfeJEoVDFCV
PvljJhbOsbQBIYkh7fLJJtWRyfFVj3n7FAsV4HGXKOopic3v22+RTvao6OaGCgHZVBcRHb/TwGI9
1n7Yl6US+wBdl+F0V2Y7B8xOzX6rPtay4DLEdx4I+m+Y9sqBAKX628s/aDxDgCgvRlAGPVqDZ+Nw
QvEmpx3pHGA9f5dhr7LMBRRxN9hwI3Q5o+IWoLbjKjTwwKZujLdDmh0A1ycREcylrQAToEpkrUpH
SSXU+wb31T+n1aDLsLeMXNWVdyoYsPoc0u83pFQpVGC7Ys40v24/mrVSUSgDo/XPXa8QU61Zog14
PsfUJK91s/UsoATNlUYU19URe2Lpdk1UR9szwHWEBDuuGHizT50sWC1/sQ1Uy39dLzThkN4T4Is1
ecOAJDKWQR3rskTC7pi0H9VJAiVYMgyMHxgUVI1HdXKsRC2VTO6dyuZr336TPDA+CkdTHrgwKUlM
Phfmi/clFAEaI+0yNPvhwCGtsum+DVc0yRwH8BfBNJ3EYNDjb91Xhz+pDJe/PLdxHSVIqaVmA9WM
BfxV1LG5eZ7JkOuDmdRfrGmrHTx+X9cPCE9diPgPFh7AsA8pLrzS5k34ZS9M6eI5yJ005I0tfeDJ
AtqoWPia9g3QHMbn2Ayb4DX2ZmpOe68uYeolmIsnczkhuRSqApwR3FQ+Zr3xGw1RRCAk0VyhVnuO
plAgqvcR6XM1OqT0pAvcrvRdl9gkQo4oL+ZGDZ1McUzk9mJ4asna6kcJZaGpvQsZnafhtQC+M0xt
g4tp3wiLScORRtvStQ8mvCHDdwiAzzShmA08KJafFtvOdW9LAlLTXUMDbUWcMx0yMw+vmWuNdZtx
m7uNmw528ynZq9MhX/kXMgoe+ikOdSq+ijpW+g6DEtNX+5b0UhhXLZ30cqeZw0v/ds8GfcoX1lJY
vxv1SVW1VxeBsgveDJb76nv3Fqj8/I8AinIWHEMDKvJAH51p/2Bk1FSa/RBIF/1/ItNMudoOzwkJ
TjhjvGAwia35u/bNBcFPME61fGD6NSndiBfnCx5PTv4N6B763w+GG/tQWMpwaWz1PiVgQEcjttis
0D5M2wNU4wbxt8Io01bEB6dYWwvxeXP1b0segNYvTrSzJDApibs1rpYuMLjDdvIjqbI0KvpbY5/g
WV5Xw5fbqxl2O1tbWHMf6FX8fZDlHH5S7Bef8jUW1fLjT4ilzPzyF5lzoDR/C0dqYsWrELgLM1/U
A0TvOuOKrKIG/1Wm0GS9XjyUCYsOzvUOw80oAK8pZeFO5aKIEVeEpv9NI0UtA1zs23XqShfqb7RF
R5AfF6+gAGNjVjuRsxW7PGr4C2WLiXBZhQPR6F35cROvsUqTDN1vjfyZTKiR7Iu6slO9ANIo749F
71SAPI5S6xtoaXOEqzqTmCjcvGvvGMhi6Y7ilQuYluOSSPjn/tRGtVugfGZi6z3+vD8P70h8oQWN
BzD5syDkaoHnWN38TKM9nmeH+xgLYvchisr0at4AQB369ZMX7RLOVh8NtIWkLgjLYi9+Y03gjZuE
hj69UGEBotHWvexxJEjRDrF/N1UowsNjI2Z9bTN7M7tScl/A78tijDKgqKeUpC8VW+6dq19vtjgu
2/q6QEz9CnlOoV2Dj+8kFahIPz58K2QflCndoce06sc7o/ERAk5OT1igjtiHpXcBoTVnnR2Stau/
btcY18k+dt/MEa22UT1LhQBJSd3x1v22A27TZO4IjPsg/uu+6kELJ1OmTluvlyE3kMXq8jNrtqiF
nedXut+5euXRM2Ab74h1/+tCfW7ow4ModolUxA+x35nFdziypfCXqAVBL3w9wAeQilt64tmVKVUY
3CtURZacHjAzh41SQ5am/PGrWjJbMB21YuAUyVUu29zl0krGuPsE50wyy1MtYIz5BFFufHrS6FRW
/VcqVmYz4ASm5A3iUBLIqYSUzHtw4C0J7CE+Q7Jp6Y2/CdD6887GRs9B3e+woN7vg1YcnLoUmPNu
HzkzA1sm43QV50pYOOmxhtidbceJfKsF2lDaX3s9fXpP9TAvdkBIrz2CxH9cAH7aredSsrnkqMao
DYgt3ex72gJ/bQX9dV9KD8fUKkDKJJb6nvLvs+GPdzNv3nsoSxzlOeUK6J6h++jRERRo7wnHp5vl
+nLlXnra8JMvmtkjEEAaJOImf4L5Y4dVyPCk3ACwVS0rLeMmi8Bit5+lToZH8Zmpr+Dra2NTqyJb
x5OPVqA3o4rbVTQgxtaG4W4j3tZ9ZRhPJaHNnJ23vDdljSsnlLS3g0uE3B3NsA01t1wUumW7XwI0
MnakiVdXibAKBeso18DoUM+V3Xjv4z33lsU0jVorpg9HDwvelyB061rty12bjiwqi1qOMuvlwn8p
5f1UPk6CxdiGMykqnVMkYufte+70sheCYUVAsHFshTutboj29RLf6yCDaPtDIjvVAIUtUIizWjPU
pAmceOg1ibhHopuRt3mQMe8tmWefsyIynbVLbwfWme0HZNbarqiuTfka9Zh7qnytdm61PjJ1LWfr
WjMLkCx3jvoQQwnPsPTg5mwThllKoEEBTCF0LNLdkd5+Qbrukn0Wq4OvWt+FiEZeGZ8fEhecO2bg
17Uqi9XQzw+L+13D5yQkKo6I2ol2YHgps3xGPHbOkfmgL6iSLV5YfQV75qkFn7wd0tpFsNxrH4qL
WemwWSyz0/Tcv3WvY7QptZXgbADxmqlTRHMbVDhthX63ZoG+NjrcQFBME21lMv9YwJA7b2yzNtr+
x/96/SfKphN/+xA5kLi2i1Vzlt6CrxsH2e0zG7p95rkrc0HZmt40gy8SvKIT1HQj0l5Bqm3XT9Q9
JDZgI5LK/amjf5nbegdgnjf1cP1UQuqS/1Yln2UCkCk6y3Z2tjrMJRwdgczRXphsbNavQvKDHm92
CV7ZMIAk/t4bnv6RoWARk4etinnt6ZdWH/DxeHF90wyFtOu+EO484dHpMiCsp0wLTTpSF6d+JbS2
ZGFpfjtQx5HlwvNh7ooXNfwRkKIV7sG7AT4eAY6EAYCAlcMwMRJg75eky+AmKsNx6sYXQ6ePmjE3
yV0JnmlaDZ5Cp/X9qexWavXcoAnubYMP3sB1ZFAee0nM6SmO/mpcQ+a0tcC7fryXR0KlrhH2TnU4
jnpOi2L5+e8Djx9qFqXRMzGVRzkQCNoJHOobqfCz7peoHwe84WeRxV0fpC4/nRgk4qZVpwk7vlZ+
s2UxTU0EXP18ij+QSonUtv/xhK01qo3N6AYej3hwSkK/KtaUkuI/DjguCiyQXFBDlW177X9BdU0k
QbikbaZPtz5UFls/4CHcPVqGp91fwQIxvmgMRA7DKx5RjuHdsSakDZcGnbQf6WXbfZgvhH4tGTEA
zBTUq3rjLJbspP979nRHY/HYfAyvwfRPoQYxbCtm+bei3zy9G8s63gqpzzDzmpdMAefFHsleV6tQ
/J16TMTwy2runFxBcLvSI7yv/jHSk1e52GSOG5pkc3X7Tq+PEgm2asr5S+RCjk2P0AV/itG0wO2q
XOdl5Qk64megvdQ/KXML3lvUnzMkS5YfioPvBUG4PpmJHZedhI9N+FJZLlNEBAB+4iJR+kQKP8bu
CwgCvdx4EuVT74XDMvKlN+R0OmROBYoKU1Y2yBkhMepsIYHO1N8FrXDWPheCIG+RVf87++9sJBu+
pSfpr+89BYkgHiYTohuu6tK4mcaxnbKZowiLg1Ul3IP1SC4+hgIlw9OeQ9gwLGE8Eg/fe/ZZnxk2
NRGG4TyfdPbSBm/jmL3f7KHXMAQuWxM/hgV7KRcH9C8Fr4WMSbbi/1Xqzatv3n374lpoRgZ6f+6x
vcbWdelAPi0WmyNZhXjYzSlOceHchoGtDoA04iKnRbKOgxnOIo+tQixqg3nehf4m77EUyTLlyfXi
0HLM7nzGYzXY0YfcLvDTaooECcMRwYyAMPF01rHisd3w4y/ySanz09x9ADjrfiomLCll+NP1oV6k
J9Ul5C3Hn08LRMjoIWaJ9wNXCTBCpsjOMZZDkeSY4TYOvbMw48N8Xnz3+p8XBurCp3C6Jj4CkWXe
hVWo6iHHRoX2bbCmQW+Fkg79r1ncQqQ24N8mcO3w1fb9Qvme1uquHlBp6vLxD8NV5sJr4lALqWt8
N2zai5/3+GR5450obChjT6NtxvMnjB3LdZRYjTREAMZib+a+2Ma2vZDg4UCeCVpo2s+B5mcM0GA0
Oz3BFR6EG3VHvJfNW8CEmFOHusafS6xLDDGeDvBRmcIrwRXKuwBGgh3REKLZlPB/Gba0rs2T1Hxl
8u7SDD8+ajenDLo0cHFDUe2HW5jQcT/6ZH24I8JmocWfOcsRlsypuw6N+5G2K/HSBAFzGCA9jx3s
GgYO3gi8ELkvzOxe9YcepE6zqIFeFWKMVNK89NtkTb6yDUQR+IUIR0q3HUA7jqnAL3nWmCT5Fg6h
AESzzuXGZNeEgsh/6ATjco7mx+HFa+CcBf14xRaVNqvcAAKHYj0oejv0TGpFu/S1Mja5i9ZAsuvY
cHWen3j2+IbWJdXk7kKFTPYzGgnHBQ7SdMX6axMEOzYuSYcmjjcSObUkrP2fM562f+JBn8zmO35k
5edblhIFcyyJNDpJ2tU0Pvj8L6gQnuhOC0eo/Ba40CIUNV9lIeuen1RzXTNCkvfxk6crskm5VcRg
v3X9himjGCtWszfWi9o2ezS/lY0DDP+b4nUF7tiI6aoISIjYMMgXBmuJXtK6v3qHwANYZCzWwinu
9BUZkZ52/ytMC7E5V/2uv1QEQr/0s6KEIxs25UQGQ3U85aSqeYMZ8Ikjfvf/fofJtiQGsvXZMqnE
kufClHbNMOc7jtCcd9mtpAH8Z4tGoOW5ARuBUB3MmJEoa4XdqoFhh/HGy1WwSDDpclj6sEOoyUwD
Ei6Yoi7kH+RR9KYKpJq90/LbjE0gaFUgJMQT+5qYfH0LuYVqQrP7L6upTJMdMq6p+NZvANYfJmSs
xdmHSBztgiMCfPUJocWeMnVJ7zrOf3HHHCRoVyuhnxdXdR7ngJ7f2j/D0yYvVbLolWN3GJbZIyAW
k07V70U2f4esF6+t8y4ltfmklyaHMGJQi4HrtNCDVxQZRf9WULJSxsn1u3sXFETaHuHjZKl7xeRf
OxvrqCDvrbuCLofL/mRYGcuUkd4dErVneaYYKW1tMuxTk5+XQTX5E7BtCpamzZxbmF5sQ9T3TFSi
sxULR6BUAwEtKPTcsG4UlZYrqSTansi76UlnpvXTsDi2jk8qOPp16M7ztmtZ5QI+DNcPuq5TR5//
XLFDhVO2uz3vJeL4xW+w43tYLEniANz8GRE942P/ciBfdGxJC9AiojkuN4lB4bGgsAA+bDNPPpgX
VIwN3N8a0cpINatPdUZZYqFUDJn9XnEK593vGHDc7VGWC/vf3rfBanoFARnE6oBHPrHDAewz2lb/
LeW/187UQQ4IjNJb8NGCXTpNLaniwWdWceaCwu3lqm4EpcgjrXul0RlQYjYOpCq5oFelvFB66lUM
uWHcNno+iJLwNLZZPX1HVr2c7ynKA02im8GE4FiDlcAApGczM6VDJB/wWG46y2tgwNQF6pYcVFDg
VV9IbD5aP7a8fiwDs3gTJtGaVkU6J/0r6iMDOhmh/R/EhELC0nsUNoxr2Yy47GON3YKq+4Z3HAW/
PGuf7hJgeDfFrqZr47z4JX7AOUEPSJ1jjI9p21IlKU7af6CVfS1bAQbCShbI1vUT4p40+Dv7qQ8d
NQRHZtJqVNgW0Cz6W4AdR7yI9kDtvsJqMLwBYboTcxFXy4iRPf7nKSlaGOLtYqX7KUapqiZTsJJp
OMfQIf34Itxm2mun6z2LRf1TmTo7GINI+a8yaw9VSZ2rJ5TG0tccLpgijj/aNRw3TJzo8ghk99e1
7Z1SNj8UBTQRQyA3dsKUGfrex/GZy5fGaJWayjUw4UzwWfel9JilhtpaszidatW5zLdcB5xpRnPF
ctmkNucVLo1A5MTUjwGZXNAxc1NQsTWI5QgQlmlCs07beQ4xouuVi5FB3D1OXdjO6KSNp022z2Q8
dteAEZFZ26H7vdcvE1QV6AEu3BuVRubOlSTYR9fU6IqeqM8UaHvU7d+V0CXSKo6cxHLyCzL/sWyH
XIsFJ1gIc9oBvlOFcqzJNMAzHJi+VCBszQkBCA7+biJ5fGVjOuAmXfmV9vWCkdNK0OldXGcq+f4B
l+FwxUShOzm6zousj1qi9mf8nHxaYs1l0QCvNq1SqkmKrvBo3VmZUifF1Pknk3i56OxUi4fqG1ou
GrNXkFIWTWY2aMXnd2Moe5dtP+nH2SqBS9u8IOXTXfNtfGClaTOLFCh9MEyLUi/1ZNN7vlN7TZck
4kNAPa7Gc7lbXghdmvCamuLv3HBmDtS0+NgNQ+1eNtsLC5o0cexu6ZQ9scrNs037up/fT3QRg3uz
DbOH1CJuYomITYR6Wd7ItsYAQSS16PvvRz08RxXQWfXFu0Z9SRVGJ1vujaKLCRk3N8bNLUhWOiGO
lvsAmKkD3FS6mgpmkQqIB6XsKVeUkc4amHidw27aFBeoFMbDld792vPh26GlKX3dAluxYApyYDz4
7OFkfCZLSuMR1IOym+4Aj0DV0prKNeMpPptIcCqe0axtI3YESGiC9ZnJogVlMvsDVjsttcy/6A2/
1RsTV3HZ3S7lNqQWdYPrJd0+2wtW9gMGRZgrRRes6+kVSJvLRSFqwj5PeVxsGJaNps41twTI8/ei
qC6mrLK1Ed40Yf/yozrgEALsgTdU3s0vFk3rJ93xz+RItmzaxeSbCQc9BVx5QI/3sCU5EJaqSiR6
e3HD8ZxsMhCNqLkNWyqPX69torTl7CQISdx/33WsLrrn/MU0WthFUVOUYouMwNC1V4A+oSBOQwnQ
Wo7HgrWjTdxBk/leLKlH2m5AMMMtkl0zKf/G+Fi4/dLXSs7VrTua67XJCGnfRc9i3TfQtN222chN
8HeAbl4oCIos11B+90gbZnabU505nWkKiHuGzjqPzK0Dqg5TTiDUHIwnyslcUa6LG0Eusca/xqXU
wxh/Cz6hDcE2xhkjyE5P/Ki/pMU2jWpntFiFIyYRb5cRBL3A0V6bf4BM1MynC2kdESy8qXnTLyny
BcRuNkiePkTr7KAVxzqD2Opl3BYA5FlGuHnfY4Umthite58VLw/zb6iDtq28e6Ns0xGdrpWlaIPS
hmtiMQvSnMogBlzV1ZuMmDu4qCMdFl5QGS7CSjOwgXO5mpY1Ug+XVaCbMnYISn8ItHyfxzq//XYZ
XheXn+5mySCiH1gIvl/pMOX4TgSzBnkdev6WwEZNaMmyQ1dOjTdeKFLWxb2S9GQCge0GX/hn2Y6x
G8+lBG8VEtqLKHpk0m897kCfOqhttFDFQgw8pVE+I8q3B42W2RpjWGCiCXjLoAojyWzBaqHl1Zvv
GhmxZYerSvbpR1OjvPJ4h0FXN1IUEd4TY83G+et8c24sgdavebb/pJD2YMhEJWaPcewKCDefCBZz
GY5JRaWrcP83YBDFZ9Yns4WFx5+LHPV4IvPoTr+3UueQCWUf0ZGf21NfqLH+n27sVsV6hZJYgqjz
6NpTXlNPiHzbuszUFJeg1LfzR1BMJfbI2+IoA01ampbd3cfImy9RAufovmj/u66oves5jGSiiNqX
CyZ6jTaU1LDpN/y1p43hLhpKPOy5x/A0rhIPGqtBPIHyH51wAnq4xhAkvbNtzemoJ8z9FTyNAZQ1
pPxrNiZhu6JQ/SjrYLdxT1GySFM44JUM7tNtEjSQlj/kzOtKtVJ4VgyIazTvwiFfi/yhOrBT6yex
+DqNBco79LghW+MuZSVTwLHpH+6QfdxjHsCKj4JUTrjaVrK3QMVmWDaQZGVMKt6Km7Y3+kWtLuSA
Z1M35mzQJ1X50sPvYdy0JvXHt5sgXJJh6Sj2r1g7cHxFnaPWcKBekt8H8hkE5YYo/bfmIqfPAsCG
VP7UMKPlL7dI1AYOHhCbdH3HKdlImy5jNEhRKcgx5Fq59+DygoeNdm/APCv6d9C5wqdYiiRQ1dic
qU+1uUY1de2+2LAdMlzlflp2rScuZNXEGdXs3aWRfCeeC2ieF0tw9B0xR5GF9bwzS5OE8eO0fOQ/
XAmCEPyQCeLF4QoQju41RInwKxak0vCDL+473ai1/9xSoY73Yg6WxgAo4tJhipQFhyIHHCLr0/iv
9nuU8oRTGy302SszaxeWKvQYjzI0HhoC7sTunOcFEE/NXtcTrwPJ28TExUmSwJKJHsY5hKtPzac3
vYw+3+Hx2k5bhj5C+HaXEpLC3oIebMEFxXzlktbPsd8xCSsOMtccdsa7H8M6dM4l1pcOcQR+wz2q
7ge1lxem5+IcvSjxmuP2rFNfSdchUpzhxPUEcaPDeWFDFY9tQqE30uc4pEAT5ai8rI0bMPmVZDVn
BDYuShVVdmQ5kqTp+L7UF31fTDHzJiUwA75vjlkRWDLn/iYGrmOVpSDM9Nu+BM5utXpyoNIR4jVj
IjO79YDtfzS6CtziIZS7/RAseL5R4Y4WmRIwN1m9nE/U44qg25FRUBogDylcycW43+xM6QxYZzLz
X+7U81FZMsirUtQY6E1zfmmCqXl9/9MfpCKd5hiimowKrwvD1PvSDSvMcNh+TKLWgeLdneFFbQZy
3UpIDsDlnycVxvIx7/0cPm+VAVx8YJj32dCp55PqxnE0xLNdSZtoZampy9mlzpQ+rfVqrs5ZO1Gw
lh8P3R9uckzaY2Z8rrPzeebo/MGYCAPEWIZUEAXG9c50qC8H0wd1zTMPuh63mTo0+aANgapQZIjG
+Z5vD8oNSy0LtgnD7sCXvuLF60iUJlAHxqbKMpcbUjMPWRSby9eNFUEZWj8PQ/sMEwtXjQQtSuNU
SRBKb/RsvZds/z9r4oO68ShPUCQ5YmQ6ergcraJUGJAUTdlTxt3L7MzSzudn/reNukGJ2GfJpp2q
umHsjlyVF716+S12/Yru25YMnDyZ3EqBXv8XJotdiBr9QgLkCXNZW5sJ804fY3FCfRNquBr0JnAj
Bt9r1kuWDK26BagTvI7f8CN9Ai3nuMyY0PvwBFmbZM28OsopADLCtLKhMSeRkK53PfRnla277l0i
ST7471NgMZHg5YhHPWX2lmwHZJRRoUHCJcaBl7vkL7HKc2C8FbQAmkd4uTyDGypjBSQKbiPfi49F
iSbvF3K5mHKAEpoV32J8Q5LuQ4KlOT+bPTe8a2CLHtzvDPAefVMir2QUrX708RgTjbkcyIT2+MlS
RPETK7SXTMtD9sOq/4Pe8DJ4FRicwTvZjkkiz5SRtPaxEWXBeIZFKzlb1pq/JaHhJhk396b4vAWS
U3HOT8KrYuTvSDmP7XdoNnbWvd06qFRRZH3BsAMsS7ldXJEXY6fHGRPvClAEDm0GUK9+qB2tzn3o
GPGUC/aOjonzqb9t3MKoNUgcDUpYfj3rwQbbO5W2YraZJYwIYs4Cakc38VM8sGU7WgPMnbcq6RNP
3ehw7mDibB27lTzVNMgQ+4NyUY2Gudx5/rCW4WQgpVzZqv0amLQbj/SXCgO+AzEmlO+FV070xRIT
GkQTIHcf4jafZWdwXu0650g1U3KzQrTsAKwJfGRri62Papy+0M4xzgs38nFrQP7c4qFo21cXAO5r
xAZ4Yp5ZQJj86R/Li3lInjsIAS3NQwGxjzIPMJPV7x5RnHNX8t2nZqZr4iSffFTEJ/SMbFxpWjht
oR3u2cdFK9Uh/FhVsNE5iMCm6WUTXGSZZwzSWWrRKVTlfVlIXqwGmfoISnFL6+nmd6iHNh1aDY3G
cuB2gWoEZfolVvhiYSJkJbiH+d8tRzurWc1GyF008I/+D4M6YR/YBr8rfwea0vojPlDxjCq8PXJr
Uu3fNjLfWdFq6VzDiJTy/55PmvBKnavwudUXCWfvULM21F34yXNbkxRnVS3l7wuhtPn6KavDyFr/
6pfN/GwVmeZ0NGtiJkItwB4qqVsNUWbOUJrUgQAEifHlFDUSw4Jk0lZ7nUBDDVlLdrtFEgcxJy0r
PKztIDikek9nCdAVRwDhVJOM1/zoa21R/P6Swoax9thvWzHC4/G8qUnZE8H7xtl/8QosS+EvACV8
Aa/6AIoIYlwoVhHEYSP4Y0SXXosBjuAopWSZDjaxLaX//NHMj0yNDU6Vf0+je4oQMXMRCl6BwBtJ
QgET8VZ/MeHbfdK/7sOlTwHpwf7hOaTV3tHeH15i4I35AlzGVoKttzthNSUQNAdbHPd+cLuGwSzi
eCQDIMHSJfKxiA3taVjMFmT7vgUTXYzCuTjvWVyfeO7VNpKZKz2B0dC33ckX45XrJ3JMki6JDzkx
o/7VPHOBA9urjfwTqBPoi+4KOe0N/wVMSXBSVA/op/ByU9bLrlqJdZEj7+Z4fCy4ejLcaGiBsj2j
Edh1wUr+OBy23GABK9A1tU7GyCwcrRyIhKSeQGVVx/Yyg9fnYi6L0R4yt4iMBWmoWjvg1tk6Ypox
9HtAsoKhUTzlAVqP+VGe+1l9vUPLzwGxZv4nt96kbUIFLYIEFowSprY6N0Frg2WpOHiOg8ejYzVW
c5hp0vyUj/9Yzjc0ZvIyyTAZtiaFcHQcZ2MY17c0zocNiekLJw44dOsu9k6MSh3P3Th08rgnNO+k
S2+jOch3/kgS+kwbPCtJIfy9nTO/ghZQd1lXVm7BScMDmhLWoUiJjilKA1dg5/0+r8cHsHJbUktB
oiX8hxJgUj7EPZQoRsskqTmG5CaLdh4MJc239W7ZlZTD0sFf4TIsjQkXYO7NjEeFxtMLMyrP5KIW
REk8ycsuVj+1+PgmuQHtfZBFrxXBUMgZG3wOgVDtUs/g9k77TFSs9jTTzczUYED3Ud5IkNPG5Pe7
wlGs6htzrQlNcVve4eTYv82xYoBdloagweT0mqC9nClFXaPD+sg3BHdjIzc8Tk1YSmWlXuv4/IzQ
1nDo9oljeBVovmdIXeEztH1/QKzi1crxz/u7h1ACLWwOuO2pPkvAoDNomrRgDNr8W+mLRGmmJz9M
syUEsNOlLa9C8ORwNrm0uOgf7UZoN8ZTQKhTd1LOJqkqPdJDbbUt2rCnwnYAgJZ9wthxD7TDe8nj
Ai7XBHY3P8rDjW5aNmyFZt6ExMGg9r9L/Zwii/4a4DoQO+gPXxBaGAls/rSYnBn+r52drbLvgUK/
Q7eJysGzz6G6P80BztvXqNTvL67gQHhhOVfm6SjHRtVAQUnay16+WL8SAzFn1L/6CMxS3I3K64jp
RqLRDYNQl6lgcVX+ijQtPgQdZrI793Wclu7CdW/etQEMcUUCc8GGUwYjow1Zkd4K2v3NDKCvtYEZ
Itm7HHnSALZrRKXFIddEPhALMmTjl6vzuCIA00CMzS8q7WTh9BX4+lobJOgihUVDJ7lVjejlTHbd
rYL2J6UDId7LkkPSL6JsuyRMGNlgaKFNQN1luA0oOf+gvNblcNJ+SIgIL8YkL5tdbRb9A7WRxBko
EPSdrmCX6LlWFC5ZDht7Fydcj/gS8YMLvfSJxzfcKq9nIcMqLoCHdYpynGs8bOqsaBi+8txdf3jc
rgUMOyoksELeVIymO+Zm5+9EAZGHK3v2y5Pr3hPdp0Axlwq7HTIKDyrZpxCT9gNjeHkzCGaa72IS
9laWE3vZyURnryd3WkKbzBT76dKHrdcvorf6WOJUPIE2nO9uVvQ4Psj921vel2PeSpp1GyVWfSBy
b49MdNa3Ov3pAql0WrprLMqd9cLiF76lKbbiNbjKXmLBWJV61HpbeViWhfcBNceWVvin59dUEdnE
UeuSdPpQp6wFYvGdFt1ZhRODQlGXea6e7j5z4JJ93NsjTqDV0F2AKtVfzg13Qt5NgI3SDQrUFm4h
2rwODNCZApObkAipKd8JKgDkxjKqds4gA3jrghl9O/uyWzSg+BoEEfJP5k985nQe5eFCsG2ukDo6
Dt6uQBdQrTTa3yh3LNaS0M9iyuI6mnPvV9oqCPAyA3KqMaZ9DgF/T+PzLE3o2bEW3U1pFPhMO3cQ
paFnmGJEwzxsZY4CctYUSwCJir5SJsSKdZwW1XQz/u4MRABLF51Q2wKheT0g2OL0y8Fm+xOIYrd4
r92Lyef0hJJ9Bfezcinp/tQ92rbTJkkpFbh/Rz3jd5bJIqvE3FmTX+Nr2TfpwOZW8qI447MRhhEi
L7MXvAFQyaMqhoHWaec7hLhqbszoSXskY9lU9BKefW9AHaEwPuxu7RXGy+1jq8QjRFPEEBezuRi+
6KwwXB1zmfwkk9voUAFSwgrv9t9HgrjrVG4M1pmldgUDoo3iRvc2xi/wf3lYjG7ovLgf17rx8BO4
gvWrcCnMCERw6R9WczQ55JxIijxMq6C58+MYOsX0jeVu4npQJnIfCP1gbkr7jJGPRbKWfR+wLGdt
TFZj2uGROrjTsomCQAQbWLGWlxZARbQVUG9A+kr9T5zFVBzkGQ72ZNWb5yRgKIhr5/rttzhefi3v
Kv7vLL2JQkVgumwrw1JufpMl4JnXJvY1rBjX2DIVi6tyqLAJsaMxwKDiPaQMRR2iyFBFFQOkoelf
ENhf5WZSlifef6BD0ZOXW32Fsdyh5+/kCwV1Jp9lHNfNWgbF9gpq8+2MjkCMuXp4vamcJcLnCMqR
HddoC3CXEe/frMqZAUkwUskNu5DdkYqcmop56orE8BpPRbBAjNkmvxvTcW4qaTqakd3MDuFcYuOa
rD2ODKmUnaRS56rhgxmuZjRD6zgVj43FmKiL79LgyAOVihnnBlrAw2GMvDAQc9O97MYzsKQgsmDR
mIU6hpw+ALgqw0pdpzJN/vAFBhKpe8ndF3vfukpA5P4vNxY1hnyuZ2g5nW2cAxqJtUFW6+g5SVpa
JcLCVjESk8cqZZVjGmKy/5CltOO7B3tS3SOr6YhwG0ZetW3QjA8iveffQH/Y4iExrIo/OiTqccza
ouxUqiScapyppkjgevWWKgDprcmq2JBkO1bO5vVHPXVv2hy5ENl0Ac/68jpuh0rypoa8S56eYDWI
CJYkzaoZhAytyal1w4f0H+JlOBQhRaRf9GVjsATHwXfINS2dIrpCq8PERtVhEm4Qne806Wj/QIrG
luOwyES50/54zyrN7hrLYbq9fqrPAO9kjGheXdz0w3a2j0maFm9CPTdR6MFwGUe1dXAeFEBEQeWh
z4vWKpPs/5rvnikFLB0EaZXXlCIy731NElhJNgYXCoHLdg4k4oWkVBCpw+oPmf0ankc6AWFOpnc/
Retf1zI0nv49EaDSjpgI2hxxuMtTYTiFMuwcHHPM1zXJKW6gfdAm4b//ZaSbIQKrXSlDDwiSVofk
JiqLXX8w5bVwbDcVUvLDI+th7uG2NFIseRExr9LZDkWwJDqOWBObYZPPd7PDTqKTpz09jKLqPHCp
rB14YSdtakDeU8frmT2oDO+1mdIJ95vwieCWaraQi21y6eC/pIhWAWRPsRG56vtSAXAR3XwxM17q
YgfSbhgsKvhyK9UUr5C7rpEyfCfID9eneCglP2S9XQQSUNx2MNufwk+AANgmC6zJc8+wDoN6h0t1
j6JDF5vWMv5bf+Gb0Yh5sakbT3Q7n12K7TUWtLhjvHLx5IMrJuBKxfVB/iXEslrmjw6qm9JWIwKG
R6CUmmiu3liirsDLRz0Ru9SnB2vxrYba5eWHiS25p+SHDk193kHkY3z8i85hEj9+9wxZ6sPHEk1+
suLdWwF9kcuN90YiBcp8jM9QSEb89R052Y4K25aRdJJ4LfCtESMjFP4aSoT4Jy+SovE4TOMlso5+
a4EEMto/Hj3WFNoGZmAHzVSDflYDkhur4fUEtkdxziqPR3QAKIBL424LDG6DARpXVoJcVrM8HS5y
T4G1oZhH36Pu0fPnwtcqwzepKTegjMARldqb80FcX2pPLmpcqxeuxcxMRkQ9axkZtubN2vhdM/hv
XcXg7cKTsrEh7f8yzSYOv2yUzvsBBwxX3NiFCVj34bJHvQpXl416pOVxiCzsr4tuPFJJIw0PUSqs
RN8+q5CF/DzGrrWt2TqhJctuq7etxU/UF15orrX9N7g5iv+PUGuOI45CjZE8gQ8Ob9zEdnTJG5Pd
S8C5GxD6kknUr7JQyq7u6qkrWc/bPvL5IQSiwrGiTnM0H0OFSq0QZ96WVaL3HlCgB4AFgfdY+PQ+
c1kiM0CmQaZQT88u/8gzBXhn6NqROKrO88dIX2uYfo0Nq/ChtHaNhL+uNlgUkrKrJkOV7L8kJoL7
ub/2Z+M2jY6u/Xb/mjctABFl2NFVzomR+9eCXKKQUejDZro7ET3HBK2SnxYRM7KSLTSWElG/lmrt
Kg6oIm4+gckohFXyk6inVHJRbcwUiQOdbTuBEIkEvrAWpssLZ6SRigKFdaD9tyT2diy4rcgHoFub
AzzVw0TWVAbN0iBDYglSLK5wMlrsSjlkIAyKPot1GdnpLCtHH8Rbfabm9tXYvoHPmDnoRjd/62j2
IiAfHfVri71J5O16FaTHNEIog6Caeq0Ab+xLOlqDniub6rwOaX+i74nAUjC1imOC/09RiR2VNpyv
adoGMx/kTZIFh4t/z1l5ZTvj+02V0SyRJVtsnY/S/7IUQnimvhnSekj41NeVVfrOp1EWCwVdqzC1
Cmk4Yk0MZRIai6NB729FFpeXB60VLhqFnMhpWlqo8Jiqok6OiBoaAE7v8EswFVMzDNf8FU37LHRV
1nEUaxzCyv6VOjV6zYmsSwGyUL5sDG+Y2WLQdnV7F5ljA+tay0iupXqXpy1ijTu5BDHPq0k7nvCt
pe39QeLwUt761WXtw+mFY56zjzkiToBVFxUrmC/92RIX2guj5hMnTbdeGE9bvFOObQiOre138IKx
vVpGgTnPohreHRHj+5/81FlrfTQ0oTDX6nNj4fklGc+Sr7+gUhrOouInMTAWJvSLkNWJB35bNkT/
i9GzzFHM/kL6UpDIKXBKc8xuZ5D5yQ5lEt3fTXvBs4lzQ3aGagHwHGryM+jvDQQPvyTVhm5i44Tv
cFxS89nBH0NeytFPdbCEhzrTRs9oIQUeSyHdcbYYBKqweLLctY6iVthmRgBBwEO1YReD6Qu9+t0a
vC5/AgmWBQupX2uq/jvBLVC1HcT/Uvpv8mvLhf+FCdCrAFLB/4i8QKHiCpVz4e6MW3vmsBtnx015
y621OeNS+mKFK0fOSncaaWloyDi+jQYXSYg3mwnoU3+ZbQODqp6MUvuYZIC9hvV2bw306QOfn7P5
IefXM5Mk3yUPT1NwNHS0ROiRcIOclZlFge5jPBoN48Fhn4nhkMgKrJtbwNL2DiwvYwClzUuLGjW1
KrJlh4WV9duDEayIJJXC9GW2uG33o2h6MVmzWR4m3ARS0SUnXI597dwMwt6cotpxO/Z6MjpgVKgd
WzI/NvHGzKcrpq/EGU7cNvzCqnsP1I0FUSkIPqwPz8a43SOTruNGe1TILu1l4RMDJ8Xk3p5R1JsZ
pFPtm3fSfpvjH/h0LA7ekQ1sHFRMcAw8TPpEGl7ZROftnQmb5td9f54+j9abHLOSfYK4mJSLNynB
cIOSgxkyDOwszyVvXgzoBiMVC8+r2BMewd2YGlXccyGMxAuIH25113P5FCfZ6YnbIuKgED5DrYLD
fTCBjkuiguDzohOb8hBadTJXDoBBu+b4HiHkUf/cPFQkVjYMFHRwgTzb2LhIsrsN0mmraW77HWzd
mYyetqeTBEBxvjZF/bkZTRJBr5cV/naPOAc8+7meRy28qo/DWT3M/HHy/JR26ri2yWFKeJghS4jj
vBTU2suPDFwn+CP4jRcrW3PnHu+aHspLoOmBak+sZbn47wwgEZnB/tjGl/+t8VXw9RnMuZ6i1EFx
TS3HRIjAKb7nLIDhAOFar3LAtzIdMiQHBPDmpfje5W3mt2NWU15ZO+Q5+wdOJCfI/LMSiG6XHR8Y
ySR85OxCFVvGkLSokPycEAoQ0j2N09ksvIv1BduVwUk4mCGc37LYQW4ZsPteriZSt9MWB5KxbKyI
FKlwM9uwHdajrBXIHPmoD+CC/a+J2BKaQS5IPWFfTaPHsDyQMwhLRVlk6Fs4kY2FhRg4KtgNgfM7
ChYkjoNzUwuPISldmSvOVtt0NUDNoHXFMIjtKvprLAfcLuozOHa/Wyy/3hI5e5x+JvsmosgEcE8d
yiJTTWK6fyBrKKnuF2lHVIN8mAnoPYwfxzAxvrw7Ps2BBWs1ZSwmQ/0LpX8XzimLbILCJHf7QKIP
7aftoF3CUFSknjBh+jBVzyEbXGCfPRMgxvvf3xHOYElrvRYp/YZX3xHUZQLc8A4sAPRf0h4ZM0x6
xjgG7u7of90SOKBdjL3kapmCs1Tt1dVH3Uq0h4roQjsUotjun9GyUHwB9XRq/qVSKu81XTnUcnEx
/R+AGFBt0oRDCOGm6MqVmdZ0vXMubqKCvPMCifVvg5VzfdZbpP51VeUSTKz61dDZLiFW1M/VEmVo
e90shHu9wrt2D6AXYu1M7Vi8NaVo8aR9nLoP8N2j3ufllBh7djRwSDNQcbAHgmkOyo9KxcxW5L4l
QZqvi24dm0DbsNqp12XqAp3WgHdsPJyy0p9l+9Cdii16sYxu50LMFiWrnIkWSHI17dN80oMegz2x
8aZ0I9ePKHyGKbR2/A7SQdRk1kMwcwWgNbWDncIx9XVDfYgIh29ZVPCpcwyUYDthnhh8B5cZ2wK/
/7bFYlG0o1xHPDmYMXECmFsGEKHJBUcAnagW+oHe9Fsi1XA2oPTYa/BjKtIOxLEUdJOcRUqxHzD7
s7OjdHNGMZBNzlsGauG2NUdBpJUcsEA683t7YTc98UMw4I/6W+6XTeEuJNH1gj7CJ7NzQP1njCoM
SMuRdD8H64WkcXvdTV2pnqdKkY4s71Y1uYX53+ySrcGLXLapn/DtWGYUVu334C3UUqCxaxS5446Y
LekCsjcROEUuM5q3bIYvxMZ5hS9x5flfdZKif44HGBfZKwBgmtMAW0eU6enCvnL5Qc+n8+wVA6pU
C5UN9DeIpvAK797GxcRolY51HePR3wfeLy3smfYDk65bRm1h16TQHTJWThsWFbvlcUE+6joD8EVf
kmW3Eg3QOP9wdEDAD6JXf7O4Y6DVZ1IL5TWkFOGLSB7yD//ylBRmtnAHlq71a45VU21Wqm/Y1MI4
O+F68sS9mV/WpWfSQvFBLtvP33ih0QU3nRa2nbyQTM9D7kpsm59b/l0mPKSGAIeIBZxYTtV5FdK4
LaTrZLCnqcyf9JxXTZKfQ/UyE1ZnAh9BzOB1ZTQhK5C7Nhd9//slavNIabOb+RyZH+jtvlDh9qw7
Np2btK2FoEADkrimKW11e/i72xWnGh9Vn2lQYTGypWXMK+yh5VK5B9pnWHarv4vue10YjjCY62X5
kgkojLXRq8R2maAZn792KPoFrr4yw8QZsOq9kiow+g2SrXTdZyg9GiSLnIEBLAdhNQoNJpPnXmFz
bSkheri+C6mleMIwDCPfLIwfzMvgrOm5i50ekxYIs/muzICDpC2pzxPhOFCeHJszHP2AcIU/Fkyz
XcGUKxKaOIYnu9oREJU0DmtuxrjvxFAYCEtAnvpo2g2mUJEiyRd7qN1uLQVkCI84z4miWDhhUs7w
ELp/aB6RZjAE+Lo6z1ht54beHeUEPa5H9A1RyI2RrQal83BSirY3jkuB9TMCretZtWc6YtBFp9jQ
8dv6l5hjjQMnuvDzZjOVGowgJzjRFE7Wv+gzxZHCLkzAPS6AAyI5zn5O/5MdfvJccHSwsSljN0Qm
1K1N7CteN7ApLfeLEkBwe2kinV+TJ+qkRu5ZkCd1OjKz2EXu6aPYov7IqZvCtNsykBNN6fKC/uNr
PpmgdwKo06w0cCU2ukfvXNJpYThgNPMqsXNpkPfkJJ+6ye4EyjIduJ9b/adtfd3LVP4QET6BBLZ+
IpdccbEIz6cbfr/8Uo8PDIZRiSvJyTvxlv61ss5hsFqZRjYyGUNnsvd72yZOsYxo46Q+UzCK9nFB
bBzHclqPBqdTy5h4LRr2vlXajsuvQxHuVgAIT27d9KYZES0NZkcEGTdb+l4034hCLrgmppqU3/xf
fPHdzIwXjzxxBZCihS0g9C8N9c8cN5ATHhdiyXwYy9GwnTSBnDPssY14bcVVYU92yj+18DF6vbR2
c7uUxvIRBb+tGdttpW03oeq0O/u8tJFFz18NPJ+oypTAlXGj1kYAEW5OgHXhpFWi3afScsUa0nyY
lp0kdjwnzMOw85fmQ48YuaHi7IQK3ru4ZiLhnnCuqmeZ0zgUbAOYFsqH/HlPX1hTE/RdAHd89A72
n/tC809mYoX7efjZ5U1wmlUEjydUs2aGC3AQC2Nt1XlRKTMjYwLZEmK4XqH8ufq3x71t3TlPoIzX
QdikY8/vHLYOvKzrQFypHcYPL1lGrpfyTqotmwpYUJSMythzBy6lCWPZkhMn9z5jRGvM6kNPDiM/
Pd85EYF/xYPb5EhxXb8pB0S7fm/bQ1WVG1wwlw3gtTDDCv6ZIAZHKRTNZR+eo7/oNeFMqyyHlbVr
A5tabTm3JjpTMAOpjfbBn/j91P1Lerbwo5glDTfJR4EPRf670NHj2PQxeifnitvVlREwdmaVq0mh
ZSmPjeUrBXMKopTd0fHfp1DaX0eqEeyn3GHKpXjNN1dAx5hruAXRjgtDRQxOkRIsu8xLw85HlF8W
AR0WMUZ1MyM7Nnc9WRORxp1QmKhPwnKjleBOVC4B7/41UVdSnZ/IKucZnoDOfXGZkjaYLZHVG6Hi
s1eA/hy42UAlBqMkp8dzevTQbwChOV5QVrWJgsAzF3pPMTml0mXyAB/UN6Qdbdr2r4DR3smSWqBD
ribNEZsD5/LNGwF4XBwtwvzfumCySxBa0gh0+yc5QON58aLLdfLf9BIPN7y/Wb9o5oGBKz6RP6gd
QHhqkiKQ0jq3PCzjFGYDqoXIaX5Ujeu3JaA0FMu8rqHH3Cznda/guIox+5e3/HQJDU0/LW1/fsPc
UvYgGTBDteRqzjr0/YtfuQW0q3gL8HqkSsOlQaw651bm7PF+XFBP423nFs12xrumKuX3TBRr8Llo
y1OI86S2hM8hiNX5d1Ujptn/LlHoMq8L8R9XJasiUC74SrZMYCYuSZhT5+6nbQkbWDVCgxzphJTA
BQZn4cF8BibAFNsfyI3/5jFiwWseztDvxWbHX1v+oBQPkbivOLbqbQOihRuXjhlEatKPz7rujVGn
eocnOqmHfjrUwt0YbNaqEy2hSHJUbPUbcP3Bvr3FtzjAYDoPvh0PiYdehwZd4g+dHy2ibVeSRwxH
tsabqHQ9DD06Z4k0pYGNI3uAWubAdrgfnoLCyN5Jb0dukoyMOpSrw4s0YglHaEg8PJEhr9THmucF
GQgMSB8EV1VtK4q/bJk3xMDOlGUi3WkBRo3/otkd1vyCicCWoLrbw5YkAEtKS7VJNPEfYhiNWyq0
TUMILDiQ3sLwDBwrstjDSr6g7buafwAoipK/72OCdZdDe5nZ91u9kyWuOVoy7/18fHx8pXoQkMzc
BkQFqDFs7XIogyXV05dgcFr4nViUxkzYOcx9QPYuSP8jJkXJNC04z/v9kIZaTL4BNkjFsFdlnQMQ
Oht9q7qOVwyKLCuCKQlLxQ27qvO8hxndLPBl+Pq39iuO7s390dA2ShqPEfN5qRtQmyW4c6ecWf6D
6GTEcBcsymhFChH1zWq5KuTPC0mnE2i1LcDttvbMD9zsgcmD2KQ734C3Hoof1GDisyRr61oKj58r
feUvO9cdyC2/XfWz6Xvfa8dv3CCNyFIs1IumrFG2uyYUJ0MPY1+cNWvtyHwGns2H2J0nCXi7uASw
eofGCwkQYW75+3/BfVZ51DwlCSIIQ6L3Ugcf7RnbqIRCITN5nnv9sXyeOSXQ6L0laPj/1nUX7ra3
XxAym5c+Axf5qh51P7teXtk023mQ1Yro56PFZ1/HIeF/OJeOSmDK/c61NKMrC4r1vhXSIOUH9jmT
8g5s1v4vWroh5LEQVejbdQjRZoEb7L0l9w04OnJAmUGX4WCavMGSpUFqIvxvcbXegHmGnlMaV6hA
4MfR5pJs7CTtbna5/Iyfj1SFsAkIvLttYwC7sOdraaPgWOOomOGNd1HeDvYoiryFwqVnYfV3cNnP
5kOfpRsy2UQD5EJRW4a4ISK5xdncK+yl3DBZ2Vrx8nlrtHvd2an9BxD11xNHio1wLJzy4gPhLB/6
o7Dh/nFSggkZrJvzRmEkJBMV9coFG26eHqvH2Vw5Pk71EVlxc/vZVlXoVHUdv5psRRfA0Gmla2oW
mzXikrwvTXrcWCjjNX7HTPre9SiO20GduMl/KqFirycmEiTLJdKrEfbnMQPUTEoH7hBxgvTMNVbJ
zK+gblwIo113lw/RCRIRrFJYAPAkouQNmC9uAPp1Q5og9hKT5jkAlAYn/YYAkGUV/5HV9DWkantj
I6ihURYeosHoCiIAPMGzEc5aKdNBmSE8PjC1WoROMTYRPXydNFVNZJP+/8PjAS3TOcq8KG92aDpD
IX3bKaJh5/dHJ4ZHSlunSnhRDCa1pnm+aLFOGG2NcxUWjeHtx4CzqirOiHq8aitWiz/q34Gl9dhh
RtgD4B0DmZ8TjEx0T74q85syfNTxBLNxVMf+MS/BUr2PnFZBD1JMBCA/ytvZlvsxY1rbNAD2cMvp
jxbbLXZHg8rQvfPG4bbxta5dgISKlhvXOkqsLwIT0zlKd9VZpLq1VEPpTkWBjJ564Vg5kZwGX7Ku
o7rabbv/qtFJM9UpQmRIXoAUPKoXGMkowR1V043xrbdVKmf3R7AU3Vw4d4GnDcvwejAFBV1BOPoV
gKNH7b0A+WlIwr/i3eJ6EuEk+12wnewQrb6OCoz9sMAlluF3gaLbD7WWRYsUwmDl9IhT17fItZbJ
ePutyUq3RTvLQgjj3M3hS5zitmB2eOXqwO7kHX2wrY4JSbZ/X+UYVRvt8EQetRHkTrBfMlI2c/87
UXFE5iv8dWfFWJCQvUWyYA2pkTEzPxELSXH1t3G3CuRB9+6kDss9uAc9mUNmofqFdiTL8S6mr4bd
jtd73mHdxDlkfaez3SNZ956Re5x9OHDysfzRIisvTvekfhxGq3Ivvw0oCfVa06CKl7CH2QRRRiXq
DYTN0T45/skaDSOKfme8saH8OqowOs6PkR4teh/HId6gdGvDMtm0VuRyFpIeLh5IcwYoMMsoXeeB
WT3ycZX2X5PbsWnzMogQg0mkj8UYhj5n3CR16Qamx63PAw0NHwX2X7smsp6+REsLMBZ37+luhIVJ
IBxZZdRULGOYi/xZ9jp347dUKSRJK+IDM/NU2853vDmhG8Kp2f4sB/HtvXXpB9AXdPGEBeb/Xdgn
w3qiKW4iwlhMH7rGpgjItCRLah2V7YKBWolMSMBSXXjPX/T/wdRcXLRI4ORDVCjAwmuey4h99Hqg
SoRd3IkiS0JUR2leWTj8j5+dl80b/fgHVD3gs/ltDaIQfMg2lsbVySSn81FKZTlI3jNtGDav2/lE
jaGsMgqaTOSKAG6NmQNNQ0WFlGNuFJDKrFS2R50eRRW5PeiqqGJo6ScXrgFc1MO7eUuQSIu3c4WF
xn0Xpx3XX4cvx+ipNkbEcG5M638Kc4tXMRUMsmgLuroZi90MYwN8GTk+Ay6OT8ltNEN7eYs8m8+K
K4yfCQuBuyi1R9GTrRmryMf7vEJIXWo1Ka4uEuKaXzfJcvdwpeasKgyrQj3sc2OD/0NCD4lsHUHn
NAzRQ/vg7YqotcW/H1p8l0VS4wDEE3SzjCAyMjNIz1w8kFU8XZdspAr59LXAIgJFA8OyR9tsxA9y
c+bCZhteaGPMlHSdz4lCQSRrisUdnxAL865iafXLugm0U7XBU/3LHYxWFt5YtDG3NX6D0DEhccSu
YIeY19jRpR0ILKjEpGmr82wbt0l88eTxMOM+E+MTlazN3OAfLgycUZyLgZ6w402Jr5ZD8b37F+zw
Ut9FUyqA/ACItMrVnEZEiUXO4zYeqsySLHhLw/Cf1wkimkBnVzeVEjIqVLeQLsp7hVmaT8aD1DrT
/0tSdRmqJoQiyz+ESHhpclhWeoibtZVcdxp2EzM8XJ3YkY/uU2E2UhNjCny7G0e/+8f9IYXLIgyz
H/ToxGHzmfsT6TdnWT7Z+bJKujFDb+7oS2CpoGnVWC15+z634uhZKmfkrMZ3lrxEmNRm83PK+ZxX
B/JmgpHYyqff91QwaOYkLNl42hImR6yZJTbyGKT3klJdamf6xhk7CWdD0QJFkSbhB++t7d6YhTEL
Oba9GZvXKPcA9TYWMIHjkyII5flEny6cYFEiTETSz9KdO68n+u3DwNrAMDZRA+JCv7tgFsDbUBR1
0b29gy6wR9bQZ4renM2DkoK/RDBl2HaoDNayCUaJfIkY8UTOGfZcZ7fpDShr93WK5WhtD95+gbm7
IfwwwdBpccRNnSsvz0tUXWoicLYsSWJU92NroZcXzKdn6hPrsK/3gMiXc4fqrY+fVI45T9y1V3PV
3iJ3sji+r6Bi4Pn6pt5YUCWYfAWabd/slsMMBFLmSncVOwSfB2EaCdfX1niFkhVykV9QFHvhOGKy
aUkY/u+bcPZyjDyu2cC4HVPZ5U+ntxjwTZqt6L+4FlcDj8J+6F8Il7iB+TUVXoWhnfI46x3RBtt4
gwiJ0EpQfeqSWAvwbWGUN/0r+MSH6QYs96796l7JvYoxnuaIFAEjvkf/sgNsIAh+aKgml8dfagp9
3oLDvODwTxvNvOQ/E2Z6ODmXodfcq+1ze5IPXFYef1gkfBkuM0EsoSgdsBievLBkL65a0f7T6Dyz
eIexYeE1MeJZnzSmPdV18Pby4I7odq429mI2RxJhH6s9JytouVyrFAO8pIOSEN3rqS22KjzXn37e
ztU8S+zwcmnvzLHhvc/BzyHs6QXWBaFwqDLHHtZzVC1UMs2+MR6U+z+Gn4C/FfSqXiNBuS/a21rX
+fz9l8qK39ts8MNHQjvIkP7k+Bx+FpTb1YGkrwsYRpT/J6bszjf9pCxCVQnTwKiGQGdPzkrEbUB5
WWheIakmRcfavoV3YvXygMc20BDZNEQttOLQRG9KFRyZ3lldgbZVWE1+03Al1PUr2ypBWrjv9Mlc
zeCLGIoS+/F3T6cR08AS6FzxkL7MvCST2mGN8Ozf53pxUJDBxBKGgrOv2zaq13jNLGoJ7WN39Qe8
iHaP5JjqxBi2Ipj3QzRgNNNPHXyi8HYmqD4hGd9C2QiQklrqKY3wbGjpX/OIzTZY3eIO5FtTyIop
PWPBSMBFvt0G3q4TxAopnUnA/Prpafe1nZ+Tyd222Addmx3dDKpUB/alIw0KhmwUyZFKWCvwCKah
Q6dgYJT20XDU80JjnsuGNFxBI/FBQITYZnAW2l00LMk/Q/BBkeRKzpSxkg8neXsKr2i7JjFwM86Q
52JjhJQSMdijoaoTFqgTRl3CqGND3MTJxYVxBeKinQbMfxs+U+NlEM9Hr3oq7MjnsxlUr61gmTL5
K+zKW/I6diljkVrchLVgTZmzVUJCUOnrruW65vqyx48n7rWqrO+RIXYNvj1OIK6aozuts9bOVl+B
/s3VYB+NvY8D2+BVUSfIM+i7oNSaZhlfv7wFOHEhpjn7dtKmVfS97reJuX3o9dhGk/KDpeRozEvF
MDdsiZE2J6E2gi+aMxhotR3qUmxK09fVUCLYgiNgka1a8iADq3VgbrcEGa+7kwVNxvAaulDY+jVb
Pk8XLxGckNfwxGohffnufQLPKyY8gM21ZEAgvg9Vm5+0J/rzomvNjGFmwJNsh4rc0U9739snUOYO
Z5MMn6q5ljj0EqAsjH0T5uZeQX3d8auz3IIOTIYZ5Q2Z27qmABja73qJkYMsmtJQZfh7w34NGTKI
alT4HmdG8fIeDMX8P5XRAMXTIE9UFE1jHeZ9wfhcijRzYEBpiq067hAJhmFQkhdamm6o0oPH7mr3
q0Bw4/wOsYe3twI4s1Snhq8tHVoHy+0c+IXoXHHuG07JrnYKzWAPTngyWU2M9HNhWbnnRN9/ObJU
xoCMndI/09wOn47M6uqL5Tt3h1+JRf5nh7ajRg1kZMam76v6K+r+zAGH77MVKjToV86E0Sb47L5T
QsSShh+Dz/MEjbpIjNkQpOL71fHa2gsZRN8vCc7GoMhcPNcaBB+ZedYUt1zZYPJIqjX9fM36W9eB
EXpk/vviSCLGnHqBG4po6Mk8pbJX4z8QgCPFEnItf/wbLbB1IeFYTHCtddI4aXndCFrZU6xkh+wV
fFxpqQWir9cCK9HgblpD6kctHSAyKGQpEDHIbeOrTyON5zlfWgrLmw7qrCFKhTT1LAt0NtYwLamV
Rl7khsmeHWKkdXLVJ9x/bTRKuRZZgQqxdx9H014eooIUZGZ26zo/zCEb4OGAulawgNJlL109nFQK
OwJZSg2ieQR6cKanA0aMPztIh1RptdwED2R4zBrx5mqcARE9BB3Blfj0SIlxwwRrxq1IyLNlcG2L
cW1ZNBRHiHNFJLMWNatLzGh+ok5XBdehS5tICGJ+nwqwNsgdvDGEobCjb4aT2Xhcf4Jk6lOc/dC3
bJjgOLkX0639mD56K4JUtESTqWt62Lm4QNzpt3uKuzVfqDR4KRHLbrd4ZmTjuKlKZXhgEsib5WB+
btfB13epk70FYs3AxaYTo2CyCI9votNpewtuC3c+x/+5Mmma0wxwKlsMs5l+qLQZ0cmaDLf0HjXL
aVsTvhs0gf6f55AgeaRp2mv8EOJiIcavufLqrjOXkacWpf+6a13Z2vLgp/8J6ZqXq1yUCdcXUjed
I+2yCqPhWRw0UPCfKUnBelAVkJPL45gKvgX8+pWIYaQL0z12UOq1a0UrAIhZN9A5SNV4OEXYx+m+
BRpOxcB0sXcaXw4IuZqnHJ9PGqC3Uf91DtDRxP6zgdqyxxnloO4sdOTg8Ykh5D2Hin5lQsZjoTBZ
qIce9UHwghlMgqFU4HKpvtoJXyX/jtNioyyCNtJFnwYyuXKwzLBKvP+5kiFVYziwTLE9MDZzeTsO
+jpWuG7NFUWpSp0Wg44sn/04X/woRti0n5jAIo8j2agKJ3AVaIGhaESkb7BUzqu+da/Cy4wMQRmb
Wp8JgGAtF2uSDrNWLvhZBqvRHUoelA2fsHf1O/CUW0cCqFdsO65HbMaWD7ItB/fCF7AatEeZM+tQ
92RoB4cRu1LzTDqPPvEDwD8IX7WrSyJcY8gEtuiTchfM5lEQEccO6czEQvftEvYTnx+T23EpNaNz
u0dmcJ0rk7APN4hfX9jJ1tx61Z+lnaFdnZziTPTjxacVAtTdVB8Sj89rfwKfXboY/mC5SOS4I/7H
ganIUxKv2FYVVzm7eWmZ0WHBwNZaxExCujmsICEYwt2cxjkQ1qV/qjbhjQzgLg9nkcBS1DM9Z+B3
dOCYY/3XK092ppzpC17F1OZFV0TQe2dYC9UPwv8xCOrL9/saj4619RKn4VXE5uCwIdXZ1QFs5Kac
+ciQjhafKdEHkXuuYW027hKJg08CQxOYm15UqZKvQ5qxSMM3Y3Y/8/rk9UOpXpG/tVoDLA3Kj4yD
Djy7+MQyescSg74b0yA9eMPu0K4acSA/XBiRHeUK8avQ5pKXCcJ1GGoR+pywNPyJo7tvFLcV1Xpn
H/fyILvG2STafpd87sM9Vw5o4oClamjsYzPOrwuqALWnfUWEUt17YSpAJZMTOrwrwqBZTA7REq+h
ApVimGbNOg3muTPC/modGA9G4Pe5Xf5UwAApNvpett0TyjyjvLrFMiB+cHY+M9QDeE77Z+tTyw9w
DK8o3r4NYVdR80/yvvl4JHq/6E+SWO/awXjAzFQ2TDdLMaDqJpCUDHoaM50VGHwmfPnJ1PrYxZzb
wi0XybvOonIyc8MKiemXKSoQg65NjWAqTV4mATchCXW/VyWDiho6RaYvu+52INDWA94Sh7hxXx2h
RUkf9n3Xhe9SSwDQq1lrH+pj7zrwLHQesHCfUQ8W6cQxgg4sOAsyzVS0eiouhd1n4Q1DPuQelimG
ZyEgvl/zK9ouUaL5jLD0tObPLvU9B4xNgezgfvKUiFXmaHSUd3fyKUggHjggtTnkazIfq6U3iDjW
2ANuLystc+ISSwZrE+VaDUMT5QqMTCCZVU4ipvUAhnkwNd+bhvd0xq/lWmaTbdg7R/jPHfDRkM5H
h9tzrmsMaC2N6fdr9v0mshhlz+dc7AN/CbluwInFC+QsWrE3vXTDOsTeYr8sot7hVrt2jhirDkpY
KQdj61Morul+bYe6TMUftiJ77z9rdsen2k7FvueEFVHy6i7/ee7sv3PtmFA+srN/+4xTXjQu00Db
p9o4teyn2KZpOHNormPsUWAU6TdoeGHsGFe9pq38RDSuP11NtVl3ESF+DcEkktugGLvmmr5rBE/R
4n2CdNrSs2RS4OtPIUwu5hKz0H6H0zg+zjuVhfSHkRilXvursO49wcg1tnN+PR+o99LmjrBdxIGt
8pI2WXcv/DAUQmQKwXfKPI9qQMW9KITCmbfT/f6Sfptzgfno+9WRSGZS99VPHDwTHnPMNiKEhfYM
0Weg+kFZFJR7oZOCdi7M3dvyBi2Mzm0W/q0YUXiZ0gqAK9jseyOx3nqVmCa+LvKCp0x/ar3T99rk
utQ3mZtIQ5DgGx14J1EwQiRixU9rma5x654/0Ba6++xinVJTTn/r/59y0JSz3Ift1MjYAu1iZJFq
Oc9cRs1QTNaTZVs363yRkex5aee+/qby7si4v1JeAfW9/sFlAGlCXyT/5uyGZMkujOtuASRV0967
4DXFT85xQfvorC5vRGfnem/XAyRTWh/2kRkdOWYAZiV1YIx7QRzKO6NGFKkhSKATTXWQwBNt8mKI
dgH7tmd/7RXX1dp3o75Bxga01RSf0+WoXLpBF1aJleIpd6nZXVFDxclfUe9gUPZISKIAs3/HMyv5
T5SEafTcXxxXeDjyx2OZPCxdJ0cq4/Hk95kJrDAKJUU20BGPvVSKOW/Ot2iFPTXA54Py6egUmDTU
dOu3WAK3mQvliR2WGvEuHButDiOZpKWuOFbqcHh1+23RI2zG5gC1FizeEgFEYscUouNt8STZjehk
v1p+8/r6M/dbFxSHVo3dFGPBmq5SdTFAJoZFnJWsQnPpe0ELksGKqRo9D1zyV4240ikWJ+cu3tM4
KQxKo+J1DJC6OqKUGoLPWhB5VvpL+HuGTaq6Pt81/xmpvChMDxe3gUHGK7DnUIzQVGgl5L5q5NA5
Rc6zayGcp0STI4pUURwQrz/itVh3Xo7i1qFES40jXuI6+CHPgQvba2uUwEbCOL25MLfEj+rwWVZR
veuAd6WdXiyxAp2UCKb71VNDaRGwa+uZsbL9Z4QKIWNETSMfE3xi5Wc5ZXT/PGZKHdz76WoS6yVV
3UduIEmVVorYWSdsMOOUDMcB+mjRUMz3P0P/A609OUJ4egGMcA/wVyBqDT3ZB+KP/hA12WcRt6vq
c7xR+J+2RapiZ/ZSD0KDvYXBxosmZ+NMIRdXy098qD9OcaKH71IAFVgyapUJm0ZyNvSmoCPTkkQo
tcSJFX8M/eN1kK4wV2XWLEFM0syNGbXqyIy7kjBgS3aHwu9ivTlcFXDtbcsgxvOw7s889teC7TJv
idRvmSLdOo7FTVqYJgFMo7T+JqrWX1KdZXuyxx9lgD/tgaALTJPa3FJ8wxwm8W831vuSOV9Guld7
LcqEIec7ZhHIkVSCokeRqpba06McwmEH0tJRB4NYDTp9/sqc/fOPJ8smEdUSNJLZFkrY0mOImncc
9iUdogzScNClrEbnsPnn7GdbCdcsPaOt0MCcL3chlCHqDoFVE8kQ3UJMvQ9k1S0o4bnCGyeCkDdm
mgU5RtnwYYRBRK59/5nyvoovmG/T1M8YmP+KUWaS4pVQG6ntig8PRpHmWtLV+GvOMVWQEJxdQNAz
NwO7sbxYeI61kihgvRqNYDP8TX59/oJT7A+OYgoc5W0LJGuHZqUJiiNpgdUJ1PGSqaOGZUJEQK/b
bYQtmsfRa34AWtjihxEukm/Nu+OICO96x64WOp4OptNiudNri1pivc/R6O9gwkXKr9A6bHNu8XV7
5A7w+RxyOvMS8WOxpZpBIAiFlumn84htDTAknST2pkGY6PYyJP7ATcit6PHQiAl24nBJv+JDpXuo
8/jfSTC16lunseI+Jbicmg+k2J63NOaTeK0sjdPOsdRlP/mYl7N2sUnMhq1lswbRnBI9uNXAGbbp
/NAxSRqVPTd2g/+STA8awCcJB8olW/97e+FJdEfPuxBUI9EoumHVVG8R6nxJhF+N4VNO9RVEPXwo
B3jR+PImz1A0KN4t/B0s3ANnaksJ5BDFtoRa6ykqz+yzzIHzw0DhfRWqZMZvshVql0OwOIa5Qphf
ylO6/PnYPuj5hBUlzg5G7w2gMWzB9oePg0MY/j04GVGmLTpGpadbYr7IFSo1o6PsgNRnEta/H1sr
KctnC9sh3gpwnqVVjYn0Vo5OiJGmsdmzyzFeinQj/wuNcEsx+IDPD8VtRd5uG73p33tZTQGABeXF
HOZ2vrVUBYRMs8rYIcCqt6+4IqSJsFmZLY8VCoTVvy98YJZH5tMjEju1tVgNV5QNI0mYTm0iIDxB
3ES7JAgP/QW5B3R76oOs61eYC067v2t5uXYRksIBI3KeediCS4R+ALerOZrTz7d5nn24wxDriiVI
lfSUhQ6/SeUNLLGcHcNN5cPAUeiMiFiIHbL9uPyPxTGRPybL8+t8O9VLq+2ZvoIh3uGmI9lW54I0
yw7gUhJ9/J+GRpN5ON+gVJRIYlXGJ4/Opzi7FnAa1mIU1ocQwTrVtSAxlUVIGGO7lvlX3SKisbXt
3nacuSDw3nKn1Oqxrn0bM04PUQkZhaJjPNocEu0X9NCtburtAezhCbgDHXnh1OGDCnLKGEUqtWJw
K0NuVePA+YBJsZH2+qbcWCIrtC+Lqk7AGjz3zDtXDc/anqGBIsTI7DgR+Tc+p4kK5Wf8ETcGD5wZ
VytLZy9ABhkhX2sQtmWnv0a0yQ9pL9qBXO1IXREVnt+GK7VTsfgDVht8NZjiu6Ippk995eSRqc1b
cS/vkZxrbGTVe3LRZZokmR2N9ixZflboh/v2DJvJACX8/WvvwjsAB8WnHqhBhpZYhiOYWiN7GhpR
HOjqecyroTftzRsJNnn4fF2dx9Qpjv+8mDFvZJgdv4lmsKNAhCKxzAHQlLT12Ac1p5pIlGIYu1+g
qD7VCYWtSkTRrOxHBqGRaik8yvjCL6S6vxD3iSmLucz4qNaX3OEgWWG5tNCltMhcEVWnF8gxeFpK
2CwGMLWJmTgAgFnI1VPM1rmHx4D/0OIMax7xYDBW6OAGzeir1615sbLJMh1XLgCcEZ9OSjbgLDyG
3z17BNUo8qnBKc+7361IhXQKeCt+7076ORVeNYo/g6YGbJ86LZ2JRw/c+G3XcjI+jVHWKgbqR2ji
QkkaB8vgivC4R02AhgShumdcwC3oqz8E3P9/DfpddpA6S4vLbd7idRENanb16EQ8n7WCKSImqvFJ
eBVT1xDaIQa7e1AKEUzAPUUGWsAvaamz3L9XCefrarQdxnAJR7II28u+GaBkBCf1q8uBU8V/nwqy
lu8UQ09HjLczNGB2WQ/qAdTa608wx6WBebIix8+0/OEWcmm3SmeU+GsQ+qiJ2Sk6dIZBVA5xkZhV
ZqTIN/aJRaAzjy7DGlqZ3pqQU3+cvlH5TxgbHEW4EAIKh01s1097nMZeUyBDB9lTZOW8yCWf5DxE
mxvVKMe3PsT5UXcMmKc8Q/h1pa/pV3T5FF0sF3i8tf4Gvs/KkFyp5Lmjb3gHugO9K81LZ7oXto8Q
1ek3DS6cFPgUtn8jfBurbK+0O5UDzFQa081e6UzNbhEMV/ExsydLLcmHRAoE//30qc69qcW65oRC
TMQHL90ei08+XwKEjiUUd8RYyZxGt7afgs9e+rEpmoYQmn1GOAjoSe/FQ2op3eNJn1kTKBlLU/em
IuIzuysCUacloPxEaJGVJGGI15zAwIUMzMYVF1AazowYVPJMeYC0vl/yuh/lswPcngl9KA6uiNqV
fPg+MFh0mDuIc9I9guVaJ+F26ZGG9M+HHWPjL/ffFMASxl4IvToqrYaKLvqixW04cXafLdYYi17K
el1qbyuAwCm4wfSoRHLsiZpOKMEcIIkk6FmC/8ukFOmGY5KYPD8uC0btF76AfjTI5M19tk60LDt+
bdaMulXJvWOhVHssmo2ukLxGHwI6FUIyjj1ZeFE5ivD7fmzBFcxKWANMYV4V8839RaQaWowwSnaD
886WOkzWsjv404vfMT8auB6A9iRFDqTfGf9TpRVwgk/jfxvpH/K7OgNXRyy2SqzndRfagbuARHdF
jIk6kmL4FX+vW5FU3yRPLR+OSbeN0C1u1p9qPddcSAxgn3gVr2n7KiJvdZrhvbXRTrwuygMRJKbd
8cA5bCQY5f7H0p18FidP/z8mxEKNnf/vzdaGEJFJkefHOy7zf91lZiXre/14Gww6yOIDPRoxgsg6
1nuwAjsVq+SutpOlbDVdmO5CjS1NvN3uoFF2N8zCj9CKqECz940Zv91yYuPPDtaKJZD2ebzaW4Gt
CDBQ3v9Zw0+/EmFQOL6K4R+abVL4MKoxlJASG+WM+F8c5eY+fJkNWcyWozwpeDfS4rmV3XOWQhZ9
t2KbxDhZVfQpRdnNvyeCrLNGRBN5X6G586UIpOSqQrqtnF36zaq66fZD8KU6PQJOsYFFHum2hCUw
LUEklQAExi4nXmMm8dkwsFdAXOOqxUdySmK5BlDJ5R85TQDGxyJreOM0SsbPIy8N60zTCtptSsih
ReTA9itVmbzXorRF1o8zGFdIL+VXstcXPsPDtMEPCEijLP2afYfJm/HnlqitxfNlt+iCegwu5Uw2
fuSohEJ1x4G+8jnNXbVHBu540z1euofjzUzxduD2muGHrH8JUTxbzPyIcQkC5+eCC2vwR2pS2alF
ZPXq20qfzaC+ijcJNzjKwjy7MR0FCkCblWE/iF4+it1qY3TMQQeWxxAmxtPfWAsNZSehaN43vwIe
7ctGBT5/zD8Kfi/7+8kvZcAOP1+xnEycwR+Ub/k8YxfSwf9iVD9EipEvy67mllRuWARWajhe4rKN
/VFSzawm0aT9TYPzxK2dw9vcV8X3J6Ocad/+wsiqX/g6+vJW6phJA8vqxDJXMB3FHdVpCBpWGP5p
f+5aw0X4SCA+YpO/uE+2sg8IyS7GodRj0EZHCBeVLgYtkCzf+Fkabb1tb+ciwu3H6K7vW7a/RXp5
EfV16MiIWpci4MSgYT58Ws7XNd552I9zE8+i+xEPw9v1+y7JGtBEk275Q50YZwalEBnmRG5Q/P3h
ociG8tXiex6A7/sy+yvtZwT89vvSOdCtK1ognqR0GrLw1MOOmpPi3W4dtGIolqxizuApxJwYS+id
2DJRw+NVbj4myh3hN/typO8jvJ5btOGkiwcg0WQ+iIk3X5wxdh947pX4PsaTNq/iL1BhdmKhyduU
7fI1mkE7C3PxI8MZyQSQL88OwgnIVYOPTlWkXEZrTMP2X7e8YALklY1aivJ2PPaVYs3agC+AXpSS
t6wUyYgU9mtrAY/DHfs1xE3ehfCfoZWNhrzYmQlzqWmVp0Dq6ins4dQ2rjrLFRdkqhY7AhvPWKPa
I5vUupG2WpAy6nI/j0Q6i3seFKIEjPA58tiulZCqhpIFpA5rM/N3jp2n0oXJApOdSHGwX9P4uQ9M
+O8p0i91BYSi6eVHKyU3qwWK3Ui5VaEnhLhPvaJE3B2QxJ9Jfgqo+g7M4NYaywCGz358rANLiqDr
e5TUTWl0Gp1mAQkyv3V0jtctdOi+mi3R0xQ5b7mIK60yLVHewJgMfVC9MJcYj92gvsWBKNiqGfD1
dEKr63Uh0v6VN0CNfbbIbmbpPvzcgvV5k1mGCx0DRIatm2ETWdDfgyJ2VNYnpZRP5es3moyjE0HI
GSG3TriS1b1xZLQ4rJmKN1L2uW9gZG3p3tA39hxOyWTpvuj6EPzGfk0yR7zARGUqnI1KBYIchhki
K+UtvOm6VMXtkSpg3DKDKMXHhRCABfKqNL0evk9epRrE9mUebSaOwaF4sK07VUc4eSi63JnM66Gu
T6KCBB+k4MvAmE7ER5avCqgsVXmPKeWi6jhqevNqimSI95BFPAzIzE2Du/fJAD08PcyCEUW04LKz
5fV2uJB78eyAMYCAjen2F0qHQXeyFMyzs0+QZxaOtk4Xy3R/5lvC0wucmksV9UsFBFeBDt6OlpYz
lNEoN/NozfdScyEkwO8V7zQnl536JE87epdN+sIlhag+BXZtCGicVl87zFFtgiaPxAOeeU+Fy0OQ
Usdv0ttbNyEhj3f+TFgATl4i+9k8sXSYBsP4ab2BwUk4dRiIAUFJTh0327xD4H7Oe00v9PXk5M7o
RlcVJorVvRt4J5a39XNlC2lYK+pUP2BuH5pDji4gTidi/UL9fM5h2t3RFKQZEbl69rDpJEC9Aagx
HcmGTAJsLaKEVoQPiq7v5ecyC0iNcSV4FSVfYyjMy+690b9HMmXStcw51vrilSVR5HY3Tk0a8O4j
dqSwbGufEQr9sl3ktpnFWR2azwke9pLZekM2g4KGb/B1cAPSmPy58Vt1wNS0GEkfiEccAm3qlQKx
ryzqvc1A+FR2Z+QDfY+Wt+4gg38tTjFxZMSOEmpnN4LySXr/AbStCkPGItfR3amkxc0cdj3uZA/1
HaHvSXbmF253mObp65XZkr1J/6ht5qZlWw0qWbrVKMOysnWgu9NZMyN44V+9SlwJRIKggAi1RBxu
/M7ETc9sowLZ3C9+4CUivIf0rvQJ7+p6RiZPEpvgkEUm4v2LcffYYN/Bt9SJ0QvjTTY57bEk5Ffh
GW8VfxVVBGvvHUg8eOjt2ulNM5Gql30IJj40aPQs+/TnslYoX6Amuqwrn8j3VGDe0PHMur+5nVGj
fMco4gZd+hpNDL//CFepSyfMtpUTGllqsZGp6RxmzXUs2udGjgshNEd08k2u7xy1jfPx/eAha2g5
/muaCr9k8V8YwYfA9N2COKvRUNddCuzigP2EGusz13KcEQMDHlUUW8urA0Ca9/2OQXMxlTAUM+Re
qNtsr08FvVsyhoqoyqoWIyEtPNd6GiMyDzp+tPK7qDN/lSxG6eEW9TXcyCt1V3EzIQScD+mrEvMq
+4zVykjd8cKp4H1yqWRztAZvhklEXJw1mUQgNRswM1BILMMj5l25r295uwPcvKnr3ocJrKqbt7zh
0RrJozvSs8bkznvr/pr/3PML5uVXCHSGcdFpBiSU3X1S6TkcZ+jzbxhUSiIYOXTSp3aLJISSVb8t
OWPLMZeo8sUBNjWE3EXrXWMoZ48xQmGfXWsII1MfNcKsYMMUrix1EDK7PvU9LfAhflP7EvxQNBnb
TkQrgTAPsV77j9SiDxrxIReghhrx5oMEOWlRYgA/WhURV7J+ivZjw1wokqgAjoUtcLYFKm9sELfB
+qKG78yiDMxWw4U1zIkTYANvKJwBYCee79DIQVhzjCCpUm5clqoQbw2PfWvliDyGbRFT2zVknnHG
MdVnsAVpxcQMKSi4UkthfQkZDqxnTpHYO9VjfNhHBEMuEv3NyHYL2OmWrXq4Kn+oKlPfEC/daum5
LkvFAqgycdxAY2TqtLbS9cv7bFmZuti/BqfOJg9Rj2v8QwTn7ymaApvjuf/UFfZ+0XJibt8RIIq8
H/0x8SFjMPmMNSIAOevEU5PLz96szfW2uuOOHQpbCzHWOm0CrC1XRKO6OfwXYoHBMLCciMUUsWg5
kJneXnIRo+MQCof8T3e2WZOsOcWWhiETCrCPIecgYsKhOsmUaUDbfu/1AxxalTMY+K/NVPBFWR/9
xGPfd1Mdkzty2EDGFasPORPLAOSv+cCtCWtZIpcMwLylN8zsIzoi5G01BdnCc0HXHnEKsqjTXCyS
7sQ1JacxkNz3LEroQanOXWAaAKOSDms2W848qTHQhKJYHHiD/rNINaPQ7lmXWuS0hrwR0al+t1XY
jKAgv6Pa3y2AsTd1sR0kJDAGQHMlm3h8n0jY2oj0bwV2GbSfdSvL8pZgS7TERf/5sH3kI9fBz553
WIzRniuhx/PlOqnJqsCoviNVUlQpfjk2MRk0ukSuuGv7kd8J8gxKAAdBm+DkqOdR62FATGk3MYnq
WuuyoGJgMk/37uffGl8giEnSSIZijTFDYzX65aqZI8N9TJC9Lej1gay0W+PRz4u8YrXgf9vqNef+
EThUx0emA1oU/wDlBxpM/Mf1DZ7l1nM0KCZQyOGYhpfqLuKN6xTtibB0yYYHogVJ9/5ej7+Ii52R
vhdZDNlp9BF9/RIO9z/4+sFo/q70cDCcyCbzBIJbLK0k8JeHGb0qU3Ka5tEEr2qJ3acmT36P4Wra
XdLkvDVAVG+7l266XATMZKMXJFmTya+JXvPAcqQ1n+IHhrlhbPxL/CRldEHIAVn2Wdj+1xpyOs5J
PjEOL8578vcavVp8gJ0EvFPwjiDv9v1xp4VLqeiKdFvW18DU16WPF0ktSSR/O0iiYZvgptwlymaz
c5gjDScAVvNwbYL+5hrtR3mbwld9yr6kVrNoBWEkDsjr4VjMc+ymnEH/mglqPYeUFASWhod7i7gl
sZrOMMl83+eN2ZnvRyU68W+69QDBZdDdSXMk3/CXiT0dyy6Xi3odrBU0JJRRsC2tkKO/CJNLSDrs
8kxg31uQOYcyC5yV50bbdkLSpnggLwGXRoNMZ9AXaZmktAHMifsvmwwntKUj52T5/EueAiZfli1n
y+KSBhaOuH5jWvvcYAcw0rdl3cljgiaM2UQ59wcKLyuwQDT6kuZsCmzM2iZQuXellhVRB8riSH58
+QsJTb8vJSZzdz2NyAJ8JkTfapgdIRzvscANN2q8lVxn4ZKXPhZccwoGtGDWBV9fsoiB9nnXjJ2Z
hr/tWV7TlXNNQaquElpYBVPp1ZqBFr2QC/KQKneuRP9j0lpeNTHosmDsqOLD5WQkAmJauyGuU6EW
4Gaukecq10nYZxJ6QlhC2THJpK20pIpwgyGTAoE7T8WeOXRMziyEEEreNKIQbhE/J53ITHxR4Np2
wPLSYvt3qpoHhBNeppId7SMMH3yaLjxCS+KyWq6d6MLH1i7LtcnpiktfS1KIpABysuXNG/JIHgsS
B1zg5xN6paC8Gk/HKll1Raf/KKnONaZgWE3+MJQwRAKgzhu/1X4xyVQdfzR16tX0/ZikDsuS1P7D
DoMlvDS8UOAmuqaC0lKbeIDff+7krDir2LK7K6MMAie10QB/L0ek7KQRZfgN84F85IIJlxDpyk3C
RDChOlI37Z0W9VF8NrSVVL/Kwk2zJjXH+Jgc3yAS+9myb4hiVY1eHuHy7c/vZukODfmqwaTcLsF2
R0py3iMD9Vrj7ZWyc8jTaNhr2nA6EcLFeRWrsyo8ruchx2zkjNcJnQzeORDKOot+SH9UlvZywBWg
qSLsGByZitoHNP5CSwAFGO3nL08reSoIRM+Pe5X/yUFxt1w7ckVCqXzggT5kWG8pshL9DgwR5VF1
90CQyEPUw9tCP5wtqLVEBFWRKXHqb1+xsYXKw+UqyFYWNhfpd7AyKjhXUh0doSHZKfIN2fLJzZxw
hiuP04Sfw1JL+MTQ3rWNWahyJUUwYg2BcIPthWo18q9sGYzViQtAgbP8QvNa4s3D5GCrAPci6j0I
e2Xqz1cTOrFACghqldrVAN8iHJg1nO3JEhasm0O7hXuhKPB4BE7jcvBF/g8xKJxWPgS75AuLOGBP
pgPnrQfCPdko2LmYHxsdJojx/uv3HEobkhCgeiWEmd1OatjoGLQcVo+MhMe7DmDCn23KJlsXynHB
vz46wxoi6jxXdK231Wkb+rRIArW5OblpW20YoR38vR3zK73d8k55YF7kcAV6JlXNQYD4oVHVSONb
1LDBXNZsNePcmz0UXDVC7pphwAHa4a4/jpybv8PboevjpsAKmpo4wB58Niee7A9+vN7UHHbx8lcP
A5omIOhFjBOYb4OUjWM/tGbPC1HVa6oWk5Jfqb+HEiYa0GRhyaVst7tlFNfODWG3bUDov8bqxPTR
vMX2MQxcF4g/2qYJMUx9le6TKe1m40C9CFN0yRL092sxKKUVdFQvn8wg+vgtJAFOXKxsJmBtR1vY
ZCX7ZVv1XSPlJ99nYFcDJpB1kNCZmrbgd6t65hMmQybXRMvilPNyDvrapENerpa+qqTCi8yuvzKI
GULvrnd9bL5ZFNpfjfoRCoxwUhd+oq+wXYB/UE27ptgv62gzRxnNVtlk31Cj6ZUZQXx5f+3tjk9M
um0STFgPcidxm+jbMqjDDIi8xrKXCuZrw/5rOgLWxu8AdZurZhzoe/gL2FbW+8pYHonzWjLf8b/9
QlXMyQN30kOQRfzl7BDqnYLE0DLe8e+TZuO4z9ohCDE+3Fii51/Wt0mh0eUp/Cz26OfHNMjb78pc
McEEhnv5ePPDM+nhbTBHzvLXK4KAsoFRU9usaG3cWZr/qqnw16jSKIzWFO2czeUcs/yWoVvtceGQ
bb4gS8r+vnNq5T2zLKBqlcsOwnjjRBpjoi/cYNKQuYaPLHi7y8bTk/tSInkniKbM2/Y4YgbuKJCV
XzfFcYRYxBnBlFP6Fv/rV4vhmaJ/YvEhcEtqwvlpqBDJg0GqRKTdKrs0vJO94T21hHZrfy97xJfK
aq9XiGGI1qUuGOQnST19CEZNcJ0/BYpzhdoZ11FsagtK+VbRCtmXq96zhm/f+G/TIfda+A/YWgdR
8UK2zeM6Iiz/GPbgdtMgq8PYDJjVgPbMg5IMZzw9eU5Hi8FsC2lv0WlarfuUI5Ho41faR/tNCnCK
B/GW0nxCELb0O5IYlDQUjVbCfHPXZOGa4aU0N/R44o3NNXIcj+dz2ANlHNUXfsf7H//dzrqhhLCO
lz9CspNcKAz9AWjc2hTrchEZj6tCRaP0uYXaoYfkvsk8tXcg/JFc7JVsNc2ssJOQjpIjk8zH9aL9
He4ODgK+RqK9H2caMueWjII348sfqwjxBYbMhTj/N/4SuVL9Jn8v8D+w9MnFwJFaX9JZbPpk/aOE
+TwWwnjKeRyjmvqvwNgaIByEi2Ea+DyUE503VFdMHr8YjPyWdMtKW6JKlLiFRSM7oB3xQTZ1cUOe
Prjfifnnzcc91cXzefS7Li7HWNcHtoIkbxfzbHel5ZwU2PaRFHl++zhdBYvvYa+83uMeM0+1L9Ly
PbbeULajj0MSbnbHamzCxv9Cv7TgHDXJIvJupNQ63yFkcRax96o7GT0mYU7nUcuFqz5F5W+beQ22
eb7d0dDNGRRaR4fiV90xa0U54Q/cZw0+6Kq+ZQXZbda1dUj5jwyUcILWMrWtivGYhLIwHrN+8O0X
2aytQUCr5CIAtOQRP6aSf9sjja+7hCwIUPfVXh8F7vGuNpBDd+5Q8xOi66KO4MQyXmxNlOBYALpr
gSv/VQqv05ORQEJCGgfwaHozN4oUO8NNpva+8elXUrShrcXJhOYyFVzu2JSISK347WWvGS0qNP0r
YwXN6CDvjX5IyW9Ec0Mtg4S24YFPh5JmQvNYnBfd3FwzgcQzqk9mvmeecN3sifAqzK6V2aQfcPWG
JvdIgg6AMXFip4q5KAdKlnvE/HwcRtksyyzDvDiYMLGMEakJCKyBera8SVKsEv6oHQg9QKF59Ujw
t7bT9MfpH8wQ5QoCpRId8BVMAdDhH2v+7eHvKZWhpxow0Z9hW25r7K561NZNtFIy9TGanPCBqSZc
3A2BYM5D11tZ1X05ddkynmQK8rIoO8KJjkuGQtG19+3eXcUih7IwMVWT+ARp8SM7Qng6INTYr9q1
lf9bGUoQ5SOVrI96+wrBi6arMQ5ZlFYULgYgVpCGIv4oMdFnmQDX9DaSDiYGa5yK2bM/m3pvz3b5
OOktT+ZvG6NutFrhdPkSAxfAVVgibTE8F09G+LoDYMXfrUtyHazhL9zvFZ0bMtCCjqqm+wNPWRfp
LYwmj2J6SKjo+dhjJ2NH2v8MPh3ru4s5F0FWWR+eDCixsOO6PV60O4NckSKFjZ+fbLC5p+xrZQLm
vCEstNrGwieOdSkQsjIlF9wPRICwbRUbhRdbymjtOSFZotQ3Rj9VUaMZKmskp+Fpp6PooZGhmqIf
0H+HGc86JW/EXXULxvks5ori/ISO6aKEO6tHBjV8qQW10Inf5AQPIX81BvirvGEWryal2tPQGrkH
fOI+cEPWxIkKy2ys5Vq6snXNNZ17sbMD7AYfTrOpJT8BFjJq7GuvtT7H8g3UGuf4zBCfu0y4+WWg
DZfzB9fxmG0hdClZ62ibKZkYKl7vaRe9wByIPVqmgRMBI0vjpbMt7WoUlBHX3WzvcHYa1zl3efSK
VCTi4Nlf/dMJcWPgqC41R6LuTey0KiSWn94d921UgYQROTIvrYxbMwB2Js1u8omE3vDaX9x1pNde
7Mpb/JsxNq0MMOgydgKy60X6/Fc0CPUT0QDLxwGEW283MjuqVshc5gKzIdc9vXp1EjhjJFt3Gpt6
trxf1eK170IrcSmrfxWarHbzI79XbAsLja2PYWIPp+6jTWuBTHBFP4EYtlf+9vPYhdftjuvM0KuE
BCCbK58WnkvWxrFYmCMerb/r/uMaOzkbv768T3t1/maiDXsbDksOweWVSXIfELATChHQ00Aj/lt8
TTgNsiixmbBdLgHs5TwUJzb+dPkW/CpD4JcDEJxNBPvQSB1ZLlGvs6kf5Nov4i0gkQPTNsdd0avC
f2RY6sHSq4iVwW4RdC4bFvti4XP3tWo+xMtWROvKLoIt5nIZ4oAhNEinT0vgYeTLvZ3ZCc3Gexlt
zmG9ohLPvzROpDabN1dEceQUY0XJdxcCBrVDaAgYDOVyZFtj0P1GM6l1VqKKasG6xbLHSPTYMxXg
uN33dlnZ22uLeB+NC/OTejTz/rdHSBSTdMi/4VCxvefj6bd6KsMgat1cRKG9Vt5HFbYVL61c0FKj
oirq5KL5KQ/OhNJsX6j9jBO7AdRVwmBI/r1gLmkLiWY9z3z5P+y9h//va8EzQj7BuxHhzSkJAU2v
eCmvSwgqUT79ta/eYRUKbDoqAzZZz9ogPVJcbMjvK+4AsOc4A6oJH0O4BgonUDf3GcixOW/RYB8Z
JGkDQleuNcA2pj4nNeJdT0UfzW3/bZeHQdCEAc0hOee2i/vEGXkUTSvuYJxBWK+Em9nGDZHuDHYR
DJa+cKf0NoiYhOvhOpme+tbNPk5D8wcnmwKWSDCQ+36byZh1sYPs9naKTa6RPUECThVBQYBIXT6D
cEKFx7ldbVjR8tXYPks3eT3VyT7Z5XP4BwNDKa7I72+lFudMO7kw7pazLwbdoRAplZU8oqNWmsOo
3SP4L59K33SsR/qkjMa8dz6W96u8nR0eLuh70VJ3OtshcX8Zf+rzvk961AJtfoMdVmEyr818Q33v
JR7iT/KYWNj+9KbMN0R7CxheImw5x+cIO76R+246+oChUM8tp8yQpEAYGOTYc+mvN1QMcikjkKN0
D006/MGbDIkVy1F9b90u3C3jesr2K4bBXxkahu3iRTYG/t1RnmdlPOkJ7ACX/sxZpdprggid9iFZ
4kivdMR354zxWSp2aS0GZQD8nKY0Ze/FMjNicuMSxlGMkYC6puPpnnOyeaXab6Go3BwhI8eyWlFH
i+JYo5Od+53Bo0e8aDl409QSZjD17c8w61BCPae4cWlokySgIIATCZRBNqWLVqPz8TfWzzr5dbWb
Zq1KAWX5IYSVTDBa7yKIBRGEIR/6nl5270snV0YIxag9P3Zzwf8oYLx/1Z8i1UJPLKiDYTNL7/Dv
pqQGuLUgCCN6qwNo4CIy8TllBaTEdp18szngJ3vRVLCljchbKtJr5HntXAIS15Jc1aQAVr9DANhh
yd2UAEIev7LhfxwZOD0t/7Q9zCKj/VIdrsUDy/ju+TCquSsp+hfLuCIQqi2ScwUgByQt7/okUXuD
gkrOAEpyC/8lJ7nqmhkZ/Ylx5TfBZti4y+yZwAkFQ4cXYwGDGfwl0TiiUNxFjUl3yuL1fU+2CGND
E7tEoNchy+SiqcXC7UuFuKc4DR/DKHfF23ZOFnIhZ81NSPqvPiWtyqqgNmRFyBiy7ZxtcYasSjrM
A57HKhDL0qP8LHxl/RxipRjqD+/OLg8AimGncRq1OvIFe8HA+G2d6Tp4SZLMdeS5lNyEr0rQ08Bp
LKYkLOb5/Nk/8Tx2BP8CC8u3ktAGQO3DfHWHIPS3vtCeHBXQ0eQ+Ew7NWYBBLcVEAbDXBlsvac9b
NOdG5Dd7h5vUiBGqHVN7H3dQM5KHj7w34Kv2gSgOxdAD4uFOQD2G/XZWF6qiZBMDrYaYt2SVgHCP
IC4TVCtF7B4EibeC3SuIYoiF7VRxycx4YWk4dwx+2fLJ0jw/OfCt3VdJoCMiHicFlXkLUxgjsp8H
z/o2VREVAeEblbuoui6da75pyxoISSDOJn3UJWKpTGWkgzcvPIFVDVzr4L6BLL5pDs0xVuvdBu4S
k7V1XgTNSIx4DlWfjXzgFSQEcbaR1/gBjI7BhDBHQ6VGPuGRE6GNqwkXi6La7tnUVKzUyUWs/LpZ
781EU9UnOYGiuhLw/Kxo9Iy4zMKM/5CIL2YqFki3KwsHtVBYAy7qfHJTaKcvVt4M7zDbpcnlSZPw
9d/BvPhhai2lgAP1PVCwSuG4IbrGvxFNuvKZTF0ZMTElS/EKWoP2GoU6Yx9Z5CZQs3AWT1pqWLGx
cNIp4mfFjKBVKuvWvT2yi0pZ3XBSvTYTk20vJuRBlgKg2rNkc7Bxx6liupVDRZ2WViaUp9lrO0ll
YqQtE3WLUvSKJB+SCPnhkPbOeNwElLzWZ3ufAnmdDCL8hWo7YldFL9mS1CQhf2KAXT7D9gNRC9XA
cLYuXkzSwqYBA6e62ASaoG2IJYQoRfQkFQpd0QcDKLlbNsrkwv1Je4+nfx7aZMspI/PLVQtAOHKP
iDeZaAqR4EuoC36vTtmcICRDAU9hXqO49GukQLh+Gu9pAt8PCyLnhsvOThnzgsC04MALyafYGs0X
KGdya58ZaoEuZFwDYfuqvYTEX4wFVv2R8Z2PEOM0HLZP0QfMWzAjc4AbBcdU7sVAF0a0YprxccgV
LtDh49KYY7MLXvJn/Vx0ioOUOq5wvm4lF6vc+l/CET1OoyoxOYnsh7FMpDg3lm0AkSdUiMnL0rv+
SrUreO7OsAlZAnJvGA77Irc4ALKMBZWE1PeePS6gc17zsJstsZEocc/od/GruzzvnnzXmNqyNKod
nc6Ml95WwerYKuo7IrYQYFNaW5iEux5Tg2pVJAMqwWYeTd+hX7OyreN6GNVGfaN6p6Ib78k7jha/
UvvXTuyrXYq4vaSYjyjw6Hww5v4qCWKfeLL85fz/ySKeq3AQx69yKiB+m/8UI1/GZuVb6XlJjAZd
eMkY0dvSDVASAXCCryiEMESTOAJMUMy42Cpiqod4Vb3hmvRFoTlTpruQqlwhRH2H8l/dJ83UxmC1
LXUL/4HeTpmTw5WDDe3acxtiSRdprVh6CD+urr31zJzuq8yyb5+h6epCNNs5C929YoR9dvuHXRrH
qi+gL3g1vhnXjH/Stk4vqB46bGWV4ux71/DS2imF6om8sO7GoUD+jXYEVPqIp/Qqx+2FZ3mIhgDx
rOvN9Ss4kcY/T9heCRhe8bIOvtb+c/vhjN9SjBt0xIyrZh6cAhule2XPYxBgcYw+uA9VSmHucbiN
MaYWHS2gu4tcvNF0ulSJQxteKOHzJMgm+PWbO1sBeo+byC6gyKmzeZFzHlGmzrJSd18SL6yAbDvk
wnfB3M8sop2yJa7LE5MCnXBYK3nejPLKFUWOpj34eQwxZBISwBYmoR3ox/RBMSD3rhfF+WjorSP5
DuV1nibFWvS++AN7C0sISK3U+6bg7dFHuBqe/HoFPy9X4t3GqK9kaaPrLWJRWkjDSiMSJEeQB5P9
MTf1P0uTfti/yN0vLImt77e8qZTK+G8myfZWL4EhIejeXw6g+iCDjYYDDV1dqlhFnnDrvD1jEwb2
9GdS6I4ZCBYQbomvTIRWe+evGfnfr1vm+r72gmrkdPKJYoaMyrhqcyn+hzImRPsVKwIoEwnIMf6i
UcC61qIlicdHP+eil7Yy77OKIRPcKjbXbEoMQo+wIvQSNv8loZ5Xe0KiZZMADrd7TkyliTuXP4bG
JPCfA9YsmhPK28dj/SX+8dW/FDLba9+uBaIN3Rhu6H1ZbWq3Twao162idrd2v9xWcu63aYzmgIC7
zTWtvPzCzdDHDRLZE78/4oi0t4EgBGvkpHdoIRswln9bBdzYvE0Futy+MEZBsNxpE/uvR2QFZ2tW
A223GMwgUWOv2Gof+MAS4uCcMbEUTANG5J3NVHlBmXPYPjrsRl1p+wbwcL/rFKzckA7WEOJDBs52
FwGIPxN6dwbM4iNRHibn4jpvCb0BLCGGu5CrcpHca2fjtSMlkx49tj7PmPgfodq7UTZ4HysV2VZK
E7bRsrSB9i8BFhXZGfB8420H8OWDZ+tZ8VN3PQtfBA4WXjDUnEEUJ/vlL2M2p7rUNAhclqPCHPzg
qcXP0XMcMPSVE2tClI2XWlABCE5lq0IRJygqKan1jeZHrieb1QSOzkyTI0HpFXvAuRIj2edtnA/t
Gqr3BOpwDaom4WBC+yF+I/XRbdktL/sS45mXlx7p9G5RNSWL8/aK4vlXc82QXUwze7JSHH08ct4r
d26CPcSgNYKREV31nNcyOBXC7IRxIXXax9UkotzkfXJeehHTAzH+SlM7hwFZnsRkXGxw0A5D0jTi
/dprTj6rXbQzAn1KMQ+a/rpZ7KsCGtbVGrLnj5BaUUze0kL8oDezH+DOaqG94uca8FqwfLKnctkq
/IuqdMk2ziVD1qVlnAmQGNVKSD/jR3DGj8qRhLSFL1Yh1oCHUBbN9qy38NdyvXtVhHHxF3h8agnQ
nFa+3D+gMfh9IG1ORYqSc59PEmLKGypM3KStNwnuuMn9pumsQxculQwwf0VRKG/hoYM9cpaXw7CL
1jwTqm1xcfI/gDhzk2pjpKb0vAbsoLjw5Fi62A+8qoqnFGI/WPignGizuFdi6a8uR28II11ggw/r
Es5f4Owd3uFbSvnRWXSQyheDc4uPmkmymUnlrVNnVENHouRHqH0tNKks6kSX1o51z0dG5koaTsPa
olWZIpp0DRVTpQF/7YjMw/n+XrD4x8v3haSaa1piwzZ6zpeaL/yJYuGOy0zBYqKi4qmU9/LjMrnG
ZaBINOPleItZu2iqbycZ0LaYfT/rXON+OHyfF+nSrddqV3Urp3glKTgjnMD3rt1zY5K0O465OzLz
WbbJBZqAviclGMUxdF+/v/HX2PPB1nadaSvBDr4pQ47BZGQLYhO3cNfeOe9lK/rEVzZJiRt1ZHSa
ljFHRTfvaRLYN9nEuNSatOr8k2UHLFupnXVtmmkTnUt8t+fFj37ygWOag/dmMj9cRegsSASlClVZ
RLlc8vtj1TW7CmRYxxs6IcGyP7dA6uWnF7RtQieuPIdHtqXnNcAvp+dp+4mgcQIQovcCMzYTYelh
b3YKhLt8Ty/1VfC4yW0u5VYUvphrhOSDtc8jX9Ml0O0J++w+GbCeW3NjhWL7wwxNHD/5ANihzFCZ
0dwjpv1qsQEU3AzdafxW4towaqpHSAChs08tTaASEyn1BwCUZ1u2wnoAi6pISG89Icmo0AU2xlnc
wtG7FJsdtBpV4Tj5NaurA+o/rVIEBNSNJUfu/Hmc+lQG9oOePTQ7a2mDZ0PpUynmZiXv+qxS1/iZ
QJvbz65f9aVt8y8PCtUmGPhEK4e3o7TX4y7MEJyESWTyl8QoYl5ASz8Z5keU17GBclPLZit2dIpK
03+LiK9wj1pzOz0LASps37tOP+zIXEYtDuX3i7KPwNks5yIY2/c6x6/6M24KCabS3+j5H458I7pX
t18oeGVEADtxq0d68nxDOawcNIzCorB7lEYHCd2YU5+Uf7F8Ij7N4SyYYg/6CizRg/mnNEp5Tfd6
+QIkB8COa/HkZiDR6ZfduxF68FV7aM1jeNM1ScmJR4rK9GSPhhNEMYSeuBKFpxGD1e8j7/EVNt3y
/95lz7/VR5xm55dnKz+pKnF8eHQZuIxKzCjHbU+1FUrvdXMB4OjHInNLfZLoObApD4HFEk38T/pa
nY0jHo5fbWx2OWh+aRrvh2kebtg3/GtXjAzRj3uJ6IUEnLnWjnuINNjzmyS/K1GVDolgqcZYzUrF
l2KFEDq7F/5S09m88B7fjG3o57P/SbLcSF4S6jYJLVakj+v44e8tjiq1ow4ABLotJ5trOl7THVAt
cV1YuUZMI3l7vTlwhVWsrPDytOmGqiMTvHkfo+cr/+gSz2c4r8VN4gNgm9lj8wIigOr4UFmrCQHB
B8C8Lm8cTEaGM/3BKF/WBbabh50gLafrAc6swDpnialcM8kk7CfMOmazK0T42WrRJ0ggifAudnJQ
2ViEdWSOn7tw6bZuEbDUd7B5wFKxJhLi9zYuV456NqffpsTEGU6S/C0fzerNIsygKWyiGNIVyAT+
sXMqu/8aiFBoZvuCJ/vTuwd7RWmLcCk/WP1RTT/pTkEwQvu8v1er38A8ocxkO/UcPJ366YzW85i4
vzZGkII5LV6QQGKNXmL3nbHlnlqzL8DF/cRuMNdFjTnCVHxBkS7bVerzSdFvPoWP+Nvk5ZaQBOER
e+mtA8K1z+0HewoYnJrtLoBHupjVwmDdRr9HjGvQ5RGY4XkZhYC1UmsuQXGyz7DGMkRA/p9L0tBx
3+DKFxxs1A4KJJZrHnw0Ot0ZLFXATYnUu9oX7zP4SBPnIlgh87x5nQ+cBRkkjeOLA+mcA2avAyn6
QqLV8sh3c58Th7sMUmsHwjZ2ziIVCTPw5k2ihgBYbrFzuLs+cSc2BKgJj10dCpsds280eax23Wv6
SIEX+RaQM1BMNJ8iQLIbN6Iwyza5erscWxNWDjb6JvfRV7o+SrBqrlvU9YpX+e0KvveqgQRnu/ot
RnuYOhRFXl5XhQvvBN/qXfp10N3fKemNMFb/fHUbAbR92fn9+cluSC8PRLfxeu3mwjgy4TNucQTJ
UPxHi4XesxVKdiztlUDogve97GghSeRdi4e0yZ8nxVFLBf55a8f6U7BhG4HUVwM/ix4cTkOcDZpz
/2x+XWWZk1KNQjp2DHhXwiTnD95CQvNY4QXyOcBqGQIYpsG9r+dFJB9+xQRSeWlCc9GGXgO4pach
+bcgHS0a1CiBckABdgnSCfE9EWab1hkRRB3u4oycBsMBmDn/oTvJ0WHEbfDfi4YIBoXH8NaaVrTV
evtU9q7yrreS2k+iLzAL9JqXkrLXvelrlxQrOhc7wBILjWxGe3LD7TizAaFoR5W5lLyzvYSWgVMI
LL7T2ut1tCllUY/AJ+knVNOgKC0m8sVkOBY2PvNxoZaPN0q20E9ZuGcQaApnUcFVLm/csC0GPxLO
UxsyY4+KcX35MEh6qMQ8VWx9N6F+i7KSa8q38a5Ykt03zUHKPXtcd8vjg+p6cdhQTA/gqQ6e+cg8
KXoQxSAKfnLYYqNvzJ2QrmSMTDWbutjO6YFrQM7J6u/FpdKGynB3sKTm/ZPks/FoT9/5mCI8Qd7b
IInfv+uTcZ1j1dgsq2Dy+PkIqeWhaivenyuFAzIB54R63PFBc3z4HMMgqH9vPcNNEpIxw4jAwl8n
yL2KVr2UZhOCrNJRyIkcNrAJp7OJ/6Ul1vImUX4Hv+NFazFRUeC2g3crthdHnXpcxyrdzjHIyAEI
czjble1iXOFauty/NGSwcvNgq24EvMyBpVuVbUv5PnZhH7pCMHn38ULystI3/THM37Z61Z2By51J
KxH0Y4W+EWwsAySHQoCRrl6FOEGUCDeeudlBPQ5+1Pe5g8wdPnN9qKQTqSq8KMtICtcLz63JX2I8
7jA+DRXT2V0TTcXZ1hQBEzMlNxF85SjDhPeszscop2J8pEqHlz9iGwXc7ZmrvkKmPnQmb6AYMNXn
eApM/jJfEVI3yLjhG/E81XBWlFxMcPtlNrA2YE8fP+7Njq44+vfvzcb7TSqwU+N8a06PCH/lY6Zy
opozC7KiN99McyoFR85RQJO+DgaExBO3b4rKifEUlBAsYrtoHS/Sq8vderkUAxGB46Uqshg07bKo
9PUY2XjNx4RoZme66gS1dODUe8CsXb7VvtmPc5ad7lw+DFbP1v9jBHnWgVml6vysr8VlpxqpFpGh
GNZBDHv65up2RPfzmTY+iCcL9fveoaFBWTH8rjUJC1300BNuqwtRb+MpUjzPfjUogo6PoHxeEKGX
ajPXOPqTj/SIfyMZlhQybnGo3nLwNDw3sZBCXSmZPsIbxWiJmYRVeyAw+wkfjXisnokQtNhNehWD
csjWExlWvnms9fLk0juLu4N69Y8+lPxyALfHTHGl5DrucvufiqF1JTGYXkRpiSZjLJmTlRJYGnwS
8cSc0RD56TA/cGlzeXp0J8uIL0xHTbnmckiHGbOErenqCeZcwEq3OHNPec66RivV1F6b3LBWDSSk
xjdw2KX7R+oY/NYxmcRfjdUVlOoHbJCaV8o3BZLnN7pptDwDomepjcYHPSIiMnnM9phdtYgaxH6m
C7hgPU4dCqURfkYZpEMvOXdtPzgKPeoPZGKfterKcmKOj2+Co7UzsAIn2tYD2/e8AuZijNv8v3yI
wtXj2KL7K4rR3NdTMPz9gKdxIWOBia733mapdXa+6sbuM5U4mBmZ80IYwUWQNYyWTcWFaP2OGKfT
fzXEeM6JOaLU3DTH9VH5WWgwZnwWUxlKY/gCzeouATu52ExLQCDU077JNG0bxRryPkB+/5HCIiJw
xsK5izKSGH7L2pwntfHvO6Zlh11AM+oZY1RBnjXWdybEemAvF9UthOPlbNs8PDh3bR4T+VF7qQDo
ML54/gIRKnZOgN/U2jqDPeEaM6LDya22klzGx0o9WPgmAPbhJUyzpt+Rcav52pqyJJI/BckuP73h
l1t8441lvlSkZyhtUFG5LWsQjfvqpzpQyS+on0TJMEZGv9c8X6o+2lXaGPBmwSz+ZNTHaWrtLJMX
41uPdDb8ToE7CIgPsYCmg+e65fDdDbtvcrcGOrwX3wAZ7LJ6N25jQceRKEiu7/8LY30OCt1TATxy
76VdWnfM9iuzyzzIFY3MBS72I6YdsFAXa0sP+CuwqXQgQ131caMtaUVZsc2+S55dGUCdi/kiDaqH
xDx9FxNBP1eAP1js8KUrDpDJmXuzlmo8QCjB8tV+BF9l+F9qsFWV8y0vIg2djaTbSOrKJ56e+LKv
OaG7ZnakjCUJSxIGHzLECU2KT3wz9eMhFNmghO0maYXcNi6bA3HoUhgQ4IIDt6lIk8zbgOarQdYz
tred8vWdasDiWT8LMLAO+HLMyOTuivN6azgucVy7KHhqHGQI3HrRbcbtNeW6Lc6xtfMGIfvppVcS
yKyhBCYWyZ+rKidVJx2EeUQwaxZO2vPUJZkSq6tqYk+fAro55ZpwTX+dcD4Xdv6NTz6mke5zFWrk
H8ulooK38Fkcxat2cjSm52VOK+c4VATnyb1Kdj7zrEOQ6AZiyrmJ5N6Ei9luX/+rUIPtnsPgKF0M
pyY5kmpGQKWuNRi5SJZYYaU2SQMtZFHhnqvC+6VKQNMI798OK6s5dFx7Ns+ejxaljtm6eN5NAQjM
EU3/UKX78WvSoCtnnmaMlWLJ418aob1zTZbPQ8Hfo7Asy/6/TTqsQEWoo4KHHczQ02H309/AUOcq
zjSzIj9v+SpPFfTHrdvIHgX91AtcfQ+fBbrI2JW07XKiGK+UV3x5x/DKp2z+wOcarO3PTq41twTv
4TYp1yRW6Ca0wrc1COjSjnyMqx21czN+UC67c7QdynpJ/mKXKUA43Kw01TmPnts8zbuVq7bGWVak
IJtfSLLit+4WQZ4BGgvmQj0Pq5/zxs+ky1OcMdzYdzA3BVuGR8LzUtS/0xBFk2oUsdoF8rOB8wCM
b4JxWYpksPROIJPDNeB70X2bA84KGmx3RBK0fCE+NAOCa19nVIQHTGuHGWIQ3xgyqZXyBcAFnDAa
D7Xp3b6TFI4Hy645uVTkpp26T2d+8oPTdYHk+ZdCq/DEjSALtX9MP3gRykJQJAdnIv+Wg8Nl4DQ6
qBouwkK/ZsU7arDKgMT5179j+/LmopSdZi/aivsk/6OZeD7YWRoJIDqfQu/mXMVLnqOgw3DLZ199
9RAtfGSVdjkvboCrEvYxaocMaJEKt5nJIGJbYHngPqg70hPWHNUnfv3k3CIHJeGcS7sZpqpViv2p
xEKiHkvyRJl/Er4DucC/WWpMcE9apnl1KOtjlylT8ET2ofTtZnbJz8B8mXSVr1Q9NAXJ7tpqw+CK
ZySBcuPR4z7P3A1KYk2mKJTA443olnyEI1czO8L35yvIXZ0vlGe//qieH+Nj4rlzSGi5WW4Djzo3
Q/gQHOVppnpToh36HJdBs5+9pjfpaa9lLWtlbaI0su6kEgyVwKeBKyJ6ymf704txVZg36k5OPxHP
vfe0at6uYOJt4e9/gQJoj4O7xytO52zP3SFwD1wk5x17bZmDX2m8RQ+6uZOd6CI9pDfEbouzlWm9
AeNYLXyH2sfgtGSq/IFiMf9MpeRw+Cg8+U0JdB1H3fpQGlijLJoZMR4hHo8Ea/fLR6qn9UKrndlW
SjCtpCUZs3vJb966Cq5zBIECvlICj1Hf1tF8tZNvn7coIRaXgduS8J6yT8dwlpjVH1MUhUjk1P/o
1zxeqMUAv5DJCT1eI9kUzjFzGM18X6+PJK0e4fCn4ZJZFccJBbMnqxE2eEIQTZghUrpBLLK3/u05
HCtyFeDrHfukyr6uFFrbxcY5uEyKhvEQcurGmRTZ4Iv4yIxwftrQWQ61W015mzU2RDG1uRvR54tT
BuAKmbNkWvuX1UxEOWufT4Gkk3pm8avtppDAK/mWUuTGnKhgAOvrAz+J3JJNpJcMl4z7wn7fyBJv
49qu4fF9wv0s5lxvOQU196kywa49i2+dif25Rv+mOYA2G3b5cw11UrYjHsQa8qTcJiYUwZkFxDlw
HgRRi4YlMhwjvxOLSQ4DpHWtSyF3bXOADz2zAOgRVY/IiOXKjn0OKE+useQrfpY+REUntoQr0sG5
TIrRGtC2cmhLo0p1X4O1jU/bs+LO829YxO/VBeBbkthnsj1R2WhjpA61TeCe6mPsi9JS7SuCKxr5
YqVTmHxkXJid1VRgFFjG4URG13Qtyg9QfzJG17EnxZqF6NJBmwaYBuLZv0BvRt0TdmYL0TSI8Pe+
ALWzKFJghsj+2obzG4/7nYUPKpbdSD/bZ3w/D5VUKSuaGejJ9ZnMKDZSKJ27/KahExPo5B3GYb5P
lS5tXFc02eujd66whn+zQRwy2WLaf9HgO/t5OPKJJlxNt/uPLTtlKzCCt6G1213rtke7IjIHuas1
uGnlVSNra1Und1EoCXQ7W7iXhC+1B0pQw7IpfgTCXWSo40/LshzokwOmt5q23WNaZVRCw6/hL2A6
fgYKGwa4xpgt1EEhjrIR9j74wSIfGDqeLp2cd7+Z+rxrQoAiRVz10rf6Di+N4m7uTRXw5gseX3/Z
jFUw2hAFsHP/zVvAO2T49jXktb7gbOodeCqXotCYl3v7r05BTpUZVwVyQLIZh5T52nh5+tTgshs9
1Ym7+9fv3W9o+O9ZOPTyKwgUaFvy20S/rDM/ceoWf7uVN80MhSFT3sv1sCX6yYI/wv2YVk4F4jWo
iKqvNMOXBYICrqO8zV2JMNxaY4Xr6jB/ho6kZT4/5srOI47TthNMX7rEimvowrDBGRMR+b6Rmd48
V1ZcndFxOfzPkbPLSkF9eglIvLSdLTCRjiQLajMSd0QHxn5OSz5bBdPbzIlEmyQw2BwIeJg3LzSc
BH40VZpG33RNtOgttLOMnKKFauqB8hWIxVVkLaepVoA/oZX+5Tr31vIBhxOhNI/cpD7jPYGH5m/P
WDYLg5fGi8Ry3aeHyEK5opV1BNvZFhkrS1RVZ+ijLv52QU9/hwQKecLE8kyu1FLJZwzGD/5b3P8e
FWToz0dQ8BewbeVWoXLcp2PI0i0xJA/kMpAET3GoOCBTH75iLjcNlvZb0fJ9dkIWzwnmQ+X+szkS
Xd4KDWbwEXono9yT0sda1hZ+RAbi8pK8CvC0grop5aDHXe7SuI6d+9IdZcoRv35TwXkOL+6FCijk
6PzqrQGf3dRU+vuEn4+WnVqsWjR3KS+l84CGkfcQRB3BhcVnXHcAvoJVpxauL8ZfYRv3ccZP7cKG
/QqITXmWx4MKGq7XXQ0NFSdtyONgRm1AViTTYZyTvpkLSL/JbGVq42w3JrYbOWe0sRl8dimuWRWv
OKm4jleHToX9wD4OBrGp5ApFMF8utLB2soSCBWLIcQl+1JuxeK9tvBzAnSM+yMhYDG124UBwMzhh
cpMJRL/i+RrWl2LfZ31D+0RHhf09VL9URPQIzdyoxPjl5mRXH3oQ+nvMjenfvw4ZHthBTdJ0WrrK
dYcEoGGMxeI2j0FUFZOYkSBQJ+5mnR77DxSLdP90+y/sIAJoQurjh8AFJJ4Gff8gcHZVoDWjtF2b
XjNezd8Zs4q6F5/7IbnOYKlTx2Y9aScZvDk+rHCFue801lAC2+tQnSjLTfJ01rRLEBtDhmSP1vMw
/KvQ/yTFJ9sWwo4F0/6QpDsulCg6uYBSvpomoLF6LW2txol55Q3xh0cYRoUFsdA05hiKzzr2D/X0
b7JAATt1lmcHzewAXAnzaVK76CznaEIkUuYpmu1zU+12mSMC/70tBvXmpvTMFbOqqh+TfiV4Amin
UNZ/Xo8yPf5j0igAEYoFYAODpqBK1dolxZ+EqNZxsNlrqUX3KXH8wnCVur1geCQ5EK85CUoAD1oE
7c/D7DQQcHxbrnJoqeMqUeMbBdYODXBmIP3tpQr9gj4xzi6j2cX/EzA/3YfNzYkLlJJSjrDwOrfj
0o1HoIFPe/uFgrfRwghYZYt4nYkDN70CJbXSSItL5Ml29n3Xpm+SmV0yIN2naRd23j6a8p8IkqvZ
c39gSdtOAQkQYCNBKLOGUXn4wivRZx2N++zk0NkcUo7JiRAaGi3+PC6hV9v7K902q/8Urm0wAtPu
kWzoOP4umaUO1sJKoDipiLy5augum2+C2ZOEFlMseXarmmtZ0nJMKR/MYuQkICrYPZZi3gwM6DyH
IaGRLDVJW/GCb6xq6PY/zUXjMj/VrmN0CF3omgX2TvDiUtDKx1cVaie0rISVhPCOaqwTHgn39zYT
RgU++pGj/OHbL1C5/Khqr6ScYgLmhWVo+JZD6NUVOc1SjZ/MAZQ5Xbz1rosbLRjey6klxRWYigpp
Aib625pKQMAqWMF1PRPtYQC7PZq7kyORIhcy6dJOKhid8a3WvXPsk85AJiX1CdYUr0LE5f60TNR4
tUZbQYCMaL1w9Fy8fKfrbNkuo4e5JCxPVBFGQKyyGAydj5glTqzuO+Q9BY2/Kp2Ms/2lOtF0uPfX
vuMFinc7SZF8M6Hvt1xlLwvraoCEv24znCSSh3zYKa0tcXDIkINSzGpHcnXKlLSsR0QKBi9oXdd4
FOcTvJOJJWv1aOXciemPHMVo2uGxXhx5rRy4/UsAaEjXPFVn1VzrZvzaQwJn/oGAK+Ptcv/9Ts4n
7MAHAV5vE3n9BERU04RSAchwccN/jVBHm71agQL5xP0i8ILb/mspImlPef7ZOwn9nh1pnU58iWMK
eE3O4pa1gHrmwxMmaeG9MhcblfnKhqF9bqIMl8X2pEZsG8VDE8s2wpHns97CCxV8/Csg/TRxD5xx
6Ptj0sIUvaiilE5XPpkMdQ4BBNnT5y7cI8+iPue9P/y7+p6m+jYpZb0rebAXD4lThARKMyEbaiQV
kLUhBm4fTv9qV7wMzc9jJ0Tuo4jXutcws75XH/coCOgPKfSa++a3CPNvCCYuzk6M+z/uNJPic1m4
XXzCgbefQ0uSBq4mSj0E1OBdJXAaPwlLu2EMcCuhNEZ9NExzHJ9z6UiDDhJbh19O9xbK+TnpReFW
xY7UyRwbZeRP61Lt6zLs/5EgZyV4zz7LbnuyLriq+TfJH7XRNIifQKdC/6ACp7g6JTVWj725I3ll
o8KudLThuXRVFSmrgih5VUqwFz4bniwNtpKbcAo7ezwAvgywBWsMqfsTiWvaZodxDQlu2YEoO5J0
OWjLvCtjSjtK8eFwzsgUKHvUEEi0AVy3adk5iak/W4D7dgc9ynUfRxuGK/m8YB0foXcD2gPAVx84
YUfmQtQpHuiKP4Qdo0b+zNQBKiVeEQ+Tx7OGNEofMRQpgHweBl+Dd8CvPg9bMUkX6HI5Ies6KcnP
2RbCdH87r7nx7Sv4KhvmKHP1urt9m1uIyfaBUp/GIabtShkGQfWrhzt6PIBI7Ds9bUHseX3hCvyd
+U23L8tzhBmp/OytAxJ6Di8vekCyY9bzBI8JGiWyHDHkWkUR3MuPg1XwVLN7vKh7nh1zOUoWslqG
UeBv/lUCHGQEfuebYphJx3Is4GttLvEtOAS1VjkIArVcLcrLTtcYPrSFpINF0VUE3xPbQMoJ7+ik
ERRFhOs60lHK6qFcmxQG8DHBUdmVGNWvL9eBNmByXEw6h/OZGKQmySgy+v2uqUjH+3JIQKv+gVDL
AjWJiuVe8s2vLl6w9nB7iBlHZOqRjlEk0HVHjfRtK8oYyWKfCgdOM9A8W+9Wevf5CTIRYaJ2nyID
mfBmF37DV9LAfuwmY3AJhkhxwmVPe0Gp1nF7kkCEob3kuBor1s57ylBjXyI6BXIJLYCe217wNrSH
32v9uzUu8TelnSuc583oWlMW9kBb63NSs6aao7kz7JAfSNnFX2snY4MZ/MSxTakBGr3lQdLnrQhY
QsMzGvuxHo01usNm/Zh67tqXGtg6bj3OUbR7QpW+pWxtI770GPh0HCCryS6fCJmcybH17BCkV346
/bEd8eQbWRcsLli0QpZV6ZHkYzIiy58AfctelGglqqvXf48bFhVEqmoutrrBlfMZspmV20Ayc5jV
1N7uxIp8HZ/CMzdJnOKRXi5luM+FscuDpIKsmH2tqrhVG/Q7X9SrvgXyZxj/UR6m/ahzPqXQDhSc
X+9yvEdrb/h137dnNCSAtr/ayQ1WiDeQ1Mi+VKWGJg1lbxPBeuRhyhxLQ1PbUDSP+xiS7f9cnJ1J
3RHBxXZoeC4NDaaoJ0evOzFo9N0xE1EBJanK7Mv0eXHPPqNiziy3KmbjX0hkDUUBMc9njCqjlAR9
3npfQaHc4hNmWPWBotS+nL6xhP5Qx504XMxrsjrXNLnh7h69wPjrSoQhWV5xgccj1AZtb8EJFD1x
I3TTxxy20QxKLBmLCJ348FJ8O9p9qXBWZ0NmAcMgtk/kfWR152eL1ZpFtmcVT8Aw5vttifatRnp3
HBcB+7FsF5BqsI/X2O4HI26WoXtJl6jxnAW+XYdA4/26nY9IGHB8sym1y3PGuJ8s3Nq63uW1ysaN
Zeoges+epMmIzvbO2hFsFYtes2qxxoSa1sfbSO1nMHh8rioh9VCcMKKjcM+3cUTmagSmFneF75I+
O7MjJg3JQB3SSzPyw7O1FXwuRv+r3ViZyKhTICYuMMTkQvxDZC8U7gSs5RO7QTghA2zucbw7jTYk
vEVimiEqAwXhilsHAuNu8YzCDDRnn2Ty0BDXKRhWJIfE4CD33lp8DH84D+g1IIDIioKZ7/BKzSGL
ZZBAuvwGMH+rdnHXyimvPY9aDC0o7qnTsV4Q0WcvduT/U83pc0QqNvqYYXtEZ3cosyw/tgAwzwK8
OwrDCEVVGbxg0o1sg0p9AUEiSV6ABNcXjN7giOTNQxtOaBK61P1y3PjCquNkqai2Y6KvRBlaJskI
NdQ7OQzagvtwIR+NJjTNSqwyo+ovqwKgTjxtddm/udnmPFt9AZ+0axWEy5z6kXxrcZUbBnIBsJWi
oeF32TXrq47YgpnxYsFYZq1qAXSKXiXkRsRpkM/a5Bk54HXoQLPwVYG6WBizyXEaavGT6TrgFqgB
0zCwfFTzTrlRaoyu/ojiTBXu4AyHisM8kfVotUVhJrERT2dl+I/kDxedXt1DSfBkOnO0IZVkxTuk
LF+1L5AkNoPSnCXpll28l9pLLO/wdv2mhPOzFTxh0BCyXkmGEyAJJfE9S07rOKzamukloXhrTlrQ
r4j3gteNfQ0rjDmb+9z8CxGd848R8guirmzpcG+lu8bq3FK2Ow2OmaKEvtxMxuAFrKQnIUQsYBEi
VpUgl+8Z4EAEdfAMeKOvcuUy8gDZfUjCTdt+TQ9r0uvLFcksKZKAkzDyIdJHMRXE1l9T2DwrJJDP
QCVEkbEnSqHIX+5elqiRs9Sl0vjOIxsPb4eymA8R9PUrepfclMj3I4iVahEydAvgUvY9uAFK+flt
qLHQ9CDL/eLaE+MGTRG6GUz6fm3c2ctK9ZGLvsHufbxWHLvR2Qe6T/02zFALoib30cdpbd5jOoHy
D0kvJtUWRKBuNdjexR0HbBKxOwSoWWtPVae89eFXCR7t4jv1z5dxRk4tSC3ytuY6MeKy0CA7sp5Z
v8PDoBuet2liXblp/gjC4amTey7dmdy7M/PgbDJmNuqM6hBfBYCvgTuF1EmFtfzSFN4F/7YJISR3
JpBjG+vNzw8RSFbI2hhpY1hgAiVIWcDtTIF2+Pn4FAhOEHY1AFJPQBZtIjx2t8xX6NzhsqokV2x+
XRtfFPDZYgHrdTK/cMxVR3hy5SQwFm4wSKCxdk5/OBxGVuyki5eL9qbtr0n8Y7t1qi2fE8+lwt9/
bfdY80Dzb82hF3cTe9c9BB4DhNEkTPhJay83Xsr/oeg3BTtUiwZ5aveZ+6P49Q3UxQ6Xq9QB3idP
alM2e8aM0YJNW3VwW1ZAYcsI7DP2FvH/IZYqAyq6JkV9sjQpWn6Faf5eoQpI4rtcASGu4b1fJzO2
JGtR0//pSFTv2Ao3RBqPxi6dEKdwy+16BcGvU/3D+/kwHl+1Cq5uiXoRo6ES6w9MJiQzNDcaUiYZ
tbJJMX8vIWgPRYdRru5y6ZVeNNbM6yzc8E7su6AGJ8ieso+MCrZIidd2jVvh5Ya3luhFC5AKU23D
P3m0Udk7xB6iuwf761Z6C9OLe0gJCuU1JHMwoN5u6RQkCaEj3AcDxuTOSeL4Y2CWSYxiojvqbRtB
S+QN/SEwBxoc+d0qI+/anWG0jvsU946IGORNU6+RrHR5ig7DglhjuyIaV7zYMbkDa9Ndx4gzSAZC
plXzk5NjouDqBQPV51iOnOavUZsAX2Hk+a64x8dnTn3dHe1RpyXysfh+xVxM8DY/XBRTWZCQNUec
I0Z23GFWhHhi+/VKrrYaBkpz3EhUw/aLgf5uraf0PK6VPmUD6ARYDeAJcb2aNcBXbZ8eFjC/vZQb
75UKwjNE/YJo7IgKIug5npGgIgqU9gdG4T79f6yCuVtWcCD7eUHDx2GSKNutEdCLBYGi7C2s7MKs
V+kLXmYkcJUuk/6jaPsnhjljWgvflczowDTZ7lYNpNGQeEVrrsdV6Ld7qxzUG1dWl3/L2CGfzS1W
Yj9fX81gsuNe8O1X+1sf6DqYuC+qkVsUr0DmYUbX6BZQKfiH5zPJUzC+dQZsqmBUP+e8rsMLwckk
SV3fBj2V3fINW6uBtoAX+CQp02nK2FCf79baMEng/XxcSo+YRjs2NTJ52bNoaoZOYw3kdx4rsJg0
arMT1crPND1jKQG9gT6oRS9SI9gWCezZEfqSgrbdp4qTnteu0OeTftX61AITcZrr60Emu4SJaETt
23SqvqgcATDvpOoIN4dnaOWFBDyPI2IEEqGrIQl0lqNLEypvUWV8SZd9DCc9s0aCl17Ra5sIu+R9
vGPwYvAf9/v/3KcLSOi4oQSvFECSZvF+2ZdW68hDl6UdLOEi680jgEC2OcA5+NMcKYC1V7kIDPhq
VGxuPh69SiSPSze1eC3zQgrZ1Zin3DuI1TTGkx5RMZK8o9nkXBQf8ynIlZ0lvg5IJA6fmOpgO5rX
i4ii617HkO4+tfH+DzIBp3JnoTMSz448WK+S3bJHq/uLK9+X0vM5AFV3oYcO0yEcrrsnrezdfQ9N
JqYjR2jO1jAezxLDdE44Us7ScndNsnilTxWu8pMsfrQMlffVByF5IB1Ul685RKZJTpiD641NNufP
amYb5sk3Kps3t/zvrPDrKl6c2xtbcmxV+LgliwNostGWFz2DfHuBITYVRO3u4UpzjoiHBIjJeZKr
TWjnbuCN5QxWODrwaEYxk92B9ipir6fklIHvd/UsHbVqL1whrX1FjNMOmrKtzdIvc8YU7dwE3G56
+Z8FCCJtMy1LpJjHqRkPGfgcE5IgzfDl6hj3CgllefZk77QwpMM8c4A0rE3pB/BDl/W/2xaRmoYf
wafxjmd6JC8z98XLkFQ1ZQO7ZA71Kix7Qmoa2gnFdyLW5HDtUiMN4W4vw/zdus3UK2kQ48iFPIt5
x3SJM5CFONrNypRr6H6/0jM9hXvbDrYdTA1NzaBnotoYgzqK2SP8KTYT3nINbd+7YcsrO1RCWMpA
V9W1Re8ozCxx11R1KYWunFl9lwBRjZ1Okrv2IoM9+X2avjJZJnI/fpEAT93x9STVinCh6IilpgvK
Ymjy0+rB8oWGtaWmiZx3F+UGyaqtR5ToozfBVbewzfvFjsCIcA+rhLtOVXwGUmPhCVc2Qt+LI+TI
GTUsfZX3AiavsJdAOFVaIXD7+3AJuZkTPPlwtrU0mwqOUoz28TOkg2t8VmubORomUkfFFGDrmdXu
A1n2hlBRikBLnX26j34ghf5XKumBRSkAgTk0W9T04xCwLA27tk9iHX4+qdmEd9FeFd178IcUbpxT
IohfHEswWLc/TxboaiJK6wC4G2poe1HUOWz++ZqXlyx+AfY+6YB4692Bre/T1gBBM0xmiE0qh8ro
ki/pmxIN80Hq+VEBLdTJREnW1mhVX2GBu/wN1s+rUq4sIBgIwobIOHvN8MJ1oyIMw58DZs7F+A9S
ufcck7rFwFXcozCL0AVSlJ7BQs4gDotJX0XVMN3lGKmO0s9O+Rrzif1IufhUFeyXfIsbkz79wBa5
15+hwlQnt3elXWcxOSeCyk3xgnPaRhIgPPGlOcvO2x5JoLN7/EHmuBHyHSxWTGrL+djr6/pOjY8x
XOYKlD4Sd7UN1Tar49yb9XPlNu7BtgtxxmyuiMCgZqDa2zDsqqROLNghFqeoTXeS2/P++S1Jyioa
9s1eIpevfnbWKrO9oOThBFlXCpCFwoTsj9LMi6V0/C3hMdRM7/WloMNy2oHapLj02sOSrVjxTXKL
3jPDf3y+9Co75rm0hDN0t+ySBf13TeXSvib8cJpPuloCbtwMpq3tbBpmIi0E2+AMUXtLAGx+R+7J
B0YB0xt4WMUQL1QTORgtcdBZpI4dy0lqqGQemNQRmdhU3ryZFMFmK4fUCN24NIaUajPw3Pvv6+Hf
9hA8aeFZO05M4iEzarkxoXr6LyoVSTLw28S2l5LugQeH1EUIgB+sh8QTlmzytD0drBtjWRrcT3B9
UwWW5QMkYFJVjAcZuwSlXTELXlexjO813silOEQlMdxmJ2sYZx4Vbe7Vi0P3tdPxBumE2nhVCFVB
HVvcHwkIFEQcJ/WO6LsU0jA3IIetzjGfNKLy5ndozBLXBsCO76YWFB7Dxj+Le2o0rOobOLvlf5MA
KCx5blIhpjn1lRZy6azgt5Bp83tEagRlCFjyrfJbe42SeTGjDvGmVK+sle00CU9QitnmEObAWVBW
KHiC1Narz7gsvMrMy1synpqxIIwTqejETuU7s+pzPKV1vo71Gsu37OYBG91dIhPgFUMDeqqNSB0Y
DcOlyqHVjiquticF1DdT1fHZiXUyFYC/x907ALtdMOIzTZEHzrEbXnUQFTrFMkksvFhKMMKAkVRJ
/X9jyMo+k9bnYNbgenkSDCtTYOINut0N5Wmj4u0gLacLJg/u+c2viUOeyrYdvd7Na/AzFif1FcvG
lQei8RaGN7TMvHuuZ5FhyreYNaexx1kYS6OGFBZcOXHSy65UcvEteQJyiZz3z+76punvgia8VuS8
gsbniwhndazeE4SMPd0OMhZ6LpJGyK7S8/9iUylw6w3eKAEB/bt7TNlVRbLPvJrh5Dtln0zHa+uJ
1RdYjCE4Ah8+wbS52MSGJpcGCofLGJwuxQnkzond5+GX3TiBVxiMMZQnODq6LFIDehAY+uqYYOw/
1S5Sue68Qjjz1GADjHKAHosEBLQPpb0wNzds7QuzGIfwcZUuHhnUYzGfi6vuo9G2owTnEAkbR6eE
MKwAconxJ5M765MlPEFo0wCyVEnxznnZCPFkucdglp7/LoGqs8UNeI7V+NjBYEdAZhL8JO73iwYY
69fQYAFpZHwMnK2G2JgMO4cdjOkF2+5xWb0hqNePjc6FPDFPKVg1GXSRVHZzEBH4s+Y9IL85yfWq
K1AkpsEcTtWeoFxLczlgOiRfNm48+oFgdx7eO3+NphEgeo/vSuuGwd2TmCpk6MAGMZRF+M/HFuKI
0Af8OEVVkJX17+UH7xfeoB5dWHpsf2jf3F9+6L+Jae7ttodhSKolxhSTdKB9kVkPdAdfTh5dj10G
SiqYfJasp/d3vfg02Pbh9DuF/XwGv0VWkGV5EsJwXjEofdVYzgjy7N1NtO5tiU5BwYC01vEjlCXi
o6hy9h3eypMw/bwWBAr3NarYfHR2wzbQQWFUybKJypb4P+brS9L+4nacZn8f2ZB0/KAvhMQmnafZ
rfh1jBPvoMkNkofSqXVJBAWbB4qgfThEZLroB++3OHg7RMXIDeE+9QMr6WqOOStaQRcc3PfEdOpH
ptASg0t8xArIK4RnR9Yxf90wJ6rmZhqRAFdHE5U3rn7dzv89PbdK+JqP2AVcU9omU3zDA9FhOXmi
EL4oIGad7eXWOV51cXniffrRKbeW7cIhwgH7MxzJ0UVia7M8n5HpuszcLkx2VIwyeNt30zmtX0Vm
KHiofSDB1Qea993foxAoOM/yWuHtniOa0TDUxaglW529KqU02X7yzAYwWYZugupTWTj3L1vGcrKY
VPAPIwnWgpa9hQYSkOeEkexIOmSZ1++QAz0c37IZfNF35WriskdBoDKcaWPBz45c8/lbDiTLu2MR
ov4odj/UZ4eIc9bhq4ZEhIQdlGVhPUPewMUzpoU3MtyFvV7AEQwuhZSPe7PBjAUWJLdHzP0rxsJ2
oQ3efSLytUV3Df+Mkibmt0wtCKeAJLQ4yWVxF5GJaeNrRNQcdox7NvCMPnZAQQ8+sNaSGxLc8Cry
Iz11c2iTPLzmRkGgU3jwfM8lXz3mKyKpjT8qa/46ScYD/k6fN7Sqz4TBDzT0Ab6LcE6ceNYjn4um
cnACipzn3KfBAJ3RHX9XZjsciZlhgksxOVVV9lXpgSIlo2J0QUbeUl0Ccsmo02/kqcoj4I5IsTJY
7VpjJHsnOxwATWpoSY1LTRSQQdHl1kuUjX2r+hFHa++ZuNL8/aAQFQ0lg77y6pQm060v+24C3CeX
5hALpExBYPttpJSwQPLSLoYjbMai8PU0a0m7MvDJ2SaeU3AMM2TGj3jJHY9JmpPpDAW7fNAXpCk2
liznpPE4iHp3DroBH0C1c794pi/MBs6WHEfN/tueBeEWhFnf62nnIM9XD2boqoBigB7moUHsyWnu
DNC4XmtZRK8yv8oKQfdkewMIamArNNWOZ5wTHcbfoPTWdZQhXjWRXEr1+zyGj6zq/RqSbcBgaDiN
76bxfUbH/215mlqbdFG0+FeJFfJAxqUg9owKF7+1yKm0HtrbDeqqYSdINrx1ku3qcPYfgS6iSj/j
c5h1hLb4+Xd344D9L5/6vUa41QCJ17Me3it2cZrccOW5x5OGa22h4+kVqsT//lKkHI4Eqii2GQ5C
i/1qESqKx7CvU7shJALvKs/H/9etDmFKmatmSN6l2HuwymCMx2lExu4h/lzav92Ezfmk0Aq9zbgX
RY0vevaMADMCzgvjrSbdWPGzWG0phpcLt0kEjUoRJS9mDXHg9byTYSRUPvGC7uuPO8oTp5SUjZrh
tnJSlQbjI9A//GuUO25k+xVK5RtjQI4/e9S7mdJd9eoIS28LqG0I4itG5ASi+rBkf3yEU4DojHXW
hT2KXZXl4vfU53BlcwZ6bSAuWORNfR4WK9dhmRw8sckwNCSbjtotMuo7Bx7M1G/0JjqkXN4jx93v
hAXrLFcnUTJWfiKK2DU3nkf2q0s7n3ZYVe+fZOF51NUmLe9fOJMbSOjy9Nh1LK68HWZJmfIPz22q
VXy1HJ1Xmg0s6vJh2T/RH3GaF1pWE8/ocwSCKMOr/pAXcq0KIlEcoE5iofoVMXE0AykeNSZ13jFr
D+bK9aaRf7hi0JFHVqMv78UJetWx4W30iwVErK93CNB4cTOSHEPx1PN9UpEzqcPGYoBmLKfZDCa8
S2K7o3DpC/n1ytqXWxJ6FpuVVwwGcJL6aPxlGgJ7/Ug289X0UCQ7HGHVNvy0EKtgOEl1bMaHq47p
dHd2xxrBENNq2bu6a8F7qtHdH4EMkgpEEYgHmhlnM+NVYfL4sxJS+Lea6AKe2yLpC9SuDaxpiazd
7RXDtK1/jCuG+xrlFOUPXycUBxrAM+bC/XsMwBekbsr2BRMfBTWKs4eTo0V3m8Lc0wDfSm7G5ygg
zGM0j/IksiO+7m1kzK69Q0rEF6quMfw2z5HDs5YWJV3286CYsX7HJA5VWsAKnvk+VUXtPUwTykkw
TAbR7U3Hm50+e31e01Pm+ud0iN0yyhSpDrapA5LXbczcsjKOmS8Vc1wZhcRktAI/FEw3/KsuzEVI
YIIifSc16nsIWeUhI1UNJIRm2/s3439w8+9GV+lkaRFL3zwHssmSZROM2bF/S5PXKCR0V0eY/DOl
nqOLxfe9UFrRTA88Jm8ohO7jVB70a41YBa5GkDkprSF/sEBQKNJqDKuZNMcvgTh4MQU0fIRnPO01
1+SLEiyEE8U4cKq/nikl9z8zDiXBRqz7MitirzIaNxUXTQfZfHYmQTmLTVzaQLe/QsBUuiVUZ12W
k64Tu9eFTPakA2wcF1kIJ45IWNqy49m6NaI7CS5ADRMwJeNVsRfd/Oo6DZ6as1pb2ZOhSjIj9p/b
kjA4YEvJyOdFmIsFY/Q74gNdJZ879pHU4iZe+KdXaADtVw6EAhBWl/qi4gxb302MBEDNsR3ssFPE
Z94XWexhGnFKE5LyfoODmOBvwsR8+XH4AiKDeVH+hNIE1rA7bGHVUI97ToAiFgG4Nq5yriC0EHgk
6r251jnUVTW1J81w2oBpT+FgA9OyBGsN5fHWf0hzm6NRonl7fnBl5tfiF3cBpv0TIWnCBBgBqt2V
oUI5fP17ZPNzdtrshcdTeNdqO0L9wCaD0nFZi2pOBNnxoY4FQv31rKAF3soMAEyb/D5OzHaFWnPc
ctMt3AMvtmtR7N1R7oMnCJEnH+ZhvgWordJggPdEUDHXwGyB1FkBwWIlxVieMbD96gIB4Go9E+HP
xZ5CMS8YzhD4bRtyj3wdCUW32qP7bKrSUkRnTW1xICD92Wj/bZXTcOzynHcdZl9gd+/dxVF7SS63
5qNnMRoUmQOe2bm8MzP4xBqEWeUthzyafvELRJyYXI0dtjCHHL1edskEeqE49jzluskKApZV/QXz
dUE9v53/x2x8AtAZZPgLr8Ka09FHVYy23wWUW/o4Jnqxa6v0kSwzas6+RpeKNq5QwjHmEQKx3JTv
YU9JuNZJqpJ8zVblx6LekLG6AEogpmqphANA25kwVBXXlNucR7e0dqv94G/Oua8kTFgVhjuNVmFn
QoMbL1zvNQg86xe5hRG9IkonSQb91l6DQ1+liwQ92mIC4EGP8GrVdBbyAQqZMh3x68yPx3VC5rFN
eJx/Qwm9mf1rDtLX9e3en5xQT/kX4Tm8oaheTdhbC4kETiRDC+xnAd8YMr6KpRBVU60vzuzKj9Xb
JX3VxC204W6jT/kDV9TRudZN/qdsVVCbj51nmc+KNnC1FXYACZ2VljYlKJaMneLmMiIA4Sde8xTy
YWE/CQYzpetJkjvD1icADSKSODgyNjBj9BHxA+VANDQS5IzK4vwE3Q2OZnNrPxWPFSF/ZJc6v+c/
53bZDbsXJ5ElGS5rtfnBzcjnn8gkewua5fVWeIOdSLImPQRWUVcDhZJe/opXzijs8EhtK9ZisbeE
sPnX/CDyah3FCldqWtgIQkl1HviMwiVKGTU6KqJsbxD0HafZyZKdUOGmlizSdXpbWGyiRx8UzucP
b9Thbh7Z9MFm+1g5JzrviS8lyaLRtc7LjWKgJQV9e4PB+Qcj+TdqQcu/lbqRynRqudJhV96zUbvI
VVwjFPgNZOtBXM+erIkYYSyLCp+2OiA+h723Q8tJbXClxsJDnoMq690wmUr/EbIBmdDkpoBAFiMk
q8RBzUbD5poSwx2YG4P4SPgkdGr4FSOXri8EtM0fbdCW44LBBSO/9FQ/yT3QjmKA2YM84o3fUjv7
387xdjG3Se56m6TA9VlYonWk+Xi2TBX2odUAlO3QS5m3n/gkIvlpl7otgZuK2V6zcMHF93HUEEq7
6LImDmpA/c1XzXmMJNKLhuSCQvuT8jyTiTfZLxLmXK4qxSYHU8jPDym9jQ0lHNRok+8wdXEDWeMI
QV///R7AjG835ntNkk5wQEeCLbYJKrKTyjnAs/xynVVyjv0xc9kSottNwMZrDiSRQPz7sWWd9GPE
iNGzHZCO4CkfxqpUbFFBfsA+dQFP2MTaSgD8WeEZtBJh1lCGPCiezhTWx+630xU2yU4lt71eepoS
Xo6Zs3pFJiQUdXY1OKw820dalUe+8OKb6pD3ZeCo+Zr7J3R0qjSWn29IJ5BIjuEu4kDI9Mp5P/Qj
yKVM8NsZr8dhN1gxwJ+34wesDD9d79fAlrMr0+ObwaM7uVMoJFxxnukqRQQOD8oM0B/T7/lHguw3
uKgw0LNdic8qAUx5V68N8iRskWKEIefinU9wOUc1H6Be77Gop5DcuveQQeen9WfbjgCIV1O0KljO
AutQFqFT9ABNip1hU74I7SChpc+NuXqDymR3XtwIqniMSdP7y+TkVkFU2l3vc2J8lMfLAqubyXc2
W5kall9sEiEUl6ij447nbhHSdZkYeRBX6JloogBAFTkQtlCJtyHG/+Nq6qbj6g5D9UWPxsQ2K0wV
LuTDmeb8krLV7hv7VtzM6o8rQyqDA+MwX1/xz676H99XDAQhqxlkStNWIbQKnPE+LnyF/fRe2/vD
BomWMrtA3dXOj/N6MO3DEnyPPNspLTxlVUhVEYM+mld4zhIdaONhs4BV55zWVfaCURr0m81+dpNM
jGhHako/XcItQrPaf9HVqgNqsZnOkTCETcPAApf8QeAJvclGvAl6BJyaFqiC+ck1FHn5jCYpPSm0
zotlj+/U8PVZEq49ykBRU/1EQEbGvmikLK/SrOIWwOxxdPUFmpArSykjpTYAr1uO2uCRVOKZTgBP
vPXcI/jVA8b1SfvyC+/2lolv9xSPcobBntzf0nxbVk6ZpGJZd2iWBWIzYpiLOfzo3IWzlxV98O25
8dsnfBv4o2p0fOeki8pJ888CfNz5b1sRt56DAgJLtZD3rfMgS4vQ1SIT/NZtyjG5JEzg+zrjh4F4
/Y0vAQezlhpe0h76trXj6L83DkAVNtfYDgZeow/Amgb+FjyVNfUeSllpl/dpgoRiJ2JU+b3SyXW0
sUqPf3EBRza7AKT3tGRGStTOp2emOts+7NNIyScs5BRpJJpltjDW2dNIdNVPcF43HInjLBD1qa1A
6g/DEtS8Z0JfvZ7SXLd/a8z6a/he9JeyXCBLRzRFgmlnQW1b9scvPXN+I6B1YucEHIOzkyE/geeH
mA9mXWxdPTdAZWFgm0i7+exkhumkrMom8wI2Z0+QPku1L230+iEg5d0yDA0VIaedXYpQ0v20vq6C
wuQocpHjpcGs01aeyoJWX619hwsAHKdIla0mIsD6JuA8nhctAajVSAjujsD+Q8X+nEYOUSD9a774
6Hfn4m+W16HuTBURM/DuPB3rOw8tbVrIf2ytmLbuPJC7bcfdoDJmBCI9HTAh5YMhr5oIZVvobrv5
eXWoBTa3vmjBFbBHdiujcOwciEVR6LYim8VCwLX7nt9d2c0b4sCIZ5kX3oL4YQ4ch/boP3NYD+KH
LwzbFu4hyDzZNZxDRquh3kGD37EQeMQp6CBEJTCblnABLHgTHX282GIJQG1tDoq7J9jnCUjHmEaT
hg9hBAc1B4VR68o3FvKMKnMiCq0XMDyqEN91yeqR7oWl+79M0Z7oYCpmGlyctAcQ3mR1Tf7s+4/b
iYCqOqFfaUBNYrZzqqSs6GmdudRwoAJCNumMqHyQRhjw5o0qi4qPsDHUqAEufNFyMFIPv3f3L6N1
hecfi6YXukKKjfFIfweJzsxsUooZ8kesYJebNP/IWxtIDHGjPFh4XQzTLpQHwCoHbT7W0yFECTL8
LspFUZwSRe6v3bHTc+vKI/zUrm1hQcz0B3X5yHZl+FvjclhgPdfQY6vxXawWW3SOOa/LPIlsh2Qb
NxBwizBu7OUjUJUl06h73aP/VdhtwljZt3PhY6/Drku4roSYLqMblUcxDruMGmkYws+a23arY5tt
52NjZfYlxXPL0uYPG43XVbhlqkA2SYSn/lsdGNRUEnylk2OBCeALUQtU86cr35JHJFBh7lnurfO5
8MlMQz5EXsIPlgYHhX+oiawPrlEExOl6vzoFO9zw5OpkHbI5RP9W7oTkcqOhn6N85CAgA+BmpL71
MuSInjsT/sd/LQge17qEWw1/JjmgCcJP7Y/YtwreCoO03iyiwqCZsDPD1GzG72YvL/7G1XxNA8ZF
4iA5PrKrbwwg4o7orQgw6uO2tts4eYzA04SObu4ptrPiM+mT1GNQvDD3DTghFFd7gpBqR4I8jKAQ
RwJGLPbbrt1r+wkOrj4vev/hFXUdBhslIdxTbGI+b/Tw3TjzvBiN+JCa7OxyWSSgpkTtP2J2boR3
sdSOy2whf3VHNnMMetTyy0U+rID/A04CUFhoYGdiNMEZemUUZgVs4eDllEjd742mlRCi2NYH8GLo
Rk4xj032ZZid+nG1CsMfKTbjkjBa7EcK5uJh4EdJbHpobeR57SXbxYhM4nOeYqgZ1Kod16jKea03
0QJEo9IBXiuyDuKugBLWny2XPkWSwxv2V7HXd/87y0UGrnWoSKzvdIHaIfwdi4Oe9mpJej7Eb7GC
EVHTLzt9CHsuIcN6I/UwoGCvZmjiE98vOmA5b6z3x0MGv8kCYGeg/bcaP0fuVQWk1SiBXIJ8ykXi
NFhTEIcIFNzVO2ZkK42Bf0fNbnqQbh5WfCwjqAz6e30N5ewD2BpqWLLKUhc0dAZoUWmmImIIfKTg
f2vlaHcos4TYHWgvP62tYJQ6uos7jDA+ogZT06lPDqyw0cSn2aDxcvS7h7H+WDRvZlBjS1loymVj
JA2lxyjZEPld4GlcDqGIFc2t6sPSLBokg7K82Ut+rE0+tRAZF0A6P582Pa8ULqnBVeZuqsy+9UQp
merhEKDarmPClqL4gVEjpLt+xq1w2Z4QBu+GNSJSg/FhBRL2gFjsf6eQwJTUO1wAcvHRFaowKBB/
BUTGyOn4T9+fbO/tmvE9zWf2bBPv1JHTLO0RUID8oRhDOmp1/lZesBnIqIO2H90LsRM/lv4SOPlP
zYsaskOaJxS8IZnb7V4Aa8z+mJp65yl+XDB4YfCT2i3QvB0pcAWCYPHou1rwAIMxaDgDPKTtDVCZ
f8IC8Gb2pfnmcPNXkZZELvtClYJvMXLZnR54MIIAYy92kWsCJbY+ktvz5CYsSayy5Cu0sJ8YktD7
Z25BGo1eataiAueMmeTBPeOHtv7ToDiCq128QosAbHhT4Zxjf3qNbIRjqhjqb3NXMXhMzFtpwOq4
lDkqSqQc0vVHJLmJMUv9xeplvQCdo+145X5tOFuzR3/f/y/4xYyvASfYg5+zUslHrrQ5WTJrMo0H
2GtkYvjrizmZhtslSUi/0e3d5KKT1+J3mCcN8HV1KxIxowwe/kOvOspvVcNOVUstsO1/j+c1Cb6g
aBKDIM8Y2onyuykOQMaM6dIKjVoSpSANry1vt7RckEnspfKj4zin0IFf25DPHUgw6XWDhdFCAMk/
Ayd5Jco4ZhmnSyVTu3aL3wWy0a7W/8oM5OU2TwZFzEHhZQmcncD3S9P7xXT0KiCAZmND7YzYWl0/
EN8zxN4C1iFOnxo1mtCC3VJZbefcS0DOnsecOXcivxW3jnw25fWRdOxiHFM1qm6L4gXSBDPeDiqT
prq6EMlS9kPjmn5u5nSyHHj4/PPU1JNVHWpg8074VpQL+fFZrIF6zyf9ldPzHzmm0ICBTLRzYghR
gOKG7bPwxqV0iCRrBVH3BzevhnIDnoRhwCqTOvAQiw2P1+jVmbgKRlEn83C0IsJUD57TPE4jDZsh
VhMaC7VuYcPpuD+bWtswWS/r5uCT8YKVaZVdPYeRJXIfJaRL08g2Xc5nrYL0Q1xJQViEfSa3lCSZ
ZY0dMj9G1E3JUX3TCMM6mOOnN0ouEPntNJk9Ac86o67QykRXWF+MTH1qEWWSjbnnIUpI8YfDjP4n
h87CJyNlJmoOtFRqAfJq5AQM9yMlYUFT9tCh2hFRYPQVN7H337/Pc1URXshC9RGGKYDGlmJKgDfD
2DX7eC7DWpQLcGesB5llzD7bU219z1de9cUQEgn9tNxzHBAybH6ZrdngZcua4Jx9utIVZ+Zptd0p
p9ugE7lPD2fBcJoKM+CEG5OWbl+6HRRDRioUASFis+K2ftc9e2a9e4F41ZZL5FX9W3EaP6flda0f
NIPF4MPJIv/u1Td3Db9vkdm5k04paJxQTGAe9vI3Ij+Ika3+TDNyiTyZ3aUdxbsoPhuisQKQDxfN
kZxFkj0acv/1sKeywo144u6miYtlkJkLv/m4frTJZXo9DYccoPAhZhVSLqgM5fcVzi2LxZ/K77M0
o+gVAf+wfMp35fbkc/NbWtTr0s2/F1bsDMU8EOsFsg9Jk/wogWz2Kk7P8sZJ2cLmVbJ0wsROlAjd
bN2C9VkcABNQs8NV6lWMlEBIInfBqcFdsRgp/yERalGRjgUMuFUETV/bmhftj25LHygirLGm6wlq
WRziz8mnuXiLZ/Qjy+J1fmoD7dywO8KSvL6X+T0IygzM2RL0Og6v4IxPKqPX9u6YPZ3g8zLBiLu5
REelKr6ZPWyTIGIGlJrZ6g9+NtfqIceElfkWUAmgUww2GDDPuQYChu3/MQFRp7WN/jy7ELaIB2sw
l5I7RjQ+c7Y9n2UzkNMuolhqciYufrbG6yF1gIg72aAXOA9EJsM84g2LjS7ccqDOlFh5Xdxutksp
9CsQqlqwXVbPRBQ7eZDnaPiiP53bDXbmUTdk7NFGc+eLsUeaFFcVcfty7z9HMoqkPz+k1d5oLTc4
pIQqejKJjp+jLPyeCiixRCYHeoxYmJ8m1wVjrxDrYv+yUO/TcMOSrKBoagpV5l1PyWYh4e1jYESA
fTivkwxj7XK5jzjQjZZ9A0V2GYusRV32kM83I17NuviQ0n3X93NymlJ8zDKtUcMrlXVwaJU/MOzE
ivN4330srB1bTqWPGg2ufJBySYcD2UG5h1N6y43r78Zz9VRpxJKFzfjXg1CggjQxIoVm+8ssOEuI
uN7V3UJHqGqfeiDMCsH7Zt5bqaOi0nkhZA127zLZbTbV4KDor2QM7W+bIxVODIO6DaTrEeo4/iiu
DT7IBOY4kZ0qSzJ1eBMvj1r5FLWUhJbSpi0y7rMETN83wbpcsm4c27K4y+sicVhRxeNHCT8qnLOQ
zhVRSWVDxB/rjMijFLI1mT+Ji2HbIXbL9Vu8ssx9CTr+7QQVTmyB/9/yYwNBn3NJ2Uztfuv/eo4N
ggCR9tTkRJs8L0ndqMWC0Szez3cvEccvuv04+fO4SO8Gm1zK6I9COhY43mtK179w8sIvxuuvTN6T
GU1cik0jiONJ4OGcHBuylW8db6KxHZoF3UHkqFqzax8Q/XXF1e31uoTIP+bQkDfLc8sWL3J7rSRS
g+YMqjpa8Cp/E50caRBsybhSjFN1GmhR/IhS0taSW51fV2bHMiE9cIxUnZNkCjeQ9I1bm7VKsBOE
+SBeODT+kHdVWD7wU3NsjETm8EKZ/eVHku072mybid2aNoyNd9/biq2/UYwqkxJaHd7NqxCbXvVi
YOaI2rS6pyfeRich655Cg1w/gAaa7NucBg2Mo/GnxHFe2L+T+ZRf5gXkugEQePwwXJnlKOFR4kG2
fGIngOACeduEZRqnB18JSOLHiM8Djh/A8Dv4uA7uZPNLnpOuXqd+iEJjxtSvQY4MK8OEi/GNZ0h0
bO88m4vDA6FgB1tGUXBT4Cp2JTv5q0Mh09aOaX+rJ7FOmuo39jeaJY932SEq/0iSFAaVURCGVIOv
SHU1xb4TUcRo2NlTQ24q4Nr9Si3U+7PxPjBoDoWTNOxjgAdm6EQyhp7vP6qfvSOnX0g+Q9RFPDXp
KQtziLp/y69sbAglD24CeGPlh+u6KwSdsXKu59MsPoWauRBqXriYxZfcrplbQVysG4kK7hCEdY/O
1d37gaIUuZF5hMl2Bu8qF+XTWd5meZv6OCZNmTlu3OBWQeYj9N3Hb7M7JDwZJztTrTvskmgWRleP
3+F8JfemXHehFDbO1WRvXvTsE3kwIymvq4EFfwgObUxjC6mWQqtwiDloPr5bm8IW6D6ohahPjzSY
OSiaBFH4t69aToxC2Dax4zpgeaHmqTLvzphcUAZjUcmntOxBL/E4YGxvDjfBWnSxduk90tIpM2RQ
zTFnToY60TAWTMeSdnFWdYp72jGxCRgNeACl1/lnK4lo2l75Pk0c0VR4XgEYPxdrmcoUnM30w+LU
mdtFL54XJnJKPk1AqpLGU+vpWEd79rFhvCz6DTR+IHyqgehzhnozeZ84xEXkwolvlz4vpeJ/ZE7G
zMPCp4SKzENFQ9vEkxka2xz5NA6hW6lkh79en6porpXn1qdPwHJOWHk4Kme8lEqNetBXE/y6SdG0
pbiyzYQeH/0IS/CPzsZwpAXMMuBZ7yDurPld5DWyNCA39laMPUITnXBCP8hRPYufwoVsZTUXN0S3
rUQ9YrCezJBp2GI80FiIgPwuea5Crg00waN4mpdTrj2Ydz4ipzJjwO0A97+bW2WJ9d2UtDDVI2rB
iHWarQ2LYvw0e6lHG6i6LP6rOq7A6IAvK8w9Y8um3jg/X+b/V+JHTdReSmbwDNnNZRTMfhVwSuBx
7Qt14JLjApYt4QYJy223yqXPihyWDnFjpgvtUbTMhC5PEB94Rc5OhR9uSayJWminYl8GoPG/KBiv
V5uw+5qVL7B46O9JyDfJl+Ngx0NMtSMAFeyAR5ZKAlFvlZfg0hQw5KH60iftyBuCu6f1nJ1U5k+9
8tTVG1LEYBiOgWHRcaaCNxP2TdAlUoP0qGVaXWo/WeAncmPETzOQUtLnzl+pvJL4/oQOberwpGwO
IJ3EUxg3W8I5ldX1qbekLWVY3HEX043d4PHr7bn7CAGKKIX+LbejCfF8G6z0BYQ/oQJe+JvSLdak
ySxUIyBjeXLs3WXzzhfwqVUxxkSiNBbidFEAU/use90zoC9tN83Cckg7fvxtaRMNjpj8V00Gz7r+
u8B/KG3LQPir/P88RzJfMqOm1JFAkeD9vs9f9FUjzv9y6PU5cfIcD+gaZkT2fT2g3bbqb2Mvyahj
+agRzfAdp/k4Bhrq/0knRuiGm7X4k8gHrvYzY91vAmbEvYkBJdSRZLyGllCgQw6f2uYjDLJRKzVP
1ajt4dCkaxKxReofXRbiNeqDOTdBeQdt12D4F6x1AR4AFkE8DBJdXnGKlKD+W9a9kZqxw3Wg8aJm
6DjtPPjJjmrlWuVJrNtGJdUx97G4OpIzs7sq1Zjz/kh6jV4p2DHqG7EfuxthAkI+Y8B7yrAH1dUn
iLjGOr8srPeCginSrkDcrdPDbLjDnpQQUkJC8P/BEfXpovV4O30w2AumwxvgQ/LzSgtwqr8CrQI+
wUH7MKFagl6xMHUIE/0+LsHCQM+9QSVrzgV/dBGYITeeUbve2N89WhPTKHf4Rnr5h27SDlQqCNgR
YMVXKRGXLYOIMQ6zJEw0L5NfM62exp/4RkhqNO2DyMrB2Wnkx3cQXCpi1ojAWGA36b53V91IdPQg
DRRzCrOSeYWoAooY5lwEUI92jVOFHmSesG/XdkyiFabEhajGuEhR0qLwElAdq9cwvUfLyCS4TCPl
MUzEwC1wlgak+zzA+2mp21pNp/WzfTz3kjdj9n650x1sQLGPraXTyP+0Xhwpo0kHpFxSa4ueqP/G
7k9Rt4QMkNxkcNlVfZrH8HKYDemQrryD14rCwWFEg329nlAYaBjO5qztzP18HOP2sG6/Tc7V7vtE
aJX79rQDfBHj1hXkbJZg4adenomz16o5ww5RCuW/HMrtEII7zSBg+pwIcmVZ96wwe/bxgFqVdmBa
TF5F0ldseJPIsoX7oMqEiX3tNh3COvEFIItcYSjjSmBsYrU2ZOnImSYL8z1/LjPDRaH54WRw55gr
B4kDkLwPu5mygdZ8ztnva1/sNxTV9iBdaqa/Rdr8/PXuN8MwTDoS5zaoAuykyBivlIKnDlkX4/le
gB7xyulCwUePs67zzruHFt4DSZf8KO4fiV81ahVW9sTN0fvisFXEKu7It6Nwc6Ji48o6VVnVVcUy
XGmS6fy2B0IST83fnQiHH5VcEPMF8iIx4sCxGHQOV1nyDbXQ/KFTjQFgo05gq1rA/KFsGwY32L6p
gwuZsXgb2V0MxCpKnMnRCwR0WozW6FetDyaFiWK+csjP9FBJG3qma1srRPinFSG55RqpvDXcyKfs
z8XzTGUgeaSEk13lViNkk/7I5gm/uLBQE/gN9mdRPj1dvc2ov7Glp678xTutxGQcrKUiyYrr77hH
bKlCSYRWUnkVpimLuyINUOatNVnbbjmKmnkveQe4znAhCxTGBmMpRRyl5UcCvAqupJiG3ipOCZDX
VJS44QC4ECDihoM+NnHPoxOyw+9eGqYyUJo8J9In1lgbvcRhC/LPP2DrpJAAELfBO0pr68pcyeK2
tOe5Mn8xuTo6Ra9V2TwXBXlInLGGgMwcfeeaA0UOPidx6RSwXZ5fgFDiAxDOILQYCZqC1z9V390a
ycuoBYwfeZYnD5CtUqq9onVhFaIV0Ko1Yv5iAPhPBWwXRYtGvKgAFyrgIEOkSMhTYfFuKXdSKtGr
Bk3ypIUPuwl0d3IsoOD3TBgF4ltbyumKK3wyTBussaW+vsp2OOazEHX2bbgPv2u7W4a27UhIc5ho
8kBjnyawxhQH/yaiYgzBKQSHf+OBIlijne+QnM/WzO0M1FXEmQghT6CeMfXZ/T2SPtx37N9gn2DB
EoDTcD7zltK7FimjhHy6GW8hgvXdbmvyber7ZMnZBCmlHLLwRjZmJhvXmCTpwMSMuN7Hsjw5F2F4
toA4a78cGfA4/T5GJVIOoErhUiQOhsEQcWlBNeg8cavrKAhCMl1htFfsK7uqxYx3uoLORFIQ0Agw
F732IaYYNo3bdclF8qJWEOmZbbYw16VX0wG18rb/R9mIb9pjRSWpZz2etuCh6mXc+Nh+LqDue1kq
DhmeXJXR/RaEyaXOV+f7DzgKWdn/huLPWQxEnzk66LTZ/IR8W6qIYFTbYe+40ttIdTv1R42eh9NH
tUVGDDE2JQz7CIRCMHlJJJ2ckgdb+wqht3BY2tjRRyz3ms6s4fOp9oyO30psRmS1TuX74/2Z3dfy
R1yumsCoGMM1VWAGPdWH1dqvPaYbQpK7lJVq3WcUINoRcCcgJC+3lfvhH9cJtjYlNNj3z8WEsgZp
3kHfPgfRt1U73UialWBJ2TvssD/ysR7WG1xiPxisMyAdJexBLM8FKibY0WjehfFFsD7At2+SRRNO
EeOFdAe+Azis2kgoKWMngGU+w6D0L4EhHPTmvuCNFgEdX8u+DCKXKD4l7JNJnedF+fQN8nEVvUZj
QYqVhk2IsrFHQqyEeTZgtHu4HSPypo+vaeXWNC0j/eG2rsJvhDSmzuf1//r+tQwMLX0vHapnoX1u
xlndRq/rp8yFFrzkf3Ja00LcxjvY7wNQHI5Yu/rWw2aOaAe2VcIBIW6KlpUHvAmkDAvStL9Byiuk
/n2+hsoL6ibUMwgKo53q3gxAyUcY5bceErXm5uaqshWEdm4gS8GJcJxFqEzXmc9udE8GNOHOCWAK
2T2F5dFssz3BhzQNBMRd8vwD+gZTQsroTF6Didv5Kwy+SCdSunUdJqE6C4hZ/wca1rnqPMFMoiZh
HIyOtdJ2fyo7EaOhJpejaQpcBdPDA5M8PHOOHqqR+ruGBipabl0J4Jxgwcpyxvph6EpDJ3Cci4MY
ZHVlR2A7Z+FoGa0WEwn89+qYOTzP83x/6J+t1k0Wqpgl3ygQF5MFvA7nzfALUsJ8bozm+y6DVcfQ
6bBM2LFBHR6yB7Dl2NtX7zKgzszdCU06uJGxSw/dcC2kce0dapoGBhgcZBw2cpRyvuZhyG3jVk36
e+Rkqf428CxubE6SCUc3aiSVnF2oWFzk2kROd/orAzZ5sxdwZ5xtBEXR8vh4KgThTkUJtW4MYUwy
rBU204hJcf2vG310l3gZzpWR8vFviJlf3aRH17QcuPzFbUiNwX3OTC5QoFhJb3QnzhwDPP6f4LPe
a4W6Ph21DfWlE23PyECrt/fSXoFbLrwHaBTmPAzR6APnfmvaXLC4QJ6h/FU5BvzYDAI7cE1lPdd2
Ieq+ETBvj96vJ1KC/OtU2BBd62vT0tkbYxoZn9iGOzAr1zGIWNRJyymgEbZVCNvhN7Ukykzmhj9/
GUlz5MfhbjwQWFRwc8+gJyojYMQsPkhGDPUVv5fHVIT36gr+vx4ktiuUm1rd4ggcKlYQU/TrzRpF
nW1M4Gj5gx42Pjq9fkm5aPi1tVDg0NE9LW1PsR4raT50iXJrtU9TNixJZ37th76s0T6qkzliS0EZ
QqsMG083WcbGOIaW3cX06W2jlqfHjbVTQQ15QqnSz5c3ay5OP+XfB2eoLQQV8VOSxkuXbbJKVVW3
5Jn/DD15dHny/hMDal0kDEvl8bPGR6PeiBr6upfQZ+hcX8IqJkO6UPy7dmP4Ybwod+lA15nDz6p1
prT32KOI8J+VVyAL1YWf+U5xok51bjrRjAQ+xk+QPvaJ9+LaBLuZiO6dHhAfVu1awsOtnVT/JgyN
5QqQi28Kbzc5VkOUMLI4N96+FFnUGIcEBBFqHx9XQjjITY1LWLxvGsQhZUiOlblrKv2wmUXzYLJx
ayZnINoO42RqpQ5XT8vWY41AbSS+UmCuTGlKopfpwMIB9tAEgErDM9ftPV7kEbOAHU0uaVUKXLoM
oRQnjPv0P+WFH9HaAtExz4WGFtmvsSGaKQv2t+SwDrH0KIIsAucAaIwi4z0qgm7xbrFlhr18NRFf
2bqhk9iXVKkCmawRrK0BJbfm/xYnO1UHFfIgeTJrltWtUZGFZS5bcbCd4HV0huyxnQdQSFsF/oi5
28+u3Uq5v1Shr9uakMAMctNQMYRs6269+TNDJ0Igvwh1wLR0Bn/K9ipZsyW5RQ9UonG7hMNzu6K8
ctop4vqVDzX/fYjKnZoLd6oXXhO7Ba0HmKki1mbQwhdiQeSGp1OnnEFk/64yAy9EpZWCxaE7om8N
I24tXaozSr8lMEYkVbDM09GAmqQpEzTswpBFAnYDXLukas0yWfG6h7FBOhvrUQ/SCWhe0kBYQOD7
lylmhM11Mjetd9LP0LWUXAd8W1OykZYKBNxep55Qb5IY+tT6TKAoOtCorCjZVC+6RY9GKSfK6kZ9
AED4T8wAaLU/gfT9+fyDAvQ9XHCYv7ETim9os/wy6Xvl+EYe5e0odHniOx/gDV6mQa/mHhKz6OM+
h1aWnmSnO57iYxbRpFEaQICqDz1ON2xGe2haY6bYvtpJ8FvKuN/fP5q+RUQolAjh8Yj8Q5IFf/su
+JRfGErn1IDjivj6BhsotpaUD55IH+SHdqm8mNm1qo8WFtuhQeC7x+7ztv68uTKGtz7nU1f/Wuec
kGrvAcl/aAF9BR15cZEib+M0vSDecAkeyQY5m9Vz7vy2xnZpgeuErlFWYXcuJvB/THzFKaU7rAF+
f/XNjIW69WB+ojqOOyfzweG0+z2FV3u8nAJCzHJBHMmpqhMjr/5p+WYBzPi2DycJa+HuR5x0eeht
XyUST3ZcpzRpLhfbbJ7xHdx9KTXSPtBC29Ek6PdQ7320rSZQjgDaJjyFa3MaRTfniT19A6jfautu
AFp0aIOMiVQFHhAoyX3U+laBcXjO4uEDFsRPTlNdQTww56I6FI2Kd5lcys7ptapox/vK3NvrEq93
Py77JAfJRij9eQbiXim1lcKsxVWux4WtphNbSnxAf7RovPb6pKj4xM9KBA1TgbKTDuA+UvfarzLY
neUYIEES9JVnktDpA6fsHC15cAzm6wEuV1l1Pu0QDCWkNwTGsYEU4122Q0S9G72cUstyOMxamG1g
ux1a0twrR35RosdoXO8/jjX0EL3TIgP8GTsMaEvl9F7a9wwOMkn9unLZpzXq1hvmBcOVjxRGSzU/
WmgSsS1/wx54GVifH6wWW1tThD4bU9OVz8dOCkfotUV6l/hcKR6VHiFS6GcEuiWh9XBrK+q9/xms
uuJsLE6XykDe8l38FqWiRHPnGc+3f0a111/7xhGbXeGP1hZ6hp9NzES+Bup43Zmgjzqau7Dar8E9
BohCjZ7iN5+60awUtwOC3N+ZzszMiZR3FMlk18PqHPgSTY9QHrdAKR+1GetO8iub9GR+c1vTLvMX
Xmz4N3u1vSWsYVX9r8W/JKohxazSe35Zi1mytTZcJMZO1x3A6RYx0fvlzXh5+iEIkt/v9E2u7Rh6
Zv0lcdf3dbE8yttOhrYIj0OTfx67EkQ3ABzNwbjsLgUcj09HnwH0m3QWxjzL+qynU3xZTIVK/2oZ
Ti+9s0sOm0OtNpky8Gm076/kLv1jl9QuiH/tIY+INd1E6c46g04BpwpvwSfYffp4kQwKnm2wUr/H
1iLcHo/IFpBE64ckZvnVmUL29W3SWrtinU85OBBRMg8+e/OZsl9OF3TWUomnNscVonxQVW0cxfgf
eEPSBnBLLsSY7bjtrEZypiZAya+7hrwg6C/kfRqZuYdsKJhIydbjEuVvVEfqGZeQd8UJ7MKGhq8D
FoxBNu7QWb2DqBin2jNkVdrhJS69o7u/FYW8QYBbyNvzfonrPRGjxiG6lNCG+upbufAqZazBAFgM
YkG/oPSBPYu1f2XKKhNFTErhBEZZ9mBKppqRHlS1nvbFB7S7NteouvuCj++yyH9zkJgVObP9y5Ii
Yk2duNhbZoh3HjQQKz4d6uwRPNC+A4Nj+8CJIJX+zytko9qQt3FVlYKbK6gm8yf29C1lcQHpLTlM
+2ENPPfKTPcXRJvPAQGNA5jMTPwEwTqbm7eHMpSYQew23f/l0yio6PtPctl0VE/TrTJ8SkeLDJh5
rFJt6qrj1qkdyCJZbhS9EqoJxv0h1IXaVCnhxluV8QS2mGL1d8CORRNM5JOlQixezfTpqgt9NzyT
xWhlYPjA9bBlwdGEkuE+w9uKeFF16B9qxTrE+JtDWYWFSqY09aMv/xoVA1YBxrl+3Rq0kYa+N4Q2
CRzIz/WL/Cdor7YKrtL8VvkCH9vZiOvm0ZaD0loiEIxCPptQaX7J7kV2VlgHDSQQZiainpDe1X6s
JtIGAG2cBrb0rnN1c894oZj0n2b2shmYh4w1IGvBcoYaR3kuOl5ItrQ/+dH7m0Lh9GgBM9YlifOo
vH0hTZhZgKmW5AVo7SSX+yPqfK/NtS7IfrSBe9m2noTvX+Wd8IwkyfyshbAy9ZlnkhAi+8kU1Rcz
LW3DM89eA9W540bek+mCbXiyO2UHn2zTSKnHdhAT/Rq/Yj1ntYl8E+MCcKbUAXm3bW2UY7fNK4L6
ji6GAR6OWsOjhluGwpMttbnFBulWEICq6p01MAcFWcoN40i5E6ytcqYBsMEL6JoXbiSoqZNelKiB
knPQHwECbQsk0UP4HqzYgWJraCgiGhYN1pP1xeLWYx4ZarSQQoSct653Y8YyIYuXm6iP+90UwrW8
C527tQ0AwLaX0+PoLWbes8KlxsfRHW03ekmNBAN88DRa1U0XHjKT72t+ieh7cJR2mIiw2t6PPOCw
La7GKWp/2J56NCWn1SMTkUn7L9lbuGTssElxPKF9qH7R8JI/pTzgohi2g7JfO5pwJnu/wShYutUz
0Li8kU+Jd3b/juFkstZsb99o6gRei8gjf1Bp+K8U4a5F5t08ov/0dZvZjnNxTvZWiXyRm4IrE1qw
p5f1L2ABHeDciWP/3PbaAfIQ7CUhuOpDfSpwrKTujBerDo74AsY+GAoYJJf6q25YWzlkL07Q+9Js
+1DBC0lxw7j63OxLjp9WL+XDkpvAbvoJJyKdiPcdIwYupG2NoWQjrJBn4aNxoebjs1F3K4B/vdRq
QSpRTF7Xc2PQyW0VSg8nuy9uJmbE7qqbTFo8kPvy45VURqvI3T8NTdvSHvW4HW5jt2SOezdiTOt/
v4Q5cQBj2Hk5NF2neAQDS/ec2DFTR96T2irHG41jC+cNXCSh2bJFHINpEMaXKh02CNYOWT6Qmby6
7hPo25GUCWs1Io8HqqixEzkfp49mV2YaFvU+aEZmusa2mMkVYqkP0xbP4L8e80ir4j/DNdy4586m
IZnJWLSQgytVzjW33M0r2aBVq6l2ws2oQLeO51deDn+aOwo5OZTrLZGIlpRrNc/92BMubA2whnJ8
QtfBWq3Y/8FoH+hY85/MRi6NxixXK05UXey/PapqDmPlK51MQAXeYZ+BCydUjSwXJU/FtBJXqMyQ
ua93peH9DWDBr+mcdGhV6nkKB3HwYqrbAbdztRmF2gRZaA24taNuc75cSd+ytSeBv2xjL9kzShfU
nX/BxMthOvIwSwLUvX45zhAp283bISVPmNFqZYLyYybJ7zgUQeUTeWbq0vbI7koHLndMCORaQcsS
V5qtPtCioWs8aniXMeT2TkAig0Lrh2WQSC5C0xTeUsAZnBFA189/wIHW6fGJ/V/KZMD7IRveu2KB
yLT8V6eGoR+a/p7/rlTI2ca4sMae0lW0WD0Jmlu9zAodvHjJMnxvt1qlUGKEJgdA78faHpHuaoSG
vwJ96EbphkMcml83A76LQ6DeY3dOJrrbtUr4oRnRT9p6Z8oWDKfxIlNtkGBCH6xWTgIxWtKvZkn8
xqjy9uZ3noQQ7Rckx/Ed97wwT4Q2QFcvDNDgBBWufngqac9UplJRgfR6wzC7LRNbWOVz6olhvBYd
76hiWXDpdBgTEW+Jpwfeww4W3Wu+rddfe7GD+xVrHvQYnuz6b3H9GQvp50F/A/i/ZFH/oC/EwR4w
r2WgdFOTJ62bCYLOvQxMWLDZ/3v7emVbra2AuhkzRzFajsO/WpgAx4XSsEWO2o13eXvxjwKMZqRa
wwmPhVAbORo3OMksjD7yBSbbtu5fKUZAO4LGUPGmGwkoZMk+OcC50/1H9mahdV+4TNhSvnguw5Ls
aNInZzupcHOCORCCTo7JKASViBj31efDszZaZN2G4qpb379FpP/64FabZemXab4d8u5xUuBJLYk1
QQAe42EXbj8VsH/gj7CaXYgllquUcG3WevcLL9e8I4WMkY+BrjpC+bk+Vc10/b1p162LZ7k7H6Qa
o+hKjRMoYW+S3JKFZFP2vZ9cOH+2BoGsfT0RF/UrSpM5HdM+gBvGFStDfL1RavdYMzwNfwK0kT2A
rUniSAsFmTsiFNkZmd8IxS8Q4uLH5A5DTI3DnsfGBNQhdQx2Mu7g4EPAcopRpOj/pxHYAoWF6FtE
FPh0f16cp7NGw6c7PZxXAC9mByvFtMfIibNan54qD4PY82+4C7+wUw2urti8YpoeC1n/A/q25nb+
+cswXa78uyko8EyFIBHMqSXle4vl5RirWp9DX/TNpbbwE0nRIoPtJbqDL57LVyxe4GISJyopGOG9
IUcIBvN3mhi5pQeTY6NcgeWQLZ6tIHCCVXYcwPBQM8H0aQcwDUXl1R/znGMUEB+JZ2ngYE2Ns8Ir
6tUTUTk41zsER0UqLh2XsUEeZAIrM59wd5L+lTeTnVyDICcBNigdT3cJ9hgGvRiJ4XHFCeCrFbhJ
RL9bWjPvz7cabglfDIEQsehZClyMX+Us4+3lWxEW5n39ThFZ4S7Q8nNY01/BYUAx4NHclwPwSDLr
SVs1xYfk2JcrcuYtHSQbmOzB4HU+aztVrvRHSu8i1j0gmr4sBd45WymREtzrRnULTGJmGeyz99Ta
urov+oyHMiL6nKHJ4a46ANP+qCH2/CYaqEDxuzKYwpODvXVheOyvwqsz+A6oYbIFSvlESbkEPv/J
K1L+9JhIqs1lbjjzzs2pTe+mhP/Rz5915HU6vwWcjW8Qk0KZgnU4+JLnunv4WaqGx62qrjB/p7V7
tdOciOEvSqWwHNivis00f3NJzcxscUyxQC5FaRbrmZkSxqvGaPPEcfELb5NfJDmN8VAih+B9sTSD
O6wIv5LR5bEy066mVOZuAFHZw5SkpCQtPKLZ9IkC7YgqCo2XEnLHn9ifB/bqVj0+qc7qJ0oTPI6Y
vpws6GNVlC8V9+XKeCmDsr2w9gFbHtMJaugZyJz9XP9REcBjxgpo4TnwC+rVlKt56RuyR+H3SxGl
VI2lNA3jk80dTFICaHYDYUnAsYOvP5RnGzychbInWopYSmi9xaQ22j36HpSVE/DP6COEnwxW5B1Q
eRXiTlfpHyBWIeUcj6+AODau18xd1THAJRP4XDH6WySyOS4EwDmy4dwVK+/M6ZyMd/IJ36XYRQAf
UyHUMBG/dhwuPvKNAO64Gqei2iAn6QHtDK1wCIgiRxmiDkhwwjuvYBbHjSc7ETeW4HrGmuqgOHzV
ZWmFpabNElSwDmZHtPVb3xrUn+IMHA/8cyM3pUKy+tr0cAYSG5mI9lu8Bv6O73GpNT4uN7jlE725
abd0SZgn3f4Vz+Pt/n0xlt0/dpsV2WDYL5vNp3AehPU5A2bRJKsWlIxJs/3rPfrbi3AlUGXidYWe
rn0Ny8Uy0mu07brMYQ7pk9StsQi93Dje4+rdDLOxMPRDI+cQtOSpz9j8O9wEAs1BWie+tSQLMFH0
+7lh1h45vP8VL2xnwJkdOlrirbeTdC5pDXofdsE/9yMgSQxWg73edxIP7n7/i7HEjEi70L8qipt/
gokNsYBPXuZyQfZaOEgSnFnjqvlTKTTn23pQBJPa5ejaiQn9sKviqG1j51gIOqA3ozBI2xeBDX38
9GlkNM8tci656P4BlgcIytteSRS53VCMmAnUN0I7XwqA0FxUBgJG/bxYeZLr8XXWvBEVRfSrjT/P
K2Zcbnfu+cQepJgvDI/gZy++hpdxCVYqRBuxEkUSh8Xy1kRIkTn2ufCgLYSBIL/+oJFwG7X9MZ56
Uwrr6dUcT2iDpjnlk9gvy+jGMgURyboj0XIR4FNMl2eChrVODJzKyxLWiMWbl0Jf8EZU8m+MgV4P
45IrNy3Gt4iLSZJvTwLV6ZFDq+EGdANn2VewUnPoTvHr2flDHcAWY2E8ZeYb3uZi5DyrdN2cySi+
PzIPwnKzkTCxZHno974N7tpyGw12bSKzBhN1hEgczw6OftBOlvc3eAkMuhKOKyAvwdJ6uXiEt46K
csOTFqrTqiJM9KEzXFCX5YGoYAJ7HQ7kxtoIYbL4zmsspHhuILktpvdnx1CUxAcVxrMeRXsNbXxO
aTM9/aEZJDNaaxaLJPflV2KgMOVcukE2mfXG4Cpvjpy/eTfKq+hqmqUtYrIhNljqDkdSz61o30ts
9xZ8vyrpVtnczjrv4hLZ7sGv2zeB4nu9t4zg1IELsnCe7uc4537Yh0Zqo+O/bXLbC3zkHs5kz71l
4gWJjGcH3qJlZ4+EuQKyCMazrvIvQGRS1RhE+Kx/ygZqzqauGcPDnVT4kIWgTxjKb/l+wrgfxG9v
v6VeCV7cxeC2/+gaqbTtTcXr5zQUCvjuss2lq1luROdpkqS9eta9QqKZID3gVcF+EO2hp3UPfZd6
/U8NXWPQ4WhyT1eKxnWG1L1nnd78VCJ60oF95IfKvfO35iNIryzE3EVrbTp/fiwtZo6OslCUl/KI
O2U2guZvguk0resCZSkaCkY4fvdbKordNVVjq45QLmgMV/9MdLZ6DF7o68ywglZZhhWRG0NQsoHx
wyG7Jq2ltgQUCzY/QsbLe4reFw5MjLeFrJGWTxGi0lps4QDm3LFLXvHQneaqK5BlmWGxahcdrIOY
nxuO+id3pibeEJLal57Xnqdqrj6NU6PjXsmI9IjUFG8GoJA2bpLUVKwk2/jzp52dOpb0O5YOGTcF
B3eSjmSNgZJtXt6u2CN1YzLdKwK/VRX0OZKrotB7ILAaYVOOcsnQU+GikS/r8Yt3B6Hl1G0aSLqV
MdsCK3Eo+mckm3fEsSqpiMdxKQwuOtNEgVlQLj1Fdgk/c3AlDB1JUNWTV9bMJEhEweEKl1/Syr4W
hbKJkrZCRhx5A6EqtO0A4zHLik8vQZefdnaTMFoz8BoZFCLSeKdUkLWvs8EAi7nV8HCshKKoKtHn
1/WQq+jAoYkpepwj53rbciu1Mhh0dUBI+IB8AlT1t0nBX5sHxQPgQA+0vktPR1zZFqbSZy00Hd7Y
SP+xytwJtSjmh5Rxs6kcPolVZzbH02b5+Ud9V6oKqQg/wHO6790pXirgQ0zvC5rOeYz2d/nXl5Lo
DEYURqiVdz/PSe8N2fNGhYtaxNJm+iMCh4SIKGNMsS/0kB2bwLLeTGbROuDUfWtk4rlEgG5L9nnQ
a38mrnT+bRa/99nogjFWv6uoBDMDg/iLrmSu06cPfDrJalWEtEdGkqKhqQAoWkcnqwC+ejfNY5yt
8VTUwGBO7257aLInILnsqjFZKJJ/DQ1LSutMxNC8H8+/53V79x2J4pZFlvEou4hC6f9vi6nEcYV7
Z3BnFfVNaXowBPqMqmRu7HtiX4GzGDZV+eTCD8BtIP2YL1P1L2hm8kEneHp3zIX6s0Sr+Ix0HZgp
P0uDa11GYgGejdUhhGdoZO1wvEpjEG92Hx1bA0bBny+6hOgCZEhLpZ2EGCY0vysry6MxwqWarXWY
YzBXzcnx8yZyyIpdkDtTMNHs9ka0l909glGvXSNi9lyB/8iKXDzBrHEFwF2TzPm6oftva1AWjBhg
2yW/cXM2LNspo7K1PHx8aqIm6X7OJYxtm79oCpQXjUURv444MONvNbrDtGBnN92BFScu3VtqUjz/
7hOuGyCkcGqSEU2VSBA2ZZgvQM9SGPjVeAyEEVMcBo1U2fxaoCL28oUtmWke1PecTPqvF798BwS8
lXe4cOb65TOmZ1CF6lXm6a1Hp45S12ep7jihslgwFcoNfNxTioexwvpEWvDgJMGzJmO1z7T8utKK
ZZrA2VW8R68qLABet2EAIRFGTSkjUgXCJp94NVt6O6PmoNq2520x1Di9gKjafZYJlVY+p/ZB2vhO
aaB/uz56HOOiUl5UVObXK/rIYlkYj5FoomIisC3xwqvGaQakd3AtZ8PmX/CTjsjMULlfdduP5WoW
c2BRyPjTFVPCu42rYemjl/WnvYHNyqwo2KddMW26SpUP0F7p7Y46+QWTEqG9dlWXo/SAMIh4YweS
CfIFLFvE7iyaE4qAk8R2cZRoW0cLdMId/OFQS47d3U+ayfKKwjyDetwnljTsR/6+26CRFX/WZIRt
WFx7Z1k2lN9nFZNHvRKl2xX7xRttAbPwC+12Bme9huiJIg3KMbWbJx2EL48pgXd2NjgiAXFMe9Fb
ZhCjRwPu+Y29Edvg8/qsk7hM6cXLjeoX2YSRRECyTARdgdTyg8mg18FM85eu+zNVAnlonmVQIPzz
BUJpgysnx/gRGuH09Uup9U4jypC/DYvCMAvynapsARUiTRzGQJD04zAX0a/pt/MngZrqcc2NrRXI
hTRbPnSIH91VIrRm12SuKziaYNqoo5hMApQlSau3Z/gQp2IgXqNuYHHaETm8eMxOvhpGgmNb/65a
FToe/s/UCF8Pn0n5NMEZ+QSRyatEopI+EBf9bxuOkO+H8I9ysUwGYU2saEActgtWjaRyCC77IrcZ
eh48+liiXccdqUsAOHWkA9o/OKNdAavqJLg8GTPDpS4cVzDJMfNFWJycJHA3En6dLMRKH7fsdirC
9lfA3ELiz85JtiQwGpa6kdzpIYbKTT7egQHy/D28exBtRrLcqlo/UK0KmwZc7YMmR2fC9H/EjrM6
Wl13av5Jk+5VOYdJmYaZzo7tBw2wSXQ37hmOXb8Ckv8BzlWL9KKLWpinW7O5HclGpx2nGSlh4Ph+
ixKnKE8ysOt6fTIw4YSLj13GZlX+LxPBynYKzmQwuKLLrp8Ew4Y5F+30zxAVrwZDw7g3I/Z+XyUK
mw6cZpiqk9mCX3FEYcyqFb3fMc8TdikTdER7a4zxec3uBOZHcxapZ2fpqBtlNYEm0ktcf9d6Q2fe
4IqUa18nyw1wdp5yvU2FWhkyO2mpv9NpLle3n867gbrPUslY6zUynr2nNoe2UhMc2Ji+/ocjzO6n
1jAnwJu16RFPrS8HIjE7E4cQbudHEDqK69A5Ta4b/KLr5uOvs9kQnxd/ddz/qJhwft8nKSgKKptY
wRDdPzrFZ1dTDjgLB9D8x9BDdvpi2NBASMYdpsuuxD2Gk46ZQot5tlkN8MMgzEBne1Lz4a+WPkmB
jb87iNGQ39vCn85dVxklQrQ46MKyBqc2tufOkyrQfuCK7mo6ksQ5h65afxqi9YwKdlHoukyXkfWy
VNogB5yumKnOuvYk+XDV2q4DuI4NIuCKiP/Vx7nL11KH7bd5g7kMPd/BRcNGeysKOLx1HHkrzj+r
sg0pXR4+/F0qmMwg1hOFOtHC5DCWYX8qknS+sUEyf6qS8lkjJuXiMS/H1y2WgZDHqSfY7ZOHI+3z
D2sp8YpC9yeSrmVEN70ygg7uzPJ3cCDGe6erUMovZ3OhSarp+JeYCDF3psQM23YMDawlB39GgAG5
2+6AuohKcAqZK1IAN+dPp5EULero+6doFh1POLIDd8tibsNXNAPzHzTRUjv5WWuB7BhxdtZtBty2
/8AIvyCf0lpOWvDPqhAf7lk9V56lbNSoEvadb2T4Nk3yklwe7n7hh625B4S8S136JFoIRjxXJyak
23ArAughrtQymnZWUKTGEtj6Ll56byMdOOsiOPtIC1pyj4vnEi8RqZsK6Udp3sAphnKOaE1ZzcHL
Hcc6W2XBk8nf3JHHJbqooRou0YthQAt45AtoIoCnnptIAYJTA3n5OTFZamIsf5/b4nyiuCDcYK7F
UAa2kU9+89fCje+Ak2VYXS+yo7z5oBZyrjdqBhtzI4ZryNb5LTj+Nc0A/l1ZPXAiDN1hlfpZEuB4
vpxB6hwE98y1BCSalfMCbSs63ciZPiZYnp2htN+k7xnJnA3kNBuTWOFK4mjAv5eerSM4UvuFM7mm
9TBh4MC36GLcDhUkwtHV6+wZ0b+ycjdCEIGiW2+MFnQfNEr9lG6uFlhTisLaVVbS60k++P79owNU
9PGsfL4cnxlontIn1XHwolTzkrC8r8dzo9TbshivNM9x/15Kdd7zr2PojPRe6jZMq+A5Vv0nplBr
u5Lp6lCWBvWwkQR0nBG6kGCaK02POcshQxzIaY4WCJepMvYjycdX31/9YO3RwwNfYVTdlNIbkc6C
8Bg2c2duKCZzUVBB3FzCgao4JJCWAsGGgI/cYP22EXN6s7olB19gB3u4QvCxFIa3Mj9Y3pRsH1IY
2dAB89uQIc0Y26cHjcSpqU4mkqUDF/l45EjuJwXY3QiLz9dXAFPENhJwNK4qvt0DCoF0rfQ1qcIn
55v4000MnjOyFbfSklge3UbZIfKHIpPXAPNI+U0OqR6t03hUi2WGZMKFE7RfUQ3jcR/K1QsWEZkZ
q8HBB0WKUGo+6aAbIUcJh18k3FnOkDUJEf5kv+hEwr9dUo3lwAP4y+4zB7EB5EgucEujDHEPrKIb
BNd2uwEDqW2eBAetvx6ZpXVCcVRD+BrkBpAaAmNB7ddK1TQZYN/UWgWtuM1EPEUACGmzLH5G3Qln
qmkB+qmegQEV8dxuh7U+QaBypLOexzMKYKCMNgRqmrTcoxqrx9TRFgJt1edDHMnvPsilaLVmR2Up
fGQpolkVxcEXv0/z/7FKP/2t2XbYiSzJn0sNTi/aWygnttJpkI863Y+DOnVyiLeLwL9Km8zfXsZ9
hbcimz6bdrpMO+jY/WLyoOdQFJws/fCiqfzBu5qaeS4jXcMTCRIB2GX8FIJdol+cxj5FX0Cycewl
4EE5sLPgCcKmVHGHFq7oPIy+vX8H3P3V72J1nuadJ7R+QjShuzERAwm4r/FKCVZOpG5f2iAzgoge
+rNmtv+KwMr9V65fR5sbw+/j33aMf6pn1CGfofOhZh8K7HAZ8Q5npaz5jqhgYQXGGF2ZzS0YSr8l
xilXQBunAD9eCw3M1S57JtshcIkx6KQalmSYbkCB/n6XeteT1FeT5DSU6jXEZMPUyDav58YXWgkV
esj9+k6PdsLAmiNrVDDcfE7pjimd1kKE95QaUSZFM7qe1RiC562r1FFsedrXXs5XVtBB9vAmfyEd
GBzhKgePH2X+0460O0jOJ4CFu6Dg0e4mS2TbEKLG9MwWR7f5405T/ExQCARPYwWIPEOH6BGRjCmV
Y6VcdK5OanHjnZZVwmz4CkCcB4gV/1M4Y52IGFzrrr4Rb1MABbjeNtVgBFMSHxvW4UyeedrH5ON5
F6dJVcoCWohJDptj9gSgHTz0e4xAahZ0EYIObgFYTjVfvwmYmtKaQjraF5bRoq8F6dgP5BpnM57R
dhoanUUdHn/Xmi4yTu6aXbhnc8m5F3GhfeZzmcqO9JFi4P9GCU7v15Tc+BMPAwWEboB76WGYDOV8
SJjDuzMde5xJH1BDepEccsZ9D5hYyKx/xE5sqf4MxFQroFS6f3ggZ8fJob5BikNcWvctV9Xnzr5x
6qnp3ndFwIhRSu/A1PF6pTnr7Mvh4yAuppbxzl8OTqyRU+41no6zN/v8nBY85WRzlji578CPB4L5
7GePSSVPoVDJYuRSJQtD41FL+pr05Wqlv8CmOAonMGm87Se652+APwIwyu7khE85rpH/0wbvvMuC
BnTtXdjFW8WO3jMT6YQIvR0zAdPhCBDojdKf1IEUU8lgs+824ROEGKqalfwsF+HgmtsT1TEjsQ8B
R8m8pmG/+UFz6NcQahywK8xd3HOPJ/Y4/YE4RDPfDC1/kBoNFdfd4/XUz8QS5mAJFYIO5h1Q7h4t
p2tPGsq89J/o6NXGfD2VbyKzPcYYxsJsAnMJMgA1zIDdUpmjQ1CEsKuuTeF4w1T4BsHxDwRcctO4
hGIa8rAAKgFT61Au9NM4D6X+hhaaro4VUjgC0d/TT8RhYnG8E3QID2JB5izMTlrXHKDk/ol1Shrs
l5IkI0+dPNVNmkDwhgCAUfVV7/H3CObLm4IxgARTv0+csUjexwnIUfSanEyGHdmIHYyG0MqqUSMB
yQSM3b90I4OO8749+CdzRneE/Ltw0blUpnTSOsVXg/S0ErNAiAFfXRbQFtMxT//DsjL8chicKguD
vaCHUWazfHyQJXOr3qjh3Vm5/7Y8feiKzsQkk8UKWkuxGMq7VWT4D3b6Qg0JRWDrY6p2c9AL0Dp2
JQHVltwb5tQO7fpjBPcPaoAT2wR+Nm/DLAYkqFhL31eaNb6uXcolleQuUyCB+AaO9zMSPsap+Yx3
Wrtgq7ROLXGhhvh6Nj2cEYFDrnyGdjBM0HnTD/cWz1ikYg91yn3hXOQd2CdcQr/mMGHSH6J3l2Cs
HlUR4VrBB1Qy00zHWXKN9zGdQ7dVGJcnxfkjvhGa5im699vS4YuwuqH4vvScuEmxJj3o/7t86X1P
prKWZFGujdHq6Lcqd2Q9Kl5oLiAnxqJ7cvwc4FiKxYtb2M5q7HjViQHUoshQXrFkDOYb2edmPih3
4ZS/ecdpvhjHLf+9eTJCw8evvEMlSSNkelkESDmK07f8i2HYLfcIjHm/ycYyWtyMpsBHfFiqIohr
teVIA2S3jVRAkFu2LLA96QNOmmv3BmMkSQWEdFYj0A7XAQxzFQ79DXIYHXuBX1asoiUzd+9kWbkp
jKNa0ji6WfYEZ3UgdVMigLb5PT+D5sojJZv/k6x9g5J8VbHHnTIZbCONGMVUJVsnYXSFuVa1cmLT
0NFPDc08xfd5gMSwSPqUssSohq5fl3VxaccwNYKzMWZkOxavDBIziC+37pgIn4qkORjCv8kSTiVN
wrLK8EVG9vrGuKoI+1x2zNY6bpqvUYZ/QGcSMHzR+Oe8beqsfedBYlVgEiLTCLX6RS1sARcUne4a
yxZIslAsRVQuZFty1e8l5CxTzm75chJAKR2iKzEuBU/XOzYQJ8aY4LtY4RWpbElv6zoLUWVwJUHa
PwDWLyCbeZgkQw9CCUKmpwW9lr7zud4vjyfSZwt2AcoUjl/qdcCQNWLW733aQKAe6/rkgEcV5jeg
hK+lLT974cTGsbbsuftOqD6dRy07TaT1NTfq0aU13AtVjD+zclqff7eA3OtWrqTa1psNgGAF6lYF
Qrwu5yT78FIraElsQwoQWITs4q34efogp0INxMBE79wMxnO3OpmyBGg88NOLZ4o7htpoN1bSuaL+
riieB0K7xX/uDZsujc4LM3kaJBtVaugBZgPHBGXO9rdVGa0xs9EjcKqBUbVktiLFxIVw+jxvM51g
FZ3Nr8DAEqWkqF07YpcrjT+L3KJOB1+hefuFrIAsGGKuwT5yEWljdIeUV6AylBwAsbWLIvsj4PTY
R5byzt0mDayl5WIWIp6k2VFeQmCwcZ41GC7mL02VX8fxGHT2Ybhyi9EEHNCKd8AANPx0NufcRqwx
PDKUN8qLkN9wI8RRLc9CjR3EjdAi06uGzndXsWhJqL+mh8NHrof6aMZ+bM6+E+scaS4CpHZAp1a8
oZoPMczpvQHGjtRdVi50lx3Rhq6QvpK/b5/jVQpOSCRjvy7sEBO/MGMn6UPX75p3S0wV881FY2PV
RU2efwrbjP3aou5Ey9Eiy9kc8pew+H9hXP/OP8uPTj/Jy5IVQh7ZiYpqM/F2320wHS8VXE927FSE
uvR97Z3HXQiRFCVuJy+ceASQ2q6vx3y7tl9oH1KHe0SVmCG7KClfEBwSiqiV0dswDpdJ4W40xOMS
vloW8pJEhvd/SZ+f8o2KSZMtAhl+DjqTbUDDkizItKGbeZSTcF042NWcjsQiVLitaVVJGO6wMkEB
Y8wUov2GG0JbRe+dmQeE8Dk/Z3x2TQkVt0iaR7oHMApKjBF2Xqg9CFCFKYMu9pbIhi2EV7yWLzM3
I4I47NrXZK1t2aBNUpCL5E6fpcalV6sN4+lwoX9FXga08s0LmuL/Ixl8VXE+A9FJZaQg9pAospSO
wAwhcAeZwbYbtiFSmxiAVrY78B8filkktCL0KOsFso4dGhZXO1E0cP7UKs3SFzLcVKkw9GRUjy0Y
5BRYd388Yi5uU0eD2RG76cO7h4DDY1Dph/tRltiDZ2j/zvLO70zLvWQ+WNGKNq6dLjuxLpfhDDDc
C7kb9IrZ533Xi4neWNWgIyX+rVXYoEZsMUIGsNYCWCEYGFIuD7Foxs5NizYxldZiGuZSF2UEgM9k
LiU8VrJJY7vIRdOOkvAmNmpx66Qoa4D0MPJSNvzme2YI28+HmZ0pz863JeRs1U2HUwGT7TIN8T95
9gO58vs0mAhsW33NFAFHsfLFoCdenzryj2nmqjXVXWmbyQRkKq82U1Ga78zTJMGBAv8sqO1NWa/c
9uR7IKr5xQbWJlGnMfRKZkmWPFW762BJw0ghHyz2YXt2G5+5C3Ce1FEibPsldpb++QNrGMaaXYAp
Z23IwDCKH0/9lekSEu55k2RA2L1o1lBjmKO7URAqSlAC+o6xNjpUR0617UTwypRiETw/ZXAOrNGh
IRA7ecK6EECKfNQ/4sB1qGzfZ68ZOhwcbfHeVWKKsoS7E0eHuEjChf83CDnggLLg8FIioEpp95db
iP/AGzy80ai4NkJTNGF8aXJBrN0imOGNV/fWFncQuPgdtwFPYjaNeP/glLum6tx2Gm37SSypFfzq
JEP3DoBg24BoSChCLiEEeXjBFSyS+FC7wwbfXn+dfAh0mfwWbKCynFJBmijOblmc49N8VBjy17Gx
YOgusbBQx+fwaeQ4+SKUjgLqetKqhlvad5TlO/FIY+qq4Qev39Wv8XibOqKdDKj/wjYKCPK7QFgz
czgI22RrR34bNc6glcdN8GJo1tvroAHnFMHr2bqHBAKFJW9lfbU0Btjqai3GatuBylqqf/Ngg5d5
ZYog8ghLS1GyNzUDaacJu52QypOOhY8hi7Q0bzkX71PahmPU9pRxXz6Tg77kbhy9qOiw7wal2HXe
z8qbeTMyEiB2YTNA/7399hCnLwngIgN3lC+zV/xCDSaH1yg7GK47gOFwN4ELcTn7ip3UOABW/yIW
gqqJzFdtGQ+kmSibTUOC56VCXfrELRseDFiqOVRdCQY0Fyt/aC/y/lPl0nxjK8pe0SAOObg262ED
KusxqHD1TOFusf3VMZsHlWv4IXJR/t+6TjTF7izw7oMKH6l7VqZT6g9E5FGHLQSzL9jYO+dJHDIa
EEeb+EWLNpzadvZfv80ZJjZRliNrobd1Xb02SO/1Y3E3laCJK47BMsa8hxH/yWQUEtBX9oOovmC3
mmv5w+zt+bIDZfaemFM8r9QI14LBB7nH8VPbbtIP6Wu79GZtO5WB0TIBWdmAd2lvalXFRuPKEIGj
V6L29NhXt1m8MuPwQXDj6XsX9z2N7qvEoOZEExS0dNS0mM1j0j+xGTL4p7vCa+tsjfAIWOEdpCwd
lbVleS5CTPUAK0+RfRmRwOqHlh36JuyvkopZSoHfsfNm3pVqao9sHKOKeo4d4TjdfOaboaLsmqWd
kILrMI0Br/YI46P4D42BCP9fj4KuCnb9ovHZ56w+4WleuV1W8MQUuKe5LzaHDjP6pwovjwnBV6NJ
R4n7KZ2DsmIdvHtqGxyWZpqW8pShC+u2FJNExbEcQ7zipyMJJfmTuvE8FUQkEaU5ZcoO3fb901I0
eIyhxzFPQCKY+FgCK1hDwmjpOKJg0DXPpv5LbrABAROAxsFJmkwmLOj3nIoulvPwtlVAAh2CRwUs
ZDWTf5/bEsL3/ghRI0Hy5LFd0dqXGxb0fMsi6IJFni335b4NthLnm1mjyR2QjHiRpQSrEeEj9CLU
qDwmYRYyZwpecQPLhb94OGnFP2bKvt0jkObyrYKd7D2UHaIf4dl2OxyB0Cd5BwwXKsoQktRSPTxU
QugZVPDk+I5PqXKbWtLz07uQU9w37bjRhKF4O5u9AGe4z4hOIVgqres87DA/Q0LIYKHAdcTMR9hU
CrfsynsJgx7lHH43SlrcmNyKegcTd1yNRcKQ10f606kJKij8cDEeEsyRIrO21llqAJL2GP2NVwPZ
qZlrULUDt+01Qudps87KNGEbTjGlG3cWuc8D+mI4+Rs/DXA4jdBtjY8ZKLh6gr3gwhQClbF5YBGK
lJ5bqK7dtmQZe93ZCMzq3hslrZB4AlMo1yZuR0+0Kgl2ptXrb0y50FDpCxRllOFgRkT4y/MXKFEz
jCv6OgFdxObNR28liBIT5txUd+zTlFFN/8hF3kDBT6X/cABeGqdltamIXfIh/2X0/uFT8bNlLdfS
Yxbtz4S/NBCPX519kiR4yCxMlTbwQ2wQIdUeFfpxnw2LB1UInK9uhCXYeYR9E7FZ4hoeFoP3xj2Q
2NxFvNMCQLvk45tDoSDsPutECX8N6F41h1VwOost2BqF70gvHD8RdLj+mr/dWHX7TcmJ1QJBO89Z
zVaI3bdL4t59juKvltLNHp0hBdcD87G0yLUynJ5nWjx+I+j1sbEa1ZGIacVlRLW9k9FyDLUHE224
B8XFaRL6T4fmVlcMUiDojgT2IaxACtpbJ7TTh+vDjUJab+dsZ331VCduBYbiW9bzLWFoMj9Bq10W
r8nkUTo7v6847WsBNPsoFH23CXgBDKEeLZPFNa2MIqjTxRywcmbAwtDzWhTH8R4dG9HUBDgCbCqg
7PxRVwiZatOK+1LDVwjFrjV/xQRhxg8HtjL81h+fZNCoVlmYvjdf3or4MeJ55+05hhGlMoR3EAv5
XpaNQgQ8bo+kPAYD09SNXr/OyZsZIdF7EzAbMHvsCk5qH1hA7Zk7QuNEkRYVZVsMjCy9IAJECpOG
KCOsyHsGPdinGMZ43XUui6AGzwdbO+DxH3Aeiyw1ihCokOQ28q7oc2rOh4DCMD43B8M3xEby3ukG
hNGgVXLpn9w11a/3hbFFAW5vIP6U1+N/qknu7byzNDsX49BMD56yKnCuL8b7gJAzewYqj5aTVJhg
8wQ4A3jw+hEZG6nzXop9Y3u1HFBWvdtOp/+0erDp/pe6qennDlLa7/+EUQk/kNqRBYEBLnskzHqs
pMJrd7hXyvwusTTv1RKErB1DE4T+lz0+EfkeM6xqFY0nH42rtLFzEFwqn63mjEOjhcTJ/FLwd7Mk
jU+CMK0bIHxJAcXAYnm6M3Pxg4k/6jZjGMNgL06/wouvBLm6qnhXKEvbiD07xCjZSTymBUv6mCzy
l19HrRcPmMc48H6ZiOs/me9UgBNe8TXuZ7RMYhLQoGdX2wKaFTahmQtbD2oJpUwXvS0BFTgm6GPt
lLjT0E6wmUNGHl9Rym+WVqx1ehqicKYn051/0rW3a7Z6fG82atJPLZG+EVyZorymM2VSROyeNQDC
7qkYNvrVElzI8f/CYjdcpUibW5pecyYzor5v+w7eAURZ1sL+JqmOO9bKyeab0JT2XpGV6avGGX4w
+1Nxh0wPe/ijbfBdfN1JSz8SJn2d+lb4+45YGY1b8QqiqFXF/w1onA6beSUq9Kwsn507k7ReLV+u
TsaOJgjyzErbsx5DWBnR/eOezkrhzkn2lvn+Cse6T7kx0H4+830dnG+VdAYnBjOQPz2nwO1VtjlT
+Z3xGV1nfyoYEigNn2Kfh/4c6ZQCNigi721qNWnNuHUUqgCfHxLBeilg1/Mv8EwR9MURO8NKrVZh
pUUxW400lV4G/hSx+kP5qKVrWarr5uc2eS3BzjY61ZJkZfCk3znuoFcRVh6t2+U770TcuBgH1UvX
jV9fzE5/aIDKt/fEmUjgTqjujusRdkrKMzzyBi6/GbgK6Q9f4oIh/cNxODHTTIqnsQG8/7dIs/t/
6/+QzSWnE1URJmvmPuBUl1EZin0yCM+aDsXp9tcO/O/+6FlWiL6/7FfYdpd7xw51+AOqgb5SPAF+
UpRFWUM7Jwng4dzGUwymtIcbzs2t4xbqKqnjbk+YqrkPOHs0nooP+vCCfGApgqKBY8yyPosuoWIU
l418wNOoEzuGIEMrkO6hyDTVehB7ttiiyaN1/YUSW0xmLJPim4Fj8fFeq9qqtdUgWvftO2VAw3NF
LddzpiwkSyqwCTy2flEeHLDaihTYyYBKZOHht7iJM4uTJMPBTsHzSZBM+qzaw2oeFXFFLNApc9sp
yHjMuIy+IMTZ6iRVP4qeo0JCvaeEhDPd68mPZyZsrS1OnIeFzBbUTB4x3psvaR6wRuRk5HnOZxvI
PegWOh6kzePN4u+bZ/fZ4fs/WAOKsND9oWl3wfGgAACVkZW42VlilmWjimXE59XdUNoDKMlK2l+M
JHf5Q65iVahCdIQNiK5pRbtWgZ4uLlUq2mUANmEeZKuuqTPzyvSB57lxwJzumoUL+FrlMWjBb4cT
R8xPuE0bwfSoRL8HhwyJ4Vv2VX/lYKI62Tu4sMV0u9rRmQEni/eVvtQFjvDT/dez8cLLjdCkmj2Z
zoXIPw460veJECN9+as0FtnICgR3mqJyEz68z+Yc3FSJIvTe1QjlGsSM1IjnCGRV57eSycCzAx0b
J86Z1BaTw/zgeqOFkGgbF4FYyIG6NBAXVgOxQF4C4728DSeoKe4sdoNxIDliSoTyIInCWPG8WNHM
LhLX7yDFLPuDhXBzl620bWPW6ZDt1LUtH58yNf3sRxX9k7ySNyobIdSiCtCCyS/qDVmnvAg6JBWx
9KXMIfxdRtnNd9abJFGvoqgSSpIVoG6nrbws1+5JHAwIojG3MFygKtU1z72ycE4Y+vqlBYbFRl+Z
onojXkPohhrUm3r1Jwx5HsDWtBsYwyTo1MukCPtpXaovVY8eA7K2tgOF8yZVqvL++iA4qAcZRfFT
xmwcHnAZRGIOG9/ccjHiGjDe3+aQO/jaSog1xX/SpumgaNwL7C9zwSD4CKjgT/DOrKFYf4wFKcIz
UCWUkWaPre5naxMzTN5GSy9y4lEXjrt+g5rJHKAzOGuSkwUrRAwPQW0EZpfCwfNC/oxn4EiXrJOu
FYEFopdpZfQOTvIr7t+Qd1SlrqmJRwsj6GrkAa/vPJUR2cgjq59oj9o4WVPlxth7xo8qdR+s8oEG
bQV3oEqd7Ud9i1gdK++iLC0irvlmOjZsiraFJP+8byya47CIRV/ySm0E1lHzVOu6v6WO3bBwvMP3
Dr1qAeod+cPdwf4UR/Qzo3tzTg/OaY0rPS4j1sVpBAwh4ozGS3UzB98ylwRU4lH0GirMKf9JQKF4
nD7EgblraHAjdbaGTVz4532qnhrgnvyi1u3bNFO8vAkpU5P8DNQHSDxHV8S1Pr6Zb4gbljAuLTy+
bWdSyKpu912zIG7pgE/qMCpu8Rr9tn20tTEnCnrtrQcVS5WkJEVfVNj5TTSEx04CqTXY0GsUOLpW
zD7ib0EkSVcvqPE0WDzv9NLPnft8t7ck2n085otB0+d6TWn0aHrKcNpzQV5i76HNrZC2bgfh+HRs
6w+daD4QmosPaeCQAa2BC2C/lNwMCfA1AKLHBRMMBn1HKrsdFrCPkICZbcbl/2sNFLUm5Qrm0sfv
yJBSXamj3+AcfRhXk8O57I3LtAqLv9PeCIsklgANTXTp0r6PEuIofWR2lJvP+wG1Ny7xJG2GF5j6
mBFUm0Pu9CnU2OTotBHlZrHyJipP3EEYdmiLo+gzwRwdv4TQc75D3I+ue0sWyFm07xESIW7uspZo
wpOPPLgIzgNRyFTN9spBF1ILvS3Eu4kwfykufZfjYzuIg+MkIGFqjgzfcq2el5ME3PNrC4dNmllp
7FBSFz+R6hDVG6fwBqVVg5Id6GCuzf85s0sUHvfGm1vLgVKc3rWvrEI63CPRmEjJ28r5GP5/7ZyK
jYv+GEfykgJral91Sz2gJM5J9xEdZ4fhlJDRhpiQiexaAcj1PATZR/GurP3QCtV+iIkjgboBZ0Nq
fVxXRN5RJe6D9LDgNknjBcLyNBN+2MHA9KisckhU6YvnWwYBy9ZKLfhAxe6PtCTmwi6va1rPh7Q7
R8seIiTrfsR5ov16cJknFkfssoYr6k3j9esLfz2O6zO5iAi1WFxgifjIpAQaR7Slcn8C/os6i0OV
le1cwEDcKusvfoMtrnm9iwK6PW2/sL6KwoM8MDjGPhLl2gQS6G9GmliXBloNiAkDjIB3FclcnHr9
DWqWbeJCMfemI6EU8yyiNO2pL2E+6hPuD2DMGSyS1Akv24FaruavRoaJY5GZOepT2aQ+7NtS+Y1+
LEmrUIxfw0TfMHCB+d/g3rP/6ewLXzAsekcAzUmvaPAfEurAmdhq/iXvtc9+OVZL/CK21yJK/QZ+
3bWfYKdKJ2eJz/O2vUNh6Bo4N9N0oczV1mPThQHWy12NfuGOOYrYWJehpN5wLqQTQeXIZycnTeSb
f0/vJxoY3HcogdrcKHdSllEjL+5GKU8jMBJl/NuaELtbHhrv1NJjNfTUFZqsYtQGQrVINR5f9+JI
kUVc3Avsk3as5t+ywmDGp0ob4w16cJXqzQez4F8RZ+8/ODN051zwBU51SLjFkTDkyAGOmvCMESLp
wkwxwAyf7DL0jr3DoEAxTA9P6c+8YNHYh0DC5ovyg4b69uJ4BJ8Kocm6I1wbJi16JCeGhkbVVy/7
cOtol2V8rBT7KJwdbI2L1qqCOmLh8IsMneQRNs0+qsPJvLoOyFY0mz0/CztuEhnlX43bcr/ZyBwG
Pe8uNkarGVePVbRMcG745L/I9QidMqIqEX30M23oLjq+wYIerD8mU7wysz1JnzgkkjmJYwqS8qvP
uyQ8r7co/yhqZG5D7OS8Y/uNaJUhZOvit+eMwfdFDWgsWJDttOzJS8sooDc6qTTIqS3fF/EDNVd9
hA5zesm6YepTYLOAHvDqZhQ8k/h6001Uj1jYb1ZqS5gp/OhLNmeDA0d6IcsEIDrz4Lk8X9T9ImHh
AGHGWM9Rb+7e1J7QoA28F64aAARWVsi/qvsX3vKzDXu4EF/RpiVVdDDGAkjDeQ51lzn/8wrxuDZN
lTT760dD5FEVVpUe0sjWHTkPxYXA4G/jdbV0cCa6O/GZq/vONf2OHhbYOROLtGL4eRyI24V+Uju8
zisY2G/6lIcrtN8JgybQNhI/UlSLj47YBxTR8gbMWphchKIv88D6LPB+PM6vLrrZdDvb9z5rcfLl
6wy4oSN2w7kkpVfhdSePHUWrNX56EsjLOBFqUIbNGqo/uvLFXh0l4Sypl+M7s6nBGE64mpX325G5
mNkzS21XS1AaTirBuDgqlqffx7tgetjMc4GBHgUNKB8xd+yEgQpfx99PJ/IgiNG61uC2qSdpKiMb
uUMrPADQ7UeFDhyyecXHAjImD13tlCNz0LDTipM4VC2sFS8koGymnsfARDkpk/01xhFSjT4odOlw
k27rJshGP0Xluz3UigP1F3dWBnYD2BmzwaBaxPiESM/uERX4bxCKmzvZ6l0jGKjgK+4ZQz/CxST2
tZ86gCHZ3YGDzEvSn2SSG1jkTMQhM92K/0A9xE1mZOwHqZgb0P48VghbG5mzqZYadE/35/5+24Hs
pQcDl+rSR9HG8/ACp29XQSDdUX8+rkgdc+3H7nFjDSeLV916EPfUQwgQ/ZGPOKSSlDk5uTBOOtnh
fhPi4N3zg7EVkPf7Z5qFISLjc157JxayzEdEYDBWb3W+7pfy86VavZ7+xdB6dPq8tvd7k3WLAhMQ
YfrIyG89NUi5hcaBfPK2+YxvoEt1lNvA2iWwPRqGYwGjqAMGIGT3Lu1TjtqwB5an5hDook3zYlSV
HTveaYX7K8zNqTTTy1oeZEajvCr7m+JnqGB7o01rjKzaMxoUoQjIU34xJmsESV3wFSGd/2p352qA
MSjjE7n2JsVY8CtOg122tGWFp6vs0Oi+t1UtOB/xNWksqq3ZVn/Dv9yHJ/YsfW6beAr25ytqWuNt
kXfVKPLiTazbonA98a6ipfJls9VPytjGjfaC7lGAhBZCz/ds8gp8qV2OdVonf5nZ2hwpUroiHDT2
VnFZCmpTiJyqpbBFXRAl7ZRTE25emdye6YBZU4mPNMpjMGW4pp7CfR9MWmjTurel+zfv78PrBF8i
qa4cVlPI/0EsWVN8PFaEgE3YU0SX41o42miuA2WqSrmpHiZs3obrd57SIoWkY/BZS3JbgL9XRjQ1
yTx4E9JjxlrF0b7f/kk7mA7THxRwbcpKVha/Tqzdy+WHiZX0yk8NvA98CHgV2eKD14rouTLbp/tU
xyfz3+uL/hKKuflA3fdHLZICMidWhKt7mlolk82gmMUG7n6PSh8+fxfiFz64O997M+YJRjEtlt9O
shQ/XMtLpyjnBpnvoln0wKq8S02RwM4mu7cxBbp7qTfXs18ZtqjIR8JM5gfDyH+EYX/Mk6wFum8I
dcRKW7maTqWaZnOovuVwfMOf5YdXjjO2hhzPcXdWyWPS9rll9aIVLNzXze0QoWY164Tf6/2E6+yY
6OByYNwfEJVI009rh2+UOJyZDdNtJbM1+7tkWmt4/MYvbRX8Omrf2BhO65GYOGDPElmSZoM6EirU
l7ximawdjC4Hqu2aiIIuIm1S1IlewSwRq1I+wisq7Ki6hJACyXb9fHBlx/uaq60VwIQ/+lkp7v3S
L+xjUynngLsBMnksb8/XYt26t8d297YVRMNkxPVSpiyd/cTgJLoPMe/UTkKsGpHEwYDf+PoAPNKt
j9O0CRXZPQx1NaYL8hi3kpyvuKQpnYlXlgYSlnIRZoJAkUL4516O/FC7Gv0xDZILBDWgbAq/QyPh
SgWy2SQFgRc+CMXaCWvS+F5lWHnls8ZmzfusIbzZCWd/YNBpgjXD2y4KqO3IykgemVmr5cTREqLk
BAhu/aG9iWj4Y85tlTD0Y7p35kJ/YEYfRZUruU81O3N52+i6XrvZUU4CVqEtMW2Q1viii6sfhX2d
8v1k6yIwpG+RDUMSb1wNWHqfecOAKTS1gcL6VWPn2MzE8NCfIBXVxgtSoxgSvYqxwoqMO7dzvgyq
l63gjN2dqT2S/yuEkJl/63x3JrTE0GagOXmT8IjNoP0r8j6gjqtLVSwnFTUs4vd/tKSATEzXVl19
bXWDgmNcIZK4PyLFoa6xLgMn63a9/uGzZ9T9Gru/n44KQ3A14Sz4bh+UdGl90Qs4XMLMm+FWA4bJ
t68hbyg0OeuB2HPQqIJq9ZQQvH4qzb2BfqWJ2p1bnP/DrWrCL0MMEHHNMDfaD8Sm++p5jA+qZVLS
wA51CAxOLCWqRavwyBqwMevYZQObSJLIfNAyuhdjxy+tCHAMICMQ0/gcum2ZQl5j9m65TPCOOyGF
a+6By5CRCIdIxTMYQBelpXrmAbKFJQqDdEYWKHuAbRdqC6kAl92WjifWTECnRGHK14bQxWtN8GtU
w3Ky2MManLEvLX0IbDCWGYORSXJkZn0sKbco6GrTNYKuAVa8CxABpVj018HnkQSxLc5Pxi4UmXAN
CJ2W5suvoTescUsVUvQZCfhTMSqrAx2Sc3mYoSzmMatQntQP+AOr/roQ2VLV7Lsfr3hLfrnVvDri
jDGkMih7Cro13K87i/Q3YhMFumEf7usNC7afHasJqgOEIqeyPqrhqDU4Ot+ivKjAUvTlBSSenY2Y
UdgqXx76WhFdmcpRlMtcWyT/RxWt1rspB5HwaYnVgV5itmQ7wswyhDYEPiQ1r8nIUECZnHMXKOLi
KfYjpF+azmGmZb/BMfPiwONht4raokupwPZBSslngW8RwnlTQEzfqca3bmyhqphX6Y6/hJWUkdDY
GoHF481SAaHZVV2Q+Ei5Miro17LBVkB/NgMX0OZVvCKFJTK4p9wogTteozU8hrJ0xTWyR3xuEgEP
FwGatMLBe4WrnjlSnEHxr5mkUhilvoRdCg5eKrSkgAYl/h0BfzVgOpcL+5EOpwFbt4s9sPEnRoi3
rRPoAg9KUsf3WD80yGhSFr7kFOWDowESOw7y4RRB7FMRPgpgm0XSBp9WZnGEfUFAwfqTPElHhoRh
lXCJ5vEWRgm5tmlY+816wTNdaPl0JcnrEUHLKRPD+azpTmdlQ+0OE25XM06MuBbXOnwPpjxcVhcM
OonObBOZ1/+128NNf/RByf9/9islCqwIYa2X/AkU3IRgF9vCw/uhKmO9TQSMcGBYIPt/Mw3VlWJ1
c0EgtsEtFbru0HC/IuuhUenq6W63ik6I09AgtojbWmq+mYFiAZ0Jr92ZOFfRIUvRmKbWLi9JOMha
/TVsv5Y4rSGDJGVf5LOGlGcO1mqjsDTyYktfTS4CtElx+qehQPzIztoDTUxm77oEBq1AkPyZjDLI
sRconussLT3li19UWqbApQHa+g18GRQN/Zf9UBSXF6i7cDnPfVjmVHdquxX6Jq7xPKx5ue2+sAlT
ooLFmxlBo7HdkI6j91guwVNWYknvjIKNnEaQcpndbdlPBFpCORDBNCqcdl+X5/ypVhHtEO3dW5dx
9Z4fvpEixmvcRXBLBjkQR784yMENROPXtWddQmZ0IWaKy7l9/jEk4+crR1mHxM5BHwJ5s+QKBFZx
SEhs5AuHyQqafQNJ+2gEcqyCzfJS1/mN0TEOJxsAkr0gD3SI2NNAXgrcRDXjzIWOlofBhIAuTKVS
jOeH+kT9eED9p8VHElW6xnl4rJPAwWjtsXtljRpFWXeMNBThylLmqhwFeU2DcA3GbRG6eSNNNCfI
3w+EuacClYJhlHxe6lKECW1nELQuf06CM8bIHGXKLs14UM1PIrCg5/dYQg75Xfn3QtkOhpCrE8SQ
vm/izyGpm27p2lT4XBVP7lPhcyUo2mJGzkBBtAApCQdTefd5ThX4yVwm63RZaVTAn/SAYs1HURVL
ARmlEumzPHD5eRBSpCxfIAIurSYp9QND/5l6OczJTji9mcPAeLD7td5XfSWMSo8kem8p1LfIDtpU
9F3amqcc3CDzlzFXTwem6Mnp/jQrAjYdDDLNh6r4RVlnrzA4FVVTecoRSYyB6a7Q+z39v+X1moIK
2EyseaOoam4G0MK/kY06qpMLLQZTE/alGC+HgrFif47E4ijESAz7CpPI0M4BsDDzicccIvRdFkDk
Wz7Zysm7XWXao+gt4d9H24EKUkLP2YWd/p/xyewOs1JiABv+a5ReUlJLVaLHIBkb6hEPBaMbzn4u
RyC5v9lA4zVQPuSV3SyQMzAlChpjbrpXNIUqDYhePmFEYtQsQl1lBF4a5ZXTrM4L+KIcKi60/MyQ
iBpHkkNImVehLog5Istqn1w3EZC/aBvl2x52CKP/M6pi8r2LdJOMjTvei33ZW1csMpboPe8NOysO
txM60q2H4vk3sBnjhG5dURYGrMsCIa976ZGUA4BjxL7OBoNvftmfbqgNVOdx49n1snIJSvLnOoVV
xbwV4/LiHatt5Z59ICADnPpB2hiC8X1uxlccezFvR7eAFOO31A0RiwZysGbR0FJqzgPAndzPQG+C
8OFuPaHmGb8s4pd/UgzctMPTbuY2fC9jIIQbxhDrxGqjnqQYf01qmh3RLdHzc3IVk4xY0uK6x9bD
ROaYwVPdxwr3BMCyhPt/RsKhwgm5yoMiB/bAzTnkE5PDkVlGYdJa/2f1YWMWP9OeSygDgOp7Cyhn
4CUHD7X3hnC6ts0znyea/52Jw+j15QjRHLDozRS5yMOKlqahCHZMVyTmLiLFfcPeB+YzJnIsKop7
/d3XSy0cTadH+wyR2ew1n2MRz6GUlJ+1nnt+4xRXR7+RgtUzBQySmeJGRxKQqspEc+/B3SF7jqiD
V3RLM4SHQj/Ta+FCygXJT8PHt/JNfmugOszXKD5OjmN/zxumysYjAycQdcSQlP3qNh6Obbk1eHVT
42ERabBst/trz7Q+lqOPapBxiY1IWULvGxEvJCFgF9FqO8kjNkG5AVarDGWC8n15Ad7eUr5xip3d
jA/FLOq7DpvgGWFgoXhuD8Wzh9BvqPYOqHvLPbNksDSvBCnmvJqr1CaOe2zB5+TEKoFc8B5p6zTm
uUCRaiE/CaFqT9gDfsAttD/1LZrtUmYT9iL/9apfsJ68NbUvqE/r8plwOiE1qwJOkkOxWPOG7d+P
ALBnPBHfjPogTHevwiBa/xxIfplUyr+OR5/vN417JW/qRddWYH9FatQPm/F6fdmTAvYVOxjNSp/P
TcQs0iAAu7FufUO45L1o+zC9upN185lOAkajIHK68kSxWK15TxYKT2ejruHfSa8hoB9wrxkjnUgV
XafUiuDq+lpswE7e79rJWRzRdIa1VwTxcPBH+lUEIV1NzQVVcMBtMRFWd7gIPS52T0HSpHsreGpy
jvIIXiduij3zsrzj6DzV4rvCRl7PQkeN74oaDGrQ8axnS3taOoYZ+ZCGk+PzLXuu2elpG7VAOyay
iUmPLGPpz75O6b3s19WP9YE/k/+PMIHtdR5eP+LS5JgpdGIFEiVvAUyKTPi3QBmYnyE6DJtnuPGc
Lv9b66vrnZ255m4L+mNAk0m7rAclPx3AKncH6spjMksDdA6T6ipyCQ11qFtPQBlaaTjUs6aaGa6q
azKk+cPIB67/Ire3/tBY0qqmUr7ODAJQBDDdn+1BRTHHssiD/VjUwCE4mynDktJ6Da20wDJMCP42
Sx22Yl9JdxZOSnwmYYbyi3KfK2vV7UVc4ncr7wf7VQLf7Vh0xusXmNy3YjJ502uAO2uWRk9E3wWM
5Wpxql2F5Txt8m/XNmvaXCTJdGAlBrEo+kCCt+NsiiUj3OT+i9pyCpJtZS0BCdxDdn0ouwHMGD4z
wCqOMS3bie9j+Tmyx2mokPbhPu7tZeeyteCQkzPOiYRO94zooABtvGwcqZCCv5GGvGHXp64UG3OK
fTAJCbsjdTl+W/lxna0IWGwAaD36oCZr7pP7M9n5YeKyTyXRsCaU+xV40DUL2BfF8NUBc2dj4PSM
NrOMsLT6m2WWN6TeWDFSnpSThfsJqXIxbo+jrCSgKFT3yi6L/WkUzS4CHIS0V3YkDxnPIm9Y9XwT
Fsp+0bWOnIS0mQmwTdL414yUi9JSvdTZN9UidEV+zNX/6lPIsKrYPAB8OorFmAxoh87H+TNm5P9p
tdb4WgLdnN3G9s/HMojSox2F/Td11dbrcUttKDL4YIW12TSXhPAcoxjsrDmxHPCx1l2HL5cMY1Yg
rCW8ioPFicGyt7sm62M1xIPCquIDzdRwXgrFnbqnp1ZFadbJ5kAprZC6UVLX2qy90FEp4Pny9vwQ
qjqRmjYcVFGVxfwXa/bMWm2L84EBHv7iPF9gAA+lz0e+ZNB5Nq8dqfjPcB6sWl6OcbOnlBvpturE
jRo/JMQ2AniNPhVLqWWFk8yulWjOFt8gMBkuo9eoFaZ6ZR7AwTj2ETd/4ugljrL6Yp0unB0Fmrly
16cTh7JtW6DdXdllDWV+fOoMNK/Y4A9A7Zkj72s9wCM0OVbGL8zkYZ1FsFWwoIYbs8YZsAanp7aj
zNDkx7jSU30UcVAVZhUls5ah3kYQUAr1qCcYzcd15/HkmcD/n/VPas9DgtN9MYG8RqMfgYVkugOe
c4oaqElZNnPXV4m4zWf8EDMbb4g4Fm3tiZcbg5+OFyHqpOj/9QmmOqRvON3T20lhFZPn9jKpRZal
5TKtY7V+kGQ8BqhM5JPSnXO6/eeA/FjfGRKKr56J1Kok1zqKnGGP2m6xD7oPCipexrU2TUka27Jj
K5vKcQiqVLWqYpuoGNHwirby+zkIjXaYm9p19vymOTX6ezfTDv3KHCx0vBZzXFM0TRhcjXWcemM7
d+jldB02/OxX3xt6mensVimwOuU0poxN7iAAntfQsKgrLNQ8f4LSb7kuNq8P/Qf8GYGKhNODJULZ
trSOzgUxJAnPax033o3FMAhC8af/vItq47hEdrFl7MTX01Ur5Ag6iym1eA7RjN9oOugKDSc2SJlL
3dD/7qEsrby+Y467EDHwCawBgGxoyxKFY5UNYAr9sVz7yxaA0hs7tghPKu74qlh94zo9d6ZvtNUi
nv6RINpVmsnfBcByZnnLtGNwplf/5BZRkfiJ5R+AncAtsP+TKj850mpqZqToGA71A8kdXZIgK3c4
9TqCa6ZGL60QWgctAn/7/oIx6FSdbSaupKNPquPJ5eZADCD8OilOmQIDw6V4ZDD36NZpYrBsMY+/
lPkuoEjpZFLKV5drBFBttkQHcmHuG6iEG4lpPRBgLhpBMsMXRESOc2Pc/Thrjm/sg3xN5rNyeEyQ
zCRqWYgneSslFlVCMqWTzs8nhOQONXFkobk9G1kizg0aBNlxw0zJAvt9YtmTBQOIjT3c6wqOpoYn
bknfIqMN26R4Pi3eW+6UoeMkm/tBXmGN/7AaFTR2K5ndNONGnkthTiaWqqcbgF2JB32rQPllTefN
zZU4EjS9iM4lqAe6VE/TzXuLufMoCHaySQywgsY1NJolriJ6Ms0KkTKz24/6Yj4qs47GajYOrsSN
wm+O5mjlQzbgjSS833Ee36avV29A3Kxv8tFe+QLAH9z/mscGryScr82evgJ8n+M6epM8knto488c
1DSTM6e9mhluuDCoS6zrvNkQFLdJ6G07ScoxnOErjPhTE84wRRdI/q7yLg5ceyB0O7v2soL3jzs3
+bEcZ203qfdAJCf9rgRe77ky/zlkioEdX633BlQdXvePK/KXcO2I/6JbMUv4uM7+sxpXOqrIKQjO
vv063kCL+gmBDPLq29eJeowm2Ukuyto5cV0kcx5dD5ePiMW/0hl3JIPFKiHZzJkVkCECmv38lsp7
UB1XeRTj1yIRcdiRlk9zcr+pFEX1BYCth04L9oI8dzLUcByWcNkZmT51B9aRoYkTEwi4r9zf7YDz
uXkSQm3C7N3w2smZGnDHJDJofvs46eF2PPIkuGfNm2hBVhNI/NCEnqgMJh5aCQHLWVFlLaanp2/J
HgeK5GffNtUrb6k0kqycCEepsfNdeUF7Y60GtyZE6//1pbEw7OhQ1X+yEe6rG1GUo+GiHS/MrcMS
ZCBmcroR8hhj73dMdNSlN0uasvgbji9knqtrxl4XtM2v0CiiGXsLI97gQcowVNnKjVFJsdlw5G9d
y+y9Vy7srNqonXr8kw7JPesYZvYyqICmdBY9rKK7Is7g+Vh3uQ3j9dp/8JnA5sm37thpWxC0KnyT
IMBslNMe4KfvKL+DLPDE4n837VqIGy9ZnrxCaiRVkhNvtvts6pJme4Im9z/z6AsfcEyvCNsLGRZM
l6NzMNIPf0j8c9xOlBhUiotGOsidr7ltFDwpyYjJ/QY0n+MPSn1VfghTw2j/ywkQBCkTOv05YPDP
Bjb+VCBJND56h/XL0T7NwFot11g8MN+YVbBlbaWKkIPQ8xPRPloq59cTKOZYCQXC1QoXgf4/MuOD
o2oG/Ts4HpLNjgABqANfsFjsIFM3UFXNTQUFeFCMCr/JSXiLlHHigPx4Ealbiqio8SpiEPX9JxjP
5lAQ0j5TI6l16o6OfdWfrRN49NiqlnQf700rWmV6X3PvznXR3WoZZ7gU5D1d5NwjQ4nSZ5ihy+Kb
GmckYLmgqrHgjMCuU0lm+Faiwv/EzX7CyX9xyrJagsaldVHhnx3ygsPWwj9idX+OHj8UJuBKQr6W
gNn4TjFrMNpF7v/Bx7F4bx+d650ThQVZ/lrHZYmG9o+tkpNujXHkkG/jggLZoGNe9e0JqN+2KPIB
6jKL1vIbOaSNgQW5zO5KWfNx2ExyiV09D85AE1ySpf6X9UaKv1/6EV60R8BFywAjpsAKgRAgDt5B
8iEGLpDAD6IgUOdR+EN4jPdwyTRs8z7HOht1n6JDaOfaZntz5NVmov9u11ANbRB6/Jz+S+A363Cc
aNWJB3ea/RuZ30RtvL9/EcxI1BKuELmN4tCTM3RvwKP5j6Hk6qIEjda2cswSRZm3MCi1QG25S+4X
Xlv5NtrtrXW7kITvt6bjus+CPy5hd9tgUxtukKDdYolMlW8cG3AAR/FvtqopWyc3hvjKXLB1SE4E
zfiJ73J5fWDDuzqeK/n7ZyfCcewctgG4aplJmynuJMTuvGZiqdUp01282ymCdPVHoRxvEobWVMGi
o/luG8f3wtbZsHOqU+ewFu8/7jvlmp3vrOBJ73Mr0dkgxzyUWo7iNorZ6pqdiGhIcl37z5UTjAwI
MsH5M5GRnvqiSc05Y2xt1rPgexph8Q3BXDbYM0oNRjqcEesOFnN7LB0lzXv2rWARoNcjzBXwV1G2
s2GaRV6LuMDOKazBTblqEG9F08mtBc89lTVGmWxu6oMAukjITWVPesPXY4AbvelUkiOrCt3HR6aO
PBPzStpaYDMNIGHJW4VcLRgmXt78pWHyRHwynUxfVyrs8cHkp9r99CAReSQmvEhp/bLpqf8uQ4Xt
iL1A8OLUGUInTtjWFFoIf7WUH0tSfYybyQcMJ/myhfmezXZ6fHUkzworqBLY9R8NAkx3eLrmKsPX
3k19PgArkDxPOUcrXeeuPwWz3j0DHfV+IoVwxacZG6vEY6ukMpyuqa/kJQ8Z/u0aO4kAFXyMj3ET
1XPlXhFPg3O0KtAdkwyYKH+LSYqQ9eL6IRuQGG7OEumeLU/vIpoI7/2QyxFZhuLoiledUXGCItJm
kfHssxdhrtd/BjFKLt4nOzTX3dyj0RbFAXO6iAcie0c8a5pDX6gDEOULGohNdmJKHaZP1kTfJ2WJ
Z8z7ZBkIkvCORha4fviV+kqRR05vUk0xESxUTtIVE8uq36o3cSo5v4lFBNVncD2uOyhM6cVcGx/h
80zF0EwpBMvpaJXk6XI0bUJ1lU+LAeGsXAHHJlz2IbKSA4kwE+DI9fHomsuS5+lUvgzHQS49r9jY
PglsBu+dNK5Wpm6i2FALRb49lqgkGoD+XjIn2K9jZ7y+lezrl9Ykhx7v7fbitvH/2HY5TPzTHvn1
g6BVH/JImm8awxO2VhOt8VSirSKVevuPJC0wVwQS9FvfpBfUuxyr0eZtPjtxWwgoMG/n8ppsEUYy
M06zjQHihIt38s9iAzHdNVEvEygnZH0xCw6jFYvvq0mTpXw1PjWYra826Y+SYH6Tby7cfmMDi3LO
E7gf47srLq2LTQ8lpb+Z/5kp0FYNL2PNseshsu5B4Sz1KB1PtCXVh627lapMa4t6X1824xvLgyoU
vB9eYG/N+pAJnKi7qiOf0tKNsA3FkrY7Sn5+lWMc3/68MtFrXZr4Y0lIKLy2uKmhxS8Y7AA4VQTo
RjmJyCJHA5A1iWwiUrPnt3JWVNLIvphmhGBSd/IL7YCtbYmy3Gnhpyusd9ghSqc7e/sIPkExckW/
Y9yGWo7KKs0zdVWyTuHJ9sAUxJLXsPeP5ZKhsYl7ja4T6bn7drYaXIpaAAnHeWeG92Zckxp1MN0O
WlAtp0G79ZQKF22Fm8Lsjmi0Pd4qw0RbjP+6ipNReZZix0K8YbKQIptcWO6PQvsY2Tf9zOzqxOgW
hM6L++SciavCRwnMbB1894W7KoOLTGZZN5OLhvFddThbW2OBOlVrWhpoALf7yi4dj1Fj4d3pfSqH
MosWQ6oy3bqy2M2FxXZk5A1wKM/kuk1RxtA+cnctIK5ahzL5T9YfYzeJmnflLiKT0mMRpHTvgFpU
t0wlloano0nekD/4k90vfcOhJGCG7mAnv2f+eArJ4ReF2Fdl6DKL6+5VE9fSyH2STlvuvQGZ4+xO
rcpg2Vfp8SQmzzF2rO1DxUAj9TG/ZCJm40Ug3iKh08NIanWMeXOf6xyq7DeZalFKyRniV2eN9YcC
xkw8kJ2Xg2uFa//MANl+8aB3HaYTOvqzQD0eaLCIDWQyf2ZwUpTIlV7oj/ayCI9MTIBKM+kN5n+t
wqlryQ/vf+l2/fzmwg4xU++Pb1nF2P8pmR95FWPgQ+14DxXJGGYSqZEXCIBFmY6qpM8sZ6Cb2DHl
+fRyOD0bZj0KPIwWq61b4LUM25Bc7ZsHdiqFyJ4B9PucWvSyRW/TNM2914C2srIwjKTwHIglsJg9
+lpu6jEbXtmir30MlnsFR44rkMsWPrt/3wSExcP0Tv3WzY15jo3pydQVhGh7qt+tLO3QOWAEv7gy
hu9ss5KO6UseNnteC7x54JFhvFYmi/J+e/REee+3H7fOOvCNER7MlbFcCsr3CDF/hzXQnsrpmzyg
e/Qnmy2IqMlgXDeLflKcCwalq3b/bHSDb9Eqy4DyaBAYWrzn1lqyf7IQoBxeArQmm9x/CTNjTiQ2
cWJPr+EqzHA5F19UjsLEZ/I3ggMRUQCj5Zp+bTOQ1VeK1D17Ol1u3sbCa0TxgknvmLK58pHtkemu
RHrGsM6/4CpVSnSod4/9SFvcHyMsAFUQQ3T/XaPlZaIT1kdAckQPriNPezN8zgNkuHQZ8JXnUa+O
fLwnPLu4NeA8TD4b9wraHma+V6gD/UnCui2PK13SB0tgrUu4nLxUd2X11Jpt9w6XvR+8acosnOt5
1MfPSPD/6j358F7rzG4+1ntEITTSQfj/A0ISG8dM//5Mz8qAia/EWLr9AL9I4M5Us1FuoNrJLrxi
KJbASbZYR5UYHDuIOA2GlbCsqyOVesR5A8j5J3cfmiNMs+WdhhiX7RG/ai/ncbJr4wTZFjKZvEs0
FmSmxMQGtc1OHACDpBFs30tUaIeLDTGZK3zA18t2HBUrJbJyzxiIimnf91nWOzRVks1qTycVujBt
ZzcORK955Uoh1uuXkxw8V8qucFFIAZPzn2v6z412+t3JLU8hCIc3Qhtbg6EcuATMeyM0lWaZXrUo
fu+GHqan1poIG+/i2jh8jq5HhFbJ2Od9B1ef2o/WXkbmM44p8L4ch64aMLhu9rtJ7W0XPmldg2bH
6PUFxf7C5M8YMwB2voKkxTfal3vaJBgWreRHLQrqCsOmTGFlsLlHWefot06pkMaywIWLBKT7qgAs
nnK45oH3ePIA3vBNUk8p2UVWcv0GbttDAB6nJzeOOcOBgLi2S7WLItvGuj7yC62LkMkA/3kdRUnl
j8G59Fg89Ba2od3BTGE1Ig2i3rL2eW+o9JEESRwEj7caGz8dg+y7QpNtjYI30TtbIKq+imtgACdR
aIo8ho69uRuRkdMdW9nHJyD/5ZpQBvUdHYNSoFoiLIdbndDtKCSMo1yPdhT3T8/82/+Nk4Xz3C+l
ORK+OJp9MYz4s0Feo21I5fOos11epQXu6L76cJ5QJlKEZUmVStYka18tba1ntK058ial9cnvbOay
YTsjZ3isw+QYh/EULRu7inr8gTjLQmWA5wT1yx06x8lz+AKIRWYrf2M6wbQ/Ly8QHrBz5kyMV93m
KUSbVjnNKFPxOr2TumRwcjliKW3uE0vWSZmSr6LL9lcQFX2eBA4ASdzDv+Q1ARQpGTdSDWJimf2h
rdDMIODj3Jru+hN0fumg5E/noEKUqYIpRFBtS6QtD6H625wyvRXYyZFNUTdJ6a/Q8Bjr7AGcGZo2
HXL6LtFjv9IJiKFpEXam+HCHy/OARSbiz28wcQH9aLj9A6YbABqGXcJ0q7w+K80SRgjYfczNdjx5
ws4rv+PZoSyoj8TTpCIC4weaw/FdUwJJu1lA4JBHrmm6tbaNXMUI2BkrCX9eJHBirbWkILE7K9sE
sp3Euy2r2ntUjEE+Ow2yKhlY4GkQ8wpXvBfwubEHqdcIDIyU6dR+5sIOfe5sB3KjDacLMrkeouuh
b3oCN08nKW2BtROt3RjkJIo1eF1AdqcRD61LmTQf+wRK11EZoLzlqN959kkJDbxAdUTAZmr0ryXx
cQ8WDBgi1TyTTVUsNvh7flluD7NW1MG8wOwziGn3w4ioiPl2JuLGB7EAspttVNwAnO72s/e/hoPg
Zt19uqXxm/whX/WjEanZQ6sAyY+bwPyJPexUQ0jwBA0rc3tdO7X0RpP8xv9qws0MD76OCphTN4nC
B3BZnV7IZlmPZz1mCxoj6DW8/3zHosVwc8tEUkXHq9mLtePLcKAdPrZWN3VvchoZqsOHu73t4Zqy
X2VWNP5ozTKIMMRu8mhW7U1ZGnu1385cLK2JPpFS0aOBp0CYO55HyJDk+aWcQfilXBT329CYpwv8
CmKihPBCtTr6eQH5cmqcNreVzhIrBKoxsF2uAycg27mqRw0IahP11NpA8xaqaKRzaWi0LVYJrSoU
6sjNSxx4FqQ0p7bfP7P7j/U2OXZf6cPDw2kNXMbvItu1NSyq6eUNOXneFbRLQKT2HQR7VxE/CRYp
wLiVJPemnG0Hi/i/SCmvKB3dW1op777JoQaNGec/w4W0UbDM5Mo7elIjza6X0m96QGaRp8Gy2O9h
XYzK/Z4ds3159jy1L01f72t3C9NaZFsskXwtRQdeVrujlrTXvBCsct+fUb3uvTc5rNaPrI1LCHw/
S+azmslZrgN6tVMy6Yrgggbrb5e7QxvMf8hCKxsdwWtNHLg0mTLf7r3CRJEW87rf2WkNRoF+LslW
fGx/gkS9+wDpSvmyp9eUPIvQvlwkFn1u3UyIrVp8RiLgaux2SVViJRcCBU2xLbYsI6GMGbmO8qwR
PiuhTSs/TEPLluubmppiNPOK0TjjHYOvd0xzap8yyIlgmHE+5Jd4oByDKwoA4E/yfATq3JWfhAqK
6M/mqv3vYAHgF/ME/d333QHm2I+/AZ33yCKI6wL/ka8bLLHKIBuEKFaf/mQpevPCNq7RZ4yGPCxK
27rnjLm8bo/dLtOl4CpbFGCldrviWF1V55bD60fOzOJjlQD6a0CG0WAGt4XfbCou25snJ+2CXe6i
CpZ00do3SSqwFwNBcfKW4MGGUpWsCxx6YO6emfv6VUMWf4O/y8nRgHpgoQS6bEa0sjXhTe2UZjYo
WklUGcqh7/MzfSdektxA9PBvwwGEJnh9JMTzGbzZs4++/F3ZI0RAFO79RC3uS/0fZy7vZqC1ssF0
CphGz+OXHXSdzBjlchhGQNGSySg2JIfkQhwNyAZE2JjoV55/FFygm+cp0PhgtLn56UU9iR2SxdpU
7hy1tVg5XxLLzRKwpsXVz/ZC/SRU1AVsG4Y/9PC/LeEyqO4OA+zY6ScqsvSqiSnccubybIMlG2Ir
MPDQ4A6KTZyiNZa6yS9sH6TqFJTIfIeWdk9LyVgQGD4VyWntHLaUBshsfmhTgfRjbbA348NfijkF
1xA7nNUbWCQlQAyhQ3P925SZVxDyvSX+aGq+Y0EZ9DKqYfFBizXn7/Iln2oTmBdyQQtqih1kQb7n
mqrnWizrb9IusyQ4SjKkxdfYpvbauRCHVbFx2z3yp0Rycn0fyGe/a3zodDLclcSfT6OCGFU18JXX
7LUrdi1056zRS7Fbk5OSWWiC2ifHZELLowzXdkEIsm6WkVxvwZYGe8SAe1UWp0qFOLHFy4Iofp22
ZY5I5LSu/UYo1fOuLWHFFqMn9UfWuWJuUlnDZILiPtoRIlLwDpQgOnKQ4va+Y+6ACmV5CjG7tnXK
odE+6k8CaWdJclpgxKeFGXZtevdYnkr9bqpiWg0dnMjiUbvW5KzEvtgcU3qhHfyK2RiBvLqzJUai
qXKvZhNG6ohqcQb9GkOioqqgIo2wreNDSeZKm6cMq61G1Rgau6b7TzWZ+y8Yoioe4QqTT/2scXZ/
tS/cbET2E0IOJBlpCQA2vLh+tFHLwbx89U7I/FJ44Nkx6oxB87v6Sv6+jRCzuzCW1AgmAm5tHc3j
VdYndVV7GAoK4pIcRheBRePcVFT0XIp7WahxGc4k1i0cz64o/bffdC4LovclnqxAND647kVbl53m
FDCgEgas/OikY4ylRTq32vqGYmYi8qQdcK+VIz8nTQ6VEhcyjDA4MktRbfEhzPay+ld2wg5E9b17
1vMnOVtpqkB0MqWNE20eyOMTk7q1NVlD7uxUcHcfC8U3qeJBpU8n4CClEd9R4FvmnXkYlr7SzqlQ
WbHHuoic/v8J/8UHQ3ol7pvFHJLYE7Qs5jdc8F73UNmH7H5agQZYKFlly0ubkK70blOSvM4Pje13
U9uyNveifidaHOpGEcMNJVbu8FjncFIgautXncn8MpsaulQJQOgIOUTnNSgGb0caAVsBqfLgeqUE
NQCybBB/2d7cZAxUguxsIi45B2X3HGXj6SQfCnjppNZOznT3ZFHzCqLEz60pRoEDnwAV0gMlH/vX
ppnoPuiWpU+i3Tsz/62/SNbC6TxB/8nPMkaY0iCe4oWSifS7CY3yTYcQH+IlVp7i2jArY/zXRO92
zJbVooWUZyU7FQBwtUE1TqfmTii7zKuHnHj4jp6HD9rje71qGCzXf0lEJLr7UEXLuyZAa0VsiOch
h3qfwkTKqOxY6fwXx/W8B/nNtMC3MWQ4MBturlEIMhLDkLJ2Ju79ace/Uqa/1HawQgdGEhc4B57l
bBUAhXG4BUCUdCXgkL9m1humORyOlEdMYaI/Ocg2qTXdMT++vdYL9Q0Fm9WqfDTFIg0ZwyF74tze
fL0wqQ8Xsxu5Y4kaCsThg2JpIEhq/PBzbZKdtcQiWQJ0ylSLrK/edlTFxrqBCi6g11rkKhNdqB3G
bXoNJSikQIMlV98LSY/GXPs0hYVjgJb9sPa/qh3d9xdbocHS/smehwH5cLSs7wrazLhThzHZBkQ/
B2ro5xsLZebw62B2YXpG9T3GPQ56ZSEQIv7p8X1zAx1XPUuAdBGOtwE832zkqr52fbTLqQG8lo9q
EPTKKaNkc3ZWX7B7T89cogLYH0uXLpOPu39h57smNTIjtSuI2ADkBV47+y9tDRpkPP9eBNi0cMlH
hD8l8B722C+Ot2cQ3cOZaqkUELROCPKtRWaEyF/An7HfKfPIl5RfiVwRoFdpxk2lnH/cWLJ9pgQ7
YiR24VDHcygRh5WBseFCijFXvesWytg7aU92Ek3yz4OkyqkxMV4sxLUoFtY7O0yZw3tmg9wdr+AJ
fxzjkJiYMABP1i9Rkoff12eWRfcVPnEq+SIeEqZ2sXtlN71hdbfBJ5fjTKTSaMdroOI0pjN59mrd
owqj+0F0HlTHI9aG4GZOjCoHtGOzWBXITGt8V/qcmxtUFaQN3yvM9CW0OaesC6Nk+NIol7P4jCWc
kBZUKQJ2UwNGzfXcP9MJyphRWoMUTsFertyE6lP0jpMCbE1iE8vg7OdNqrm0nCmipKf+kmneYM9T
hIHhceVXRK1W+6+tpO4Ju3KTvyvcndFnxDahEdpJEMG2w99ugkl6jyxh4FeZ/B9Sz6g60IqUYVR4
EknepcDjb3zP+LzPto4X4yd7Mx+HSm0QdIi8xRJpvgnJSAuUgdK3IKwSmZHhtqTInDgX+32ZvIyW
2qHjFv265FcUaGH61dUa+NyFNZNQlZuJP9kbIAluYnrPOjs+4bjz4WpZjZHLhWkXHS+nqzcLRAAZ
rmIhRiu2OCQv92CkEysqvr5AmQk31D05+hJlpQ2Ghv0khzGMn+CCQCmKU0Vxw7mrqfzSTWva5nj3
Ts9A/s9RQVxAueSNz0YC5i/4jnJwM/BjOfNRKAHXB52BQaxsh4sMpTgMRak0fWhPJpXSdfNvCdwh
ageB8Whoo6TXEq2SyDgEKViDoYATwTjIw+tDk2fmJFZtKsIIJqT9A2a0STW2BlihI1DwgKgCW8BZ
Fm1cDZ+BfqErXff0+zRCRnQ/cw81f8K0ueQzt8p0t0+3rT4KbVAbtzv9ikPsh3aKc/UXsDBgwOiz
kTyZO59u4VNgtztMJ+KSs53un4GmkixYubUYdtYbzeRr9au5iDERFmJPyhLHPBAxezzA5mZLKOD1
lp1N2T/ZXV6pCPgQ+bjcVI3Ho5XfahjumYd2HOE+r4DbwSW2M5cuBeZQZeKr18c+YYVn97fGQL7P
6Z3iXwFI2XPXmEqjA/WXrfNm69SSoMDnCUYcWPx0XURCPljynTstPCjuxDiLzPLMVox2D/pyleMn
fhKaCb7e4f7HExKS/RbqB3vrJ1R43lhbV/mZBufcmgI2SZOliHKL4eb6045pbt3rDtamAO7j0dRn
bs02tk+/JvEO2B2qSrILk1lF+enEcgHAIBEtcn30gM8yi5XYdAsA3N+zMPa3OwUb5RMS1i1aNZG4
LU9vLn73clCB/DDFID7487iA42Z5Tvk2RaOqx+7XQJdU26zYT0BzF/3TyYEVbqvpuCJtZuNGGzvH
bn7j6p6hGMHZ8USQNXLv+FK3HUmdBSERNPe0v9pTnyTbdTJPUCY4JuHbpwaIfIOPMlQqd46bjbPU
KNm5iEZVnf3cWOcRlzt5RUyrXoajQK+klrcqzM+DJWO8gzWf6Qy6cFriweG8asFkyft/07i8Mvf3
qlkAIHfuUXR0Z8OuARLG6ZaBTjYbvtscANtl1wVDTxvBoCS7+0JcT8E5fjiSIQ50moCINdsXErz6
ZwxxWa7WiafOldz3IQyrZmtE7oAENMKDNcqE5f4iSXuEct0zoXu2ipxfC8uH1DEaECJd83SAmFOg
l5QKfcarWnGjEU43xXWtAgo7J6s1JrQWhe97m6FdlNJZtX/xZRMvZ70cjM1LB7AxliGcwGlIRbNM
1hXxglOB8/u/A2jL1Hi/P+1rdyIoDIfo3FyXX34kYo95bI5wDwBalZlkFxK3MYBdgz9VGUciBBKv
wLkpphlhiT16EjQZIHHME0oqZNt53ej5l3Grs6gi1Tc5yAF9MXnqhqA+JfuvOHx+hRGKIzNSYhdS
BSrtRxy37RXjegb6UB9dPh3f9zjMOVraS4mPKST9hMnXJSeilihUK8bSSUxwne2Qgy+9X6ZRtjEv
RPfeyRhZmpJor5LsEAKo9CyDYClB1afyg0Ob9HvhUgdVHsmKpKJn1xbQ/GIkpauHjfe9NC6eCvx+
l67D3/Z0nL7uAaGcxn54dINHcfo5lG4If69dP5bMvHeeCTCJ7ZHE0/oUBl2pcdA2pr40kUJSlv09
ni2wxHCx+terDqAFSHCKOVA+zV+duA7lKGfWY59MGDyixP6AY0472wb41ibayN0iW3DKfomA4UUb
0XQu+hgs8qYuMuKmP7oKXN7vrLqdLY+eXpGNM3IZ4bWUGa1E/TgpVBeEFVw7vced7YGBsVe/eKfw
SJCO00cqz3XskV4y5uS2vpjsdK+R6ZNV4tbaxkyypnWRo89h3gVKgywIOOE2NCux2U+wmxesGSvq
x077TDwpT5ss7QkUQ80fHHeDbbN1X+RSTHDiuBxqMMo9Zn4Uvu6whxp1ZhzS8vcNt+GFHcQge6DV
M+gzkbXF5cAX+VdymmVFIagj9RZ2v/P6qa7GyfawNqmyDN65l7WACziPqo46Gu8E4XIJoqoKpknJ
mW0IdeBqDkgeqXf+gBf6zHYuRfdbDUXXOPU+JotwaUIvIL0r3ERS/W+taZeEUoluTkwvyPTJteuP
ZCPGxIPokjPELLpeXEISdRqQZjY5PXwoM7WYbcm4g5aCc7HLM49LVm1eq8MlV9bNNJmyB5gjj3cV
0HBu3v2TkyuLdwqBh33kLQAh9B6nC1B3UUxvcwHWfv7R0zeUcw8rVdr67khTnu7ZNI0CGpGUAuaj
N+9kL2zi4MS2wAEzN3qqX+bL0QdvwQu8MXdl1DSg/PdH23EHvZJRICkbldA6osp8na5OToLP7FXO
fVoPkV22xm56KSxhf5+U/9sRbc8fRLsfLeJu4gV+TkgQnATzpYekH/vQoTtu6AfjQvt+GVAonC+n
rWTcYWkwzok7K7fj46iqKkqEFS6Yi4Oqro34bYa4tpX3ZOEzbrbDEYJAnU51vn0tJrfjV2Q/pP95
P3AIVamX9u6fIkDnKnCOGjMvLEW/JP5/HS/mNPDaNvHq33c2hvq4EZTfLmYwTUopNBcjEgmxE5j2
0dZ10/DwnLT1vNY/Bgn2MBp2vpmsvz6Sd0hnvvZ5UBWUzhNeTXQABJjzQkvddChrE+BzZ1sErJSD
sZH0dxLI33JKHsrgpdopbnlPMjT0+Nblog1CzGktCPr8pauvynJ6nm2MULJEVgnm8a9yS7EUqswZ
sgmfkjwQcjEulppjp7C40L7c5k0vIV+feGKZ9XskT04ScDTrpZFXZw02C4fFCKIYTMvlUPtP+zjh
Rs6rBwHTkm1cGorCBbCEZGvjKOWuxGx8HAv1dYweNLWMjPE9lO/6nSLOpAnnTHSqaa47XvDVDQaH
USm+Nb7nLjbz4704oczFG6hxow4mRg97ttjulVwdyGXQSapsTB54szXV2FjXEuZ/ri9EazI9W/Et
5/IfN+1jBIlUGW37AYrPlVX1rBEd4fc+xGAHHi9cycr+3PxMbISamChonQrhguC9vYNrhHE3+RgY
6J4HyDwPWdBaCKffWPogyNainifSVzvzSc1lL+00iBzdNOt+/2siKLL4j3NDrYs8BhohCyKifwvl
IIwQFCgoMTeVNtffNZV9cjSExJtFdFgLtn6QmjpoWgNX4np33MlvFbtWFq/HE8XtXYtMo4IC1hS3
ech1tBULOH7/M7DwhzQX2y9bIF1Edymhr8AaS4W4FxgyfWEl64kaUeScKyVNVFd9ef8CJ126rPzo
LhOUaxcRmzD1dqq4T6DJOo2v1RJLo281xtjQQVFELJRDo6fO103twD81HdW1tCkKFqXUsT5V2I0X
pYFEarAQHnoXKyBPbIOO5vZ6/sjeK1uyFdwfGqm+CQKN5/9HNOc7fAivS1o3CeHEiilv3pZp4ESP
wQxB39OfaPwv+MtPtRXie5Hw8z88vL2o9XuH7wdgZgIeE9Qyad1j0kYA9bnYufWMXWe8/KAI7jNF
evgY+VfioXEbEkLnV6a7DkyEbaPLJaN5amtIX5cmpBPG6JzqvMpftJ3hsdp59DsTtBC75b9+xV4H
jE+UpRkDG/bilU/jTypKY/r7YRgl5LlPm9Aqg/QsdbsIPT767m1iShGZLtWDH08PGNojtEYU9WDF
zv+j/wo8rdwZaH+3PECVsGCEiJ5SvhgR+0NoSF766mEAltrmdY53uigjbTD7r9paEhIJUoeuRmgr
tHeonINqsQ1XHkhCDjlwYMxq76AvZKNN7lwm8QZQ54TajfYM5jdBHvTm1HUlMxZaxcPglI30PFL0
h2adTjvSoaM2EdGNfTV39WbGBLJOpkuzdX7HtE6z1r2K6pJjxGhBZdgwB0hHuxA4pm6LFnSMV5CA
/yNid1UUaREN6vmgogn47mOQM9nYVleOa+rtcT6LHD1c6Fw1jhFI36292okYCi7ct0ltrgx4nzIY
3reQ8R8iHAB5VXwv+Q/VIfqOLBntpPPYgiikJsnNlMvILO2XPYfzT5SrP0yT0+mBFBxcdC+wcq/k
XY5QRPs8vCOvyOXkUgVz6B3L0lmPe0IzUGWuShBy+J+8iRvILn4ym7m9kcM9s3plOm2WlBsRNRNB
CSOYnRwZZJtnhZ5ZRgBBRhwMAetGyAUgqsFfFX4PC7jc1mRWUKbum4eAF3hwejMDrV0qr4+0meeH
6B3aLJi4RuoAOnSjsWJIWecv1gSUhHJ6sWmVRFVm1QZpnpjB0ORW+NcwrLH9Bi6zITCGPk+f8Lh2
hUMU4B+IanbVVxCG1OlO89b1gCnH7Xjen+sGHXvEqXQYGEV2r4qTHZp5WszpXTSsqruUEwQkcwdw
KjBbAfa514XGkMs+dVnUFCntuJQl9FFhvBPFIgzXeBApxGEEnIFLFXxDSsce1dKZTW58LAUupUZF
7ZubqGeV7rvjohZGTrFgku4Tx6ncpWaco0u4gSE06UrznMx9cNF/46l01B5ZcmF/dcMY54xUSc0N
P07Pb1YMKg77kfPdVZyC1aHJ2iOGpBvFz8ySKuWg4LS43vSzaBoBPqBRCE9xfO2xCN+kwHkpYgNW
0AZL6ZPoOLIjMgn7u0st9maIydOOZ+Qp33A7Nm8YRQhpGUP/k5zK19C40N2wI6mzJlpdu6XVKgyG
E3rvdxm071dRhUVquHAWM8tmxR9cG9IubcCUvnecjlFckghjp8NP6HO9cy75QsUZicvTxzGTeLZC
ub5w7+pdo60Wx9bhxt9Y3I5OpHpK+6uZHP8K4h9Ipn1/KwZnbvWM6daLo/UDXpd19HBW1aA0hnXy
0W8PfIUL11nM4r1LtvZ1Ps2GibttWTLRnQHkwliuWkLdIqwtXnUdDh+3j83xI5k5IfQpF/JP6tj5
hDmYqgzYr4wnI70X2qkxkjh1BsAUotRYlYw43s1Gp5Ih9PTeIVYCctCY31LjtifQ4p1mHnbd85mP
5tkua3dKcIvOOBEmCTvdLpobVJ1zXcOfvTsDgRV++uWlhKnAq+5qUf+5xNYCoIVSODbZYMEEEDiY
8xpG1CbDi3OIEXdIgcJBYrLpxvW+jSK9RSCuaMu0cdZbT/ERXYMEJB5xSVwzkJ0gm0x2L6bOAYDV
y8WxyPRK4i+ndkJTImXBQK++drRmrN6jAJLl4S7MfJi+uNAa+rHi/5g26TN2JG2F0dIKHVh1FaST
rlh5SVq/eRDQ9s8Ud3ReJ0K4Z0Ar7kBhS91RWDJhXcI2/1vCdsXWcaOtlhDMq7yguROh2ALwEs3/
kOsjP5JvHZKG2b7zvFwRTiXC8N8G6S7JGMRfF82XuP81O/vdyQ99Wb8GUv9z4wDOrPOCfyYNvATB
RlT8/SS87M0kkjDfxf0mry4sILgrMxNejDHKW6sMeJu108CscCIwxff8ENjf2jVL+Xgd8SmFsumo
gF6GkoJuRvT1hJOARbpDEjk63YFwGh+ua7lLyiBKWTVKD5NU3RoljCgcGTdJdHPzbSeT1O0w6Esg
PP/sOPmD3sWFpjRW4BoYt5md33iHdf9B1IeXc4Dt5WLDPrQTdMdqJK2nJMalgZElM5QPVTe5+jqa
9wtFuhusA0+UrgqiwOr8S0dePcmaQfsdHin+2GPOLgAcweq1J0mOUKwlhlzlNqlw35luKYazMGdi
Imszgd7gBimxgviVWDEI+pqO75lEfrFf9ckA74FBQMiZiURK9UT0lEbsGc9hhMV2alQM1ce1HvTF
MRLNNYbebksUPQNfpjMWRr5NkmNxTuVgagxEGKPIASj1wIM0yjhcK7/27i3YVoqZx21XaCxn3keq
GXDoJs724FwGdFt65mAoZ1JHGbNcuPc6XcsoD3XkdaN2s+OSEakv2cJj+3qjypwHwkSW/zdjEG9h
CGXvdm5pDjiJ08D5gwl//F8UY7TD3DhIWt0EbsWuRg6SQPgaOaAQ0jN4LxpENRl4BaAgh2OdKvSr
YxS92BQBFHAEkHsTcMNQwK1AD+nkFzrWdicnPPUB0seTFEeGn5IaiuGNS20JZv4a5Uh+OZALlUo4
fT5iOqDUoMDBeGrAUudiE239FyDDK35mpJUbrWSd7+9CbGVoBgRS2etrKB/GaaAgVXUsUKBXs+dZ
Gz/4sB3kO+Xh+A0xyqibpouzLjIeS6Gq5ClvWjz9EDNvjB5Y4heMca0lshdJowOk66cRI4d6c6je
uZ9GrcUnCYQkp8X8O7aw2zcmL7z1A3qjQblzmhOSr+mQAuru2EM1DsSuktIEqm5UDtaj5581zMKC
3eX2xJKrgk5XsaDCHCZ44AD1BffM6eOIytyeiLjuiJWMg69yYKEPfAWvFJPV9GpOa6CbQb9XNCOh
yLU36R4VoPjspY8yCGaHoV0MYjrXtLtnpFJZNZDpDvx5YKT28ZFcxsT15YwbP4ogyWkJ78Ryxs5B
/ArxL/El4SzuwvM8QFZfrMJ2WZ7vwuR106p4PA0YM0csV1cmkCW4C6T3KcxkFH1oQbLqvjupDE3h
/g0D0e0+1LWkd527c2daTbBoxicqrD+nvr6B8bpOvPSqX+1eQnNYa7/rHKjgetC/vs5b2zAed9Ee
lTijktvPbI2lI/WWlPuTq0V6aeogs/J1yJw5CsXA67fnDmXU/WlzTAvI7GWGXnHw7Gj5nRmarXFz
YTHstdTdBRUk5w96LZvf77q9/JRNfD465KPIo/qQvGpo/ljvAIGFiLgYHZNKZIkgc38AQsZjMhEy
tis1BQUkeXmNXqHoqNJeE7DgJbaHYOpEMHBw3nCAvKSb3OVlSk8ypUBNY3ZiBSbVHTcFZRX0wq8V
AMLcXwmu9MyUOdoCwdNCC75YnX3+AARvjDJc5wwP4C8M8YQvZqXToXw6SNUDIi8xDMpvmaluaxJx
g/eSVrYlOuEiTcbzxk2bao4wmSlCzX5cn/t3zNn89LkWB6RVqNWFNgiCtqZk5oyf4YV4+5qzDV9G
K26A05TcNkwRSQQhrvf5BW4AmFqy++cgGitBpD8CNFa3wjfMAdmByhJNN8JF+BzjBZGZ/pxaJEmF
FW9UZba2wn6O3LUTWb78u89Rm2F4NBruWA2FOEH/WumpeOUwc3gKcTE4t7dZUaZO+9CwGvNtd74v
F79RqIRqPEdAiYnzT9fkj7ngWT9MBpV1tuwQD/lhdAcUipX8GZjz3VhS99wbwi+ZXqz3mGpydKLo
qx0SD2tUYc0o5X2L9QDwSq2wBSBz4hBhXXvPFsVTGswzxkeADCLpj/I/RwAxJY1PEpcXmAsC4eSE
2RgJACClMMPHXZVDLCEqZqb7/sfQi4lzMJEdNtdu4XFsF2Bk39c/TJEThGrL6hG1DzLS4PJHWsbJ
bK4DAbFyXahsLLis/4+HSn2icRQNdBJiPSoJJ05CrO3WP7kG+U/bcXit4GZfd7+35YhSRkSladDq
eIk3pVLyCFFO1sKiQJdJtAlduE+iPNCtR/MJrTChjBxPiziesdT6uUSeSMrLAPmedLuPOTyCpBHS
Cw3SJgIcsyGL00LL00k8o4ywFKN5A90yI+2p1rGObtcUQxsAZ/8okcq9JicuyN2s1m0AeLRkhIWY
XgYx9h47jPM3ir0btY5UU1qGlnHDq70YICsrOagssUvCeAJGgjO+BbRXBkJcj2yw75d1RvfR+dT2
tDwMwZxLFwP8tcemsyDfxgXuxZzCqEUuE7jMZBnB9wybY2/Jb02yJf+922UqA0UB8+cmiAMPho9x
fKWtf3zjsihoefhIxTjX+XNs/UvutLT3iB42iY7r89wnVmwjM1Hz1Ei9CuLHuA9tvGkR1d8+rHO0
oQrBaG2QIcqj2mHz07tmVu7Mt2W91DW0bEITH+VfNBGeFrTbc+y5FcWW9S4UgmOrUBJknPj7fUVy
JjtdCqEaymr9CY3qM5IwezAr2iKcouXcomdANnxo7YURcaaQ7GNlbxlSzezqvYFo8RtsxstDRKVg
1fUPWOI/oqAXsiTIExD7fayJWCyAFiJ4hB5hscKCc7Vg5OiKQ0SQkvpPpD++DpD4Nr54jAyXwdSm
0rWoaAQuBZAIdmKCr7X68qidTFwJWy3hC3ja2UwDq/3C3qvTxaDBcDLAPEe4lXy1/MhVLJCXiqqa
z68TPdbaqc4tmN8OlT6HEPohCMX2uPyAdEa9dvmFVxyx7HpVoyM4ANMx3sK3ZVeRed7bBZPbKP+g
tLpxENvVrZ+/cEk/SSJIONvMttjDl5w/wf4SnNgeRQQpUlMhLKsiXh+miehMZbftv/0s1QdOUBMs
ucNZhHwZdQS5ZxFHi4/4CZB9xT/IbXhULrQRgnTqyVcztZvM2laEnHrdYxlbjoGaqEbjIei/gcXd
bWAHvsslsV2pt45UTAtJJ4v+/iMWw+TiK0IXbY1CF0YSXlOtNFgbn/XW8W78g3M5oleq8/5prsut
Nfld6ty7rsm2ARY2r3VjhJOIvrHR+4OYRwIjyOxugA+u/fwhp3X0t1bPYGx50WXrSWObBaFi28K/
71JHSaCv6yCsCMrreN8DEovx0G+RghhFRkPKXbw8MP1Wk9gMFZv8Zx+4C7amUX3G6sdT6dG5vuyI
N+43MjeLQJvPgJtSrxxe4dsgNp5lA8x94FogRAjXbSu1j73jwMrffVGN5F3gjBfE7PN4Ofs5C71h
ZF6B9md0oBS0BX3sIZWRnroflnKdlGRYn7dDO8TVFaZbTx7rcm6ka36J8j5XGyXjZNHE76LoxDp0
crsHVJIqp8HHEIG7rOkvtEBFSCg7pCTAz7kro3i5AamdKSjO4W3u8x0BdpPXp12Kz4PAPzVbdc4Y
KLKGzkkEjo51NPyFSKGlvnD/SNq77TwGQY9CzMCDxHgnVOPlt3n+7RHPb4Wvj9owDvyn5KRuibxE
QKNMiuEYLnqVlPrN8Ieb3q6WA/Im4UhkDnXYd9vUmTqMqvHxHrTXIARP61ViwCwX0a6hcJ6G+IPA
D9JA3VIpVfw7HEk/caqayTqkq/qNfXTQDEObhSYhyXy/1WwDFmdMpGUU8cIAqhuX6f0wcTcw7G+9
LJwGSxUNvVnuUnzlVW0PChthFf8Uxd1eAYU8l9gVm14hKEmiUTa9fftjWMbnBO6H98bGlgPb2B5t
wii1uSONOjr+BEebksyC5C1NZ61lda5Z8KprLW7yiheYUFVlvrRdXYKI8+dnIpLxnuIa5/e0Wo7O
OczUXjRJ+Nt3zFH0YgIC5t3AjcxArnr0ogZ+zCtV/psEL60XzXeVOxnqKvI6bE3+JH+DD8XIJ0ua
74reN9LIqoG+2A54EeKn/oBST23LsJwUDM3Scz7TNjevaCHWXjSuJrn5O4OaXyUuoByvB1ZhSEAq
tfmB0u286/qFTqKvulipeR3A/7IpN/Fj/fsng3HoeTQYOKUNxQJtLcpkWlKKpk+NMfJ8m0QQQIuR
zOIdne4xwrthHHlzLLCQWQ1jqz4rf6iI/C2ZC7u8HBrOKM1n3fXQqTKbfspp4Fdzzc6PZjqa7aOK
ddcdo7jx+Oi43byVA0/guvOk3d2Xk0G332ZCio37j1SolbFlz8Snw98jXXet3+0PYvOhzayed7J3
Eo2HTYi1kWPPDIgPLqz5oa4KiNPU1yZf0oH1kdIhTX3QXJM5EiHmiOnlMAIh3zTacilvQB8t/7Yj
/GxOFOd2zl5y6TJ2nGxm4c3LiGfgV30F3oyla1HPTGOUs+Eas2MztxUZCkFBrqsNsqraem34lW0e
QC/WLFo60WqY5qZTPPjdT4v6IeybLWZ/pcmSoufE8sjWUWNXlxvBv6NNNs0LoKiwT7tcic7rvNiO
sQpGr1npaVuO6YFBvxSFCZ0+po4EL67F3KCimZP70P4AnJReLlH0nUs0EPkp520IUsSAHiGk/Qpt
zPmEwDu/2ZHieh8NnQt3GaDIZ/15Bvk4rJ7L1M7U3HMU+360WcNEmMj1qspMXlb7vj1Ay1K/TruT
Km5BQO+MAjqUc962UT39rRrunNe78BCJbtrXmkecbnGWTE5qI5A3AZpXeFo6CB0APItWnwavcAmV
kOTsrAOgpni0mOtSz++c4uc3gC5bGhaKv1Dc5TO96RduLZQr0LeP1gwHp9nAkgbbWmbG6d3+R6Bf
lKWF9xTAKG4CvyqphWoIHoHOmvbHQYaiw+1UqeFj87x/+O3xjb/8FhewhqtsR00KklaYaxh4vk/W
JcJWfPSugeXlJA+t2Bf6IxAyn2/d5rLz1QK/bbg1V/ulP3f8Bfl6QSHAoMar9JqjmaE6nfGWL+gT
HurNoOVK7z3/wWszKQPNXoGOl1/wpEzvrwbWYC/cZx8XI+Hz8hFyYSsAJ+0X+hZK8RviB/owZpaK
VGXAdftDFfQj2OIgeiXwWP9rN7EGIDe1vCVNBzsg/tkuZ7mfQNkSYOEQyXw0Y3n5v/Y8VkAP0dqy
YruILzsgd9Ez4lonrhmc+ECACA/eU7n20IU+uabaZwlrPqA7nuW2lnv3b1OzXD8iRVtrjtFyojLw
i9k6KrRvpI1PUrpiCall68opBpQFaw0DX0oCXRST4Ms6bO06aeZHvLBM+dYssPZiDzAhFqBL2srl
wV9CYNlq9Lwjw7L2IgBOkd6zDTOCPiCBD8zKJ8fmJR+f2eq1JtDMhlV2fOLi7BhcUg1bodd5LCwH
7XcwCUvEJZTHhzIWC2FCOXwB3RpG36MeyITDrHOfyApUcJT3d3/av2GYCDMCJh3svMEBZOGq9DX8
ERH0fe3rNYegEL7a5aQY+NuO4VqNMXltUUBg7hPkd49uTNUmEOhOQzGMsbpDkUu9yXg1VgNvSgxu
2uROYcbpU78vjWKAPSKa7pr6rdn6rWGmh0rDtg9BdI85YBAQ0eKolbSOYijssu7FLMCS/kJFemcb
bmWTAQ3Awvg2Zaan4M6GyrxJty1/6HehtkxeJDg1pZwjI2Xlo1L1de6kF25+NEV3rqcTNIIhv0J7
cqqvVbqzMoBObipJXWQ6UE5U/1RaX2/82129g+uGoZndyq+nvLu0fX0jfgRD3lw5qOQLMPV+agjV
tLEm0THlMA1023LQ1ZSJwi6hIe80j4xvqbJbnl//IdLytf6jCHsDHY2Wdj+C7QjknbMI9pTbLIUJ
WS7v/SYEH7e18dIQPnYWSD9CQmB41yYYOUYB3LanUTtKsG/TEXB1LFZw6wXXRgNqZWm3Y2iSMNE/
7L+Am5Ge1j6ObKMXYzBLZ+uCmJvt5uujkl4Z+/gKcSLsBxim36/6t85Xk6CRadf/lBYNlq/cWmt4
QWYeS8dE27H5Sf7y3Kqa++I7daVXLng8bbyuZcOMoN71XQ9Q8iN8al8fK5XvXKSwgbkTJeoeO/Qc
bDBbMi0ICL1mmDc1I/WG2jZZzJXyw7deDuDD/xaNW0NaY4j51Dc4JCGPWTf86mZUCOJct7hyncLk
R+5HXn7yISeLUPv1hovypvNwlgE17Vu8aQ8PVi5Ah5byD/e9GCLnCmzFvTfYXTQ7JnKfwPUI+MIv
hvMX0wxcVOoIYPHl9gDGHeYkpBLSJNEjD1Bxy1paDT/j8eSB/jZ8z3cWyZdSB6ikgilsEFnUet89
axEXPT9oh+fhkhXol5PILTzFXhry6/FErrMZFGHqB9Xii9GAvbjiLxVOy/hXItlL5x33cfZbyO/E
NX8cBNHc/F/rhuu33mBIglSNTki42XeqSdOvUC9rNuxxoob3gD9vCTwnvF8OTKC/1iJbTmzo1iue
oF/3D7DlBAeAhvUuoJA+Kd5+aGYinD//1PzW6k5hEg4pMNtjsUfBVn22POXbt18x1n1UueFP6mH4
VmQlNXO+TeNuU2gAV0/mMyDYQUht7G1cvRVzYhOJXyWS3wJMu3eva9aWxRjWI5akP4z6H7FqjuJA
HzwzhmZb7xFFHvN2tEKgo6nBdDcZg+Ub5t1olxqDqjHhxI1d0V6c4Lwd73k4uEBAz7e9VrPAtKPc
44Yxm2ojr9AYQPZ2R/BVa1QgHdsY1M6ayD5LJT70mGc3Cy8plIiMQlICZXZnDxIztdyUOjriN+GM
z7Nd/01Sgw22PKtEBmm/7AJfS8SAzIWVI6Cl3nmLgaxQwM8vIIQBp6H3RBmh3WGstBezgyPBpRrM
3C7Uzp/Yy5tBJD+NpoL6D19e8SJGy1I2pwuU0CG67YnCYCjhqU0440X6kF81VFOYmuAFk6atfPLn
LQiVQurE0FkX+O35UP9o7MWW0Y5Aq1Lqs5iZSAUUOOWnnXUYTZNxrkEb94JDD55QR3mROe+qGSen
FDDh1x5s0MZ5G3TmfakJeikke6RifgZ/Un+u9WycKrX7hXEPS1tMPgiZUwvmpufkBg3+pbuLbt4r
qSEAzbyadlt/gF53ZflktNshw126ZtFDhztoyUVCWGXxvRnEqOf53MvUKQEBfzVdnmH0jZmVwHJg
mq5oAlvfdUvHCbfXa5+LNsO+F9i6k0uDvYf5s9Q7qv9XpDvDq+sHZeIaody8yYjhWuTIf86F6ulQ
yYJF+mi7Jxh2RbQeksCe8ijw/6rsthyize4t6+tzCq7KQ3kCSTU3jHQQA+4Le1U60odVnds7FJF4
p5bQihML0iWkp9r3m379wnzKwaEjeNgiga4YxoJMpBjiobAzG3lvfnTb09f1/E1ZMFTt/EOfSQNp
IqUriZcvF81DO8nyB42z7V1idRPt4zYENd5rzhOBwq77YbK8GzoVLVkaePQn+rJxuseRnDsoD0o5
OVULkMDX+fRBwUhLB/q4OMSSp3s9vkvz7A9Y+ZIF4mAhbczCzD/EQYLHf8vIKJA/Yfo0ICNVkPp1
qyqC1BQLrqYk2nICOcJzbrDpH7aRthOfBPEvkyKKYVy5v16wOzoTPt4xGrBZuXCSmKWV8X9pd9HN
YR7zleU1F+ojavsDaf40SjF4rqzMrpoLysSjxzxt5jSKPNzuBMvJKFr2dg/DWb/kEDvz92Pfp+ZB
CstEMOjq4ZOzuk/CdRk9K1RnYmu39cz7mYPGTBrgRlJ+08O5tJPM9aQrje50xDWhE3AFPx6DYbll
JAepVA2bjIR512z75VI0oYCoik55kg124T7j3PSv5uoCJwKVL7b73Q/IYj8ZWlUx5lILmwyUEjs5
3rZ1N+RZFidpNr8XFKGpjWKy6GUmhVSuMONPXqRgz+0cZ7tCxdLjZVMtTIKISX1AZQoLqbvpRLpy
4dqIXU8ofNeJAdHhFvO83DzKqm8DyXde8Lk8rDS4TuqPi4lMmK/xOTPyvh41h19FT5WWdDyaTTTu
ZgnyzDj3S39slW2EOtZhOiJtFxOxGXzu9PbeQIWdRsW/l/8AZZE+4iq6qq/PljJgKaeaKeX9VYIT
a8pVeHlf4lldRcG2+KY9x26I4dXsByK+L7zXpTUWh7Eu06eee20+iBMZZtW8vg+PBbxv0ncHTQmX
Fsar14+IAXDscFWhdX7qh7zcSmvjmMmCOs5PRnWsRdIwoOsmo8IS6BK3Fcer/oTHEPEV5D+p0hfg
0L4ximqzDyEtpeUNKBUcrgjaMh5LdoyiXu1lSdFGcgrVwbHqSUe5Usi3JJQV+WJ+tZSj6tBMJhfS
v/QutRI2Vxqy4Ts0L9AFF5flMM+QbFA+VxEPajcwI9ugeBqE6VZPcXyFHZdq9X6ZTeFy4A7zcXt7
pAZheeWK2ONjPQDyFcfPVInfYOqDAs1kbf7jbNP8/SQOaI/il1L0ZVSdeCpT69JfA3uI5C5vk4Zi
fOIRV2mnDvBq1D2n/iz324xFk/04Y14HurrjySsP/LLUuAaUQZerIpopvNG9tW46UhyyXAMGFzlv
rhFwAf6ls6GtwlSQfv+b2VT0SFd05b3+1d2G4UbycyGauG3OW9wwbp6v2+6KB0qadPFapDMTbQRb
nKSX8QVtwTsoXV8YkhjSPxWC781vwusUvR4TOchkYVlvbr4+G0a5MUhk1w9u5W2Fb/YevhsBLXU1
2K4a0Yh+grAAWMOHcKZDi5ap9TLCvC45ugcsEFWo7pdyG8SG89ippVha3kmHw0EjV8I2lIRQpQfr
IZHLZz+MlWIdT928rS9oyD6T2evsNdQc7tRRrb4fUFeG42C63kdGynPg3XlggMnc8zEYuzVcnxbS
1a1jP0XYZyUI593LVnip26yINFUiRVqFJg+ZCOSNZusFzFDv4qRmDzayXXhqY7goQhXUH+hjay8T
k0I3lZqBOUPHsXA07iijkrxBqlrueZHnRqEMjCAh+2F1Tvi6sDd2cOygahnxB1Nw8InUCNN40Hil
VxOqcfO/hSgVhkqiAAnC9p0L8et9bxzFcKzArbp2W2Nq6MWuYA47xGXmXngAQ0GRS2/0j/PpUpUJ
FDtUx7fd+YY36KQyye7rVkguxTyFJMCH8MaQcgpEtQcNDIwSH5W87ZLDEdtk+gwzVcAYrGHRulyx
waZLqlnwxGx1ewnvoOnZONAz2QmsexS6fuSozvgn5f0zlvuW1BiyYSbcB/R+AJVFISfBukutaw1b
VnCWxSh7A2yPsqG3GOSH1dZRpwVGrZWQwL47aeFzKrT9dHPeQrU3ZsZ2fPP6wgTSK9nKTCzQGbAs
jc2Nld0KfvMR+U5lnOjas62IRIi0aOx/ASvUbBWBEdmbe/naG+MGjzISg/Fylxg3JTUdNKJSe1gU
y/HoAAr6JGCemFtcMMg82tBhQDgNf2hJRz5WnMy/TfRAgXvey2pF3LeKF1GYtGTIBEIsMibg7ySi
q95NcEy9S4wxZuDWn0mbupAaaa0UD0vyfLAOHK4hQTFH7ddNuFSzsI5GE0dCil71GzKz3CdHEshq
XyGVha6EpBkKFWiZ2ifC+oSkON1qBODbrWzTh77LSQuJIl6xl7gegGke69ITzBfm+D4CbDP+pU3u
GGIt7mrg9iS8ji2adadrMw4XGoTF8h255vMaNzQm+kzknG4jtUweKAJ/L4XIlZ6p1ws7jmds/9vW
Lj+ODMFbOtMadIT29H06zhQamHxshsxnZkodbR7JT/J5YjDxVmOm9Hg83s4m12BAHkoJnRBWcwPD
ftYFL3ExDCptmhrDk7RKg45mNB7j6ntE8ljGBUiB2JQSLiTwnYOrUa6vNgdepO/tTG9CvdKUafjU
7PENDu/Nih0Z20wHvu1MkipCXtcC6UvIhj22xsBY2T953nE1IecadlBt+cfQz+mFhUftxg/j8qaz
hQ33ocUtQDsotAgaC2vUZIZH8yRCZm29M3H2ANuBZAHlgi0eW6qvfxUQqs1Dx7ZrEvVLVZgNlwMU
1MGzzQUugKqVNd30st24WZXZmll8nGqO0OYrsmeiD6H2QefFEWxr6xiUBzeLdXK/gUuDW8UXNWCc
rpeVaRKWzqU96dQ5Hn568KJFj0IUR/vx4xPvZqStetyX2I3QQa8nj7hfmKVNwr1/N49hWgJpEdY+
1yIwAPHuhCET/ZDUWDxW7EIRAI9DlzQcXKYr15FDqOdZXkIJvozkzIM4OjAc8UhyJ5CXx7nA8xz0
b6XhtNdjuhrIrDXL9F9oY3Xn3kEUeg9kIgt4rwNnme26QGaRbDEPJwzs6WTwwLq+huRKJHVjE0Ff
K4JcfAEYPejPleRV/HGWloNmCD48Uc/jQBbqSleIgAgSK7JzV0wk8Q5LaR0wI6rOUYGQihiztHAV
7cb9FoaF3lQ00UUw43F7sq0+eChweETGJA66bKvJZAlzH9t4qdlIV6m3vowlgPjVvqWl/x9v8NYV
C7J8BQhSBWwUDxvoUsnr6oMMkBFfmiVw/N4TPnEb5FzMsyHK/bmuA5AM3VVwIDG2ADKkHXu5Wp6E
Mo/XjJsJPcRyGU+GBxBXvUv7w/rCS3EMpJmb2r+W2HdSBXLH3ibnjWEKOaC9d6JLJyeqQAEap9Dw
yCWyWIC1ogLh2APMDG4/Px4oul9TznwXeV4jbkh5K0kzRR4HbBdeEAywg9R21Z7ywyQa37nalJAM
Ba7xv9lne96qEQ3b+AaEGR6Noal6H1bYu/7IwtzApUeBa9fzJd2zbOnCfWCQX/AQGlAj4rqNYQ+U
/d9N7smjxO7mtrssXclNjShvOlpsLckgtEZh5l3FL1LqpN5dhdzV73/4R+Z6eDH9RkTzwxvcGvJr
7C+SEzii8dDK1kYNkqK1c04+UftTECFRbD8FONoolr1y2HWwfbLzAlnNYjmTBDXeL+yHxDuMHDhj
Lc89kzMhRBD+NrvcOGfum/cIzCc9fAr15BhC+xkNqo+cO+jcvUywqqZ7yvGA9CI0fdahTRdch96b
AUGbdJJ4t1tMVhKOeIPpPKekY3VAwXLR0Y7xG8mk+EtyGCqBQhXA+3lfZ7utJq9vgchVOlk3cUN2
RF2pLGOlZzNiSsd4l27pgjUOPFQhT89+BiY8qvbMxb+7gVluF7wsuLxVTaPzr8uoHb5QhrSazl3S
hWlI5woRGOfoCG6pwu6b4QWlmjF+hsZ5/xqBPq6ngHlBA3jOfbiKqNYWwHItNTOw2J4d0AmcE6JC
wWea72Y+vnR6Ya3vH/vfG8Wxh2DbhEBXs+NiigAZI+o4MBh86P4Ho2yy03dVSnYHEc+s02R8HN84
WLSYrbUG1hR0InSnWxCoxbmL/kWf62IYvlakS9KsSm4FH3TYM3ajXZaqjz6alYKZscA7zFEbELSx
fAHiPfqLxbJw0/rUQ41bjbZKdjV8zYWAxcA5bDpeJfZLMDKE5XFXPvtzot/fwAc2hZOb+/xPUwmt
lqGW3YDaBnl3R75cg/bgdidTKL9xV01sEjFUCYeqUTUf4MOwVZc7XfjCWgwadBKOSm/yV24io485
VkarApN97AU4xbABDALIcYbYM7ZHfWPuunu3n8LbxkxmNj95VNsK7BFd0zCq0VyIx4M9N2XAEgfe
g6WWZYpBI99zq0nU59Y439RodG5AnSfB22WzOWS5YE3K6soKmkMAAmkorrBDdQvh4xmKBsUPxqTr
wjHka5fcFMHHs5JLKQ3rBI45XMhPOBxPptUFFvMuPwCeUQCWDDS7+IKsT8T143l3mBFhjKrWSt0X
fYoP+5dkZLE9MYgRS3j41/H86/tB0KbiEFmtPYpmiOlfMUN9JIQmKGUiC+jpkim6hhVupXzX9uKJ
EV3+KBxuvm6WTdQRrRID+RsR95iSr9nZYUN3wRZ/NXKTVtI/i51z6F25qp9QEpSQNcLmJsRXcJpw
x+qFS6U2NDrS1PdwI0nm5VlIaD/usBQ8TwMKucEawAQjHc3YuFn614LCrCNDpf8PjIHeCaa3tzT+
bY7ku+fgdecsqIYs756wNCpdCc9MR7pYuPD1khrP/jsg/R5XwkPFHwRBsFIKsal5KgqQSNn9eTih
kZSiYKJv1pBoBsCBM92YRO7v+JNmhqNdsJb4M3IILS0rTALPkv0eZHPn3eBUpJypPQBJu2ql+b4u
2t9HI/d4W7zIxBvIGT8fo2A4oBXHffR4yBkOu83z6W60DfoEU9YKc1tvnX0ZMNXJTEKFUX9Xr8dZ
FKAIPaVIefev72AX/AOF+hODSIYLv1Ovcj/wcbrNCYA4sCSKLGzHRi1Jo7qbaIkXETOJZ+d7kPOP
4kbqokFf9xAllFkvtM35hYkZu6gITWBkp76LNnxe2mC+pvdZmV1AzqsLQ/mpwSwg6fPDhKCRiZIu
czaV9be5ur095CsemSZ3N6ILwb1/jVsY/WiXW5Ig+radJD1hjwERguCe+W3s2FXCybiN63OK8zAw
OU8REkS3zQBMYgDVBimj4UB7djFEGbgbfrgCtfN0//hxfNBSqwxAd0D6PfTGfLWbqRs7ShDdIllf
Vm1VPYZf9lwoPCyfh3HkIoGNlLvigUWpw2AZXw2qvJkfqcf0WpVm528QHL+EB4zi/7EM8bIy2VKr
1hGJNQ2Lpzr3R5qVGsduzWydhzCVy/BpalX02frh5SsnxPXj3qOm3EXTMjm/iLnD9r322yrEjiTm
LNlYcypaKBEvcgfBbTgaGR9YJpDiVla0Ib3ZcojJYNhnva90Q5ZKH0Nu4mCXns/SzyP9g1ZmJfpv
u1pgtJsS94JuIYpkLfHRWKMVP+S3Ao1zjc5zwPbEPxmHVZFExhrpVG3yDXyJRXE4pcnX7PI09mBe
BGC8XsqKfecTL+WsBHWjsRU7MZCbHHpUIvgnjvcuLOAkRcNvwovsnLVziTS0Qe4RE+EPemwlGQrf
u8iNJROo+aZAN93wrgCva6ceNfxvJosLv6e+DqeHbbqBgik8ihRnOyg59/eRz7C6bRqB0zi62SLp
pUPOT9YT2qBrd79VuaaY2oHzv9vMyxpBKVr/lzkBGN5gMaxG9xYufjv7JtueHSvex8kukQTjogGn
xWeyOI/jdNNoTyO0ddmclyubltTwUWzKIbKloxydGQAMBnGjUmsT5ZTDohWrjwgwTjjxWgmQ43Lj
+tn7mjU8pJ0sy4X60PPI1vUkU2JA3s7Kn3SoEd4jWFk+ID4coQ+H9R7KPzEbPnVlO1iKAuT8a1R+
kTQcZQuI4jwloP8zoJAazBUmFb9VY+qaMPRUNaIxhz/Tp6SpQCET3aXAhjYdaAJ+UDPx4WwFnYr1
vwrtaL4iFxKtBlrqUblP8I1l+ajO3wcp53vRWHOcBWAiDPrPkFqNdPH0U9iL5xsnAavoKxCCe0C8
021hcWnZRUuVBkb71yH8W3L6BBfIYZ20R5O1Jcanq2cPjRfQdgPJrvgjyhPD4qKXMfktl0UYywHN
S6z3k1nOLb1z6F7LNd3Yjf/ytG32yyaErIhNij44ZdIxmTEz+Ec9iLA3tTROhg3E5jQnTTfTgjkW
WGQzQkcAcEVB4xhrdLeEDXXoBkJ3K/b5gYY0Yh4L41CmkA+kffgMd7HmpZ5ik3lk4diN7vn293g+
kQA1XQD3IK48aZBivhMYkYRCJvZBFhea9/Vt1w3cDU3KFK0O9UfgMBKCJx9oINBZmmS8K/Cu+6nb
8XMqZrct+z+ut9GdTvvF6r/fCSUIi3SbcS1adwA4IxxqCKTtf/qhmndoRZ4SB68t/3jxhQ+HNMp8
IiPPvxpkkfD0SW2f5LjA5m7ov65XJn0opiXtr+JJ3QmasqLYPDQyrY/IGhPKV/Ct6ACJXQHljNXV
7TRy5vmsPdz9+pBX5ZGtHf4dBJg45LfT+12xcmSZoucDUdUVoQmcwmKk6ek2gJc5sQWBm8BCqdHC
WiDfK5O+VF7ma3hRb6My9L+0PMKcDHCmpPCkhevnP0L7G8Y/1Bu1QNkR25qdAsVv4rQMQJ6SwibD
QZllfDL6K3K1LalDftDKRv3L+4/yUF78ke67xDceh3fX6ivH4ScFW6VeD6q11Eij7LSdMCwMDJYJ
mtVCnfVJeOGGGST3Fh98EyGdzV6pkcFy1JCw1VtwlSuS8x8cGe9cRg/A0LyVAQQeQrWr5GEyCCNp
zmfCzD2pyN1WW/EHxa/e5jSMW4ukLHD2nmFyh5CC7aXs4u0Kdh8wruuXBOpGM13YFHm2CPQuTx1/
pLSYbRylQ7XplVV2FuwB54UueeOWbqMr4GTqQKSnYzzCtuNJuVopKgCRocXZMUUYjXhk7DZpeU+u
03FJMrUz4YzoGGooBJs6MeCTbx+QaJmhJmhtsuMMzcJB1ohJ+sJGI0VMaEphto7hkV/06Hwus+5q
q6Y3qkp6FKJRZB5qvMK3SZKZ+Lok8tWqi8xkmkR61k3FhJ5djvQmz5LVu2ZQ9eo9VnlcqP7il+ri
5EnE7YzDfsdzeJZsrxBJnDGHSvUtFk/FzkAWaQUTgMt9Rzrd0qgOqxk909DzG3r+2yVbqHKQf82V
oaGD032sleaLJGRuDlA07W6pxmyR9gXH71G73YkPKfLygCeP5opoTlxv0l7UXsilfgyeoR0pXseT
RmzpjrMgC/fXS0QDdXXIRwupSMiffXXrlIWzPCcIFubV6VWP/P/7u1AQiEDCEBzwrEXoll1Oy10Y
pwWN1kYDaN3GY8XklyNQTATxE+m7Qmxbpr4Z3Yx7EIVNjKEicUHvi8jBW38TP2p4+CpDFfQFLO3m
C/eGVrLjWDjaji2G/OMeFHP4KPR4JIr26G9+/dqJPxRf8XZR/KX7RPFgXB7Yen/yGjtg4Enm9j0w
5myKc7vFrVNxkK+s0t1xtJU72ZH4MHp72EwsEF7WUWsHJvDc6zhFPJHGakNK4zFunI/J1q82NF6m
p3xpJJfJjhxKVrvPhfMCwMdYfXESFYGC/uK6uzSJKq51zw1EGClpNyo/61balveA2hJH9WYobtyH
9+bPGmrRYXuzgJuHP84PgKkqQfJGzgtvEl8fc66Lw1odDCKyUEh1nfkm+rfK8RGzLIGIUack47d0
jG+TaR6PeY3ApcVEcL+x+eM2z1b86oAq3+K495jPfQH3C2FZYaWXX2kG1jdnnW2vV+6+jAbIvMKs
snDRC5tnBoEUwYb0e9xGywxLA5OaTdFrl1jJoA9X0Nurq2grG9hWS7ZGNtjZaoLs4ltlthBfb26L
MrCz2/ARzY1ovw0xhOdwHvsX4BnnXRn9WczTOiZlLySKUjjKcFgqq8miFaSiUPwdMAxAac2v5l/0
trpNWrQtLJ28kX3OP+5Av+lpXxEpX3RYVf9/aTIe74SerjjO68/aQB0mpyP0MTfoxzNSicMyF3Lg
yFGVcy3kf4D4/heEMF+DtdFmvH3TdeEeAWO7Yf8Lj2DqCVZyKqOpSfktWadTOOqcii3PPZdIyf9L
bhOIF/NgoxHxoAkWxbNKbXD2jlbwhRW/Le8MyUy7VLtvX9G1fR9chmoAYTOy03SN5LcKz6XDORp2
PsbR79LVbFVHZHdopEaB6yZFgPQA7PEYH3RAxyw3btyyU3f0HWJE92UffW8O4gkcR3DRALJm21mp
US9/Juu6cptnuEoORQ1ad5VIWShngnxtoVSdAj6Rsp9vlcZnpdAY8IWo/JRRHM17N0R+ar8gMKt6
sT2/W4shpptWFjFBFHSqYp+TRjQ134IImMHoSCo7z6sPEePOpRoJtWtx8ehOFflS1Tm/VWErNQ36
3YKQ1t9UCfEigJGyHqa7THleJ2zht9M4fGjSVgsNMWzzzGQelCvXrE52RmKk2DVU6L1K7r/K4PWM
n661ZHwuzbJ+YrsSIVcEG9ZUHY91Sbwt2iD2nn3uk7RVe+Peb34pY/+KW8qKyuqko3MGJwCuB+Rv
H2E9zbbLSD2km1JKqJWCb3+iCGZbA19hlQrhirDq3QZnjwArVBiK/XZoBWqpBbhLIGZeZg+pncAO
Qf79VgvRUJWfeD/yqZgu+bPlf6QNSDkVmz6YO9anrHSX1Y8rOWuDKKlKP7HQqZe1j0Zx+of8S7L/
hs453pi5VX6XYfP9g4WuKKzQM2h4ai+9UzE4CPtY/fmZfF+XbUQQE+aUwOb9jK7DQrLVfUYvo7Mu
nOzSjThozptKOtFDAX2kygMk3hh8WaT6Nb4J5emMmufad29J9fFfPR60/fk9NRmIeBQtOS96MbsV
/P1Y5OoRJWljH73Mduy78W7ZjsnuaiekgxN8NRFtKcgFsJBpqwpNeJQ1ah7BlNEacz9J3XSmmso9
Z/vEXkyKlPM6fo8lieqkXeP4Opji5rmXWkv7p3ICaYuqhqTMOcc1HvZV7ox9UOUgVq8twD/IEcGo
7N/jepQ3yE4CSyp0P6sOvNPhGEGVxLkO+jnaxibniArklVMEayn4C4W89nuw4PDaLplyzziKA+dM
VX5Jn/S2nzFAP3IVMPTY+l3FgX+JaqEs96iMwN9uj5T50N4i0utNdesUAPIkUTF+JLV/0cX6zDG1
wURL/4m7YN03hb+IEdS68eoK9ZziK6fqwgSiaGB5qUI7i+Ks8kjQ8LR0jXt7obxQehITG1nsUNPs
78TdrLXcAMwfUIV22Y1uxX+WDbbj6n1AZk68UgQraPDvjSaHA3BfoPN7jTKHmEyuVvbl1jxZtqKj
xF0KTzH+30dC7YmjCVA+SAy0vednM54kEzzPSWtwVplZ5q9HYHBg3+JmcYgaqf+43VIH70kZ1f8V
KFCL3Yhdjkj+pELkPbGuv8lefro0J+Xc1e0nhSTM5o2SHYEuPnCIWzJHceE0pS5WEeNXjGJN/SLn
KKR/vAfwWJWyvDUKshq87DlZbT72/wYoICbTksu3tY0BG3ywxIPZsBpoA3bt/6XxUnqhAxZuVqe5
1i0mkhmNllurn8zaCAIQkAmlgRVSZ/O6KocS6hGeHyKDX3fsGcXstAEw7wcAcZwoe72AY3kFtQQR
N/fQTMnB9alaHGaPjuqNM9slT+hymmm9SxUNaRrqcZHW1uFSRH5bdp6gX4zg62Bs87jdymYpPwqF
5W9NIXeHVa1A1t95DMTia8CVTmc4aYWJ7ost8ZbGr07Bp3X8p22NZNxNzkLutq/weNZ8mPZoWtJA
uRY+dh3q0PI2zJAz9PiU0SVuhp59OXuZz7JdS4XpuwDz0VqcdT77BdNXfW3lFn7fyIE/kM5pFFIW
W5v69sHiBuV0Me3hsTEqLPIeZ9ONuru+Zlnp9jG5lNT9qh5Jp2SRnQMIBoNTlzhiBfo0Ye+Mwhjj
irzIgBTDbvtRVkmxpveVY/Sh1j1cKytoCPD8In0phkPxfsjURXPD99J4M+GEIfyFaCCQgxFIuPZw
7G8nAHDg/6DzPP9vYn2ETZZJbzB8e6RQkbsGuMi2YbwphyHQFDupCf1oYyPALi5gNFzKxEndsrWC
qQdO/IylwsI11SQZJSEX7Ko4JL6ZY0G3eVbgEP4F/euA6p35SOwmAkWjFiwJpA7ac+QFtkGf17iH
NfbLutzjJsS87yCo4uWqjGwFcFQD2chhQhg3k9AFeq7wldiChLfjy9nTMpXBXKtR42Le2FWhDMPZ
hGsNMFiAsQFRrq3QH0r24mabDTijfRGSN3X5LW2YfTamQ66xUU2rInZqOp+u8WIk5wBYTCWsluPz
w0O2rbSeCvQeQaUlhGMMcoQECHgj1kei1FTqkwmnNhyvX0ft6E0P7fZAGLEs8aB8zq/oo0MAr17r
0hJoraT8vZo5hvK9qHbg9XfRZOXPktuz9BJP5wYTL6mYv8+mJGNcOG8POAhn311uG6cU8MqGLP2O
JGahHbft6E5u4H1pMCBOzXBnCfxvYKiqRII58nokVBJ8iyrIDZZ6XU0n65Z/6cHaZX2avHxBMV1b
J4q/LMFtfiSMqLwCIDUVXakFtVmTkrZV/ofbuZaB2bWjIlz/ugv7HlDHCrlSmjKzP/hhCkKgturO
cMVS0jmNsyuZHKiDiV6q+gaNir1rVrrTQw2ckPHDerEvcub0dtp/Bg0xDLZlW7Yuw9aqA4+W1rgd
d0q5yZuASjdpIVaP9kVm5OJ1y4oq154RVO43618C93wukL5ae7BqMogmHGNdn6nBqKeF6SG3emMs
Ic+N7wK0OLlouZX/ZO93eLB9N2eQ+KZ56jilv8GJaxVB01yExf3TqNCp0LBYqmfhYwrgGrAkp3zP
w94dAFRlR43hlvxENY7SDl7tVTQ4vY4TXynxUECSKNeZAojpAtQ4pvR7z0SDHf4cCFtan8le9mjM
0l3s/Y2YWHfvVTsVzd2WUZfhZi+sTqCDdds4sQwXlcjmggLREzB2dLz0MtBP1zZxXuJmi0a422Fq
DuMWUeuofJh35I5ugbMjrtKDNjQRgysfUchpIUwpL5cdbLxSuF8p/wK6L6aLcQX0kPCKsPEANmwr
Vs8FZL+Cc4TjK4gboL9BFX3Z5qUMfs33hravhHkaKATmuutLJMmKeGc28sbsaBtbaRgpboXly8Sx
RC1LcI26q5h/jvTd5sF/VNsTceoH5BB85eoauevCXzS6He8BTo1nMRy0aRi4LhiZQ6X1eLIelUGM
4NeB7/rj2JvFh1/LXEEYWF9llihUteks9uqmvG3dfylJ/3HFFioAWG1mFFCQ+dRlxfu9+JoLLnHY
6B+k3CAyiFMo0M/w6r+Z5F0gJw9LeximM5SGM7+KXQ4h0BcB8q7QQW9xAUUnL2UGss/LlH3CCcuZ
kso/ReZBxbfkEajehjV/W8JwODm52od6/11vV4ql9YFVsI0LojvEqG6rcsM183/ZGuKjz+55G6C2
JFntL4lgH7jhlzCVgDUvMxD7iJqbCa0pSiIfQZpjV9J8oUM+KiFEgdTYk4PG7WPzE841NXi9Ak4c
t/K0vtHYgDSqvtrWmSEdKfEfrfRRbVEJE9ZDttVYwYxtHQO6lOIg2inpz6HwahB5sdvQTwy8RtF3
RobQRRlxTjqdG5+xDOj7tzoJUbfsQzJkCjyDHxxQQynGeryFuYPk/TV85grpw/NAdQVaGBNJOe1W
bJPqNIWtU7Z44rUNMK0Y+Ewl19YfStmashf/ilKYyqVmSvp2iyiHNZGCSxeiUEWY6UY3Q9V0niUo
KR9mRjz9FBT0HnKIXhYriliY90duGr5ITyBlSMnehkiTGeOFTOefQxuX/quG/POVGEhdjTDqKrSj
4/ZSsaIytatS2XBjhjVUhyO7H+sJgiQN85+cf8uEfVmeBNCj+YqF1ErBD80XU1DCLa+27F8m7XAZ
en0MFCw7lzZh2ddPTdBRSlzOpD4fN+uO1AL/Tr1HlhO4CkhQ+ykOK3HM/yU8477AdqW3S1fAgwn1
KPd5bpBF8/NSBfYnJbCLBhQP9pnAMdEz7E24m99CLAzAm8SxJKGtU/lZELIwGcsLm+EguDdt4kmd
4BHJc8V7MapDKqI0XaiG7pgmLZybIlfZ8cAA7zMfJAUFU74e5NsrTdH6d+KUfjGDH6scPMX8fYqB
8F8dD9bTV4uGaf5Ly6RLgC6GfK/gR7jkrTzWyJkVvUg5VKu4nwjPlMN8n/ArfPV52PSIUXWNOZM9
YJTpzbwDyT+QGqBFL/a3HwWgv2kozUvrQca3710hQOzWJu6laUunb94ZTdiVWQI3P7Fxx/Zs59hr
7Vt1VBgBiAfIQoEq0DYfRHZSh5PUZ+c57buHhGT3Xu0Pt9vpfaQ6rhQ9qF/Mto/4T16oT673/Fb8
VOsHc8IASjZXUX18kEAf3ZVq3BnGAyhVdwpQnWyBHveSA9b3tJh+kGqf9ta71vLc5R/KildVhj34
xW0ru03TNnUCUvnRDOnLV77KRQuw3HllTT+qo3TUX01J1ZF2dTm4kKHwUGXteSoG1mF0o824swwn
3AMQ0obKqurlxEMp9pRVGR2H1HfhJrNTZamZBWkdcLl7tWlUywLSg4pmQE6puFltes/2fFp09Fn9
ZqbAFxWsLkhRlgKmPeq3YJDwXGueE1wmKSOZg3wDMnshOZyeizYYfjRJ0u1Wfk9DZbd6+/RUritV
8S74s0aBPKlmmHy6p5/MtuZe71LWvk56jQjLmj0c1jsUWR3OyGTCUIO5JYevGe79eNUngd4qP6CZ
ffvqz3QcP+GnI87QTDMatX7zEudaVvX+RZ98aSISz5IeTquJpnKvpIhHvva9Xc4eeRo05AQBelvU
jp4F4ocIlJar0HZAnLKslEAzo3Zzo3zB2ApOBB1mxQQZAfXP4q15NIfFQ0ow+3bV9zvdfK48k8p9
7RHvtABmv+5C969f6Ns/h2G7WtQamwM0JuHMNU6fswlzqsW81tr7pmTEYbetChZfVsLSAoJmqvZL
KJPTeW93G0s4v+OnHZtZl44KV5bfOAh+yJI6VFzXsymvUP6itCRZEJIEbtdAJqLaaIVFLd+nx9Bb
z+5G3P+XuV7hTDX0fVIgcQqGejTyBTVXXC9gu7tnGU3iodOJw3GIMbMhjdJeuypdfy8LlA5Phk0U
3p+xK6n1yCIWfE1ofr/4SBKYIwdWGqS1udS/4B16ZdrcKZuu6S8wfLywLMa0drMxufExbt4fnc8C
JykenHQaciPlu2pojyh274lBrvnuec8xIMXsh5n/V0+MOP/ZlMot54bb7kyXiNUBrZrj9n4bMyau
dhg1uEoz8JBjlrZCMJ75k/gyY8ISH41tZviLZqlTxwxTUTwWT9rQ+SXDYUq2lKyCXOAmDICOaA5A
GUY5WvyO1goDcYiDhekyHIfWAYRoolYxvJMWLZHm52+EU6e0M6g0ZgUYbendamB/sJNKghUKdogk
G/Z3lWWSJTbN0mYyZHgUYjXkbMtfeDMMyt4HX4ru0DM+bZk2/e7DZy+YmJK/EroPGOJp3dfw1Upa
3rCAfwEl9HXwhkpdITc/wzcwhE5bPqMurRiT4QZ1fjiFnQbTrFnenglIlVpCqtOyPSn8CrlcimHR
3p7xbeeoq+weDUQ0eGqNo83D65PLLD4Xnd1YbYjHKW092X1023rW/cbVWRrLBsFw1h2xoLHCF+Y2
V6NXq5dP9NaF/1uPJttL8d74gQDrCCFto5FXJo/Nh83QlfSpEd3e6XuSB3pq3DejES8JxiN+MIc9
qeHiL89u4fBVVYtC9dsPZXiHrzM0m1/11eHVXL+2cSnuNoLL16Xs1fQohUaFnMZyCzcjy3OoUN61
JRJoui2jDxxPKP8F8Rcle5BiEfRu0NQ5NyRDiO52RxN1R7M7DBTfklXdohKNcSbK2vYB7xbv7wAN
xiyvkabCAVAxpcMM90FAbVopkMTAoiQHoGQ3mATIMTu57ixoPtB3tCaagUKzQaj8wWUvo81oSZEk
QbFPu9/LYSBvyQfSX8pQwNDNDXWgwKTuGTGxZmVy9XvUYX9HuP4oA+BBugPkBHUKNgbO8xwZy7Wn
enl48A8uegFX/7NVCNsDVRXkRTaBnxQRjSLWD3VQocD0l2ZqaHQnLZ1zEZgqWHZAEVeXWnwqkdvY
mNfP5a2Y/OL0q2ZtDJPKrZRCB5XI4yK1Yh4eWfygPpZKUr5eeGkbMc0uMtx22E9ZzWHNY24/egBq
aRTDJIlXsysGejWgH1fNPhyB4KqT5LGHMsfnr7eu/dhS7sYmjjuYZLgF1uDnvKyVLJK6A7iTaoZ+
rFyLM/RS7gK4Tjk2aljxBgLhMYInKMwHrIdgIzcL9uQZSqeK+ROqMhBi5ybr/OyKK5w1OGXQgdkC
lIVl0EuOYf5H8ofvjslvWOnmuS70qV+V4euz4kKlqmaWcVufFokGPxkOtfqhn4uaMaDkBIK3cCyK
dsAJNeRqbyy9ITzM3iQvxojAoZj+JPlUVlgSwxjAkuK1On0Vlo3u0DAVjVLKqa8WN/7XkPUVI7Ll
lYMILCrHXqGSk+Wuriu9+VawtnoqCpPWbYBATSwb5nYs+7MFPZYRuNS0fJjwAxnDivAMp3suRrgs
q7YgmRwbb4Cgpx7yzuxwOwPNKJ0Kq5R9Rr/xFopebdlTs1JGPMvVxqZ1BA/mIyZkiUUbEVud4XrR
cOmAgSSCBosxSdYjMBeF1Rx5bnCseePix/3ysJQfeQbRaQjD4dNfCUWkD1LEM8gH4MDV3eUjK0/y
ATcpUe7jOrNNjWdy0yDERUq+wwbCEqaf+UsV43PDrNtWk0WzOgmACT+He2SEvXgIPlUi8Ji+aNHy
nhJGtUtY49Lze1AyKmD06jK9K3q8YzI1vdfPHmGDjUnaCL4ALnnrdwMnfuvJRONxt7nJrwtt0su3
q7yMD8Tdm4qRgMM7jCIFl1NZE/dh7rMnp8hzCBMyYtbXtxtzZes+6hH9F4ZI2XO+ZnSpwrCI1zd6
DBJbVI36BRJCYYczdvgAPg+4BC2EXQi0nrkZleFGpYxa7/TrsIecl+SEzms9zQGVR6QR0/crDRHh
SbXu9Hi72pXEHwC5WriN4l47smg8qA6FNrJlgpeYTQ4izlVAlhdexKxrJ0UX8AE8I4JZK2kE50f9
a2QDuq47gWBftzmTsI1qWg7d+RaKWoC3Yfl9/LQOVhkk6r91RfOYpuMXUC+OWPBKN94yjxsrE7CG
uNkPYtGJE4nskiVVbqc+FDerhholffTyEVoF8Hk19u+pgxU7OHYxlIYPjvRWaIKvrE77qykUUg16
Kl4hft3MWpglS4o7TmOh4m/ppjRXkTmvSZU8dwfkRtPBbTvslDdReN3wp9jJSfFhDu7GmuJlllhd
lQJCAm/dB/cmOz5IPPYuy0eHRZnY1JWVMObEFb1ocHJ4m8dXTl0yOL1x2TPpAuh2e9kK0sN0XlPf
8meBBc2piv1A76ViLq9OmLw+m6Ows+RC4NyrvIYZ8SEgeZ4SjbAzgVn+PrV5ew14xX4q/IP+fUl/
/A6BJzMtH5qVjbI+YQfrwYEm/UIWMfUiXbjgxrXD5sxubAUgr3qKkKbpasufuZ1c7u/wxhXc2jae
DJZRWTe8GYUuGJdOLzOt40KJL9enKefJHVWuTG8oMYgha47TpQlyD5PXZblnyyvL5LN9y5rOatKd
NP79mGpylpf5bVZUnc8NI5Qm9p/38lgVj6tofZ6BAP6lJyNGUYHqw5MRXuPCFDkb5Sa7/3rpvq+C
rvrObofuq23pdrGPjnow5yWBud1DyHkEU+zKv8Gibezd2WzYnvgbaTQmMaUbD1UfxXxiOTkCQMZ5
6r/elLBVzgFJQSRE+HtvqTOv6yO5LL+GwG1gubMBTW3JOqVfsIs5WKoI8wGUNgiTGMYf6UObt55i
F4zAdAIF5uYXu83rNHYT022dPztMAjEwiU93PReQDjGvCAsHwa+VUji6NRdavAAGYHo0OMuExeW+
4rwl+jKYQjt7/DaAUz02T2KYR3H9utEaBEoNq1rtlcHiADsN4yxGL+JEYeaAswuv0asLZxS55LwU
MI5yLbnGX9EzWzoZzdTxc4MBIWcseS2JMLPzr7oB2aj4mtKAufuY4YPCtqMM6jNFOK+SFGZMKKmH
OQxzeNZOl3KOXAYAUfxCMLJ9FnURS31iPyr6htDRzuJYIy51dEVz/8ADmxqs1BC22cFtclbXyisT
ZGGX1e+gPjUdPz62tIc5GQrcIcdCHZsa+eiHA+HzrY83iGjYEkfVqtIhksrTN8q2rleGVOsI96o+
2Plw5k5dWWUBlvX0NZ8Q2XlBlN5f7eKs8YY4P/NyfXpcQFtArVKdt3i9PEdirlXbkk/F1gzfLXXm
6mzp8I6lHQxK+OSSTEF9F0/D0adzhTadVA8aBuoi6z66cqJ7W15nLuZajsQKmPhbWQBTvD46fLwA
0/JacWBnN6yg8eUAKA9MT9rGa0OBQKrtEBZ/pFhCPdUOWOolpB323c4u7ZugeXhQzl9RBt4NtFQu
dC/YqZXkI3se2E5fl6Z5UzeWoAiUtl6ESJmcDSOWX6VYteWke3ucpYx01ZPlAP3+HuWVJ/4+mgWj
zroJiIwlNtie4o23OQ9OjgAzBL4xX/u0gxb1AjCXlkSNrVrbOHek5AuV6B+SbL6z040lgbuKHOZS
8HogertL4SDOGjKgujy2gqaMWV0woCnyYYDrDQbARLDygMkjFi0gBZboA/LsxZivqPECTX5kLOSH
62HBKr2ty0WurxfY6XEQFtV/SoKQtuRnb4yY1/68mrqrj6ja3yADi7dawcDh2+3dcu/FLdUGxmm5
Z/EsywzpMqCo6iOihc3iJDcuvCUQw7g3Ox31NoeQogjH169KKpHEOZ/X3wgUqXRjP9wXgg/3HC/w
KlgExZyg9C1Vcqg+60r4L50uOcb80f04lx5q86Cj+y7MBpYExe9BmG3/rYLpDhV95u9yzl97IoW0
9fVMRURrJdXSnsHGs3X0pBsUtMRGVZD+yHBaBeP5t/avafic3D5Rn/6o7g/Rpr+at/3qg3nEqcQl
Vu7jKEQuqpHXjXTJRntxacepSAV3GGv3Av/ON+K3VTpeWDBd2kfCDIAXCaIEuwbZhSSXzeEMUjr4
6UedtN7fy0NTMrTTD78no74nF4XOaYaG+ZMIScUP32NYSK9XL5+5PJmjLORCpqGtpvInK1YSRLRi
3ef7kp05L5pQFREPBQ/ZU81YmehX95A95bD6HjHNMpBswU0gEe3ekjDwKpi5Sc7eiMaRiItzNVBv
kJ0BmtXh/DsQmN3kUIUGrl2T91QjUSPbTMAqFLzClBlu4tyKJq3Gkf0mzXXlEEOfcMwoasKVrVsn
GWTwVOO/J5rUqs+Ef4Mavui2wuBDX6iw274gGu5E8xT2mpBCuUxtXe3DRNJeEGlemKNxnJ7FEsl6
fG5wyHeLl/N6nVDdltkWNmqpK3oGR+dT36NUMEqNiyX857UzDYaZ+z/i7hsb81fpQKg3nWVHdnO/
FnFX5OGPx6Jd9x4J1OsWWl1afDax9e6+I+v9jpotJ+6i7S3GwMUydrQ8g0kmvbcvBXCIAwJajME1
PAb9NtaF4fdv3WuDBBWVHNIctftRAOYuXg9wClRSXHwWOYZx5QgHpdhGQbrWS2W7CgYES9jCYHWG
+kIQ1QAcDv69UdueOcOoi+FTG/FbB9yHTRwzbMElbjo8h39IHkq+fiiGzAuZrtltuXBD01A7n5H+
V73EKovwRq2zuiZpDLJQ/jKKjDpo5yqmrIEXH4oMTom4kTbvKgUf+DhayNe6+Nh0D1zFdFvuZ17G
ddHa4c1b345xPWZ+hNIp/KwmpVrlz3ICzmtt6RqYni0ee4R/rJEkagPNeFAqIbJiaPRRShb4cT6d
NuKS39OwnBUUI18iUmf3iY9ePQ2uyodVYKqSgAZTw01jJGYaAsXbDV19gtfgachFxXyn1q6+wR7x
RgMv1xs6FnLZRauzldgJohSCpfk7fw3Gx4UmQmgSyiU1O9Ke2fkoJEaWE/GNfT1XeW6j1wSPKHyt
q0dnMKmrc7MwE5pDFNlZm2ubqJZ0c8uDqE2/NbFxz2ZSKJuzO0qu7YVvFR4YGA1MUPt1M0GHaHSL
gN2Vt14HJPP6f1hyBIhY2ccrMIyGOMeLsi2Y4e8jWY8eMB6bjBvoByxq28jXu1mVRMAwmbxx5Gyv
Oa7vqZazjuQsadlYn4BSmIvRV8VwCF5gWCvd1POYFy6PNkVo/Eawhc2uMxColo7xMReq0YPWkrF8
HPxANnahOicGFx/yBLIDS1gnfLCVRBfgiShkh6FtV+OzvHAi0SchxnYPAFhapVJjzLOwhylYuadM
J378UqE5R+R3p6NSWYmrMxzGfmTxc6Ij0wMF3FBoXRLp38URgCO1qpM4Vk41jSpyEXq6uIv6UlIm
JlrHh9KRMLKvQDrXDp17vqQlA1/+l3h7E26lqi9SEN02iH23S+kFMpLq5KqkIFWOxw7MEQSIzXB8
l1KVbRrwD++KNtdbaA26ndmmPn8FZaPH2y7ug7bYzKkEFW6GnuL0btZM8SLkX6liZCiJIxg39B21
ly51YMqicgFrKmmCz/zvNUmdemCNnPz2OsCbDEVQwF59V1ki4vTvkTLYs8yjnYfQba4McpEFkb0p
DWWr8QQbiU9kOg5IqGnDBlnKVVAIzQFxmAOruxx0uBvo6BB+sdWge5fuoSyRfKtTTExcuTCa3OL8
GlDvK+3nWKemWlrAkGGqpvRL/vLOOSDAUgCedKfCi4K6r3U356ZRxqyhUJxbdr52XgFAqnbrYOuJ
CA10JG+3dcuFYpNVRJ6JIzaIZcczUosz2gghXr0fG20bKzjWIbwwGn13K5KSWYHOvhj2XAXNka4I
xO9WBVo/TWW4eWf260MamybhQmdiLMu07WMaDNhPAFbfx+VbVf+a3mfOYeXjUcWE/QphyJra64z/
RXA7IjMQV9+TBwjrXi77yjKqI4wac+V/tFvqsvso1h23ZPoD3zb/ODtKmMi7kLkRyK+zIAEO9Ugr
qoWePcUKSploi3lRUQuHhv7LcUdVmSPRYoAnE0eNEV6CipQdJxxzXzGAs2sefUiIlpgG7pKRi4Lx
pZX+/6w70me898gcgD3dutdChNbh+rofPoSws1ukLjTspB717cCQ4PZ7nzOyYche/OfOK2oLRt+T
+kC2u7Yl+ZmG3mhy8xQ81fvQOppdMUFkGiDP6Yip2vfjQIwj+fQBYkNS0K3LOS4FdDAhTSdulp27
8IycsfqhLfsxLhFT0ZGa2CA1spZ8wJjT5MsA7neUeG4+UyRh7oso8/4CMnlvxzIb+s8VzZeKLZc9
M6WpKPStabdWsG1URQndqfEeASPNbJu770G1NUhUIwgA/HQeY283b+sLHvCwJsUhsPzAHFLaPVIb
4KTIZlea6wbfovH2QFGAdrtWhM08ouSDPwS3Bzh7EoveOv2ngwy5N7AwaNz6lcrU/E2+pkWtKL/F
VO14fgE4cO0x2/Fze5O3mvtitwBa89aIcrX+unOJHpGPv7rUXn6u9V3X25oxArfDmW9N4tMVGZwk
fmERZcK+pucpSi06YHDTpOAniEOI/K28OaMTESK64Jqu3DxNAmdKdbzt73PVqL6Kn+7gpFpH2NPk
ZfVHQwR8xZOUONzknGg2bIsmyxXSldmhyXebKtnYPWQOtJouuz5vfLPJ/KnpFsWGHDxCmXcB4RI0
0i7NMXF1T7HI/gvFp464RCsQV1ccCjz3xl4Rhf3oVs4UNYoJ7lmb6gAgOS/XsVgsi19GHt0KTbDG
ZPll/9rZ5yYRA4EX2llBXKDrBmB+IjRglTdungipedn3QXb/BI0HrwJYuefNsNpR2YBO5RC8WCWG
WHd41lGrghoXnORxuv5H/oBgqDYsaX9xCWSz+i3hMJZYzPB0nVqa7M/FYGSECmXt4cAVRBdGGDhN
cWu1xpJt5WOJ7VHII3Y9KZEgSusfPWpCSh9SdWFpiApCkbP/8B2LyVC9gUHLW0Lb/fjqpPW7V188
b8JFD/gnnpVehoivN8nh7J6wIkXjGAFYpyb1U2Jxzlu/3i0Bb0iL4RnBgzHXY2zQ0L6+vAl+jD/r
DouKfoAIl2r9o5nTXsbBI3A4Z6ULtsXiRqK6i7wPh73JYY60IQlyrWiKgt5z+bL9svQ02e6h7POz
4PB54PZ52fWTDuxMmT4up/khcPJFr4FyC5CmqgSVtMugXYP7G3LFS9jjFx4c0yhAjIR55WLSb5t+
RIYjW7gkQgz1Q6DghzozinCNNuzGsPpnJju/cVAXOHm9hkFOgbjO4xsHv5GxAsVDLeuVkODeHLiX
fc7dOseUf+48fDMurw5lWwZZNZFLIsJYKmtvxKON4D9bxUDSt21FAIpztJo9AV/Hl2jnbV2G6u1p
KmDwwQIjcPsztq0ebJSUXWIQmyBsdXwjVU7TklWvtC1cmM/vSW7wB6axTGFRZ0bMgm0nDGGpQ4Lq
2hQ2AFFfVxAqwv4EJsipANFgrmVe1or68riLCcgQi7CnQMOfMrMwXYhWSIpgsmJRR+Pp7DgGrOPT
qirGZWHJzvyVPFmfPkLHh9zuUibCEg4HRg9t/hXNbUXxK3/HNI+zzKU58f3HAxR05yTWnusXgEls
czhBjv5Y87/1augGyIwQkqZK4FyNICDqjzrkon805iQ/C+35aia1fP/honE8hxTswe1AqstFIvS1
xMs6lZtERrfWNg10VGdRaIYSW4XSDLQRMB0pNmyZgAhp+Cxh4Go4al9LtGaHt13GA/2P93hHdXLm
6eIodAEMM9OiVy2mNul1He2WSjdLx3dixUxoPY1Es/sC304LtW4MbPD34D8uY28y+fEUIUbJNxUH
CZ98Y9jKz2ZnX/gxaIQkJZ216QFsfeGhaDDgZVjisdAIenCO0t1L9TduXrhCkMvrZk2i1fD7syRM
tfLr3XvH5H683rppoVlGD36ZRCNcfGmsdDyC0L8sLIt0tx65er5XG3J5nkvjt4CndsSW6qU3Ee8f
n8x7/+rohX47m3C84erl05CFtnNNxvVJV++4TuAwYaO3A4wYjTu2rVMT+dllA7GET+oqnA3U3cB2
g5QgdpNIjvC4NbTSlMxqQD94lH1iJYv+lwTVPOptjP1ZbqGtsxoDfYhlGLW4InE6MrMZsg3gvsVF
Dy0bb7O9PrzW5gpojtjpt9/U27vyNbJZG7yREL/+nLYTx+kggZmbqZHt6yuSzP9wJguQ4INYGI71
eYHABH+pYVd5vGhtkub05rMq9VbcH5W/iHSPQkCggZrsrN2bLH3J06zIL+GZLcy4v1WtgTwpfPyH
rH+iO5HIOsNvtuwdfjlsAJ+7rENOG7cKkmQ9ywKSV14wq74xlSSgECmLpQb0rhUu5k2RzfgQEZCZ
Bu1K+OfqDoQTrK8Lz2QS6MtRo/zDCl9ChenvubB/pCm+kLIE8zWbhWhq6qCPzGMOdofzHc/XM/Tj
vrAofOoMe+DRbBJNPvnyKp26oiWyWWGTEpuYjF2XFPHP7ObQ5fYWdlJRVbjfREIoL/PuFKnlzh5Z
w7TXzTkU1zlz3ScSaEWaUh0ldvfgwsGiWXek+alwcu34IxWgTNQ2ZfvSUNJ3k55a88Dz59KUveCf
zgHyh1bxdfKPrpRZhVnVwntuHJYZ7UMS2NaVC+8WrInR+laY9TWGejAdAVOddWj0q/v/+9ri/RKn
AgGo2TDg0nqy125YuE9c9iydX2decZBC59WaZV/DKrRT2x8rbPmr6k5eTZhp4fhixdMK7g/w3f0l
GobFV6GF74JuY/+/OtwKOHooa0PqtvVqsP/GVVS48WJGZhqbg1/pSW6k8L5dmLgwAdwQ5163eclp
xA+M+8FwBbwUGcm+X6ZPBWdkFbEwEV+Bf8mcnfKONIxzCwcw2HpwMg+0wBbzwEANKNLVSAz2RKJI
zcIJZz3gXktiAWdgtOhctwMQQMchajooPMS5o+iEplfMqA1YlOzT265c3uWVKFdIhLuJMH/fgIDq
UQE7ND/SRKxcdy3MpCF/EIuWwKUH5zETdr5cgf/jAUVQdwBNwaNM/VPF7oc9TqXo6GABV2iHghjz
aX5TNeFsN4lcB1WOV46gowAaAe2XMpGr5ODv2jOQd3ZVf4mm8Yuae3i0ptBgJthf6MsgQ94cinx8
qhQ8Chb6i8VPLh/fjzimVCvDRkP7voTwLDJOoHLhWjE9EWslhCIC3FhVvnFcBtc8Oq4hEEic2R9c
5srShq5llcBq14cT0jeynq/9nPYmKaG7SLcHNNou6sALZV3J1S8gLYa6bNVm7IkDIi0eslvuHEBh
nBPzrV4esBD+7NNWkuxydcWWbKooE4nN4uaUhoHcGrCFVYr+ROQAZFSJkm7ryLa/dpi5Y1CZUol2
JPTPxNmdxx3X5FwRwtHpUBwIF2+l/NRSb+fn4Iv2Gq7a2EeMGpdJxJb1100zt777vJLjqSfrvlF3
b0OH2X+T61j0SGQaGRRboTSfHXhXj1Evb80K8FrxC1d1QEagTOQZRFezCJriDAk0QMWzGONRgYPk
jrl+GEA4+6nfM7Nwk6Qx7tZKxkwVhb7xfu2QuCGNhNazu7Vvgu2JlLaLblu5Q5A44i5PsEGGWSBz
UBfR0wIWQkuv4EkKDRz2B0X+7RZwD76geQ+3FkHsVz/Z7r9Qxosj9hRpiTuRP71WiHZAg2CqiWUk
6w0vIfs5gaW5qxdkrYrr1AK4p5onl1SyAJ+kvHQB1K0MTZhrHfZDxaxyr2/CEACa+1YOtMdpmAfN
EjoCJ21dJgBUBY0meb4lV0/oVE46+rO2ZbjvacmqP0dEoDpcgKRv10JKBtVOeS37MxeDu6Kbbtj0
cOchcycKWz6ABRefEk29ddA2+nCdO102wqgRzOiogfw66L5b0HFwFlk6/TqnwJzzOFr/EIuV3uJm
aqNa2UWHxIzOb47jKJwhZjzdZT4ZsXk1PsQ5FsTzw5KmvfRPBw9Ls5EHz9qAFX3It6woixGJa61N
TmkrYIsapHziza8SmsTiCh8SAvSBJ2uEqg0sxBRE7h1SBTkl7Wwwlimo8/8l7a7GTOO4Hf/64yS/
5h4io3X8Cg9jZwkghKNrSEhwSF/dW5uZ3qvVQvn5CpSfln+nWzAeJRtljoO8vxloEaAaaqtyG7ep
QzGlN0jZNUCGvTNQfSNt3d8nXqAeCP7lWmsKGBklN8+ubMqLN+BceAf4eKEl3ssTC6j3b4Q9gK5k
GsaPuF7H1Jb+xnPFjIRs7sg0StDT9zQxRkRmMM6CFglreSRfyrpAXm/Ma5QFU/kNX+UB78YwCogY
R44cJAI2WjJbImMaC+toy5ZQSCRASYWvfzGNdbCmkv8qgUy/JU1Q8suG2rNGelqJRmnWiNf3frTU
mb5bZxgpB1wk3YEsoATHHQPA6Q87VDObUVa+s25Z07WVke2mHVMHfHw3+iHcBpRrt+mTMIwNX7cR
WT0ZSeIQ2xaF6WdlL+I4bVOM9W7zXg9a3pKhYneJsR32BqDdnqUfp4YzBxRB6j58ObZD7I+aQaca
UzP1LGJBwWtaRCtWJ0dhHWGjkVRi7qVIbrZBrZgP9PmrhZJGkqy9vEWhXFfOHDfsHK4LcrSoKKCo
86+kJ2N+Op6HLMlf4g/3Ku4f1DVt8ANlRZetWLd123rPFd+7nOPH6YPZ5NBMjUzT6bL7u+19czgJ
IeQp8dCyAne6K/ydCJYKyZRHtj8JkrtxqYHEQqPqYvOBhc73TH7vILpx+KhpUw+OAw2xvIRyE0lw
0YVV9yJTjic+AMxg9llq8pHcPuNDJbUst6osx0IjW0hK+pkHP9g9PPX13fUvM48pj2WL/o3uGsgm
0yXpHdYlfNvj8YQ1UJkVz+FvMxpp5qxwBRnq0CMFLN/vin/efiYKE9tvvBBEEQ+EjS2eGpzZQq3u
vklxfhtfLDyBTa3hD59FlyT3dxOXVLGwqZar5LgqyeqVtN0UyrDEZbSeIlxurMuF9xCHI5bQgRzE
IUMDUq14M8+BuycLEqr31//4s9N6o5LFF4tJWmUrpgSpOHteftUMHsJDr74Pd77s0mZTIIOWx/wi
kuWeTSQCwTIpuyT5SJDV2yhztyWvJN3AnSkRFiyMJUpgCpFuiBkFv0Lnjt7M4IbLMhvhTzBTIayF
Vs7my9AYtKn+3MgPvp4NFol37W/8CXfkgh6pUH/MdJ3MAj1sev1yF8EmkqyIQWWh7Dol5VMDacJ5
QYe49edM3LSTW+dfzoLsuKtO0dNQT8b2pngCGj7etcpwebMpkfOx1Lgy2rV6GxCtDOW+3Z6l2eaj
fUpKPLI/QXGPAB05Sl//l1GvuNDxYKBsERsx3RQrtyOjt+BXQJUHjFPCObEm3Z5Lgb5U/tc5SIvB
hgdgZigZ8pjYB5omgH8G/srvADTUkaOKXBoowBplvM/nFJuxX/nCAAjnuY1qwYFXkAeRYZg75FL+
X7/qDQf1LFC+H6JpeTYs65pG1d0r5QS0Fb/RUBSnfr6aMo75+jvVAcrlHyYs9pCsrNYN32ixo3Rh
1603k2ZgSa2cMTyhx7tNtpfFOp8vbliutZytQVuf5mttct6eYuDgy7MQBXz67EoOJ6/nhtNOtdd7
wi7lzw6oaL5gE6asgcQyX4uVh3/h+Ra2REhdLqak0IWeZcIjCshii+EQOkyiUlrQ6GDu54jiewZO
4F+oSb3ypTVFU7uKLav8oqWDs+tvQK5vP/3bvPfScut2arCAnnmTM3i8g9Ym+FMZlHch71Evcakp
gLR0MyM7Xp5BLdY/mYm7DHwCf8wt+YwFLx5AoLSGCiAqqWbN5pyLBHvGcdnq+7XQ4+bHaFkjOQkH
3ZPWjNly84mtO1C8BHiPuUJczOAs1Sw4xhxEZL8+YXL110iMsVp9dcMashWczXyaPxlZUtqHDo7E
EIrjz5nlLAIQSW3agTEHCS8YSloUpQDjDSNqceMQfwL5YRik9+OpxEMQM1O+6oIL5ef1RyyUDaEC
ehL1sU6YMgjlKegDFjinCcPk0GkoUILoF8P2yq/RRHcyIzbNZ30MMg4D7xNehDqmDugNfpBSP7+0
+j0erCljLW/EUGroHLmYuVAIrp7QtYMU6oPVvCYtDtE4w80cJr76LCFWg7/0Lzk2KG4HbuYI0jbp
0AvVmAUW01z/Roa4PCCGaijo4mcXqbVL/U15kEJjhiSj5xyouqcv7O01DtSaOi6yBL9QoPyaOW8l
UgSWUtQw5HTBmvPkWCjKLUww/dfDnrXGQmxhXzNHEemLFqx15IIw/QTk1ouLob9f792QY1IW1lq7
MNGJBjAtq3e2MIwRzZwO6oxY9jTq8E2ZbR12DuAnpqyuBrh9kQRtX0Te2kTPn6pXKgVSZIHSCvI8
e+zvBHqC9urs2idtDN33sSQZNwfyOu1XYi5SXn+A/WR+bdHUgnglEEl1AFWNZYw7SmxhO9+CsBhJ
ds8p/yoZlCKIChYxThuVWpTUOsJLj7+Wkn6hj/1xNTWFUcp38m8e6G7sVbAxqiG97svXYo93LeBX
hoRecIqEdmlUW9ZNbPkDcSX1k+UpNQqkOf1tIKZTCCY7Dc4G+mt2lOgsYKc4ud1g4RKmKbTeixQe
BROhzn7SsG6U6aayZ5Bd6UQGEdvRowQdULMQ9NQND9FcMf5HF/4uboNkky5lMZ/hnd/tEYtBLlw2
EDtbOEjKrsGysmRz3ag/rCxclHhzX9cqmw7M4koex118kR+A6GlkvwyMEKIr4eO4HIHOT92CJ6eT
NMBoGj/cgQTmWsl2z2A8AMH/s4qADoU51Ar63jELRcrWEWizl5l8+RnDkQpdoUb66DG+2zIFwqK9
S6dtAy887WYNjagvbn6WT8JN6z+wjmnOY0pCwqiZDqNHZpq5JmTPhJUlKwWCXW3cvlEF8sJsootR
JcwsFx6mlpaBAPgZXjcI2mBMcF+8KWB6jvfnpDSneUAtHsD3hebUt4+RhsqaYvuwugGYyLYthq8d
mLUFiUOAR4e10r3u/n4YhjvVGo3YCMTwJzZm5R+eJ9NbBPZyxhOdV5uXHRtz5xjCZ5NJy8lV3cNl
HQI8EWEs0yfkHRuv6nbSzgneCa6iJ6kG9JZOsljmJctCjSIA1h0j8/UoWS7w5G+2gkZOs8oIwro6
qBrTYiobOwViLxsO52haw0OezhqOt/+MQTC+U7VboXPoBAdeBz6LV9oXo8kxDLajvgNlIIx9tqp6
APKkA2YapqS82JhkdaOWZqkrCbruMHuqHKkC6WgvgSDP6QydqPAFGrGBb0YW0Q/o0FP1R1NdfeS4
tetyGAn/n2cbN7Pj/Yc5kSwZ6quAu2L93w3irCfMuwY5g0YjWwOwZTrLsA8ArGmiSGaJKaBfF0QJ
UhimxgiSd/JqNr5M5v3vjvMy0rXJtpsbF5XlH5F1bhTrWKfekeN3gGaPYd5ENvYsVkSoGLckC3S9
K6w+YsXFhb2JEdSnTj2XiYkQN0VX/MdB7XVT8ylEtPqn7KgyJfJA/49zayjywgT785rZJfvaKwVB
90AsDyaenqU7z3CbffQF9BfnPRV7tV/5kras1dNxe43dzXK6SzQjlGFJQ1gF1R9saCKOpimexKMj
N3PqZK5ngyHWGJ3MhhCLPucv18NvhRPRGrQdny3kLk6ILqkBiZJREzMUubXAf9VQ+Nuuo55LhMTf
1ULP3PRIgaK0iLktxc+WrM4LiEuCm/v7DQClLThYFES/58er4ZPqvW1xsn0G6gIm00dHAdzLMW49
yJ5JxMcXyAT82Ti3HTSLbOZpLftdGGmJaCEPLJXJ2IuOJRSKlAwlY4Au7v2mEYPka5VfBznCuTkB
mevDNY61CwjSaej4CJgkny7tTamc8zwvV1TvKDOFIcLb/wnKO7AeMH3CJNro9bsLwEgCmuFNbMob
ox4OoGz978u9BCDqXLEiynhBqw5vki5MnHJujm94wCSIE0KY1ordiwHw9Pyymt+PSPEPpTVcAoAH
itl9xHi/MtL2zcU0jXCTDC+a33U1wpI+i+5zk9PqygNzyxHmylx/5lVUYfEgpbQvB06LlDUgYxgI
ludu7l0prQjCoG3FJs+pjzr9FdBKWyBTCXSAB9NIAXPSjogKofrnjW76NsJX/arfYpi0citqQJy7
XqTt4vU4TZ72bl/GsQ1GZpIffiojGTkcfiOuKrAfwCOxgDJiaa84f80O6m60IMHldMCiPLQw0d5G
6WVtXj8hm3K6IXXl1ZTiNI3AAlCRZ5qXwcF600Q5xoniBpj62ILCIae0nsu6oDxLcyaD41dK0fp4
u/vtuo+sjAMfePuca2jVSENENLhPKs4XStCJvaTPVEyDa4OLswsHyGSyI9/9tfoeU0f/dLt+SEIC
9lsE0RE3w3Fk/27U0Km28LOHXDB2LVcTDg50DUcTMWCs381A7MvPoj6JI//pIW809QPclblmSSFK
ve8guCk3g5jLV0sTpa6GSb/O1QEwOL/qPh61yRdhwf7qb2H6INUxZGKyo3L4KDOBT2aWQCtMGsOM
FvnE/Li6iVJdejm5Wl3DyJVyTP1ByetfmDYfMnvMUUlSOhBgvTKnKbYTcH8GDlOa+OFSMSckr7dN
jan1NMg4V22HN2X87BdEhbgQ8K6UOTM1e1ygn4BBoCsSwOL68gehvh2+EYQxOd5bRIf5ABCblj+f
HHWDRIiy7UtWZd65nJ/uvkOzLszxNJzqNS0/BwOxSWPyfAF6UsCCIqXaiVT5Fba/iX0YvChFYPTm
GTv6eC4UGjVvN2Lu9GXvLAuQCwZNtySZ5g6oJd5bCKryaMy2X7XbpHq7eSKfmg1gCciKEbcL83Lm
nkWdF8OpfHaWdqnZwC22BgWqtXxM9Sygz79hrrtyJ6vMrbko8jtr9cMYtA83Fn+ARv7SXiPcvIbB
LV2poA7V5Bx75Afi4lVgYl2nNCMGeGQ8P24nymhicOghSOZQsWYZfXzhPPjddAExadcS1vSxKbYR
eUAzhcVxLOO5gLYxNWDyiXRY7joSmT32CsW6rivI0NFEzlO/U4icxN8MzTk+FPptl7nQXMtRqVbj
NDzf7FvkOlOJvqMCD0rTXOT9vnUXp6QXOY2Ma0br3xkXmHYzzILW8LQBzNz0MgtHbOgN/71UBwm1
NK3n6Ld+1U5q2S+oOBp1Ocvs4ZRchBwwc+LMJxI8s54CjTvNDVVG8YpnobtQCA4djxqFAQabFv+W
tUmaD7bSPpM2aDFNhN2mDprZJndk9HRpklqxOIZlOfnWKbW8aFJD/eLfQP2Swz6kxSD7nGLXwJ6e
bimlLpQ+FEw28i0HQOUd/0BON+z3vXD6Qu0t4V0UUgWkSYkawo4rCyFSgSOIjdGZa1vHuoUejnaW
BJFA4R7y9kb8aOfCgTiMN6cMiduUm6ZJO1oYurRM5ZulwwK6Nd4s764AHo7wGwYo3SHnsUjtQZ7x
DcJLDdI5aWxvqqs7cV+WSP93x8B8fUf/EQ+4FCmHoMKR63DEq7A58aSn29T6yczrtyXPEWIgnGgt
RLZXouGd2qNL/c/Q7ykMFPm6MlOeKKLUM55hyYZPA4gn7UoQRn1LeZpk0rVVyzcagmB9f6MtHjbX
S2oeNf5t858cqcIliI5buRlriauthDFYfPKhQyeQ4dLztl1bFynQQmfKctdPRgOIub6tMvLK5p9W
PVSnpwfsmiIqlw2Rb5mfEBeFb9cCmprqlRhEr0NHksD4X1c1aL1lxHftt2C1NfNrssEg7J34Wwtt
KVGciO84wEbU3n3lbWSXN2BHlWXoYnLUmyFX3p186ONu/kXoBC4xCtJn0xn0KEzK7L17y4oL5aHM
rkgeg1keyCff1rB5t6pdGHlRWFOOi8cw8fsGHR91LB1mJHl2m/JGhKMwrfBEMVMSpwRZ8KudSKsL
CV4uYj+PUL27NHgXWt53p4C2FleTxWOO1+4piW+Z5FrmDnMQ/Ob8evR3ldaaVOcgKL1miOmqfwyG
PeLrZPoMVriFq0Z4rMTlIzya1EsXpsQIfUJmtHyXNQRaxBDsrRafkkIo7NYGDOgQa2lrr035zVKz
e8s7PdgeJmSn8ucM2vf08K+x6RmEXFzXPet6i8KQa9gzvXOwiq3lOP6/DgDqimf3BvTlq2N5pM1h
GJaKpOUmasHCFo5gFrnhZDFLPRdqUI0sKUBg4qSv2kdY9jGwQtZBqcM63evh59u4bF2DTQGSxVh0
ZbW3Bc6qfc8xwaiGagPZ39jTZ4IzuDFLCTkCgPK9hDW0mc8u1BZCn5f4aqMBgvvCz4w/8jl7Egom
xhVSluTyA94mJt7cj6gLH649XQKzt1ZkA20ILuRfyqNeJw17QnhlFlKyytSLk4u6wG+vszUUsth1
xdLnsGG/9gDWaOLi19sNaVvxC/xu+iLXGwMDDkari4oXC202gp3mStO9alcMvKsRwoExvzMoKcPn
t0MltTQ7e3i/JufHpmxSNYOV03JnHYW1c39rm+XYDfUF7JbN/zobKE0+XpAcDMclxJGSrSM7vYAO
jFwOo1yBwdsa+R9WNh/7nJKvKHA8K63Dyltxpacd0V+1nm+QNOUA3fV4AEyejioavZ9wzzJja4BI
aDhNU0WCi4g5QfwXPYaTQZs8Uzzuhi2WZ2WCmOg9RMnh01r2kQrsCxNVt8Vb/d0iscuyEtx8WBO/
zUoc507rXj693Tl2wSUP8W7tjYxW2WszZJoV5AqflVyfLRhWHQPgusHVZWONWBXhikP99Xn7knXN
LBqPG4XGg/tnyRmgEHWidmdJ+pIBK6yPrilTcWk/APTdBVoSJ6i6t8xjWKmzwbh3u0KIvN5ITATl
lqlNzPwQzOE3mMABgaV8v0fP1UN8mfiyBfqPuEDXvzIVVVc+jvHfEiqo6FvFwvOp4xiJFz2M6UL4
FPnSK7FdxIAQdcR7ID7jNNQla0I+AySLUeqe20CnKf4cFTyMhPUDuFFe7KU1XVlLR3aYRpMMRprY
836VzFgk52pCaC7Q7+i91dNP1mvHKTqmpVyXVStM6eBrA5qzcVYB+/m5b/xa1b4GsxvCk31Y/Jee
LCjTJXyQE8n5izsfMUMifzcPUTF06giX89GeHSx+TReX65KvnvpIMAcGk2lMHhiRDq2498YacssF
RyJM5hnUN8mlE/xcjp8fpww3QLhlF4RIBd0BlNj2zmxhhL+XN6DdaLlhWdZNqKuZ3tiGV9n11oBd
PGzSi5yo59LiMm0OraIudbRNq5XKNNda4PI2Rpmmy+pIgTjjzJwYLchy78OvWpHrIZ6Cvhpg0tBR
c4uNcFG2yaHqHzWWLCwKdv4be729klv2GCOXhjzwwhtR2etHWv5goKEmrwQ5Ul0Hp8+FgM9OaBvQ
oGkjA9Fx7fEddJcMep6MoYNLvv6JBaf1sF+cfJEa+ChAGxMdrPkYR1ASr5d9dK/zy9ERzgBufoCa
FIN7iXJR1o4e2/Ye0m7DnhVJjjGO7wTTEb6Yg5uduffPwLj77nE/Yk4s21NTpr7Fw10dQX+itFME
TNiYbJyP5KvKcWahevBcNDo5QBjHCnjGagWdT8vdRW8p2oK5qQhBmCuZwIve/iPiYH1RByHHggjp
oTEdWl8sj225YaqfAnzXqXBp5gR/S6f/JmHlGliODNlASe4jGKi6BzCbDMB09/Q0wax/KC4exYbx
5AQTXSQ1nfSlhPfIVrNOJgm9nzctbtf9saPA2vC9adMWL7HzBuuv/d0zZ+PHNFFiovTM4zQM6goq
RdFy+PXFVYYk8HzPJBuMY4NLUYiv4INzxENtdxFar37i0iuE8rY4ZIbljrtCb8a15JawTSTDVuQt
efjEH7mWGlqUPuD5dMWDwuk9i6vDKN5VuRKXR0sZXw6Hex8kME+GaP1tLfAI6pLpc33fg1cVIVon
0DoA4mFj91w2Ty7FbSog1xjSKvjXC0qsP+jgqPDr3kgyiKdAWRn+8YZ0Aro+DmWi0WjOV1dEM+s6
Q+V/9ww0IzoQk5EAPlSLCsdh8Ip0iXIItB47jwXe6Fhd5plIY93MAQqsgYVe7fTCBB8mmfh8Gswr
9L3KYao80SIaZNh7JvWidN+m4pDqOLpkRVJQ4m6zSKKzOWcJri7Sn44hcupqjsj4FNiZTMnUV8ES
5rh/SgC/gpxEvIVLI5xapquumpMfIM6ogKhURswH46McKVc2XzROfAUJq5onyBtr+WLT+GK7E5/L
cKNoPEe1yd8cq034MExXQem1fSIYr005j6qz6rkQvXcpQ45AFG0qWkGGnkSiOr+ZZFwdc7FDB5L2
bcHhNBHMhh5rbH4GJKQ4Wmb1afTrVaQ64O5Mw+66s3STIrLZFmSTQ2wIEwKik/gon73LzNGEQlQP
UPBYiqLNufaToqcLW7RuQ5tzbZVSCjrPLHEc6fD5iziDOf9jasY155zJk4DaeWqvhYXC7fDCxhiG
F/qTKn6PkX0OSOOedO4ffUnqTTucmGF4hlKXC7APdEx5NZLxQChexrG71+bGEhmZZKABAvicBKC+
jCYjfdoCxsN0F9Anhmt9O1KURuR4IGMAIoENX0XnIZsRUEFp1xqQioAuy1l/GViY6PdIYExk35t9
14shKz4Kmh0zU0VwgXOZIHrQvN4TXbdQpy0r58P+FppItJ9QN9/BS82hoXKLg7o/tM6DtZCFlQSX
PPOl7X9T2xm/syppGLVM0D5vL5BlIdGsfeGTB1iEMuU90bb0PRkUovgJuaoHMRQB/M2vjopfWcQJ
CMNFXqfuvJePix9xyQHFqJeEyOz1MzYI+oCf6kSG1ImMSDYs1VSmQIoibXDcAGfWJjWYQeOiKQPp
p8faFK6z7GFLPh6GdxV5jmmNhJUMD5E4PCXdUd4RbGIh6I3nhK2Bi/CPoV1X9938O3rtcaWiS2e9
eSsgai5nCD/XGrcqEvUuDE0T0+ZSPHFqB6f3t3EOpz90Qb2eHkJ3/BUfL/FVgaSyYpttuA0dtgcq
7umnaxy7e1VDSDM2ty2RwX4246aZhLYdMaqrMAkArWUQ9Dm4kSjSacH6OVK1jXtk5eF2cIAFbfGB
KS+WG1iAZZWd42m6w9PHmE37ha/jh9RQdrIVfSvXuqPgR/8GVtlEd+GA/YY5mnRB5DOWXriitMna
+9/lutMfWyW6MzDsplM7/la3ArWlslZrE8yWiMXWm2X116OtlNbld6y0O+2GFkJq3B5Dyf1qWLyf
h+rvo1UkxcjyZvR1gwcIH82fh97B/Q9iT4AAWZf7ZQb/SYNncHGrX9lRUoHo4Miy200nvJxfw+Un
lsP4pM0Ln2FiFW7/wLxxeMHJKR1DL+op2Fyoe1JKymtLBy42R9VarP5refNEAO3ChpZThL3enMFW
exlUKhgSI1iEzKOLgyGviIIry+MQIPj3xQWm7+9cwxCgw3q+4t+OnY1dhfayECHUjWmSeHChMVAj
6svKe2uGe6aL/H146YC2kE9KOeX52Uw3ni4EkYzsPnUAv7Ltz0H7uBBkHoT/Xwuy6nstyVqYQYxS
9EXqGCs1ge1k9GDr8GeBWFwhZpOvbZBEgVzHd95x5Z3zy2mcTsAtj/UF1fd705JX+3vT8HQ7f3eh
56f6Sn0v9eniEGoM0tH9JDYpNUK5gxdQWXX9APe8ACBXWzTCUdEWF+f/t8vHit+w5U3yS7WSALdp
o5JJ7MAtjSWj82aetX4ffcal1oSEfnEJdXYwnAdlFJh/K8qtBlMLFgMCVb/g58Z5UVcR3RSg+tK2
Y6g1bgnEwz9RI8zz6vmb9K9AH91oH8UHnR8R2C0BB0pCxMnTDuOPWpoBnm/OdHaq9TWgsUkP/UXH
BpACC0XKclhpZ2OGgxuXBi4uwLaaj+8FAVqTR8uf2+Gbbhxngy8DK/NfXzRTqZD4pC1+GpDyNmkZ
FeVEMc1JZC0oc9p7XME0as0aTJjcnlkpFRUVijhiQJXfp18JX1ckH3Y3Fqq4VjAsYaPMS52qMSiH
nT/hOiKS9h5D03MtLHqANX0zrqfUGKc6mwm8gvPoUfVPqLejvlc1wNSVlamxAhDwP1Fz8bMm34FW
U0oK9dtaMFLR6MPSMu9UhrrW9fq9eBoTsQHE0FsoZEed/IBg6qSDHs3J6zrHGJRv3PghINRp2y6q
lGhkxEVEjBMgDldT+sTRpSNzA/x/fQuIqfkYxMZ1BFA3oQqaNTYsOptdzLTZJErevZHpXq9cC3eF
HqjA7vlY/BDQ5V6xc7vRUD6Rl+HbH04qqpQ1aDzmxfv7McD1LWgTE1M/ZIAqIysDr+RE2uQn/Ceo
7w0ztgZMq2H6ex/3Ch68SISyOU0pd+06l1DPmWZfTIRfB2LVQD39xOdkGXW8M+uB46m98WYAskh1
McKUea+kqq6yVQ2TpBJw/9v2LRDUrQgSBidrjWI367CFJFca9iaY0UEkkEn3MmTLnubpsvmtzfbc
90aULY7Lcx8nSor/5vZUx48/r/Sv9O5FKGK9k1TqK1YeO0zNNAzeHsG/DMcYgIQXR1tR7qHxso9k
tR6uPtBlnZGElxVHa74Ef/QWle+rFk9ef3ANJ/1KDjAsdK0qRk62bxXikEWiIsX+7FnACjOTm6W0
pAYKe2cybLlLbucuil7+P0iPeTH+Gmwh6sANMC8j0s0nyCEWpOQdCsxl06h5/1nHIu+AllSVP6bt
XjWXr5WvQa3jc+NhzcS+SOrIQWHEHh+NElahVih8w+yA632M6hMkaOAF0Ewi4U0FZWm7qP1rc1ss
A/6Eq2nCG9ZuLLaPEYXM8XnHj35S27LRAIRAGL0nlJXv5iLaFaZkPBPLfFHTxduygqngM2Yy/LHM
3BQ9tS77nUyfLnTKN3MEaY6gmCDvN9NYNy7yDlLvL5xypIIOdPAqP8dsQL1rgT5dCjNwAURDSOQk
jgY2SyQ2mQQvLJmVPQ4k8mck70/DmT7aXD7HpbH76zzwjlw84Ug7C3cZ+iJRj4+ggxLsNljRdjl/
u4WSXqBoeefrxAhu+6oY5AWXN1XSgFKTcRWjqndwViQoR2L5aKqy8sYuhW7T3LuTOIvxAOZl4mJK
aeZlZ9Phnapk5wx1lJK1I94ow84PPaIZ7HRmPOS8UjXN/+EDHrSHFn5eX1KJyNiSq4ihG7NI7IGL
+FJSU5ckFGWp1+LpgcMgg8XDQuEW7gajIHRTPQgjjfhwyBQrVyH7MWuIZz9+SR4+DK2DhIO0vTUG
hW8tnwr4FseQAR8YsYofMuasVBDsN/B0Xa2uEZ1w3VdusxYz67+szLxSXdgu7+wINr17D7vqJ3z1
HoW2jJxDmM8MB3beMDJCl6XILqat2Q1FlLjA+eB0BeZMNxlpWEpFnZWliu4ul81LhMfhS8iz1176
CBmZmDPlz8Nekxt1cF7zam51OU0x60BTq1Ifvsks06KT1LbGA/tgJyGWGi4OqVG+KyRMrtDPH1ym
X4VLz0n8SnQ9xqcUcVUjASjjHkcFuKRzB0/4CbwNQ/rfOFFgWbMNqUZK1Ag5dBIrl2GrDOoJAHgS
H1c6C6Z6qzFR6Cn2aHNrv9V/kmGaEwwMdvdpstQrOmsyGY/rfXOybMxILluF94Fw5sqHJoHi1gg+
2i0yFjj4IBwSMjfzLTMaMs4Rw+ZQDKLkODilXw68bpLekHWpAAFIUwkdEFSf3A9rSiPGWo5xPmPe
5YdG+iH4q9DP9fxX8+W/mgwvwvOJvED1aIoBC5yTF3F9tV/hL04KFYhQA3eEC0erZLapmWrw7AVA
wubD3wRoiED2PFfI2o9C1oofI/8bzdbZEuKwI2RI4bR/0SJhewx6GYYCiFMmUJ23of0dQiY+T6ZW
zauPaFrLpM3pqAQsDLdgKila4V02gatOnizN8lp00fgv8HDi8uaif0+GiRFPQAgXWO31NcKYz7PA
W/Pa0ygKKNRz/3mKnEqxCSRk6kBoXypBs31QSlQobMwPt52rSOe0hpsLrX0t1k092eM/rHiL6rIU
dSIRBts9qUdS/en+AHP3aMqVwd9/VOuiSGkoodcxMZi4ZVibfB3NrX3POIkmD8QxyI1+jrnO4slQ
KX4BE+q4ZM6NPHZjH1y0k1rsgTxXAMjhrpcPRX8/uP2JNMxIKIu2p4vRdo55iCk/kmeeDKxET8SF
mzEd7yYxnXRjYYyRyh210/LHgPxtZAQ4tYqhIxxli6R0/su+Fms0W5sZ6Qn1iQBghsVB3CaYFkPY
n1zx3SwoT+I1ZQ01Asey3gjQlbsna64IqU62u4O2nXEwjyny3dbjfadeU5CnHRxiTUURd+YAjDze
2s/qgI2RDGa0xwWWhKIUcUeOMU8v6zPbOieI5KSNBWX+z9eQPL9iXBsvLYdbnoXTzzgU7bW27AGq
Yvf7GvevcxRB74V5zaRTMyn2v7Oim6cvCzIf2Hua8z4CgIxX/Yxz2MwJZFuAJXtYCVXgBos9q6kg
lSbUKN+YYB9Osi2ifkubu7Aoljso8/2GsdVfI2agjxFsP+ubjhIvTvG4tbYO3RsErB9BB/27E7Hn
KAKWCBUiOb09HlXxEQkEe03V5feyBoLYO063JG0dt48nhIhCrXHO874fzTsaJO3t1dwy8WoKqYYw
26fC/6lZzjhkggNyCjDEH2Z3VHV1NYFzS34uX+gYUue9sEOOJy89X8tra/BQcJ0a0wei6oOEeN4t
9AiOJgzRdkUmgWk2CgbPgV4v0XmtphHsANhfaFzXOGfUgIryrClb6kmyEGZzr5cbPtEip/mL1WMa
R2K5ymqUadeZuHgc2eVNy2inzn4/7oyOSD7nfFSEDsHVpSXukx5K06uZi1sA//caSeyEj9z2O2Zr
O3qF+W3y5F3GnGD7UGWZuuPZCj0U4TzaaWfdHN18FBQX4iiomvb+/ybEWZdLvtFYDblz/GKRWzAE
xX4uXXaIZq2bpdN2dBxBNrjqx+tWT0kOx1tUtozEwtiU8Byvjr0xlWuskJdvtveEsUmuIRdnFRKb
L4CQHQZ+e4obNlrpLO7dj/7MWhYjcWR/L5nMAUc1iz+DP+hn9RELHvZ58GgCIdlBoBBQHMPef+QY
Nl3yDnsjZdOklyUmkmCHOgXM8/sSALSqPMHS7Hln887bQuuC7WtqbOWq2XEHKkrl2Z2UgZsESdMY
HvUVcu15jq6JeqB8X81SgewXQEV9tThU3nIxG1Uy3MqlxhLF1SmwjzMzuSDCbKoDNBFqsggvzNom
tliXDkzdEoSIRAzajQG0W0VruIFBNbhbVslscSeUCfEZT4374RTuCW7gJrkkK8z18LrpL7KopGuT
kR0LtSot4diSFlAHbSCpxPW+wGBMdosgDrsTa7Dtww9roOvfFYW9VPuMe5hYdSpi1mnt3UIh42Y+
BvVAkfV+2xeTSzu28fLA6qLiGJFmuWLBD6p8f47cQnp0PU8EJeL7UhKlivAHgCQLv/lzawp/G7C8
HbrNKPZIR1Wou/7BotKpzKpN7+u+D6Zu4B1ji8esXMk6yDZKBZ8AooKwGaytoV/ate7T1VsB1lq+
qiOpwkzSB5LtAUzhFkziM6Dv3uh3DUnmdmXPI2A35R4nXEVsDimjhiJF6PISV5CdK3sS14/+RnXU
ECucttO1SMPhUe+j8bwBYNCTOaLbj8QUmMnhfw3LJuVO7NUxJ54ItlO44g8N6zuL88951kuvJsRM
VBfOKpWjbDiTDgL+AVXlHqxWlXDv+/WmEkx466xLzY6GX356F6o6IXY17+dGzr7B+e+INXQHaS7d
UEzeHg9uI1YSW2liKclvEBA6PAehEs7zP4nF8fT7ZcYBlpp97kf0OXRDPePqJ06N+DSxyBk3Yygm
AuWw/cHTq4YtPexScboTQWDtpWsa1dSaB5hM3SZMA4HDVaS2XI5eydM+PxZ9VJ1DCF53r32DMi61
P8FOApOmgLrd6KBntqxIAz/AezYHPezImNwxb2YtbOGWkrCmrleSUDWhrLpWnAoSWXz1m0CicB1T
6H8V6AKUlBM+vGwx7EfDziz+3QWmNwi2MG5z1HeOnNiuCORJm4D0b5ZcMbbouiiX4T2eBIVtMC/q
uMHyWpsFWa61OdADTnlTwcmG5+rRzsx7VajgCBQX8HbbKqkcf23PsekfhE4iI+r30wo3NhcwK1Rj
2J80QBPArAbg8bvM5SvLUmojmy6DKh0CQO2qlGP2JG3n7RxRRtKT1hvPYoBItpZrQASmP3UY0zJv
9d5cBVOf0DRQP27sUqv9WsnLZcXjzJ5v/Oz5aQPLNilyQVXFYHctAvSjUEB1Qq//R6eqwR2sYfbF
aIczLgfcr3ZnHF3OJd2M/cNdWFdpbCmXPvJ0666IIhOTMORGzf/0MKn9kaSGl3myJxsFWl13vCTC
HSKXHNZ/F2uHRhCOIyZKxJu8eah2bCYcnGVbejUYrpIeT65q63OLxIRGqUbTWPqfZmMPrIuqE0u0
a6oaQ+irMdiyl56fTs1+kc5k8h/rD4r/q6xcNFV1MPQ052w2DulJVSlL72BGU5xRbtCB4Mox+Gjw
yvlOgOekQ8e44Ak5f5Ef2oqnf1Dm63SCgUce1+LVP0QmBIoECP8nhg9qjxcUgb0BHpBy+uLHa0eS
Eatd1JLXS6EqKcZq7kkzc9toDVzJ6AI6wZhzc5qePy0tvRjTsBPMsjQa0+CdITx6jF2SQytOYIC+
LeX16w2IT1Oiakmv1aBSpWzvzvSSQ2uMupsqvUiKvqkAItABmXlXztre6mObKZBKKPgZ8w11T4g0
TNktTFZRkQSKtN2pmv7KtCnRYyfDsiYalyGz2Vpn+xe+XE3x9ilQTXyzcFlQ2MuEw1VKSUG3Tamp
V+7TgtkKMiGIBVEKBfvQRz1mcByAl7kJzCnHeq+VEzzjSb9hh3HHzVRE+qc/8b76O0tcelRs3aSY
BN8XThYP3FenN0bsnZ7RM5Mn9S93diDYeEZidpJ7xgIhXXzKyzcf/wvC0xEyw4cTsXNJ4BUhkkdy
WrSmy8/w8T3oE/i9RgFx2yiCebhlYqQQwivTiwYgFR5V7IIjWqaFgZQwvz9lFk+8dpOtdpwvF0oK
VYPDq58EV0mbseAH3VDfuJA8W4ZhrGmVCF8yHHuNNvyyfQb2mUyOKbEiTgdMQjhbuGriChWtojdo
rLcUEjx1GkjpoEJC7mEqUu5o1QU/PpaXsOY+p95i0smpoxaNtiioC/piKtq3/YUXuXJ1DhmN7HZj
8vcpVOGfHriWJL9ft7yeotLShcQsBpTAFwvN6nWGnyAdkOB9uqMOoNgfRqUJacwMFDTsL8XpE8/E
d9Lbqj2rRzpYyLOR6xH0kfjXaqJEecJdemScPOlAN6AQKuO4IL5mvAJcDfn5CTdp/lf7zBfsklHd
J7wXYFBwRrGBftTmotGqzEaetpQl+loyMF88PuC469STDzF9opvDi5DJ24a6ZtCiJaAL8BIDscM0
Z8DpsXqiuvqUzj5qrJriwixXhWaxqVRBuxVvimy0ZheSmjPuDvwm62EETdvOPgC31EmPQrculokJ
ewX/XzskXAPAmADLoG9v2Pdc/9FM5PmeAyBwURB4wWsaaO6Kj3p7LEKuDkwewjkaS9r+IYHesiOD
rPo6oMB/1fzbSw4Xm4IWWlOayE4OlmOa9stt6I/8yCLomfas3XZsK49cxQ4Lv/uecplRcIJC8axl
rvMc+s8O73BZOl80bAXsjmQxzIENRD8GkDbjRf6v6Wx7R9glSB9HumqlbFfBmuSmOZr37Ro7whTt
sgob/sEZskZQAE3cFCvRNf9PWSGUPihHmecvqVmaGufhZxYUdBlqYn89HtW78Jx71InPy95exeV2
Ni65xJfLnWLLiSBw6qG1meXkJsBdbTdpIZI6nNvfg6vtBUjQTPdt1DptvcFJA8JMUswq/q81zFoV
3A6iGTlFy6DUcg0JOL1SONGoklBgN4OCku5dkQHdlqMBz2Ud10y2th0C0gKkNETVLpfscFsLDEoU
6ziPymhU/8iYO6KGwx24Ena7grYPVTWI6HgkopwB2jg6NSGnB1tFcZLnqv37p/mehcrmL9BAjsv0
RQTlrxuZ6s2kwcJX//6KJ2OOafW01S+PwkjVCgi0HzF7XFCqnpDwmpNuknY2UJhVisKQUbUyHy7C
WimzowsvcmcHarLMdGBJa8hfGa8bruuM7gYpy4VoBfUGJoBgdMUIsJ+UKBOtaJM28o4YndOgEv0j
z5RmtTSskYuYmOd75UdPdoNTdpGy9Nq08sRBFnQ3vN1Q03bLleTx463C2g6fbLAvW3DTfAd/GpqK
jo1CrClzBaWYY8aB+Gh9Qp9/v9/e035eFA5/XBt+ciB7T7vX70bSrNHmlCREs3MpHXqzFiX5/2pr
LeboNF3iOdvb+bq65qyco4TzeK0dD4br7h/OQZIiHs777Fve+Op0leWwet2NNzWSHWNsQLJQZbjx
wC25VX8OjBL92XCExf2Yul9uG5QKtEKEFlAgeI685OtFp3OirCrmPI66152ArxCNlWAAPcJnp3hm
BPzj/rDERku5Rxv1YXe8nqDvKE4ZDVEgm0GUh4xIg8QWntWA+Ot/TfAFjeAzrGrKlT/CItkg3mRi
UKmHPQzUoQzONnArilCQXT64wiyDxJHKn6s7+X5uMmYLKIlBXPyH+F3zR7swGYsQhgz6Do4SivIS
PhpckFdnrr0hOB1j92tVEVSmsYy2SbKpDXz8GDsHsSvJtOM3FSTYormiSCOirz+cyiQbD8oGdfZo
v2vXcFhYz7NKVJUHAzCXhX+KEDg1IBcUWTwJYNn44A4Pgfq0awUUpqjL1LfNkp4YCjmQIVcItVX/
iZPduTojxk6bkFjm3gMYRPXcMAmmeBokhvrBIuzUc6/1PMDAPtRkp93T9GC5YfpTmYXbSwYgnx6m
h5iStu0OA6cHqkWSiJNcN/kpYMNYuBojljEPipdqL5YtSoLoS/62QJBU7ozSgpBTmRg4jjPqHn/I
hpdiva4H9Q9eepFkyqEbwYOHccy0D4w1xPTuBlhi0hEOPoPaatMXzjPqZXIvahSdU6zRaKai6RYX
1/azm5+eWGRKX6cn04wzDG/6W4IQpjBUxf2Kbw+iEyhbaMVxZKjyEMXzbjm4laa5hgdmL0k5gemT
1Ez7DCVLQElfnNW6wYRjYSt+Ztkvd0PcUYaVLUuH56leeFw6X77qoTc+Z4DvEeRTq7j23MHCSyHm
X+iKD1vAhuiPxA62kO92k79nUz277zIJ6eOcJRg/k852UF69bGYXoatVDLCi0ecz5hV2F8JybLNd
RgKtDmbuj/IehZYcF2SfgW231Bprno70wib78uPXtgpu7/mvJzK3JgbJCw9A3eLFQXLMrAMkM6Tv
wHWKzeELK7xn4W4DIdCtrpRONHZ1Oe7vJ3mBiJni9BvSNB6FsRwIq/TA2ylaTEVqEKRsB2bom2e9
x0EU5tkCXfV5S43etfBaUQHv0qX+f10hv+MzwtoN15pF/KxnhZBw0Sowhufxr1hin9LGXXQxQIdq
fnBc5sIpzA5Sy59lApY4bO2YcZsYk8X3hZYo/ZTOZp15AO2FqtY6tcFvNp4uh1tjLDPK+EBQFqaF
7oYse0vU3I5xdRmZ6+F3SXfK6qP8dpP3s9G0Tv8ktA4f0oEDmvpc1pA4PWfIOdjklsjqQIy6PZCx
El2giaLanhfY1jDAW1IeyVyk98v3df5+M9RY+L1s9jDL0yzwaSNBjArxfHHKGzzAkpDcaXR2+pdj
ZlnCmFNcFxZZmygWeKpWdW4/21S5xMOz5zbJ5nr3kdAaGHNtNNgUzjXmK5QqwcDX3/AEDzWVL0Kw
pYcGmJPP4cjP5wH2EzM1ZPIW1rWqyOAcAwtQJEoc5D7wgtvTZZFKiQXYYGdlZrAhLiW+ahtYMhSP
X1dL+trUlFUO9Au10LPTbc48Qgh4kHdalprJdsj4aeWuS1mBoOBYdsEAE7bzfT0GdoB4qdpob9Rx
zLEN9JFNkbGhijvVNTXcYA+H+1CoILlt/BWVTewQ+QsZuBHGbqtxmNPWJeIevpfr4Y936MSlS5EE
rzNnqcTF+rXJI9f9wv6DxfU3Ys4bpdGnIow9VYoQ25e7TIcG03ff+r4zrXwsUm0fmABcUX2pw5ni
S80Fh3zlROvYOl5PTnUokYtgb34i5luFdBmqAFybZHZdl8sGktcBECZxRNe4kQTtb8aYTcPfRoqi
tm23VpDyoMfDLlHGozMFVAs5cJRE5UQeAqe0FM8xevktQWyysSBJHR2McBwhSgPlQ631o4KH8asB
CF/sA4oHaubkVzRET4eo7QW3QB8siTLiLjF87qLSTH9Gz3lzy8+lkkQ/WfmlaZbdzIvGIQm4kVAg
m18+jjOI+gglmdO9Mi7Iqt69FyndrlWRCon95u36eaNR0vihoF/h5+2cuaXMdkhvqw/PPKvNOl4p
h5gtYXdOO7Omm1oxq/2aw1LNNFlX2TvjIuVLn38cQmHTYZMsoFFtQbO2FBADekZ+KpzmMOwil1b4
fZVdD7eVKHTbc+LHOK6y7RcZw5LTufe9oUdpSpTIjoMkO3Hyv3jk8eBwZGgta2fmXqOUBknvkcwL
keem0x2WBY89mRqS3TdRmsDMdnhXjn+86CcDe6QvablfPfxrQZuKOLRFH61umhfgQYHChETWO07+
odB6GDVq/A5RJFG7iuu6rDruLsc8/RvkecdlN6ZcS4z0eXwxmSC/4zbs78YYuW5uPT4mfnUPY0yM
U+bBotRQCTdN7m91cSM+njsg0AId6TFwTOLDZRabb2Oemt9VbQwpL38FwwADSlg03CnWmfCmzFpS
d05sLEQdVlp0gNA7cYQ0oPSubVWC9sq9PZktPD/AQp67qNcwbRpr+6mzJEweCphMbIYkYvyzwjbg
AzruB+25HcfXHbeFmCKfkO8GxMtKdswoELsCQLGYJUCEo6cIIzyGv4Bd1y1tQ3HRwK+ck7pImLJo
DR2WJs/8CWNTedzfbN3XocTD8lQ2/7NoITxQyJlIHDrxHdHCjbTIbrH9a+Y+aQcZkORNgQkfAvZV
CUvQiaUIjbp99bzANozg/OEpIdSwIE7om7AsffH01iNcePOZmHsRc70OQflbCx7Ys4bqAk4yH/KG
2CpwiFmxqbTM7f+aDtdfHD+7BbA0wVggyt+JXlnxIahHepnz0J6AjMHceva7X9/CG2q6hVYeE5XK
OWwrSMqN+C7QCLZz12yNelbAabaU3+OqJxNpI4lVk0jAWrYXqC85IfBnjq1iXZgU9WbKMGzVLd4Q
69WBIU1pAK5aiXXxtQscI0UZhcgvSGXmqryd86edFVHqnm0Zsxu21WelupmlKR6A53r3lS+SCsbn
42sRNDJ/G+3P/uAIWZoq9fxtjZ3jVARNM7uXGIICqRArFVBz/bBIUyF2rPZ9ga8ArYRGM8CKdv52
BB0VpVpVVMMpPRI5tRpMZVa1rx2KZAMS4cNOe9vw23uTc6Niv5HIO2pVCYReppkT8dAbW0pddXYL
KyqzdBSF0zcX9BE87X5BdoXMSoV8qfKGsxwxqmoSRl/Olmni83hlofQDj7Sh/zxuMzcEcV2kR+if
26fFRXHUQ1T/vbjcruzN8duc8tcbMzLV57hPoWrgB0zG3Sa5Cn7sk0VNFRmmAtzBCHXMsrCXe1Wr
2XeMoQNbx3VZxPUff+mmSJbm8lOKAwwKOpGq9JgkRwIjbD3AR4tsnWCg/qQC2N/Q1FNmjOdRCEFX
FptRROBR3rNJrMitxpKIIGhZ16AKM13FGnDVqhYyslhzTgAzQGMyOjuNJRN4Oq9uLr5B+/srE/I5
5Ny6kxd44MKesnTv3RTKSulq24lMYjaT5IdKgVnqNYUkVHl6mzEIl4sX02tFISOyOD7fZYi8bqMA
CFOoPcSQxMCRnSqauxi6rJ8sNQs/SbXBGCy0E+h82JXVOaPQnLa/mgsCtVT7/9Cn327JcOr/0C9t
BNZ+NvTEX8AjSO0KfyJV9GBOqICFXnDNl2LDv/GbP9lYRJOglD3NoockgzVAawx7P2fhDaVWAMZI
DAvJ9I+17ohhlroBMZabymegriCFxuUCgPJKXRLOIZNpgCjG2hPcd9HpA3rF/cW8NYy7Y6wk0I3N
tyThpu1KnvPs1gMVyXlwt2QrgzniqTCuSP7ANCMO3vnZgEKIL1WDQcvVhRPwYBAb9fTVN/U856Rd
b+MvRODe86kte9fMDetKcWBwSwGESZk22vUc0NIgQfMQLjaCZRkJYaxFBJx6GU8dOfSvxmxiHmGa
5Xx3Y+stCMTS3rhjfkh3OV6en3wOAmAavTYOnaccSq3iJ6IMoUKx11hLNFb4tfF9f3dZUXcb1cGO
WQ84gUwldhgWckwLclbW5SN8qz/pxZ0ZXVdbM/VrebJceiWuPKO+FxCyqWfLxIsR3MX+pwr1ZA7t
HeQjJLu9I6jjj2saPrGgaJ8JIIne31Qgc3U06MpLd6x5sIz77zY4Md+loJyUz5L1SqdSRJhXE3Cv
tYLMkwAVY3JhVIfazAxAqIpNlA7BCtKu6hHXlKLggqDzcL7baGvKuPR5KkpM0l3vTEPH+7fZoQqB
akd3kLplFUQ02zlLnNJUOXCVHV1g2U0qHc1V2MgeiZc5Qh7uFEMKtexcxGvfADiy/+cchUiurJnf
lfKW1TyQZEd+yOZLHFxtdIZyd+to7MXBYSC5bxjdMg782dnbQ30X+8LtLgQ9qoePn5tiWfef/wCU
c8Y0vuB7x8hd0kuv8qcOQM3R9XCRXCe2jDPJdwqO2XNOsHHqqUKxiYIxXSYnrNkqmYFr6c5IATBQ
LLzF+Y7zaL+FZEksakCr33UypuqST+NjRYlHrrkX8IOV57KMkWmkMlk7NIEza+D4nyRBiS+TxopG
xnbwqSOMJAPh6TFbjHqInKyTP21v+DwBMUAnCO1U72yrjCE+EI2HaGiKkdNd55+gUB7v6TZuhJ8s
CZcb9SvN0YOS7rTERD/Rxpcvr/SJJ2BYrOe/LqwsZzuQfLgYx27ZE39w5Kd/xouNIQSGcra90306
OOs9f9CaD25EW/+m7JvHw+cghdGM0PSAif9UqPMmm2mTDJ9o34dJGHC0DRPFOd3bUHvIcYdHsogI
mCIZCaCJIUPYeynzeFIZ18Kmm3O4NkPLdWNcYVZQupvrcIWvYUdwSl17gz+mnxG8Jf3FJYktNxdk
cswGTwhUGGAEloRyQ95IGJN7LX4AgYYtGMYuGxLEqi7UhHWCLkGfvZU/PQ/cHPVbaLDyQEi7v8ZS
/g4CXvxLdcLJKPu86ACmupBEPHBuQv4wPcNnZN2spMVKl4j9iCbvFt0swHQyyG+AvysT9nM7ykOn
5DLZTiqT/zo4bKYnOddHN416/ukKBNEEJtv3h5ZHb94e578GOizowtEw+3HvzUqRKTNqA5Ppiw6U
eQyHsYBxVdrMVQYp+If2Uwevr2wxcDxjDy2SrFa4D2HcZnfGzfl3P5xos+r/pRr1REjfIgmfkcKJ
732EhCedds9tdx9cQN/XyGczAMsgFboEICLRGIHTRXEnnoxiR+IjwOuZ7aP/2+1Wi885kjjbuaW3
BmGK7wew5pfEsQbCj1UKkAnLsz+ksLupGVBv0uiCZ8Zrs61mmGdkTCDtyJqyQByU/vb3gN/OLiNt
Y2dX9jDkxLX9moIzEBPw42lld6c03dHw5crc2IDoyzTU2bCcf9QWR3QzpaZoUSxRwgIxsN33LWJV
tRczpAUraeAjSZC8NG6MHlqEVHocKgFWDllcRxzPufYPe61QFYnBmaBqO/wO6qcSM+O7CmzSdYY7
d/73L2k/JXXezSkdLl7m5rJKL9i5kiMCgBCos3Bbw1AhvTvMiZhIq1Q4LfcyOka6COGm7tiOH5sy
FDdahFY5wSEOdBpL3Q8OVYny8MX0tqtvHMTsy9yb26nrg4CB1yWfPrq12vtE3lXvMv3luZx2aaj8
StCG62rT1PjnDllrNLzPTQAYpwQLq4Nsc85A7A4HkqlFO32NeEJlBuIcNt3H2dJVnn7Ba8aKWxmn
PEm+tIXUyWzr6BvWEmVOzKqgFiL5h509DA2911xZrj6sMHId4U03mubBejs3itJkacblT5qqReOU
gK6VQlTf44CvBIm7o4iMyg7L4HlSeTvXsWaVBVkRPHHDuWW74oh+X3jrNNKaw5U1Sn6tkKIgkD+w
SZHJTUp5sLqe2BWyVNV4o3eUUBn4dlv60inmHpdbCtabRdYs7mMn7f3hC1h/brkXLvk2980Hjbsa
AKgGAf/JrQ+AsphsNYpMnBGHAel8iVpP2Zj0LO3lgRZphYiZaLU/FLBJ4JpSxX2cXscoDRUwp6QB
YUgcsRMCJtKzveyXQBISh1Kr5fj2ve19x4vwfsi5JAkNLIHq5zwJsy/MpwjmFiWdfsPwWMCtujK5
KiUMWIuFL0F6wr2I3I+wAdFvKkWQiQRu9YgcIOOwpRzddIS7l7omjvWGE6czx+4uXpemep7WtJt5
HJiarykyvOceGhnA11H4S9Us1a1XQsx9AUnRb3gN6NPV3OLs87OpuVIG1pcJhcgRBBw7jvbbn8pd
A/PSz6RTphsoeCHYQRhKjyALmG/F1uhqxhdhaS0vdOeZAl7YLdcPSihjPZAD+7bbM1pySdP8GdfZ
YMQqO16TwrIOfsNTI4zJEWv1bIEI85J7YeeNJVF/mNLfcV9p934aWcNG6GYqZuWs/KpgRAukbuez
m/DZQkCrK0iEn4lgKv4rd/LSNEwJIylKtx9y5hK1Oi3SNbpzxCjMy+hJMIvGVEtGqI3wS6C3HbxP
uZToe3APzp9VbndwTO/ELoQ9BUKylYukODiDcmiBXlGqAOdAm0C3a06ef1xBAlQR0T2cPfUvprsw
qB7T6A3bzpJi+y/I4FXP/Vn1157uKIOFgD/ISPW58hHCUYwsGVo8tTedVN/rF5DiWIN3IRzPkEci
ZeVvgIeGnbs+KaB7joNMchFfnh7kY/xnYQp7fzwL/rmU1IDWZocQLipFW1hCkxwS1pnSBuKhQqSN
3qeeg+3/PgVrvhj2IasuDYy/J+sr3lBy6JNugN8OMAPn2f02yGcq9rZnhWJ6lFhnXt5CyXzuU/ol
QEWs1LOqbhUHvyG/dhr9c4EyAbcPP54nMQPXxVxf7VtcpAOTuLFtwpVPw0NvKjuTF6h5nM5qXt+0
S0z/EU9ni2k0CAHd0AvUpp8BEuwU/vUzRRFVadpjaV1cFX7qaVUktM86HqZN7/GQ/u2AdwL5w1xf
u2BZkWrpaI3/ndvdzK+/z1OhQXdaRDmM52MHTony1qhrRubdAEC72YWVEUfwX6+fymspE5hgB2Vk
It9xqyNgG5u351HjLW9AFxhOFXxntUf5QM7wdgEWMdOdt6C3Ks7BO4WSsEDMgT04lSLJqVZfSd8z
hk7ZEIJr16v/1nU25F9ONtL3rwYeMSraEUl8Pxliszs/6XaQeRE7sSPYHdYlrozPbbezOeRqiMzR
AW7NDyYPycmM4FFHb/H5XdOL8pkaY05T8DZhBpcMUs4vVuwKF8+LElpKohgx1dJ0/O5sj8AvEOFA
AGImKyGQX1xK67qmxs0RGunLbHMYTBCzWSKogWTk1uCxu+xUbQJIIHquO1VaPQcKqhESzTDU+yyz
ZDX9WBSOSLtvV0vOfEu/xBkY5/0+g2al3MQkUueldgBjuFJeeror7SeRQobM/tCHIs2051KyrUYL
PHGVi3ULhXNEnp05oYCFzPoDOfQ/QS6SvDk5ZzmJlsczxSSnxiB/45HnwoqJhVhyCvCaf7swYdMb
/ciJMmQzbmZiOMKoGZGXBqj88QSu0gv9L8mZQCjLV8TTJcqZhWQHf0x6maC5VQr1iX5sTkylkzKQ
nNXJMvZVk3+nfcyAFZOJk2zR/y/+a0qDAZhRkZox/q2XhI81/nWXJSxMHdlJ1cJnx2w+fr3AYHFc
+TyhoksqRPyYF4beaZMD9QCqEpUnj4l8tXyebUdxbRe0Upw/YJgqk/HhdQ7fp3uOrCmbQmG8ite+
RYDELaOsbuDlsWpOZ7h3v0ZK+9NjMKj5RcWga7CodKxfCY9w5hGCX1wA3ea71w7yy0DRYe/InU2/
tyzdgdSuiuUojl9s975GTGqY149Qots0reJCpLzEgGudfYEBOKu0S5f12LjD6kPUkOJuEy8fZYVM
zsemDw6wS1C5L0pc5xHsEE2n2B1ihm/HavlL7hxWe6ldZEwuOHu2qZdihV5AnkL/6zlHtVCsZCF+
I8kMwy+AQPBgkEuZFKXi+cCzG4++YwJKV+YDML0lxvhw/oIZSc0SWG1vCmh91UeAwAinlC0lUUrf
eQN46Mifg2sHS6YAczGE9Gf0KFMTUyyUkNWtGxoo6yA9eajM1+BNAkO+MvUNg8O92eHDxBS3PSbC
ckvv87dIH6ddVmF7Ysbo6vy5dse58UFUtkXD2fdzlLo/G33ArhdU9LF8/HpvfofKXo/STV8oqS3X
famLLftD9ATIjbn6kawwn2LbTykEUyhDb8qJ5k2omM690ei3LkriQlqRkmcQ4HteWHGgEOiYbI3P
6CNIT7wCDOI/laVAenKYJUigP3dQt6aqqh88sn7suxmPrT4t5Efrcmo5mNX5+WYlcFmVVl1BZ8rV
GwUCHLdP5+6twGOTIkt9H9zyREzvdzTTz99ZiFYDPf/0vunCeyEL9NKiZpFK0SfIwElX2EhiY7kH
NHqx22i4ygdjvgM1q8cy0/15PcHAcTonYt9n4qtAgBbWAPm97YpYIlp90eQRm1IUrHhagZURB7y7
O+6i7YJ6ZbwEKWuPFbfoq2UvXEfpwaPbmWJGstOYuDbMoOdEGrUCnF6iNLCnx1nR0geMRT3bq7zA
5Aa9+bb6Be6N5jx6EYZMTvgGFX2l1+CmJGsmmBuOo4G3AVLFVaW7vT8yQdoXhyvzEh3hsVbOm9x/
Cppf3QXjGrevg6X5LG2n8Vjhph++QVGObCPO9dQO4PjXBcuIrFUhtGukwQn6DXyCe53nrlSBomwC
rlIXeBtGcq8whRkLWr5hHlQ/Q7FKoUq2gV1Iao3agRZSeh4JogGz6NYi6zO06yK7/v3E4inMXUM6
nNxUmyaIHahkvSD0mMFGO6wN4Stw96ZN9ivlZiMUwNUmkYECSxQwHYGkrLkjtZqpr4HwYYY/dc3l
Izx2CnD7Dvx63qfORxa2BhjRLN0ojVuGOKxoT1Y04iEKbD/h1OabxGUm3Kpd4wlIq/Ddj/goqM2u
QimfFoZ06OdpfW6lrL5Q0mzyMjGR+zUGXruN5g+DCMPjn9OzBdizT3DAJzHoTyB7OkJhWtL0BL7I
Dl3bNa/zUTyYEc9mvq5WgmiZ+Bpd0qq32lradrcQw/+jbR0atwQoy/pxZVSIXNTH9PoEnxSZgmJF
JmDzgigf58Jh70Pw2MUDyAjkJBukKIBuSmGoSx+ECgOdJgNYhyKFtlBS/pvuJPdzoHVskgHyOryO
nE5MyWwbTSF4YbgKoo0aI5oJfOTRA02Fh1ml6oPqtV6y2XTbkLinrnNnPFxeBDdgTpa4iAVvI0N7
6wtX34kCQ+lQVHA47HyOpM8EBnoEGHI7w1xv0TL8cjEC2vaDNuET8QUIqOub3klS1NATg3/EW7Pz
xquSleyFJcKMN8+NllMPZuMmkN+HhMvFLg2RUOmOw9KDMNLeVUJwp0uXFGCl2PCvrXJau1ycJgjm
Z+S+P/XrxXf5+TtI7ge5pyOlBf4YLcikkL1+D7Clc1xkXAs/2eCknh8re4s3ycEdU2tJef5IF/fa
GZ8pp1eWGbhaGQYHCNED1icgWMpwAagIi707Ew842x8fxL/WYtL74SFh7L6TyRL1WIOFY2bhiFk4
kdvcO7Gt867XmdZGOHptKjda8JmiPVYNxfqGeobMj+pz05Wtvs9LwGUnPZX2Ylss3FcBSSpfNmeP
9oBhZsoGb0XukLQH8UQgiVn2YcKfM86xg9KQWzu9w/sEnmfymwyy7pGd4JTUGF6y4u4pPe8b+Qg2
tW1EIcihcLfYkarKdfxYBgttPOobTiCPvM6z9B/tDnazBjVOK7wpC0SFVzG3xV3rX+iF2Lex6bvj
EUzbmkFe6fgOgVM7QUrRdzHnZQgH0O9a7zag51MVtjhd5dDi7xz3LbgWw2Zqwd43253ZO/+ezr6w
Spq382y0VDN0RS9k/Qyb+y1Bg4dtd4GDfPW1ICRlMDCGLGE9gI6vnTWCu+5tFCDoJfxWcMnPBUbw
uvHw7LNx9wjbPKcLZeS8VFJjD5Zo0BsyXPHCEHTJkVFZO+bcS5KRWp+mEMAYXWIqZl1rXIJm0wSH
wa3sktt0L4LFRAPJ0aV+LePfOwXAqGBbLOoIofqYLmUAWt0vu6LpHnVsqLwV1vvfs3ECa3x9CrqI
w9xvzce1+wDo4tOOFqcEB3wC/MeUV41mfAyiu0wtrAbt0ifYb3XDbvfLLBT8+C19IRgSOXidmSNx
Ks+1fgKPYvPi1pigDpOKvhlREkYqJ4jAtKA1albcduq1fWb+a8c9Y4x/TzoQyoICN8lTv9kPVXwl
3Vxlkzy6PT8mvsN8KOsX+Oeoh7oNfD/h5zQFiV3o/spgQ0amAlqac5ztmP7PLR6vENxVTq+zSV7+
Qys4sfIqc+pbdYth9y17XXwxLk+0n+uqEeQ5LeiOitrCDwWaaAOx+QVn0ujYXrsw59pcDbuVU2m0
oHp3a8C4MnqkH72YH+TblKq/ifR7VJNG0KQZCPVamMZx5GTQLbp7caAsYitIl4EG8+yinKDwoK/5
jEDpNx34kGzr8zvJcfkQ5WtZCpIpD4up5VyMQffAHz4aHdnjGT0MtHuX4J8HD9ihsYHYhMghKNk2
kkT60psZ/4FZV3VtxOn6GyeDbhUCpxLvanXdEW1x0rO4OmQVu+nqWo1ER8jK8udbTh7yv7e/jEq1
uemY7Trz6dHJ0ldGr2zLRHn68FHGdnauGk2XLV0G08abc/TF0NOr2CDcmGxL6EgmIQI1naFHZY4O
hiXpYVssI+Tdpe+ZpQ5tsHTJsPxai8nwHkdTaXHH/2oxqse6f6MWwZ+H3ue5vXFnu1MsgzIjUdIv
HEr3KYJYWV8eeeoCw2aPO+LKc9s4heWfd7MrfztAvbKhZvoJAdBGi36C0KRQmHYpH33PcY92JuJb
zSyd0Wv0fToQ8Lqz6CmsT7/CseUp42lCU+lEHgWO1+5P+ERfL8a7eWahml7CxZdHSNsZ9W7zaBev
JJ0K+kxsXbkyHqzjDlKrPkwwZLvOmZoRRl2Zi1RlUSqQrcuMgY7L3c+RVFBbwKmPore4G7tO4awi
76h5LXxzUVpfHkUkRWrMNkapZGM1opq9y1BqkDgO/f3k5YQULCd8CzR7T0Ql4bWhJa6zWtRUUzxE
lMezMerDYqH5k0x+BWSuIDzcM9PYBQsTX4R5+Cm8hHyFHXxcjPLJ62311ElWP4wycDTUy5K4S4Sy
dSyUuQGQj97COGuBuGSiIh5WAA1TOyaTbVjq8ctxRVn9Q+70Dt9h1ccMHwNEERXtf49KwI7p7NqX
9JeWGVaag8CQ9GersntgkPAew9tpLc1icI8TS2VUpLqm1n9ZYHqje9UXdkqlmjo26zZZwytCGKqp
BE/ZXEzxvFjCdIS59Z8ontXBo1pJxC5Ry3HWdcURyAfp+whMuX3dHfnXxUx+YcbJeOhYLWQgOyWT
oSF6y/AQJ12tSE92NbXmcUTLXe9P0YZmZknhvIQd1jnTDtywq9lbMl6SCU/ix/EEVgd8AB0pVpC/
PNRpL5UctfXL0+u9VsK0G+NsJnxuE+nBrHLpFdBqetSyhIIWcKxyzwvpgXSI34c4aO98gFx1J+rH
GQBf0v6+TBQtI5oKHRRiFQuS6+N7DOUv+c8X5NjSNhcDStAL6GMGdwDMCykLSrSWmyy8/IcWpaox
JJ+sZ5mQTZCadj6Ki1/Bwe4UTwxYE+EG7Y6kqhN1XTnzrXNn69PU/Ig0p02nuMRbuYJojDKFwo9A
kZnqP3wHcpJPz1WW0lmRgSzvQ1HwHkn/PTyPYH/IzP9xkqyVIIwsgEdScN9QuTptlU7APOLPrjRr
T1hTHi+IMMvJ1jrfNb9/OGqwagcy/Jc2bQnpFeUpom8e/2i00PD33FMsfDHyYzSqLGXQGG8mAuu3
VlqGm7SkqlD/KBFBFP3EeyCjIMBE19gdMKzHxB6WZI08aumU//PUyzTgApaoNR3XrPewJB4MOqml
KoX6KHHcUtqNueifaKRRDENZH/6Khh71dt+65HmEI3YkCbB1b0wpux5WhBvvuWd/5kOv3AeOVeaF
zW/WNwlLUMW4HoGnKZWfpGhjJbvRHfuONIfp6hkfo3UMpMj6v55mmIxdvb4eCCcPl9ZZ+FB8J2oa
v/O3znsARWBfv2hjIEVqDQ/qNuPFEXr2a2s0NR/ak3i0VvPPrtAe1IhwQOEf4oVHpjam71+hOlPS
1rl3cf2rllgDAZLoNkJJ5ww+XhVtmZPqXPfIgZTEUVUTy8yswdrqyxF29yVZz8R8+hz9/rH6juYH
e1sU/zihTObiN5TxLNVi5WHO73h3YHZicgLEz87+OBWGwgH7+phCANc5YRvHp409OmCGahrBDrEv
5aZLcsfKBSJyMCu6QUzJJBZdIHVfQW5Pa2Zyna758KOQj/zSg+fJvwO8yWpyu7xBWuZ5j6HiX/A9
FdbFVcO3qQykTA8aqLBkcxWn4iNvlmhy0H4inmtWvl79oap529s7h36lh9bYiXzQ8wOnxcZ+Rksf
Gmn/mqcwSQzsqrVUqh6HPsZMOfCWwa9fDZS5WJ5R4vFUsnmOE66Dwdj1l1+SJ0hZO4nD4bGilJ/J
vRGrOtXVdcoKbfCV9xCJuw8EBTNiuRGaseXOVJKGpx5lQHvcP3NNvSGiJ7XAaUU+DR7/eBrFaiEL
5MMaoQHMjKZFG66AcaeTysIIoH2o9Ab6QBvRa/PvFMMR2zKbkEtiJE0hAdRDzcSI7R1RXk9XmRRl
Ahtcd6uACqvKNetLYSCwD5TTIzHpkJcsmtMgRU49/5xyG3LyIjkK3hxeRJ6kU6ccOmCCkhFm+5sN
rBnS/IYTR4mK4bGVEbIIFUsga+1PtyyQS2D33EXAxrdZf5NOSAHy611gxGUZw0pgJ9SlRTtMaZFS
7jV/S+UJZ0/AnSXVD3KC7KuD+g5ZrPt72MIyVIhRydFpERVfnqgBN+Se+38hJN+PfwEwok/OrM+v
mZn/ON8XVX8+qMVywv4vMJvZRUJsZ/nf/+24OtiDQ+3AYTyOAxmJCFGH13PjNMQOBnBJ5zxIrn9C
nwUtZG03ifSOZtsWowM0pmMDFZ/x8f8KvqCEmX13KqjISrYelcmbNmheVvh/SHx+wa7y9WFHUmPZ
LLLQC0+upKQRDPZGYWsFOpP2mBi0BH/Qk7blioztx4FCCRvzIFSPaZmN+FK1rUvdPcpYVPwRf4Vz
6X7IVcyrjFqrXR0BC1ovdD5r1W1F7F6G48Gewa/vxf9k9tF5GO/YW55VkHoy6yuGMu87LskagT6n
BrX0cFp/9CsEWcEaCzRdYuMaNIsoZBGyluaucfl+W5XHzOlE7Idlrpbr/+aHik8VzFSV8P69qNS9
Y74lZplq8ueJd19vfwy8U4oTOXrOwOvjwPmaZDQoZkRkpsewR0G++vsVHEPaS0ljIRuA6rCkgJQ2
mNDGChnoH/yMW6IQM//mzkaxu2bcx7RqhKyXbhhAt9CqK/cYioHR99PNcjLRm6kWZ2ktyMVME0Aq
DXm/4Fd0EzQXMgLgFW8Te6IRYozXjE7zfTAgrJGJWdzrqhu47V5u7Yhh2KJ82zyrUoLW3rf7gaG3
Iu5JURzQxK6UU0gDpWc5veDftXimrK3YjWAOSXvZ21RTpqkIipHTcFGIv3mBHDOtyv/VRtaDVdKJ
N8vQFD/7ISAZc/YbMDTYxhJK3bDThxs5jyb5H7ophnXHBcsusbE6LQvnv21SUlKesgpagetM4Ps8
bVjiV7738fu3ymlcnBZ+CiGnY7FgVYndXM02133HnJPZTS6giw3TFueVKiJ+/8DLnPr2S+f0frwu
/OJGdhF3V95lKYyQMn+UWC4Yab/Mn16ZrIXIISMBU/e1bZflQXzmUSMqieayTv1dD8nYzwvb6j5K
JDJp7ekzHQu0RYjqRlE4LWALXcRwo5HA1wlXChIryY8luvpB0AblUxe3V9ipeoRjy/qBtnKf3kPw
Chu/EeJ48YWqjAlLaCotUdnVMnCXB3wJh7RYbk5jrDfr3PtXZ/8TSNt5VqJfNZjGOfEV214bn9VE
fzX0hWDhAlczqrB82TPB/NWCjouQKVefolNw504kWHtqnslQB1jOQoWljnRKUQnJAwG3ZBFPzzDf
az3Va2tM1qehpiZM2YijxFO1hUPklT30XaoULVuRtsNsqyJVwYu+chgK77Soyz0N3imeKaW/l44B
jVNcw3JXGSNi+JjE8/4BMOebU98fndA4lGhaadkdsJkByXbZV723f2hHxV5Dqj5Eq8etB6bSExTF
7CmjggI5jj5OVMYF/RlMnmGd/gbDvI9s3mbGRydQOD4MFvfq8rXH8ZG1+/7U3/aKKtpNXQVzfAlx
ujKRzHt8dplf+iSYl76SRFOlQrjM4Wxj9/ItunYj7TSBuDy79QSY+LltZNDPPmOeOFDLQztXLnba
d/ejh0KEQdNV1kCl7b5gp+E2wIr9T5E7a49BAzWSzk3rLN1HF8ro6VcVtVVHmVt6DzOQmxlRXqX6
2LKOmItakf4mi2Hf9awvN8Z+VQE445q9KyG/4lMrRHSP4o4UD2QklDKOopcEqAjVl1XIiTvqUqQh
9R1annCDD5c8CDQTTL1At5nssJOJK9Fh26j0KMcsuLvOxId1x6IQ43mSV1/UXrlZG/13/bFE1BuK
69YEdUAoJo3VOgeQu6rLKWppw50Wi8muS8WbW8udbFen6/9sjutT0yD6SDPdk78xOYQ0HO4UhYaq
HMNZC9SykFVDatbHSli9jG8wA97djcErlgCZ6E0wtvSzDHCZgjIDOKdEnztYclCmCqT6xgCr6aKl
fFkx9DR8W9fTrFOR2nQeZUAPmKMxJRgrDm+6hUxme9tBeDZqY9qqS/n8AxhOu4GPpfRYvP7vEqfI
TcZnNohPQzpl4eZb6EJLmzFGmUeH2nO3RgBd3FwWEjLl3R3elGsH/g84LcLcyIeMIHzK7QObEVfn
O/CHBJu9uD3Dnu6AIfX5/+9Pzz2JJmimWe/FZrMgsZ2e/0xnm+u9MH9s42XiA0Vt5Sm9PmtVANuQ
JDNyGBI8ZjYfMIuYQHH7qNn0xZlctYNxbUhRHxVxqgRe81kUJm/p0+P+i+Dt3UbxTdfmr/+XkMkv
3z6XR+oItkyHnricwpQTZG3o9aCH/QwPqh3oDy7kzc7oqNyC8X97742zLMK754SW9MAU9ORTMXeX
mPCRZ9/QR5nVUROfmiQw6nAa8fYPpp/T4eqfTDvXkIEbe0Dvk9siOKBb60ZazBpL8m5TzpjqD+ha
p6V1/Hmcv9EEWsp2kthw1frwzpJpHBjx825EmjL7xoEic7XX3mCyw4Y3bAFLMogqGvkbBPn3ovy+
spt446DtwtURQsG261IEcOFPXuaS/VBXKvNfZ9KdQZshAs5KK/lkAPqJm/N3fNYvgxYrwVX5pb86
b2MVCZkaJLuJV66uX+SXqXPPA64z0MDkGS60EgjexrCLU6dRHQ+N9Rwa8b1gUOytkNlUqmoV2EaT
qD/htZStghFfN+G/EO9f3VhjWCr5LEKaosdy/+jy0y/3owMGH3ccdAgz/jPDBkOpZ/gGm89PRgJt
g1rmzY2tch+VCoKrGM5fenDftIdfwHZhi9wqSbE1UROFxpfRmvMtbILIbyZ7Va693AlpCjoH+Dat
RIrKoLGRmrFtd7gN67v6L9EV8RqNWzShyeFf/GcttYqMvIUaIC6p+l+cS3EiOM0L01FKh7Nys9xi
0ZOgZfbE0GoPJroZwUhi/qLM2Jl16VaXqiYdKhKQ6LrQWhBOFzGvqGoMSU9F47ovIKY70iK3tPJe
TAzJa/7Ryhd77bBzneOLIUdjKs5XWNmD5jNnhel4goIsaR2y3ocqvEgmXRK6zZrlVlpQGPQZlTQQ
gn3JOj7NWWszY7eA7IOd7jc5VaNlpdE8dPlm/Zr0v8W9GzHL2b4EO360SEEtqrJCZRPGYjxCkbne
YLCPfTQQYen/NP8V9dNucqq82i+L4PZmcfhUgXl03RAoCFt/ut7Xh+s4iQapywJKxkqqHpXPCOvI
jr0hPfBUlatRl4Sm0UHTVi9CaMCo+Xq/pZz5n8DGPlqxXGizh4dU0ZUQVp+LeEmlu6BPJXa5ZceL
4LKRwnfr/ZEXweJj9jM/E4ORW9cyn300t7MNikcS0EicBpdeCUmsX4omKOTAZM1HZTbb/TicETdq
s98imoOwrw2n3Ykf15JmE9SpuyK8qaMVJ7vn75cuKc6lUwTJnBztM8twivXPt6k/MjZWuSKzQAXp
ZajV5zoLjq+YIhfRACfbNLdhs5CmV5b9MRSRbkrqtoU/nB32kdsm9931eOVdL+B5iV16JxbiVJ05
B2Pllz8uhPgrQVdf2i2Gk6XiMiL6lQzKITTSPGHX1L2Pk+rB9rZt/FYnxAlyzXLCFVP/wIAb8R/i
o657Z8x2y9dzNmA/lsd+uhzuOqLiAkTT3vGiB0A4NclGxKCcznYZKyPDagjMTpTkC/KXQJzBKAjB
cCpHXHVZTWWu2+FNfQqRptPsH6EnH/0CEi7bbXPtk+zvq2j9Daz+LWW04++IH1XIYhxGZAce8srb
woahk2QL6HUlpO6y1DdBW9MKQtHNYIZs1LPGuWsXh0B7pvLBMGZ3/5X1LXenA/O5T7R/zgBX68Lu
p065SaaVaEP4fZIFtPnVhQSWdIpMs0XodHHKosLmIMdREW33matl9yvODdc5J0wye7qTWATeue7O
03I8P04Q41aa13CT0cfQ7LIhjxhYBimn5rWM6ZOW3EuvKwGYe4nljcezvhn6kaWSSu1/VllEQ7Vi
G+uM9CbMjA4isFBJdW06dqg2IjVsPSaKNHPVd3kVofA/2dbKPwzHCs6zNUHnR4kaNOp6abTSnFu+
1G+eeloQl2/5D1kjg0ghPQeyqAPnduvJVkN2XLiZ8cc2SNj4wwwU5R8KTsyhBFaqhRI0nfJLjIr+
ax0Bjx4JZf9iRZl/uhhjxyLCSAaoGLuCgZ1nG+drBvdMHffnWpzeOP/AqeSsjQYt6+Fe7VoJPOSc
EBqGUfIytwEVfIwj+s6hQ1VZiq/hxPjks6LNqVyZnOMtXIQcyO+QwG6rPOYg2Abjy9vW8Mo8Gl+4
yKUOteNMB941orPHLEkCG6PhKTOCMbXrA9WIb336x2RvPnINRu2gOTHty3BlNX25TrITQLplRPIh
WjV1weSnMjTgFPkGLHEw9pWNfe4vmoGQ/Lqejfvg2r4hH7ozRcIO/s1Sm5ANxWpaMu2EgZXsB5L2
njKXSaE+qVCZLCJQeG9eReeTSqiwO6bf+6lzhDusj9rjCE/IQkuZdw05Xa+KWmea6jmVEkVksot5
qWYwINGthD6q3y7tF/Va2FV6BuNeUh/aW2xiSyHOSisrJYqhFCxxbdslQvkhqxeKeFg1sBpSYIfr
gvov+vSFKZABWUlZz+wXvBpXMNLsx+57muVoOt3yj6x5fBfEussAhxq9rOt5g1NGikAS2TDPtWtJ
SJMdjomIJw0A2EDjEqMKTjPTvwX/DIrTygl3GB5bvcXRgPrZ5Ohsdo/RIpzOslHV2mWaS61DH15I
oHX8tGY3hhhWU6OmdEH62vmvEPo6lr9F9SpHdFIjTk6guZV/hi9j2/h7bd1dDHsvf185MbtZsFQp
NCbDTl38JkL8Coqxe6fYUI6xBjUnY+d+BE+mwZbxNsYSIWwgu39MS5Qsirtd2yxtyWu6zFv+Ne5r
aiEvFoaKE1PQqi6VfqXC+Yz+qhlWXK9QeVUvuKN62Fbsrh3wmwBsjMVolZYKWeV6GX+55h9GQaZe
Ouw7KbHbSY2+2314inSj+siI5FmJoguPxb+2+FJ7tDsIpCjb6VyUH1GGnYc20p1ggUvWxIrGC+od
NoUF9MGl703XYBLmj1ZNKSgJcC9R075ptfq8YWNIZELG3DywqToI3ynP/e9+UhH445xA12JnAat1
zjV8CWah4h8wUrRZEytTRpXJMFxSe158ch9tRgCyGiHDoDSN7wGIInAW9JS1JmAtqrDh+UhTZVg0
x/YpHSFxXgZWC8/f7JhDKKWzd+zpNc6YmVgKia9Bw50Obwn/fHvoknDzIpf8RgRaRBOPthTXZQrS
lxTGVxFU2DmYwaWXCva1D45jYwhVQRQQTLncy/lOUMg1nPnYfVlmTQoLvFdZ7NE81oIlC0XcSq6g
DgwPDuFInmdvKYB6JAbzRO27xgfE9oBhFTMx+pGpe4QHIt8Fjcii8B4ppwbmnTASJD37vo1xNS8G
iqHGOZMouNNX1oONGqKqRk7hi/Jrc1+vch1dwU/aDBaFmxjO/NLsX2bo86o/pGxEzvhRfCy4ipP3
+Kr8AN7ykv06+MtWm/nFhxv4owFHk2vmxuuJxgdcrbsxrKbh0qHLYxmBiPqvcOBnQwEeAUp8q39/
E6rKiZrAqBuil/8HUzZpQ3p6GloMiF0JnKYwYVI/6atIjcteW6Hwl9PLD6yydAXhxcLXQNhMZbLn
pE+a8SKHxQj1l1XjLSNLQkmS3tmEvoz0DKoQPbpGZ+zLrsALgPI6Pt1GsxGLSo/GikFFV1EKC1nY
7wqlGtReLVkyXAKewDAhSdnEo3fnDyDAUWCP0zBQMf6YeRKXMuGdNT6l9cFIsdeXFWQUCLhUipKO
UkAkoj85pwoc4LEYlf6X5kreMcfd01RzBekfChH298mFu+OSJtPSr09Q2oFVGWlXjxniWn3kan0m
uHDBKlwu8n2xTHwaiH3eeapbnCK0mXwKvf3YdoTA56WzEKY/yt0JGYsRwgtWRX92oe4eci62lHW9
yZ2nv21TsU4t7AdwinCqytDzHaloIzZZfHH4dOQSdcSda3b6jSkK7dNQDfaIcTXjOn8mX6nTvyNI
f+Ku+h+TZa7c1aBTTSQO7Hp9r7qiXZ2TMsYqoCCBexHklsXUVKt724ISMpqQiSUwFEk5eIe/7qlf
Sz7Wt/FFXrwy5dQkyWimYHz7u6NRP/YLEH8v27aoJr8INwGU++VNqY8z38NasWxju9OUO+7eMTBN
RfE+9saYZ1gdHPIyVIRCBd5DyCpixaacA/j+SZUrmTAfXYV091xl0ILt/dwWdmpz0b4/xel1Honv
LubIjfZ9c5JCx6MgSeKmx6k5qHKE5pFDNukVCH8R9FvxhRCffE4BX0to9fAmcDUl4c+udYBP+VZo
hqBpc0gtXWkstAK+S3ty95XOHWjFUUEzmx+PAiMG6l3fWlJP8ESsDXxvWhe3oIurZfENwbq4r7rG
1/ojEH9vovT7tmiQ6agY4Ueci1kCBiYUFISPLa47gKfxnyRh85Fd4O7qD6HHk8UGNtGpDPetXvbP
DArzISRzQld+TX0UPqCt1LhaYvxCQdKcbVzuROe484wEg2zT6C75xtLrAQcWvJgBqx1eVM/96rxS
6SJjjS/zi+0hXTSdnucQ3KDxuBzTHSV1YHZHtD1nIcRBPt0fAV3EfkthOopS1tS9au2py0WZAd5i
apTrReUIwOXAU1a4cYgQ8TJ8GIpx4F5p1AfzeTWwFJOJeeQkxUWqfs2Y2/mbAHrtb6rHo+a2CMdl
K8FdyWJTjYd0PklJZ2QA/P/QcW1bhnJZYfTwyVJJeEmkXzTIy5RqcRzQumJGTnf8e7+iSFktzzHB
HRCx+sEGBZj0Ss1G+3fZoVObVg2bgyQ9SLyUQJARVo0h4C93kZpcwi9By2myRK8wTsoQF0dUNNLN
lGokhhZ7EEfZGmYZls9vRnqe3/YQQyWy7bx1egfPzBGeAlJgQJ5J+68WyfnEzu1bz+Hk6sLhwzX5
++M79cPAdu8FNWE4rRbDQY2e3d1nKU7mT8Jlwh+827fNT8haO9db0Z/BzLKUAOcyYc5kqaIcUDVF
oPVxPfQJRaYDXL/JOeHKPKjFjoaiAI2hK+r46Yo0fDZZKYwbv09cvrjoPuE7LcpaeXbmf2GunSzV
plf3nuhuK3dhvqkp6hy3d9lGJ+/13BoeHPt7O4Z1VO0sb0/s8+ll7aTU2uRjrwrNGYPSA06AsiE2
lHPxFTiVjoVQN1TNzp2Zj1irzM8dOnfRjlQKryu4NLHjNCEnIItaXJFgFLE8RRgwaOgCDNMjb9ZO
P1X3xgLqdrEgZbNDOhyEn0v4Go2JInx05msO73Ybd3NjGJtRPe9u+nsQqP/9jXJRCthj7v2CHZlO
bycwp0mf+S9BbwIOSM5B+DkzkkbJwogi8+OCjlCnB3osfgTC/iYHI56qgnjBkn3hhzfJk9m4H65B
60D2QDECNOebER+ZgsGnoGY10kr3nvjcRcjVd/4K+X9+Y+3v5WTEm1PYBlYZ7b7+bcyVTLSTqN5t
nqM2KGayEWTQggQJcoJjxU1zyj+azdxkxQYPVLsgC25GGv8izIRhqhmp7NOHIJeVxP20/DmBfEuN
gmm/nuO3QVFSGUwKINO7SxJmVCj5ZPqrXxSZZW2e3LGp34hy53z65E+3O6A1viMd2JEZHUOFmQRq
ZV/h0GO6EeBU3gfOv43FT8q05UihAACqvSVDwnOSB4MuxaTNeg7EtsHAbQiDqhj4bzfcPUJfBPjm
n+miAL2YvrgbwxL2i8odam0vNMYWsaCSvOnfMjODbKYN83BomlC0qyTq8QV/Ut13U4kY72B7vRbm
eW8DEGlEWDYMwmWnPY5SfwLmCAPqF6NK8B837eY0jkR3BJqYEEqpthqoKhhTSbOt0cKB6l5m961/
JvbNyLKhVcYCdIXdeTODlg1DwNkIGnqnzXsDGOyMmqXql6QJPf/jvaCu1bCgdSFCbopGvi4PZGPq
VS+U7pDwEL9bO1v86T402u28OMPikQUJjiqyRcWfuvfVjFehKHbApTEegVrIAMElFWjs+tBBEjfs
PD9iHbsFF6Tx4WbFF6EZTsIbrlFWleiqutDVK9ljli84H81Wsihjj+u1an+PDULdI1G+z5+//Jyh
6hjkGckVdfokQzjVKnyKSNbE0szUvsYPzAWMu2FdLlWsIVKN36L+I3yQM1jFjjJEp9ghyYba24Fa
CjgysIpfwXEpfN7izhh4jCI/1xTIFFmz3s8zC7Tw7uGpJ9okjIAmw7y8HNJH+EDdDjNbTVaxuiSM
Cq7Qdxxbi57DWH8xgMvABpQBFOBQWJU6jeVwteonKt8KvUSe7jxWkhXhJdfdtlShxZepVShsILOf
DHodeNzSt0Jqa4PwBek+dY0GKUDsXvuRtkyg9ZuGFeKIcjt3s1HCtB5JmS6QnVbiwCMTzVHhOkTZ
TQ9nNOFKnrX/ebi993YeCSC2xxX8ouTCfXFrip7qkf5tfn2XUewRe+tNPcFdg/2qJuXPGUznUeHO
Pr7EA8URSETjP3SpdsJkpJ5KK+fe3/B+V6vp1vS6eCRT/KEFAwP5K7HH3Hv0WHfv3qUZ50mg0kHd
ViK4E2UXWBX9vgnbUYxqi+genYp4u6L4jpC+CdVi8GBEl8EdjLftjlntQjxRUNZpANof910j0nNl
Ya5hmVe9K6xZfa0+J2915HaFRbAvBNTYlruYGS+5YnOmfiNvJDBvrH+SW4t9f6dBEOy10uWrrhaI
qHIy+tadB3yf1LeTvi2tP05CQRlUNdeqWT9+HGg18JDuYV3tpq782diiqd/RBI4pAjtuIWx53Ain
PaYmHrbqkOtvAsitlXIyIFWozn771sI09anoF9HbGbiUICUZLQQcy0Q6SQJHQVL5RRgHrG8N0djJ
wTm/BmD74vtsODA/m7fJXnaGgo2hMFM7B6KIfBS8gRbSZJjlf8bWrlEU8WGeMkV4znlDS5gdiFTp
wJ/DvqUmubFKTk5OGS+fxi4FtWT9rnADTpfpNbeDhX9FZfFKrx0QibO9UV5hSy9tkuJQ19CZ+U/m
Dvwk0caBKsnWSK1Aao6+vqT6L41wZ7W1gBoOzDurN+TLBo+vWN/cumLxN7mYdkiHkyCXpItcYnaE
tiTz8J8lCQ3yRTjIxUzfQzCqRytCY41U3LtSxvaXn3bb0GoA+8GWyTwEv/Pzu2H/SuFBpsoKuGn1
UCDMX1EF9NyWrzQOBzDEnvRtQbblLV9/Nv/Cqs82CiOcGSqMdnCxpedvg+ayJYHWmcCbFZsiGJ8v
vPBWC9FcIg0lYDd9UDC7ch02TF9R4LZWJqCOItvii3DHfNluFptZPvhGrg3D+4MC0k27gqN2gdu2
H701u0PTQujjslhdh1JM3T/km0t2/R0o4zoaRjCkR/S4mOm4DYXwq7FUOe5RnC9WCQJD33aky83K
tGaCuxczXH1IP0AtLGcxCuWGtAjKbJ9sCTm8gMaXlWCXgYOOWDiGCEo0ll9KmNsQ/yhdwJ34YaUa
sqTaf6HkjFP3e9hzPDyEc/8Mqie4CNbxJCB2AicZXhj6fwJ7koMiekOag8EvkdW+bZxMIH1Xg/nq
ixP4QJ0lleC7nM/GWEGAuKGQst6qyWCUF256a5lCfgNpwo0+98mGb0nP/KiYY8tW0o7GPPcWXosN
njFgQLvgL9Y8ahXEV4fRJv4feme/h3cbDzjJkHO7XZsm95lKDsL/j/qLUkiN8hu+ewsGtyqSSaAI
V8hmGSOaGdnSo44EYojjhUFduFy/xWNT2hWT8EwmErczOQgazsOCpCWgdTTGBYc5oe6Pt3uTbRIQ
BxTk1kdiseWIe4TesOJL82QsIeYEsXppihBTFdiZ3m+gUsQBOFFkYd+7QQKv7MC9WPqube+o4x64
n4w2MLKde0pLgjZpivEg/r7APQr45teg+Lnico1z5k+Dd1aGyj8Em/WGisJUZZB1Tle68Ia0mLEx
cZ+1pjMITKxDrf0CVvnWR6KdrHba+7U0mFuROSRbDSbUw5yoMQOYJfYV1qhZz6QxgwJlln60XJ3p
Rgsrl2kdZCFku7Dre9jH0NP4Ag+Eo2MKugl64xv4HLJZBBs2uixSLfVK5ceOpeKC8dWhap9vBVyc
R+g0vPDmqGjhsgC3M/X70EQVIT722dO/hOvKkEu2pNUoC/kGYznyl6CYAVTav3Bgvm2KfVxE/ns8
ODwYkRnSwvJO/XlZkiwbGU8GvpvxNV5slPm9rAVKOlWj/KFQEJX3/Xl8rlz2+uZHKNyTbqgi4vd9
BrJGA4qrtsPEy6ifrkKl/MSJtAQ+crWRbV0RXTyFZLBNrA7FnCJRy7ZVV6joSBrN91g6zmwhpvG0
1oeSiU6ijloB6M2NU72McJpbxZQy8lh5+EpwDX6DlaU6fzLmDBZKehFVh5SkpQoyRGY4pkt0fpeg
isa0bwKgO1z+lqHYQN6grDG2x//+Np9s2rzzHQdNiZUej0WT810Kyv96WiUOtUWRr6InBFB8fg0L
Lwj+oK9A9F98tt7//quD9k7R4Wzyp3hn25uyqmhHPZMbls3fiGWQeDD90lH0GA+CKWGI6zZdFyB+
g7nd5r94Kd9D4gmbs30wZ8M/yuzmVeJiFsvMjhlBgAbuMKGEfCfwruIgw7WwmxHmYLojACWURr4L
AIfmO3JKe9NuVWp1xcEe0PlBK2CVYmoi12q7TE60VJi3YTU/JzdhnhnVUPkbU1kVNRLUtjdVMV4n
rQNdsF+QhE8+ZEvsFI85KplLWhC+5Ims5yLeihbcUuLsEFSIhQ13R6oi6Bsjqy3TQq1ZIhvQH2A+
qo8YuJZ0/n+xdWyN86fFlTgRgp85bHe4xiAAzbv7CMmb3yV/ADnKIfILw7xTjOGmbRk7fSSLb5fp
ehAQDAKbQuDddYkakr9rWsV0HoCQol7Z8Hx7sekO3SEelgt+miHvHxQZ3bVSv2eGGW+wpMzUKdFD
RQVpOW3UNOnhskev6g2SujAgF2Q8baY4Lija6cRHUc7bpHLJWWtyJZ/nSY6+jBiK+skcUumfOLAO
4MpeewOC2pHGsbeLOKdHJuXz6JkW4kBtLm2SRFNJir5eOQExzNAvh3B3tcTbmDmCe2K9KrgxXmja
oKapm+JMZZTu80ISyRho26pUKUevvq6Xd2/5reKMoAItuKy4jpibaB2uIAbe+mgEr/UcYGcOFbqN
KM2fY6VA1dHIVgC53U7y8pViMxYSkllvSkMofcVtu7HUHy4wY/PWGbkAMfntmtN4ILwTMtE4VzSO
Vk7gfHgVmC0iugjHMtLOMmHtg6B5hs/joOtm3Woe2I24JJwAN7yR0ZUjhsvIuHBkNaZwffc+1Gnl
5VoaG9jeL4ZIAfyEZe2DOqalpvf5BFld17uMwICyFqjq38ZkOIRibTXrHcanVuo8E0KaeiMDynRm
ryhY+b/mlaIcnWy70xMP0UgLw6d8O8+YvEdAZgFoDj6XhT3Oj7HfSmMyhkVymrhjQ2SJw5uMEUqk
6JhA6AfxfrDm2TqSbNPArlvET39Y6ip/QVhFOHU7BpagEKKKmqM8Mx6V8rwu7RwX27vU/qgP0oZF
PBZlRa1/LcVWenU48HIMx6+ltEMbEXHDf7hp+jWIZRApYJyYwSy606UbZuaj301Bm6nynCeh0EnZ
HZFtoJcfkRr3RXkIEKi5rW0SNdcoTuVH2z4hxDhIq5abTojwp/hhKSKYy3q5yL7rFbUFW00cuesb
z0+srcN7Yz4y7d+mO4vzsO4zauWSyzfURqXQhlEMWdjnR4P3ISwcxOiSJnp6YgLGfULYV/NIbryX
1diqqlit8nlDcZsR8/Fe9rMnrZZ9ewQSrB4+ufLhi0IlGjCYfGBII14EA21DvsL2M5IferVdfsep
p9O6CsxY7zmUYv4SS/O31Y1cCDc837uMIp4BtR0RTTc6vBimd3y2CU7BDinMhuJVbJyMFNUNfI6p
kw5uvNuwnLdbsfogrHg44zTitKHVGVOqKmot34CNqsNVa0OtDhNlmjpF2yBSiouc5+EWiHgn/rVS
NbdlQ8BaKxBX30n+NpPOLSydLTjA/KU7XLEAmHU4/L0Xi1KG2+ETDnGN+woYjm/+r0qGabR742a4
iLtSuSgGsx0M9+tFm+3MUHkrfVjDdcKI/C83yv0hig1o7Y7Dlx3hhRsOrHIruBxSw1OGSNqLiNyD
NoKpM+2t3+hdkjJy0UnSJVznfyWyC0M7OK8Ivx8GJNd1Kb3VSJTLQWZgoRPxsR3thEkUabgvaBY9
9gBbNeJYW+uIHbEhMd7NqsUqk3rzcOHw5M76/YqV/lGjYDSnBQp+F81K1mmipjPy7tFpzoAXrhO0
QhfE4scQ7P2PkfXW7vm3L1mH5sNv2oZfeygAgbOjBIuD3+eieW6AntEZPitLqb6A1UquzNgC/bYr
ogsyu63a3llzGDfk7+E4Q0A7AL9e0MLw9afq8WKTBKexakHK2MXzu+IJXGX4aREWNpAgJkk6gh0u
ZlYvT+WwJaxoiRNPBRDzoc2XkPfHMUJ1aDbkGaEYdPXnheHCjZMmiMR1pUBLieB7Gs/Atgt1H2RA
xC5+1Rkbe1jxmDPgk+IYA/wMkdZCsqU47PuOJAuiy/hT/5M7BgAgwsIkMBHVBO+z2oSOb97Td/Hc
ufXhphRI82/VYXHeUiwybMrq1I90ioIsj3VE53s5OeGXkOpWuSqDsapM2M3LSo0yuFyJBLq5qORL
Yix+idhKckEgAbAtzvDjszoCfeiTG/3UJuGehf/4HkaJNDSVPWzJOdIKdW5M9m1UlBSmNXWmSVQh
E3GxH1xgUnyXyq7U+EfEDT5y30PXsnM2ZkF87x0QmJScurP0b+SORU5zlVhbXon8vsyjOqzSOE8x
jrBO4jLI+JFYyvrDy1dpaEGQmRbJ/1YsHTcUA7zUjYqkOYj4Hzu7BXrOwqXEkfSsy2upWXh6zEmb
8srH3wqx57gaE4OYhkRscROI3yivG9JsyYPvxYU4/E3oP7xvmAI2av1CZGA2w7DMpPCHDqim79gE
glNqiTN3ftKTZY/AJa0tv/hQUIUA8nQEb/ix50kYEB6OvLG9so+Z97YSBOG5hXCtzVNwMcY6SHPT
Mytco2SeqmypYtmEG1PXJou/2mxJYJgQaNaRuWeQc6ZAjcNvXq3EqykqwZo4oNEuPgeEFLakxuTx
LDIlAhrWGurBkfj2YvadHnrM2VlmxEMMTNNfBh8pUPpzfkg6Wniu90Nzh68W2H50To4n6G/TIzNF
C5C5YEuzvh6YgnDqA7FjYLyANt3Ulc9D47INbGKOQObdxyE2tFs/eRORm/gxP98DAxbNZ5tyEwmT
e37WCVOdN8ICnD2SrwPm6Sr0GJ47utjkr0VP/rc+F/a9DBTCEGp+dGycxYFPAxNUOLeVW0mUHMai
Fm3Xn+IuWD6YNxA1z3A+R4zX0ptiMG/jvpddbraquYqzChxjJfYu7vDlXRf1snaqnBlUhgmbV6gq
z02GaVcKcnTHBlN6zgXbdcxZPBMKmFt7GG7kpYW0X0Sq6fI6sV8sPr77D8R999ztIrGv7c/u463R
uXoVbI5U41vZnVrasgtUFtwtRn8MsOLt5cqo6swQF9EeGMz86CM1cJVTBDc/UfDaY8YPrDSQM0Kq
xVg1DFGGEqIxt3ZmMW+8AM7+Z87J7lGrqs6rfsW9MAUxBIt4UTZXwBJTsbuMOykp2a0Hecl+iHcR
SU2DMA5MXZRIUj8dJG3eDNrBNtMzbC/EXhfcPGpeeES4/f3QMWKsO8opPdEte8G58n1NiwDtxXKh
sf+82Sl2i5w5bjN+VQNfjisJcAAygxErb4gpezeq6mm8ZMPVjpmMqabmkpLL6CCf+Po6921p+oop
8PiYe2on3TPaU2ODkA3JgsJZp14s64EDwu6g8xf7BZJiVVmeEQmYJHfbU7ySsmLHbiDgCdyRRa7E
9PJb0uLXUF6zqVah3TTjn3dfcP4TGiAiPGETEiDYvFZHhr9z2hN2b3NihHhh2Tsfw7W3W+3ZwvCZ
EbSRRYn5kjRi26x/LNfvzrxYrNYNb3y+MgrX/6l0iGcqfBoTwJKTuNCjsd0upuh4+7WJe+mu9++f
rKvOe0njPAc2XD+iUFwra5U+iuIE539ltZnklnpUyvrxEiMGtacDJA6L0Z0TYk4O9NkVZRdWEu7Z
VhdM+fUumNtK+k3omajRKYmy/CECYRhv745A/FdSqJnoE296cLf5YKw3KPdWmG2Vc+9/AyT7xRMy
4qeN76sP0ZKbUTTG0lTzYOHTw4QP6TvLoO6yjw64nDL6VlyGeFAAQ3w58HpPKwsHiKTiCvk084TB
6beXAJ5uwgBbD38bipKXPo+PE6Z6/rMXrUZLDd281Xnn54q988Y8w8GdZ6zpxE2VJL6X1NLKUPgw
GQz3wIHITM3GyWfa783Ge+/4b7itpo8F6r/hqqdkrSMdjQVwCkGc6ZTFxNCCyxlyR3p/Bl86jIJh
LLOSubmNRWeeBh9r07FpShzP76sTXibd6DbJ7h9gMlA9qttrDo+9B4eOP5iyccPPn02gjCE1NR8i
y5FdCPsJ2cbxj38m/EIhVHa0I9+7FKQ6YDRc2/t511K3m7keDfrj6T5z2Sak3+FF6NvxZoPlIRsN
/oUWLqSQ1U9Voj2pYqcl445dfoCgdRp/Ly6fLmFx6eZBl7noETwlzODIc86l6nqWQ43BYQP//Qvc
+xrBw7eohsmmR++TZh/aWyoSGjDv+1fMOGiL8HuftwSN9nQ5d4IJo3vMqYwm4/A8FDMbCh5/xzZJ
jc52khozbqEbpJZKjiZz4mdyrNWxnAVwtPCdoEaO89k38vDR07waIyoNImkvS6FV2LL0LcBNYD/q
JACYrBEm+onsHNX6xeuBQEwiNY+iDBMYmo4GfzYdjLgUFjKLC0JcPA0bjboPoVeM78O2Ep4g1jY/
zgPxDzDctmpu9oRt+ihLTl7Nln/rWxt6N5ikyPQKK6IoJ5Nu4g1KnZaHwBOaBy7jOr2WT2q+AEmz
YIALWfgw083fAOO1QiUnlCcAF2MHsRzmJGD3eu6b70j5o/6L8dfxVjP6D2WGoutmERerQazcxASt
PEEEV2AIOyrHoigAjW20cIw8yATxRaz46HKOtBHA8SgnnXn2N2f96KitFD2KFkceGMJ02un1pfO1
nHmv8QhV28PsfGtWThQg1fvLnEx6BcIU5y1ytGLK8WABMEzT7oeJZUEiipcS8gg5mHsL9FFOe6nH
Q/Nj04ih79Kdv5NakWAQRJGsrvSnbDUvJtkahKmVaZafyz5XjmV89iWOTazvTvWstnkE2ouj1xiX
lVEa078kX62NKpl77s0yS8QR0O+Z4yP8PImcnFuhMFULgw3JDXugydw/3Q36gBzy6jEUHBg/NEE6
cUuj+EqwFHabXwzSNZzPeGBn6QXIxJTlsGwGR8A8HmQN+ErpCoZyoj7cRAebQUv+2j+JMeBgeGUT
B/8JkcjSpvv8cCQSR8P7MX/nyw4OMATS23DYanS0hS0vywkjXYC3f7r6ORmGrYo0c9tPJQ6Ubu2T
t8Rmzc4PiP51FmRRu67Pbq0Yan+HJWXWksZiFe9JTuPalIuyN/o7QYPRte7XyQ7CMCVfMzojEHko
8NpVbSR9rTByRwXB4Pa/kgvzREuINzb4G3J3htI+MBhz5npFSiaL1ilMCFDwvCfVUaFYRH0wd8kQ
HUcFzEs0kfsqgN321TAbXH3ddpaICLJCM0woITTx0qreOkP48PnLiUAyMwKqARbVXBLqZkdAb1ig
3hLXLEn4B4PNfvmTxF2BeGBAAUdQb8QmBWCNXndk9BgfZZA9mK75YOSSStnf5ynt+I0YpyhfVBzJ
skf3xzJ79hAAOHvXEtbeGIzZcuYcu3Igwz4jN+JlIn66v8xtl6KApBXihMRp9RDYXeNE/wZvEsGs
dogfahJmvK3POSCYybH96KfUDdaQohucErzkcoW4qTLKq9mVoCXP7KujEdq26zqpIC5y66Mf2p7D
g9OjL5nyxGwO98PRQgUDrJ2/ZUcKkW8wJ7t8aJi8kdj+Ai8Fg2I98eDsb3R9FPUqRzkJC9RrJE89
lgoj1FZw6YC1T/1hKJUqMIJFNYOs1k5tF8QloSZBkCExzWtYS+4f6dBejLNLD8ecEaUsyWDql+MA
Uyi6UmZnQ4dPV46YuFvqYiN62Q7svRTk5VJdHUbxTOBQTDGUOi6/V7iCCVWm+ApFZjGMtrN69a/L
O+g3bbK5I6QvMKGtdbnkEDXBevb1drQdzIkmk0QX2RkPaDrkfwX0k9XXM7AI7F0MPbaUQIS2CBCt
gCCmOHH4oYqym6Up1pDPrpjIcEzP9Py421dIOhk1fbgou96B7OGuQuc1NZhnuZ24tmx+ccqCYlsy
LB0ZznYJvX1ST6kDjiPEzL7YzUZh1pZnipbCVtUPrO1w3Ij3TrK8bmYxnqZrUZ2BMAa1HwnrBiWF
KQdct1/T79994GQ5sqzO51C9qEqNw2TU7VLloNqIBT9f2ksvqfYWWzneHgcBG0BHJlge+XRkk3b7
7GueItoZxzf9qmQszZKL4dpU7DNKWDj8W4dqXyvDL72adM/FVd7551Elqqcj2FWw9rN7/r9SMf8W
oRdx37zid0RgzdYtLKgWy0LhMDZVMcV8Fimdm469DkiwEWgOG5KOajLfuaS7N/GIg/A01rHuO0al
bwwDOMmFnnneXz+RfvvCx1wK7MsbpOXSxRFMrg+MIprLlQ/rHEQabk8dpvB+S7Em630am1Yi2Ytg
4o+yj/ea9eBrEnRlboUiHHY0uNXlD3l6PvxvyLwwi2+fbtRPuSovNU6b1UVl3dumWNpWru1WVzOc
sooe7faAcfM0asL+vEqagmOK4kaZII5VuIDp5SuCBKxt/Nt0jzVvmhzxLImhCZ+ndgH31zMnEbB7
hDUQAzWyFI6zhFuNtVhl14evRJjE6b59EoooewjnU0ZJnONJbcO9X1uP6CWVfWGejzz8DBjQJv/v
f5DwolWZFkcT+QDLdDKkZ09mEiCqAiRab0rt1icN0ZQaJ9frojjbGLTS4oOQJxxXaoXkud96x41P
UDnBe4fGj2/3rnBTLDDa5Fi19SoIXBMxGHcg0+cZK5OWLsaIq7KCp8T1lIXlB7S2EgqymltFDw+A
ZA/OETQ53YOp/YPrbmjmBLgC1jJphrv4ABfGl02kjRivqCRU2fGgDFsrpRm3ywuGPsBdl02cX+N5
pNGZvpSod+8rCt9kWTg5zaHNnc5Lyu7ei1HYlboVYLrfAavrvvP2NcDXMxosCrZzUK113GJLQI6F
TRv+13zHzg3fRxl5QlENjf6JJdSqoXk9P5wWy8sbivBDgy+T27EKDjCx04cWmqsjILdg9Zb3o4Ql
Sv+g4omRfUK511Pb9822uKv5gmo1/WenAtnnEcNxfm2g5GDggZzLpi0verbGDaY7O9T2lrVTeoFJ
sv3GDCGqDyUPArv2wHjl7cGdgadcwsZE833mx4tt2m+TzalWqNiHzkRYO22XBuTejyHAJeITIJ74
kBuRWdxhOW4Zzz+Ow3JFJq42Lppb3Fnx4aQS6/rlNWEIf5ygUn37cq0uofenTtJy8afSJqZGZ073
CCxvcIgxk8aeQsNO4w4e2LkYHpLK3LEtUs76M/AIJSA7EVTktFbLapkw888Q/vV0NYVtMmG0lMVv
OqH55allZyDqoZoc7PeWjwnfs5TKD8C3wG31CjjPrmo7rq+1m/eSmEol5WdbaGgkRqR4egfdNQ8c
W/EinYH+Vh58zxuoTGYa6Z/zOvg8YV3F14gZhKXOn0bGmlf9au3jMmFMv4OKXgLLA0CqgPdQFlTx
GZA7T6kKiqNJwUDcAvEfB7Vc+GQiwPS6QxoRDSaaFz8zC4CMXOJxZt4ACU95lc6taqJyOPIqkfdj
fP5guGwL5yKUIYZmws+anU6zPJGm7FWhW3WCPM6lTvYi/ZI7XFx5rfOvl6wA7/9M60HQdknvi96Q
H3KQgPyDKS5DdaNM7cjQoI+b0kYCxVhjyNpqszRkMbNLcnaY6vcJnMYOP78rmWySE7Nxj3+opGAy
VPC8SWCNAuKW9dgjN+nSbPugMDd7GdALu0/iyZNQ5dljwTs2JNaBnz/XlPv+gCGJ/0ZbTh4YOOxe
soSTJkmIenTJ/H7SP8kLMMd4PVjrkCkpcCxmzgnz7tVLwgR9gfKVFWeQWNscA+t0be+/nQth2qoX
SrMSI2z3HpQThqE+ihCFxkNvbN7FsZBPME+COXXYqjQ8HAVOj+YYlifItzQmfpJFremSR3UD45UH
xjnx0Qnlmie5fjvvjxx0IdcwcfLWCfD8gDUf1/1KHVbB5F+ZIVeWH3f8SZj6VFSIKBqovctb55qi
S+pCDtfBKDkA/EVHWKLWb3Ib2Wff1t1rbU6Q+C3dkdrDKfdOFrMNhRSqODTRKsnfjuM31IJbiz6c
nztw5CZIEEQSh1/OARg39MHQsT4gRCaRKeCrjo314Ak7E2Vl2c0dUgB4GKNTaPaM7RzHAbnpQt93
hWoAPIkskCKqMq1O8DYrIU4A6QWhiwcemw0w2gGVxiLrbr5iT/3XsOA17AQpT4Xhzw7WcQBfSGue
apRPZ3pMo2LyPe4jp9PfwuL/V+D4Y3A6sTXNd2r8IsVq2KIPPQz+80LGRRzCI3Exa3Eyf6Yy8ufa
STURs3ybTkzT1mAwTS2uE4srTkAOS9Rt20FWZpk0hZjPGhXbUWXWJsJyrkVdcTUd88PfMrOIwkw0
PNAvMHiIfpvAcyAUaJnu7tPenrXjOI4XkG+tTHShSbd8iWtbq1IG5QI/ZNLLS3kjOrvnFPL7p41U
yXQ+4Acy20WcaV+Q5+AA0ZSaASagfHllS7x31mNvOd8fSyx8xWPD8I7a/eB8wcIuZjfAaNpL1rvO
biM0q8VEuqVMQd6OrTaaH5Is7b3EQmkBsXM1SFiEorhtYifC9ieUZwR9x22jUI4F3lJh/vT0fFKc
83yioEbYPGhn3tmULy30Ago71AmJ85JLorwRYkL0E6R7FhbIoahQp3u6PND3Ta33P6RBOsgEO53h
TDPm2ReQUtXjw0SOG/iThyxwjRZOBvh3JpZQvuHpjYdl+qgGEO2Ts3Irz3AZ7KEFLuAaO7/cDMbp
ARLuVJ28PuEGrsJM5q5uXqp+KBSyveLIZ1hasnvoLQca9pwK+thRDRalWcmgzGBtaQcKRiv/a9Ah
T2Hwt5xmJxbUPXNpPSgnItlqPlCN7nbGyi+vnlHLCoALsDZKkklkvzBffjnHain89ZP9Jk3fSycu
lk135Y7g8Sj1db3JNvfVTYftu1A7BpWqkE7Gdd/6Xinl7xX98ZYQ4rdOvEE+Wto5hBuFCoqm9GBC
VDjT6hBsZFJbkFdnBeOo2bH/dD8lBXqgWhAfK+I5znCFSN2iZQKoJ0wVLZvTUaDtZelm1eW+ouwG
cIZgZdttG+gIDcaKB+VyyBzu3yHgddsMbvqeuwBSjh04S8XFKeNCs9LO6PTdNd9vGV89oj/g9lpF
jlL8h3NqnINRqDMBiK2uPK/K/TpMl53rWxH3lkSmAemnmgDCuTKPJXUU1rHycqiDGsY1ChRBe2BD
8JhPhfSR9Myo1q34D8zgefZAO+3cNnoJLsNjYdO2Yv5YohoOKtdthwAHRG6S0taExP+M/4p8x9x+
cmUlWIqXwvYxgnlNXrxizHY5//nKjZ+WXsxlNZNvdt7cFMvMd6N23YYKMivya/yzp+m7P3zNr2e5
N6nA2CYJKzsw17hp5azIajok6EsQCwe3D3qUWe2rRdvLHQCDEMj0Xo3Is3oKHWTQqH/ZpD5lKSI5
dZvEuYumoJ0zU6WDZqQ1ix30+ri9F4ovx+Eu5LLsv3DAUZR58WTcN/ynphmPLbsgPk7HgpAONHdM
nIU4D/iOSiDwDOGF5U8mBkyS3u3MfALjIACKob28FvTXd0/caDgylqhPw8TP7HdIno4MBe88e4on
6mTFBGpCnSiJC2/BFz1J+mjyd/TfndL+wgjBbZQJCmj/Mtuc5W/xGtoyvDEggPTR6UgATRNxdhUX
ekIkYLtfMjh5+ML6KplkJceyIWEnaqRt8pywf3kG0wD7s6aNLNn9Fc6SMdeZd966FfyZsEYN9RTX
n/BurJzPGtbF5jh2WhEDUqRFj+SZWrh0f713KtAYwTMM/79ty5axX/aN0aimAzWOaB20RX9mEV8l
h4Pbw3To4JvpLC6zMdkrSFV6unQhMM1aY7oyTuAVyGVgI4GRbf4qMHSmDmOHsv37SUhJ5/ClQuo2
umhOf3qU16RIekUScSm4KnZ1uNG1vLnr6cTgW2utCQoJdLJ79jm9RueoUZEfR3es+kUyyTOvCj+k
iWjYxtt58Hzr3FtAxciezvW+qy+sN9N315XNiRsPLEUxhSA5PiqtM2FilobBWBK6w7g3Xb7aNX05
cwTV5rSKQvdnkRETN7XtRBqpwga4gGi69Sno5JtWYt1gX2qH+v7aLJg/CeIh5uU0MKOhNfbVcpRp
GO9tcmy1JjmAqXmD80FcijmZm6tqZcyBookK2HZv1fFbtGDghm1vhBTzL/3N4Y45d+LAuy1ltn5i
5epwn5OCksR5ECP9v8J8BRN5qFfpmIlLOtcnBg3wIA1J4remTuXP+SykgK/T3j0WNKd9BDGOJagD
YGddJecilEBrraf1VEFKzQSZOeJTXKK0/SjO0dPvWWmZIZ7WadIhqS+xyfwtyxEfpBx9koJ43jaP
nK0nCb8GEdrOGl35HoOPETji9t0uvj/Le/IgVuFZrRLFVJN03pJ8+yN7+0Fxp6PUPVq2cbcEfKLu
4UwCx9bVYtniAgt+0T+fjonSaLN5CMSAZrBOHJJX6Kx/5iyTMT+KFayIDtBXP8V6tXIDOR3FR2X7
sjCfhOf5KR8v4i9bHLOBX0FbndMJDETseuhTenAiwPtiVXdKNyHrfsvHzi/nA8ih5IdDY2asA660
UQRVxUm2bxM5n8S6p8pE7U+RsT/3neXBO2gPHGU+C88/MOiYr7kAA0e6mD5RQUPve4SN2qAJZOiN
cgoR+j+7M8mHmq2QgTRWi0lAJzuje1i/dr1ItsVbdNrk0k2WVkt8JtOQCZBhBL6b9pg1qFrdOc6J
OpAMXd/MDgsboBF6ewR/jNZ6ouY3Tcop3flGnczINIT8EUVQ3C3ahlubGCE++FeqhJomJNOF4mB1
dXymYwfDhNog/fgPeCQgK6ykKU8nAwl8oOlGTzbYjdQ4KLQbtQtfOQdv4DWNF3z7siKaOnZq0ah9
ZJvcGIFL7lpC8KmoV/mzbf7/TlA8j7sozq+lKYW39RBUXb6isYaCAiJqGAoI9Z0KXORNHp1Jl0L7
1SEw7GjKvWDM0Yl9C9PrvzP2Elacd2mUO27Gar8upd6dEzm4B0wPGIdPrbi92O3DyICzjK2KnghQ
Po3DvmGf33IaYuqT5XSegzp3Srl04HjdLYH+FR+LmcQ99vj8jTB0vBVDkZJzJvBLgZPqQUFtpqCH
TVyhgly02/9OrZuvoC+Ew2K8lm1X8kwugUtlIVQY1mVUKKOeYE/8lE0Slj9/WmKlD78Gh73OiCYQ
3WVuGgndqtQaeIGW6Tyx3Z+T6RjmHyjZqbsFFZjmhiweqIG3c8t8DhQaOgBx6oWOA0fNHANBL+21
iS9PVep+ZF+fncd9cEbB8XVI/rWjKckFFLQBBgm/skiNHQjFEH8AuImTkzZV03vgo28RRRanNyHF
K7W8oaZNJmOVs1QTPuNPfjH7Bs1H/u3DGgkOphAzUhmZr2BQ0WldJpWqebmYtFa50vaWvUrETqSr
9o9b9W/ovDkHl0Js6ROKuWnCj8I2vZRG80SxUh70gtq9FgiByPFgL5caslYO+ZArVE83fbgeiVx8
ghAuuQH0440vcqUmtIYAiLhKR8SqGFpUzE1TmAiBy0v68VgTfXKK+cPs5rF+kOdi/mOg/kQLxBoc
rWEBeR7D3uYrFc98csGTIMZcLvNiE81M1Wn8yNG0VSBzkieH5FCVmivwyHSmVsWwH2pq0TIr57aC
TOJ4FGcWAilBk+Y8KTp9IJOO1xIkUc69IBd1ojf2nYhZQZ04VC8OrA8936XE2PPNvxAS8qtXqfbz
UU6+SU1kPqdJ92tRtJdtc5TgwiiMkFhO+cvSKUAIc+9dN2Ml8VFeSevIDpqsvu+ykACmIUMKAcKb
A3+j4lrgLed3jZEHkzKsgPMnmJX0CkJ7wkM/Bt+Il6lsMmlXbQtPrwzK4Q4DP+rBQHVK2mJlt8Ua
xvQCD/FNLtwiff5gs0IoIqIVxqvPaCRZ8m3p1W6f7Ad2pZGv3HwwCJqnKsTmy07gNQglJS/LxBoe
2uXyPS1qex7nqTx6U/TpkrGCS9lAG69bdc/PPda4UKkDtew7+5VglsEtEvlyB8tcxHszLwwe4h7H
wTz3qKp4rauCdxLc8sSEG4AQ+0iaQ/iXI/OpWqAyp/qEzfxNpuvwwYn8c9bNMRyrh2dzZlh3oSNf
pB7YcB7SB6LfaoeYfIZ5YYFcv5Kr+/ZbGRblFe/awNhKO+aYg8eBSDzVY9O0XSPod1W1S8qOoUJA
TlsAh952qEMBFOiJwSWo1h441a5Eb0Qeo0erEQhp6WErp5Z7qwq+c1x+nUMSKALBR67yGkt4IQle
FhDQtaDC9s4wZeBkEKfr9sWWwVaMaW2qzd417d6rtcbHO1OsRJEVGU2Fw3DYe/vx3REPkQy9Xfyg
OLv/Z8DOozRv8EuuO4Y2MDPWQ9MQDQ5jpcNvl6jGnfJR0scUXUPZUCa4ZBvASsm2gPX2HdzmvltS
S2n7TF0lxwvNZQWenU50IldlxrHonirfhAJmYxY5mv+dn7wTyt6bc68EnnJjO4kh1QN5771NrI83
JPGPyTgbL0J+5QRUnEwm12/5HO6ZrIY5HNKQGq4pDA7uqJm6eFUJaWZcJNfH+MJWsLNbGGq/I5Yb
0ulpHZYg5kSFIQc8JpI0AFtx/edVpVvXMuMcbyVCu8CcVY2JBEu3uBdU7jK4tQh5cQHecQ+wfsLM
m4pT4bega73esyvdIEcyZ1Vzn40fq6ZL2Kn28+nRE4NEoqkBvU/vdjMTycZ14TH5cQ27gMPAQpGg
7Z/uCuu9O1YxM65Ifx0K5wV32/R1oszS1L+473apz7yKUmsDeeMipqEJa3rL9aDQqmcTjw0TnH5T
NvOEjZzoFmagBo6IlFmijxIXaEyRzSGqfeWMNNwOkoymTxDJTtxpwfP8vWq2x6cHDUqliUkQ+TAj
4ulqBGjAp5Egf3r0Yul0E58LKkntEz1Jyp8b+nhagOkgxmu2Ogxni8aNBfozhj53t/VJW9bECMsh
a2JzOTHfGFkpH1Ft/dh38ERgIYDtv7Xe+WDlpP16e/f0V33Xo8q4nBS/dg2FcGUVTZOEi+/hlPg4
ItXiUGUJudK6uEn5sjIV7TJcFCjFRnQS4hj0uYjcnsnXC6RUAfZOKBzM6rxavQSYyx5pli6KRUOW
UlMXaxintdcSTUEv0xkHV2Qip7p7ePx/nA7Ne29I40QP/aTU2VSePK2d8wG0LOlcRkD4XH2IUl1j
SRUrf+TVnzXJ2ESI49s5lbxWO6/TiJlZOeQ19SKSJ2aEZGy19JM9H9sV3gtPCWreOf+sWCYT24zb
g/98lMFIbXxWf8mMXjHnLjgBzDMp6mtD5DYHnbF6IN35Qr+ZVHDNMsuY3ka8IJhysv2GO1jNpz9c
dAzCth9z7J3XmO034aovYBweDtsiV46K5FIl2+Bga7SUIA7j/CvbSVzK/8kD0bPsXur7A3LZ4S0n
t03wwe62AIlK61gOXF/SR75Dwb8Vj4/EPLIUnJ3tmMa8XRNDidIY5bQXfCKqouOAwIrR5qWqDTuE
PNJwZHOhJjGpPJ4iDdCmF96m4nBHAmNWR6Ey7y4xH8Hps33YR7Z/DStVyrSNx+KLO/d8L00UN4iO
M6TthilI6pBZB9HOejZHFzzvL3GxilSrgwlKE+C+9UynlLPGSuEuDDmL9i53TuCigzWsoBHHjhcX
IGt/uFQ4jFNYbL1/lfP5LgGjerCABcuHTegzA+ORlYF0FP80OAMErm12aaf2RTx1JobH3wlL05XM
U61yULaXCdQBB/xgtRXN+zMf4R5tcsC7SYJvfJCIfxNB12r8rP78Fr+OL6h40Mi6gxq6/965pEUm
ptcstj7cSB+ysqXoU31ghVZEO09FRiBh6uHCMBcmZCxXFjeKGechTA5OX9Wka1X0YIt9WCF7OW+2
1ixPi3ZAW7h0K+dA6/ZLnrh5qe5ajssK4HABsezTO346yUqeQAV4RfdXHTJBuM/LpI5PMQXYSD8X
zfgPGT8G3idKGcAFkpIlkC4KFXy4I3ljQU+bVY0nrS+XKNkvg0nQo9GrJUNl/VXy9NTtkriDENAX
UNqdqEzHiTrv4KH6fnwjMxpfyFM3iW+Rdl7bLLTmsqTQq1cvldvaDpfiim3fHgM88+LOxD9P6sls
FZJm7AajeFOPC57dYdzX6cDiK/+ssBoOIkjoPY7QjeEVQBwmusaPfmyoY+s+O9sID/Iuqn3k9GLb
F4XKeUL9Y5Aoq2naLBV2IAMiowq2ObIue4TMyK6UnGPZTyVMOMN7NiqbNKkT20I1CFv1iWehC9s+
OWXtc+bjhKiF9bOBem6ewigHO0M9urbH76lIkoPYNq/tEGHzPdaOMZ07b95MwJhLqPF/LraP+UD0
wvSPo3GReNwCHVH/V8HXLHX1/87/Xy32CX56rYdbTSbuXYO5hrtnYK06KfS+iGRLxw7AjXsVIOBA
ZZtY5/nH0A1/FjimNGZrV8/whRGgFtD+RqkN7ZzweURyXUnQzb9YshMzfDxOxQm5SDnKjXLRxLQs
CWllRBYlgo7ShytE9FWIuNCMiBJmoRB9NZmaF6nDyiYm5+P3u2Je9pqjxduPEdniElRTciv4T05b
IiuwklgbhewlFdoKD+Hf80QlnxrAJUbJG6+OGafCgMwRaI/vrY2C0XGhRuIuDhlDO68BzwhD6g4Y
9s6ruflhMLL9J7VIE+4CcpTU914kbuVFv9D5Si0oMF2mQCYBhary/MQowGGbQXS/X8aoefK2ptcF
mlSyh/LwB6u3Rtg7shsHDt9VJbZ9BUoj73rFMKB8fB78A99Omr+uzfga26kuxFDdmKgXrYKLao+r
1KUdwxjM6KOQwpAup9fC2wogi5WTVx2hQGJN+LQu4SI+hTbDaKxoTpAQ8OAZTS4TO5TU+YaB1F6n
U0awX3fyq2yofc+yaEvw1znywsWrErvy/8rwbzXlMr0CXA0eECT6jv+Uvfs9gB8c9gE6Mlb2lNqx
Io9LTMmD29b0a/f+8gPb2tcz4vM2wGaDUKCOD0WQdq33BS7fsleU1/6TbAa8b+MldxTJ7Ek0tQBB
a5iT5w21how9dfkh0tOoz+WuoUtY8bgEpCJGqoeQ46Q8sHpu4lXTgld8xSRCG9laURrqot21dr4m
kVm42lpwMIUpJPVXtMgDWELyvyH3DLtwegjY/Ho0jnUEkB5MYoTfTkfauRaeG0gGcO3ZjuYQACFB
HM1hLPjDVbvwPcGkq7c21MajQ3tW+0I00q2bvZcNHd6F5prU1y+0QoW66e+E83s1S4herkUVLyvO
1/h8w9MGQ1hqXnypGhfNA4yOdISaiOlhZRk7KXd77tEZe8LqQOGVqRi0qDIXBgreD+zNzcFds2kA
JcPSix7pcPKf1jY+g+UMLAeRMsCbY/NqEi3grO004xbB2czUTRWPOeL1vnuGFalrsEJ4fcy1MLT2
wb88s6ojG5eR/+rcx7jN7Mg8mNohJEyXAFlFUD6pbTp8/T3TMOitHvPJ2OSEq03vRtTHMs2htgMo
4I428VGhXCU89g3O051y5+D/cOwLbqS1JQcGIaemiNquNQbQjPbmi1py3ZjBz0MeGDuZdRchOEPL
3r5clSaoDiguVtALspJTu/TbsAzyPi0FW5EIDibLQIqL+Woz1dfw76pCS+SMzsCTmk7RejyZ/yjA
Gr8trjffr+NENWb3UPVgW0b6/6xEtiivOgQ+5MKq1KXZ2vFRrxWaKO2/AM1DWiIT6j0CVRfSWVK9
C4ZJ6jtFZVo+VeQU95qoVs4PA5DPRZo611N9YApgJn3sgWsQLO898Fhk5Ed7DcqTl3fIBZu0HD3O
ch+Mk+OBKkiiWCd0FRKeelae8pjrtcNMLkw7qI/AzbF4qtcAqVjd0/vpMcHXP2ga3ze8tFooXyt2
jm1lQkiayuOiXU6tATwEzd5IztxV7YqC8tGbl7HPmcSaCI4YSayfmI1akJtq3LyYv+77faf+sg0m
cEPD1NZJByiR2a8SBI4oaAyzKoh32uSfzmBR1h4Olxef6+hvEYhq4obVPEw/heg4+aIFJM1JKdOr
VE3NXIV1uASJeW35kcXgbB8Rh9iSuE8vka8GK/QmsoX1PwROOjmXYIhZpiamHoNyOWXhKa1eW+qv
ggMgjtxRuI+dZdS2HoGucwiil1ArNZdfsEUolUcNzIwq2OMHQ2z9WJOXIlPmHt5PRF06voDzsLIV
IfK+85Z66IBiM/2hU74QIW3YjQiRSeIwrfXSWl3Un+5DFCiySjsmyCvW4PfQOPC4/j7IS7Evi39Q
ZlqvDE4BgtghOk7JdotdeRoC7wryfNHIyAz/jIYgiZBGcIwvfmrTNJj2+jaYKOWkpiI+PwNg+LMI
IP4a13jQtmQNMJh8Hyow6mb1d2gkT+Xh7fnE2uxqINRuJtc2qZsePwGqRQec5MJWalrimxWSVWzs
mmfsekDGdVzf4mEkSVEu2sY3xoi9m9ptDX2NlkCGXCIketsC3ohLfPSo3BrLYKeudxNUEH4zjge9
J1ucpcR4/dvU21J+vewZ0S+Cw2mzeX+w7MWU/V54xpRWM0JowGRYw1pma4n4UTNKOt6N8T9F41D+
DI977isnhg24IwhjCDi1e9Y+JyZhsjBmTTDj1c2z77aU+ArdgfBPF/PKilCyBC2/+34z4ItDTOCE
XltVxj29JvLLHjW4F+UUr6hxJ4zkiIVZS2VPr1o0Gmf/lavMbpMotQMKuM8/me41jNiimMf0zde7
mNX9J1W5ZXrKWWsaavGrbVytGjKgIrXT8VNJyOkGNaVlg/sCo3lMRUKdsbCApfGXsSFbzOcF2MIF
NdwBzOZ/uOWnysz/SlqA8SE9lI7UuHmEa9uEBggNatr0IB+7MD8w8gk76znkoYgugi53ULTIx5P7
CnCbYl58S11febM+S7SR62uFqd39D/ZaOtPROJeT0KF1o1epWY7+KERov0WlL7piD8/sHAJV7TYO
+qxe2jkXBuSYtnQSfDLmEk5PTiGikbAFQsVyt6UvZbmlUN1Ki3kGB4hnXoRgnXYyVUszsPnJRglc
bDLs9p5WTvwRVA9oyIFyVnTADbgEOqxJi37EEW5+cyI1LzpfXVtXU9t8dQDlHW9RzE7Y8ZuXOZmH
mqKSFXHr97EvFb6ZpMPGuVvB3qiD7kVfzxCVb++Y9PGSmLzZ5Z0B3O5ES78W654o6usu2D5YkpPg
FtsLg9fgxOSrZl5yCHLOVd4tcowm/QWL4e3zS7L93RECHiHrdCaY3Vub6QUajNuOYVIllc59j4QS
40cc1Lrga5fRinGp88qV4srGqlaOx/JtT6ZYoG2N7ikiqkgl/mcLVfZdrOxcqz5oJQ0hV5nFu1mp
HpG+9qp17xbcCYh1Ajh9c9Z5sscL+nzfGACAbUWwcKx2FuOW0osFZgtua9KLIPTnmxOGKYkvuALV
l/rQHHX1ymDAuAffQ36jBjeKqtSUtJj51OO7bk0bDNfaH91PnrOYVzQZdZzdtKKspOEOeOidu+rq
q+d4IqSTGAlXUb67SWaNx9+t/qAi4vB7nu6RVC1kngE6RLcyQ0v5/sH0wIVsDe6gx5tGVDLBPRLb
ohJYt22h4eb0Mzq1lShb/7CggY0klSqoJ4RwMHFPiIakiGUrPOgj9PNyztxoPmqT9H4MTn/CgBTD
BRRkgvX837RmYBIoc5WA+JsNVmLIj10MfFM4o9PvR4COp2//6jtq+2q/dLMMYz/2ycox6suxvLWE
mY9WozxRmdsvZ1HFAxbESB/h7hRauSQvHk5HgO8PkKlefQdzo+GCnY/kG+ErtPMWajGcCs8Md0YS
EjO5bHOtmlZ8bPXhcN1sKouJQyeidQbY3tMnT2RHXaMPjx4sMbwQUJ7dweTHH5QWZKnbIhyRRatN
bX8C3jD/0MG70iW7cmRLQTTjtcAya/re2/azeLlXlHdJGy8GPTitt4HcQXQKRjhvHW3rDx61kkKx
QA5KKIB9yGThv53kQy5X9xOLK3U6sUeMMQeoyGJjcyqVXRvj723ghcLtIUPuZzjqNsFJhnuSgHWE
MbQKrHBxpJmIEsLsoMN6ag/8CX1oxVn4H2L+UfMcvc/8/S7Qtvq2qxo4+J+4RjNU93inPtLIC/h+
19BkF6qFgxJx1eSv9v9575w8eeN3wj/KbCVR0kcV4lQ/yCZ/o+cl2mTV/U1jbGCTnbD6R48cAf8H
kYU/96gRfTsx9z2yjsBU31egvWFzS4la92d6kZCDJI5UyGZmzwvIL1xYkhmHaZXACyKksTz0hf7c
hjlcXsuJWTsXjIaJFTu334PFJfWWWC158MfcQ6ujf3gwzoN8lKE8Vz9ZJqHshecoUVKVCGDXtAhx
d33HKouRY+KQK1JuGGZN+qWUz/uwHRrSxLMYs7wGH3oBvX0Qq8YI9ZiHXBZMqQWaQ4iRJCHhl81u
KAGE9LcZn761TTV+BuV78iXbJ4+Tc/Tqt+xAaLXipECxCZ0IXeK5iiPcg3ex9ODqtI+DF8znK6vG
viGeMsAvOjVD3zDACEgXME0ZjVasWax6DC8sPf12DZ1tDIxCGM7fDSfxcb1msPeUswW1ZgXnKXAB
JkWd4wiA122vv57VK+n5ofu5lRllnF6zjzJshWBFyqzn5sM9j+LbLYtlZm6e7M1be05Sw7AXFWvE
LytlSJQhbN8JNxp5piaYh39eTMVcwygqtzWpZLRC16O+yYM1eIpE08hyUD8s8KPfbPd4FLPTGehE
YJzybq+czpArJIb2ONfdhuWQV1rta3WADR4MxIkz22d/jX+eQgneruF8+ABE+m+DTpBXoYswzrE3
+RN16FkLda2x6xqMAGekpNRLUNrfGG28JaGfsz2YQaegwsPy67XFUDv7MQGrcDVvJRtGLjwEUwTz
aejnl4iPwl8zVqaxqfBkYEIVLCe0el5cVOl3eWmrQjVPPt5fdASmUlAm8B0p5lDyJZsjiu9kP+v6
k2uY+ioPFowEdxU82Vy166y8LuWyHMW9NdfbEoO2a0N4Q6pw/I24Cg8TPttDVkHy2rO95fVizJMg
fs8ApFCWViEQ98LfmrYXpqOYZKLXEHAbN9YkGNyHOEd7CeQHjF1g3HvW2c6MZW6bEEfaMcJnAcdM
82oZG5qth30ge4aWV4o8hSqfEkh18OH/fiyL0vedgQzEVq1tTYUzi8OY1WI4PNmIlpL6MP7UgtMU
Lhvg6MvUqVJayFgjWrOXkpLjpF1c2GKCU4sL9oDzeOh5LQzaOtuRMUOqVC3Kj9gVk8ujbT8aUeas
lD1B/cU/N/SeePVx+OIiXURPGECOQ9MZDBWg2Xf/+SuucizDe+y+uQeyx0BiJBbMqxB1on6B/MaM
drB/5eqtUK66DOdcO/zfDPZNvDBcdYB+VJyzQRzFSpSNfbMkNFWNzQsx7A4QbzudLt/oLa0ffmL0
RjDvsgwrt+A+khDBrzp3EvFFKe03j2rnUSye9UDYuvYzwIl8goHftb9JVxxb1MjPmuOn8ez/jg81
0JLH/uWRsJLREkBRb6x6vxwAofXl9Wap5JOtEiSGSL/1uzC7Cve7kQQGUvXlJNqed+AwzEiGSKPt
lYycB9fCLR1VUXLahZ2Wv6P58XHV5WYFkAaC4qnLCB3JgL4DamBiVG2bfv18WhBc+suc0Hj9lio9
hNOlf8CgAAU8b1BnMWY64P1VYwO0Sgo8Lg+/IL+vF3hfmSUXxLrzgAmgqemTwZDOxl33GcNMWVl8
vdhcjItbMxXZRT9BjmS4Hgrig8Ltl9np8rXjbWNcLafTVm7i0SGtoYWFcZ64q1KeiMymf9Ygrf+8
52+WPKm+LkBqEcfD4uo6+K6m7+R4U7/kdHQJW5MT8S8KvF5q8dTGkULpVQ0gNk9LTBtKIDDQeLkC
4OM4zoMqPT0kBK0h9+h1sBo2KJQqSH9+LqHOjjCPAVwcMjlvYPj4DtAApgzSWEC0B1rgKCwbQRZ0
5oTjLrZZYfsebqbcDblDjd1qhxkH/qFVvirKtS3Z4Xpe0CK5jACD/BktltXZ2VZevbFH9HCU4LYV
9YFGYsxJApLM7UlmelTHS1LXy0LNBjEBwxGPvyYa9o9EILD+D6AfkNZtmOlhgmWO9kC8wiZqciG1
bCZyi5EXpn+lbKjm4JGo2DhBhpdDI4TIal9SPJ4aeQ5UBt3PzvLW8FjaxXs0FkN/N3Tml2I+M12N
IERqiGHJmaKGwlmdWJ4QgDP1VWgsbbgarF3eisHq4jJbgbedQ7BjuI5LSq5M7fvP4T3cxUStgkXd
W/c3lX8stpriogBbP5cb/FcyZBCW5n0AGvYOfKS3OCys+py7gETwcoJuRLew3pZxpCxxEl4O46jw
sUCIKee5GDuWXMWY+e6utqBocRp7h+0bI2YREzIxpUwNaA31S5BA082mjU3ZO+UWW1GwwVw7LD0K
MDoD7cEe5RcdGU57dmyUsl0LCbmc5Em1GINU/QsgAZolAYQc/976qBZ7MXXn8Yrvy+h0AD94uq+l
e+T18/55hZ1uhq1Rg1JkkRgVa6TkStjT2NC72/PlM+7lrLvcpUs4xD13OJlL9Ly5C0MeMccvQmL1
wsUnOkerBPnO16NCkaLiIsjdVWtK9konPDi7vyVD85NC6RcSJ6hflRHjW9eFOrG5qTN1wR3Ck0vd
l9ZW8jB4q1fDEDmSXyxeSEHZ0tZuL4DeBkpxzTgQVo03ULGYZgDz/pE0N5IrIujanbdmZ+A/b/pY
WGmu6ll7qIRKbwyxKkebmQznB0B174S1zPs/jWaPvxjXZh+LZM8P11qjzZ+JXRB26ZdMc1uSpbCC
zEKreHcwU8sd+DovkiAV5lFgjKFwD8O5ICRYnoJifNr5s82H7ZSlK8z6O0tzrPW2JvcjvmgUJUx3
ZsYOATrzHNQ0kUy2GGsnf1KH+KOEHR++MAgnqIhBh1LNhuBrnhep5Mrq4Xt0UlRM31O9QBualeqD
nJX7h6FEcFCNDaIJIR4J5FkxxwFVE9DEPhd7z7KX4GSb14WUcmsNmqgV/ehi+j2fyWOdHbuXA1FX
QO5GSVZebjxYZ6pjYy2vOZhnzzr3n4Xmpedi2JrttBGp3AkOaK5iWIaBNzvbH/B01Bv+7JOEteKz
Edk36X5YzSEossFVmMhDdx6owOOMqWujv09ji+T8/icbgq9SHVFf9KwW5zhnngtp9M33wTZP0PIO
LrkTBGPnnn52I+SPoUM7PJsyTQf4APgS5d7p/WlsILC7e9Q+QMNb2IOHstEkbe+DkOLMN/N8BBxY
aXTHQDT/vlNnZk7Hcq/3vMrWL5A5Wjv1WRURuT6oRbrmgzsDSMy9PYk/MgE8wVM23kF9AmFi0hmj
8rGVKekicg0e1h8YQdWMu7vq8qnOY7kXbvh2RW6SK3lcn/RAxThbWSSX2pmEPJP8eNC/+qCnzJEj
WPv5S8AZ5sdZcF9dI8CYc+RQRmiETy3iw9nzN6+9i0qWOEqHpkSzIDoNHxR2Dbj7SF7sRAUNqpvG
7YWQOaQiQ1rezlfcJzTuEVACphUnMqTTHblSA/1AUvNxMU2BFGQMFACz9U1WkByZ1TUYtyvnLHpM
N43ChPWiq7ezwX+5gCe9suOxaKXpEQiyz8Xb4wmFGERtyhPslGBiAwwOncCz1E1unrdn28G3weiB
WB6+7Bq3ATR+ImL7AqvnbmfkjUpOl3Rh21hZkRGnmZofd3+XtDFn9A/Si1Mz43gHvDLR3wk6Ur2B
kgUYzLeDA+Wbc2Fg8OHktaq3JtpSwIeHdVZGNaZ1ycjxHXQ2yHvuVV5AZ4T0FGHCGDyVKboOWqKd
rDbtCmhCIxWKr1jjfmFoxPX2Xo2yQMT9c1p7673WXrmAPnNJ3INTP4bpoeyGP2imx/h25ndRup9b
pRVNlNNciP/6UF/TYiLJJMYS3JXa7u9r+yiIfhPQTIZUXGYSdzEdKtO+q1Ik/pBnyP2mAWMu0gyK
jYvrtQ6ml0IGZgG95aYYN7bg6mi9Ruouq3o6djehN04Lg2XsvkrBGhfeJu0mQ//Bagm0mGF1egYg
eurT4/+EEwnMUv4lqb/i4/sZwtGP6tbVNQw2n1NpcwaOk8GEzPk6I+DNTX+hlgTe3D9Q3rGG5uLh
TOEXnoZBGjIUIZEbOVQqo1hkWd0Z/GjGfWFvlvIqNTN933Pkq+QiOPiuxpBTY/FPM2CE1BVNKPm3
zKcCXzcXn+Ra9DA7aI31KpLZ/P8o7TVP+mdir8WfiHrir9XHP4x2Jf2W71791ydyqAn8f462MOql
0Yseqya3+8tK2jNjX5lbLvl/Pp02asqr27ANedfTD1ihrURfa1Iju0d+rV9EOXBpYuXz1trRAE/e
AdxiUXe0SKJJo1oDPFZYu9ttmfadbWYdDtWqbEP4Chni7kngtRaexIqIKWWP/opeR3nmKUoxp6d7
3K8b74zo7GF0s6zdlJwxPc1AGxkE4mbM6JGSHKwgrcoTFWI6VOH9NEpeiKwYH72v3lMPKmpugmUd
scu9m2d81h6UUgFoRnhpM/2iwTNIVjP90oJ1l8iwSDdydVP5kLxX5nhsFmrhfcYcfgmzyJj+aOrV
2foVbtZZNkZBw1B9fbWKfMNPChtQ2mQX8FacYn0rCNbVfMOPDJMTq8rPPBhRn0P1Td4xhIPkcLpd
ozj9xIEBQPCFzSLqUAjp/PVdb5zLN8AXehe9BLL0i4ZQNdIuXzFe8uiHzt63zgvuaiSNZB5x/Hqj
HhfkfQRLoJDk2HLtMXJppzT+qJ66SqrFUBwNi66mq4mHIZic9iHSTjKPC0XvkeMPgTxL7Jw93TCA
eWqJ1vLkOvcuAQytQaIN/40c98hOv7iVJUSfGpMCA9uuJ2HJwVSsOpJ28Mzftksc+6muYiKTSIpY
KGeTKDeTaARV/y+ohdkcAMy3phqOaBG2WmhsEe19WtRgChdLyJM951LMZxH4hosoPftN+rR9SnFS
U3NmYQqr9bp6pc/bCqUUlA6fRIXsZOXhYSszDlT8v3lQuzYzxrRReZHT694QTLrKz4oQlDs9M44H
SW95LJ6MKyI3ErjmYCS/euri/xR0AN3mdxglj0Z2AI4eIJhCWq3BXf47QyDOOU+kY5enTtenSps3
At8IdYq+hWnlIuqksJhhNg9e+AbOBxffnyWseelfv8RuSdK60QoWZPPZoLPTaPBXPT2WnVSek8bY
QQ51nPgSptMU0zaLAQQoX+3DyjvToiUcS52/Rkja7WR64aU+QDUPGWYJPeWcyXjRyloeuhChueP/
31Aq8N+Xg02MZW4ywVbwgZTpoeR34XRU5TEl0M9N5CSBG+g2mT97r+Db6ScxLoKjit11/xH+wNdy
SCoBsRYJPk2zcgeeP6ipVYoL2vYk0D6fPcHc/V2cdvpGsp/sF6Rrshid3J8TGn37llqSBO+T9q1r
P8RXE0ird3YkOhPDRacqjkMNbnOs97Jek9134wcGhTjUDMW6cYZRQtnX/1eXmo2Ih5ah+HZ+OyUM
UiRYOb1n7VgeQU9C1CLreaXEacWVIg9JZInVsEBDauWIwEmgMb+IpWGtQgtG2FL6F9Enwo9CTwxi
gpBp63K0emHXOE4qTpMP1O5SXR9G7MUq/+1f5Cw+DvqmP3j+DRycR4HVJ844e2Vs6gQH7Kp5JrFa
Pb/5FvhCMljRE7p2bUv0bqGEBAsGZ0qzrVEqGeXyoUeyMqLSzfg2jyQxW8q5oX+pTBZTXH41L3cA
yxXP9hcWhmNTVfr1NTR//nrFmJx7oga6y1iJSf0ObBuFODTI3+nHF7ZXP6BrxPmtE65JPWke+iSs
wUNMVTPXNSBYvj3c/K9L4pLdnhuHeZvBSTV6AvIiKhGcMv038CL+/W2YYMTMNfuDoTvR/xmwbh8j
0c42PKv4W516iZCXeN2S8UXqaDnZ63aMltmTx45VY9zo6Bmx/juhSj8/zFOJUoBcUeEDD9YzcIab
Q3rYIpUuPTAIr8sd+3AV2AruJ3aavhfAxc2cDLSiKC9ZrS9FW5BEi9zbHkQPJT247KVI6CLfRp6V
6ssxCoA87NDw4q5vhF0/GXU1IzsQ/rwldZfP6ZJubsM3NVUxHv44ap+clFx0hkEGpPIqeDK4hGqS
W1CqT+8hRLRfUKPlWBnc/0TVXknQDr11N1d6oIzkh6I+c4Jxqtxc1rjtdSjxG0QUhdnJPR5MHFiP
4dwAoKLd7OkZAn1WnTN5A+6dplZttdLpHTdWvagtvVkVSNTMLWxzyKXITHNbubzRiPzyWidjro+P
0sKPG4S8ewyvCnzCUKj0z7cUBF78boLkRkXyctqCmZDp0m2BKFJrgJ3iiYXt1vd4tc4Ijyqxw2db
D7kqtHmYmb3cpT3l09yn8xpytYL2ivEDHdL/xIWCgq8ViH30sViXJwJcobVdnjqYG1ANoG6EGlRV
Apbi+oVCwe+/ciZLpra3lEpw7sgI6luPwS9iNMWIeQ9qQi30pItqo4ZcTfrIFN+hJvuOwJRPNr7B
HXO1dKV0+mUjnlCaNCmoxHJnu/tMzrVDlIL3YuenSwnO02okO9y8q+7PCERlWVsLgnXxiHxQUuvX
kIn8r2zjOZyET8mfg/JlP87j1RXSYE1HNrrTOna3SbsEJHWdYfKrNHBp4diMxCG++wdZkaj1otKU
FcxBqJNZiZ3tV0nOv3ren4W8NyDmh09+3Co/bilNHS+6NPPS25Z/qe+/5em/mRY+X54cBJkYJi6O
bnJJb569VuXxTE2QBl3rpsJ88v9ABQkOA70wgIQe3vH/0EO/Ey2HW6vwESlTVUvBGrthZFcLe0YU
vG+v8zPaLxq38IFjja9yS06qRNeL1YXBqBlEqGpLe/VMoUFmKXHOKUyLWLOWL3PgLj1LV1wLC1Sh
l68/wE95787BPEj1tpnQVD4o5aYws9RePGLpChh5ugi7YgNwd5FAn1HND34GJV0ryb+Glk/26Hyo
PR5nNEf4BlpImur805Ph41euuaCaRyco2vDhOeEXDbQdlZIHMrRnKYxeFbgHnZMjvaUxr9EBgX5W
UBvQalTFGWvMinBKxi7Vnkisez2hUw+Fi2P5n4TVvYOCn0Ec8YWPHf26dnN0SXYHNUc3x/wZA59r
ypVJLe6gIqDYfc4pwiXKmngWY6Ruvctya1pM1LfSbRKchQ6LZ+s8++RwCwOxhcGmBhl2g3SrTV+i
WocIwHFm/tG5ipEb8YThBd90t6zSX/zMrbyaYBflAml/ocve+vT2TXtj+yxReiMrX75xrpuI+teC
BTQVqAw+yzQ+FNab+oU14d/yDdNEJEPsyZ/c+KWxh0BZ+xlVLoMLp+gKoBYru25lNKLPjRNrrIp6
DSFjPP3ONBJ/GQZcMcxP0vH6li22viUAuP4uEhDPRc909412hntwjmxAZ0ngRuT7zV2r5ORalt18
7/8NB+TV2JKi/AzsCT7Kz44v8hW23y9SSmbexKS0+ZFul1OaERYq9ysA0xgCv92iRqswTBgm4WS3
NFmeWpfUH3HX07uPGXunqlDoKeHsJ5DtiAOJjvsVFGlDMMIZ+YchvmF9bk9lj9+fExZV3Fvqn1aB
+KoGhir2+l3AqjTA/9P84oUzmwxQN9sKfMZ5RpefS9xHuRD+8ZiQGfJIvXcat4SLyuznqmagex6i
RGI/srNZYj/VzMJ2V71BffKZYVCgPn1wXmFD20ecgzfi9TGuPoS598tJCz0fP7jpy+HxspbMcXnk
nzTW/EgOz8snVC21BOyMtBqayqOYfzNgkk80U8YKE1PlOhSUzQ3ph7Ad6ZOvmou0iBvqemx0gQWp
sEXHNaGEKaG2DVWqhYo977+ZTkU3xdIB3/Q4gZ37WLDEd8vt9vLUlthW9RZZTjrXDMGFV7jA+yWf
qi7n5WV7DVGTAI5Z5GmuP6WUblQ8Y9wcImDNOjaLZFe1TGdSdlJjXc3Ut2EFVYR9b1p6hjKCdtcl
1YB5BxscYg7zL33UZS0LB/wdpc4u/eAGf37UrVkL5WhmSnyRsn0pzLDKbwtAyff/uDl9bs63JSkS
eT3eel7ttx8G+7JWjwnL61+Fw9Es1t5fpWKFDghTatE7qMc7b+lNgKzQIewWyH7Hqt1qxqdzRl6+
ir0N9HA8JC4sGkDVjYgDjzT1FI+JVyxglIBLXHDwiyeH6e8PfA+BSMpvLSBZNOIT97a/Mjo7S4Nl
l0HrkeZVlRrw0LUAx+3UtfNsKh62AEay5x3ftCqL/xCZXpXQBatn+ZvtNKtIxvlFRxZZdCidZFyE
IUtS0CPj6hVnWC1ckz+DzQJB/VOcA3d+X8X0mpHsf5DTVQo72Qgn2EeGxSpF5meKuS7m89WBXAAh
YXtPTi8QGOkvtXikh+SfqdRs7jszOctDLpWRJHhT0o0PFCUPLnKljQ0j4iTTuU9XCFUMuWRk11ts
fmFlaTQHXXdFGsQPpvHiFWRpB/QXpz9CIQxeNaMKnwoZ+lcUuhiZ9/iA43O/4FIJJkQnx8fV65lh
OjiXnUWf71+TIBnhtbM7YZMSHEh9UlAGATZ0FUldnLxmx5OBUjNZcp2ZOfBvUzxlfD3HlxmcOevg
c0tOGJEVhjp/dPZpbCY8jI66nkM+bMsIvV7fHFhxB/YqpwpEE9fD/jfpMIk8mX1X/zeTnb+ictVe
OQz9Qhgzpp3KbrV6POU1PvOMw2caUD7rnJcgpRdOYnpTX2mH7QPOZ4iQSotTBbIWPSIdD/IW7z0Z
V7H9mB8Ii2Op3z5htTXMOCaQosqyoc+UKOy+4MQ1S0tTQ/oY/sVRx9sutuwM6zzB5hh9ByrTcFSE
B/ffqtJZk4W9cqVSVhSXZ+FL3vIw9IFjLmIBI0C1qDKpoOUz+PXOWqmLRxdchUPJSx964seGjOim
pg051MCTFbCRkWidYGpquLjrX32edJkl1r8W2sKs/aRdnJ09eCdrYFWNTZeOU2/UY1YBt/Qy5gLl
R8/vE3xifOUUYezwf38CjEnE0MlaGeHD3S7Czz1ionlSGJTAt/UjVttkU4uX1/gHGXeusNe6vOsk
ivdR2k1qdoVryAG4i58OYxfNvPTcW9HJ/ivI19s8SPBhBf/A+zIllxpqNNN1lhmXFpNZrvcm/fnP
97TW20leDtEN5ucTXRQdOxJrRXftNxQGeO/Oy221h/KGsqn/dJgkSd1tKIEYKTYfqh2OInXrbCWg
8/dLDbULF5EKq51DgUdzofOamvlM/du0EZpJNG9l0jiHWvoA/o3U9S4XAbkbikY42DSvbHjgSNXM
9TjHBGCnWWwPUNoI4Zxe5nG1v2+geRp7F36I+czZvLnL9GoW9ZN7yro0S1v3fpxwKVL2r+Bn3JOj
YIexnM16F0Auqs6O8gsXtO0j4WB4/7dnNtSJs/ThRL3D6UndkybxOsJo+a2PFxCUv7RoOd7O/8xP
SZx0GVV97UmtLVDRllgPb3gU0qKQtG43L/EUeNAk5g5IHVlIKCqxtk2FnfVAaWspVQ3VAmZHxplz
AdUkib6weaSN5cLMEGXMNY/8qBD5cMmYdtUaM8JZAz1GcgoW/AkbGGTrXx1mDYp+HlstniRBJyrE
JbYixNILflEgF+5yBP7p/AQqEFHlXjGThOBmvrE6X8nJDCgUW7EGNz0UOQR8OCIAtMqf7l3H6x49
WSJ/rPwcmVtWVg6Ucb7caYWt1bmYNYTB406xqFguRq99cGOxhljiEztf6WeIOT1+pn4oVTYcab6U
IQtXJZVfV+QX+/kFscPliY8DLoRPLSoMXy1i05j0DJWRh1kjzJF7eDVfvSu66bw2cUQ18I7DwnTZ
N6cAdrQqtE3/o5Czg0rQ2ie3G0SxY713Ff1mfLANsEz+KdHC8fmRzKcRVP18MY/2+Y9qLmsxt46J
+yk8dF+hDrWDKEGHMRKguOVCPit5SnfVYwgUYL9do4uIxejBNzp0dPHWfaNs5XAs+g67i/nZIavk
f3I8UedmwM2MTfndfe5OPommwFlIcDoHSGbz6R7uA9DL1WX7Yr7w3Wx9uTmgEZzy6jcigKbw86VN
V9TRDCtTYM1C7tDGCpaYVULb5EFMec8yg4d88kUrf4MjRStDWGuQHnW4lTYItvTx93prjO6lA5Gh
igSM4VP3iSFjWEpI6kx1tjTrZZ5M1jWzyzI4hU18bB7N0i7NiHD1yOmLebwXS+yUXG0J6clgLcio
SNYU8OKhaIZM5YkCbomg2E3O4LhQ86nVGKz0WwuTF5Xrb4/eGU4ieuARNgs+xOQhXV5jNx1Y26G4
6twXod6e/FKRC+mHW9M6dpO8N2V/nCU3jzapXgua85tfht+kmbbUqUSkExX8AUHvoYr0pUnILNEL
8iIClBWK5RkXG+3RoDKKkjPmCzl1H+Vmy9QXGI3jwwnhLeU4wN1Qasea8Jf52a0I+zw8Yc7HHYQM
DXunoIXc0wRZeezbjljE9lzJDcquZokrLj6Pg9kwl7l7Nmp2ylQ/TAe4uTXg5s2/OAM/AxzpYC/E
asjL0hMsSrWzPC7MBpM6dD9Cmkuwau4cf4c/8465U2tk2gWuCVYsFpi38qync+BAvHE4bfo+klPz
BGR6C5tD0sLlmKWPcwxk6/+Hjh9+7MVbZD1hhmkoPEMh440VdL5UaIJn/u/lVM6zrPgJdxnLqLmc
MsFpy9l1LxE/JDJDscDmpA0DGLrq07Rbq5etsQWnNFPeofpJrBsc078vl2Vy4s+uLMNv5/N6jHGw
JlYRcjzQ1JdyI+v+It6XICy50T/osjK3gPw8Sw12M1QKuu0S9/BAWP0mFovCJV4xW/LKK75W7ytg
HrgKV/IeJrRtFtQGAkkIg+oVM60iBOZrsO6q4Rfr4yvPSzU7Xu1K1SkuU2CZAxobijLbjGMNFOo7
LSd5jVJ5aJjm/8hUK+aTz0DEOcm4pZJ1quK4QugAt86a+ghVxPvG7iRbqcCZXbdUlpsjQfvdOb0k
/yrsLCHUh09MvdpNXrgsSjWGC7/K3RPxlaj0zBmgZGR1vYsXf3itFwA+XLwGFI0wbete+bmjmEFH
DTRmNAkufSDdKAFn4ptidnCKpzR/lgk942qvh4jZKSqwt5EduN7k8UOcI6U/6HR7aO7pcSuKcogg
jJhVIKXsk2rBdbd979MSKnSrYLopfxN+ydlpBEBP2gKRB+kYpumboNxNtVtR1gXxkGEQx1quBbwt
gGkn2wFe3vjwl29UUr05wRvA8u0tM2tsX/aCXGOpOfGdHZ22Zx2Xv7uenKUqxmoCtu+wmjDQiQhy
rjG2wtDmhGusDwrG0aLBIEL2j7Id363QVcAPl8FnQHID+wKHWVHbwaNoO9czLp55JcG1YUV0QC+Q
YrYyGIV/uSqBxuwtbXET4bOtid3yfiTJV2J39OSeCMIzx3QIQw7JSFuCSM5mD3wCydt8EzvpXK4L
iQ9QE6hRJARniMDCRmV3UHCh6C3CQ4yNqrfOVHNmMuVxgPdrXbn1f3IZo7V8YuHDWioDWccrEntN
XNvT21hB+1k2HGSDn5KVpskPIh0Ps7z54nrmz1VnvqF554s+N7lWWpDbRm2D6/IVMbloqvNiF58t
oKlmGmSlGSVj/ErLwgpRIYgFfamtF9ENvzWBdwerLqJctvjwoWg8xz1nsLM4LdiRQY1aRQe8fc50
v13m20fRjmrgHP0ms3L4vgsuzRO9m3aBXtfs8+fQrE/FpMJmYGB+CtjL+kRw4lmVBbq8IDDwri0Q
hDuFwfOZCgC6p2yGBTCKuyhJvKDd6UyN5MTxT7cv7KFxDrIaQOlesoCYpNEA25fD/xElcHZyktdF
KGgoVm1VF82k4fV0aO7Ufi8lMqJWbtgubaMMwpWCSDhU4r4bbkiJGW5BvIQL0bX9ymnmVaqC70zv
EdYVea/Zm7LKzbR/EHGskUi+sl4Zj4tDW5mJNJZ4MguJqAmV69ok5ci8+KYK1i21mukp3I1bEHdy
DWgsqDuSRDRejyif0iZNJZLmZJlFD14VtbYGurDD2cc3gm7tCuA/bHVDckxrcXPrr4r4wYhlRjL9
0rsuoSsTCUTkS/TDQGhFVYji7xjpaUOcia1U5c+17Fr/FckyPPYJRdxj12B18Pwe9pYyC8kpH56j
rIa1C08aC0UMtZscPrKBdCSiFlEqFArFV9vqTutWeofYxf6WK0mymtCYctN3qKyMDQ3KgcfsyeSR
FUGljMeef/3VIHOh8N0Z7qQ8ByLI/kZuIflXZKnTPMCtgAcZFYGAOLdGslTgNpMYbAmTvaUSNXNb
QwA2NnHG0ezZEK+c4Dm0BH68BXUbD7kgfV3Hu+tSCo0BKzk1DJ7C8BioG4MizjG1TOSBpRCIEsZ/
TiFk8Svw7f4B6TOKsmROBn1mmUfVZBvfn7vxtKVhj+OIlXcyi9l0lH8zL4syRxDgQzYcwHqrwnmC
lAillhzIaQ3H++LZIiO0Os3kS+pHYzreE85FONf4YQA4G3mbnVQGcHNgcCfMFtkILaM35+8ZLwZ5
ZGSkUM8brpbBaqK/gc3xrzAaUIHUifC5eWCAt1Upyh0Op5wYbHyRhyIBTaQiF84HQh86YwjGx92W
CxgNuPLgFM3hDu9FJWM+KXHN18v8KoiSARnMGTf37EB6H+Ty++4zxkBXlAB9+67UGJCa0FffRriK
vfFzjn7MF5TV33wDMZOV3rSKSXd+XqwIGVr0nta3QERRI49Kkcn5kf1KOpuO5UBD6p3H//mv6HPX
mKex040vPsLhJgR+dwQws7rwU+pRr8VLJHW0eQ6NSApP7VSPOiWGECl1m/N14HYZOM8HKxDqN3b4
vdqnPGLk7XrSY+BKxw9Y7Ux6okoRcXIVSHZA6NCqlYkXGQyzr1hrvh118IZds9IFwpVzItgqfu7B
8FgysdUPJjfUu72KlWP6fqUtULxgT4ok8zwPdXXBv59iiT+WLQYQV5xXkm+BXx0K0gNgMcsIZ2ar
UUIaNl0aL5xdN2eNZ+08FuUWAQaPdnAkHybEPpkKNz5PgTUDspkdxAtBdEW8jPROBcHWKWJCFB5A
CpmpZhdB35XwYwZW2KWn6GSjcado1yyrlB+Uz/w4yLJROMvUNNzMf1tJP4Go7y0oKp8lMQNVahlt
vjtXDmGNRnYKUcxWsIJ8kyVja+VXq5rdVS2p84+4oZn3LWqavUzSqpkeG7FTvFszm029nqUuKhcv
Xa29/o3m7rA22Gvf3D6M3FbzFClb7LY9goaRAgKjnAg0/3/T611pZO8lm7uCcrYMxF2tSYjREvGW
X+aJJJYUNKd9Go20cDgkXb23Pd/p+Js5xt4J4NAh+qRAAInqxBmuHkriR2APn/kEUGujRPdLmpw3
t+gAlZJeWSfpLXuN0zeZe7cIefKnV1wKt6V1MRv1QyJZZHjE+Xi5C/5YnxhPUveesPDcfvlcFfqQ
FPPCawAOxUpN2ILxhj9s0iuC/lb8/QwAIDBftFbridqyJ4RLGnZZsMo4mtFhLnFu4sS6k2pZg6Py
a/3JqYpclskGGRXFWjf4uCKDoZoy82EVmUzPCRiiqSVWHVjLM3/CSJr1qOMNTIwQZlusNPXgczTG
vXl60RkfpeggajEh0miQ7jojknJRKkqO4k/DXV1SqSnrUd6WeCxgFlSGDyPGeNOK8MINiMOkDVFk
R3/p3jBwI3dk4lvuW367z6faxdlxbrX0XkAzQxZsbvtV8v8UxeoKlnvbTu97EPOtpLMRxN5UddR6
mMUYfR2D3JVWZg3c+7FBJ31iUTYltP6oeMC+EOJNc3r5q5FL9pYj6eSt1S7QGFJYOCH3/pLebODp
WStKhb7rSv+CJkVJNmJWiOtWrDSxuoPfHJ5ywTF54ds9J8j8lqzCI3hv3XPog6iZZODxDec4ZXzd
sa6iDcHW7i8wpluWoquxJ8lPBsBpNFqqRvudi5y+JFWpAaFOr6UGQfwxSbuecE+ahyAL/hN1Rr5c
3yl7d+MLoi+xpWq7trrkRTJnYgGBuWf+2+9gVIW6RYNoFnjO2SijhOwXVtZSXEZaWKhQm8NRg2un
vYimFhCzFO7h9PvNlGSVv+/w8Dvy2rvtgKfDWI0zX+clRJtrZLF3u1tP+2Hd5V7BRGBaodLxqSBY
V7KgK7T/K3Lt5bqSKGIo4nueptpuKWDTHfvWUedDDcRn6Sx3ZeKkpSAEwQ9gM9Zs02TCHVep9OYD
pJh65V6p07iswAFsAAwIy23uJnEtQlE1zIrcbInKzU67ff8FfGW434Ix0jYbvp1U7JUTIYC9vnB2
HUsmIRJrAr5ILBxjZkVS+Ps7b7PY4HgxsL2EqouuBOUGospFyA6+M5CRX2kjc7LA9hNikfaVLm1H
eZUz7U4HfvwJVKzMBSiEGmUTguoWWlRR5GkKT4xkZb3hBB65EjUfZh5TsV0iiFK/j3KInb2PSkEs
t0Jq7OHPeBui3dL6GeJKOy6zvWdkNjpZKYf9GjtMSmlGecTKI5+l/8KplXxuGkuk2HbU3KeIJ6KU
b6rS+7vyB+3tNa9JDU8JGKD4Qt/+w4VIFOQvog/wFcXC0xOrq7Hya95niOYF6FD2oCweT7k/yAHv
V9qkt+CP98Xf+Ro4Z8Qdlx7WFqgUw7XZIVCWlDH0vS64e9J9IaOLFnQwBN+nLSbOXYkyu0Znfsxi
qtjDLpWOufqsRMaEbA2JCtJgEysw40fOobomUWUzqDQ/9G8hYJUa2p+APEV9Hjko0CdVTyv9VgM1
0x/ZrHWuBtg5gdhsfG9tByKCwcVMYnDMoNhNN3Lgf2qIviBbY0MUol5pAQ6VmxZJfDdLNr0OtsnD
PaXGV9hNddiEB6DvOPO28fgceyFGXUoStKx0Iz1CuF3qiT5xV3VFwKPLQ0F+ppg1i56PBqBkAh9T
W+io6tEM+aQZQZxODblHBBYrW9Uq6k88O9NcReAdEj7UhKH5Qt1F9fw48+K/BdB2x4bRYG4jUOO2
mSkwsonvua2FLbTy8VRshzl+Thq5dsdtEhLti3sLoIYM59flg17QiXBmA8JQT5J5WMfS8x33CYfY
2KqmFgI2j9OJLm1Bbavk5yvu7Wk50wsU9OIeAkdAs/UB5MK3fh4FkxbvvnS55sPduVUzgBbdtIN2
9ptmZVlDRjQvifaZboRozBAfPHif/u85jCYiUpq+cOLCyUAvsGtktILm48Y/TghvQ2WMlgR7znu9
iZX+Tyvtru7a/3+GNI8T39Okxfdoq4J2pihj3ntBZu19b5W0L+L837LLjfUZRyQVADJK2LZ1VGx9
DtjbSJWjKTw2GkgVMGDljgZlq2bb/jigOMUIllQF3KoPCozxbba5uAs+GmpKFJyUrfjlnhL3jEW7
TbaHL14/0M/GGST0wuXio0FQaxV0XVNreYvwpvVOaIJeWK2YWvFMl4uKqp869ZDZRnFeqH8YEWgm
JCYDLXlb5J+4SWNSXmmWHlzninFzTRi2qqhNt3FVoaV6arIADXugSioZIFnTx6uszoRcfTVc9LZi
i1YTLMQY2zGs5boh3m6JNmUfuRumdY5a339Zv/TNnztAAQjpwjs+Nt/wD0oSM4MslCPNDXpanD6d
HdlCFBOCzcEUg0KAzPmZGjgkLFCeVU0N4dvkNmakHEb0YuBs+vB4q1Atg1x72gxtGfME0CB24138
5c1Jjv+FA/bjmL0TPqL0qtZPAVh130lF92TJkg0O8JBZHjXr8h44jRJVY/Bt/DvwvFPEk3cKdOPN
7Lx67lWfVb9Owh3iVPi+fT7EZDxZm0jP+h8h6/DWCJs1rxc9Cd0gyrrMll0l4UQg96Za0cQ6g3dc
O9WxgCtNMPeRyHkk0NZhBDpecjrS3NhA0ebBCuj0bPcrVxsQ3Pao2c95TlE8JDezWAqa59UED6i5
vjm10lBn7Sy4qlAXfWfUJv6ANvdWgjOyFkBIcmNHNLPCjC6ZE75CTxinLU2f/e6uA+hyWSj9zLM1
s5RwgmrIKM+JG7IZO0zPUdcGkiDIFX6xCFjPHRCw3+9xV9zyjzZw9jzA7bXzOfGPeZ/4479mdLry
UtiQMDtCS+ey3pSSOw7sRZhiJvEHhgts08bdwmutT6YxeMl4cI6rLaBQNCIjgDaPqJRCtsbR5pj+
NUwy9nJbdGdwFC79FRab1Md3KCKQzVI17a+yIGEukbaZjIy34Yj63dh0Xg/CZ41HzeLAO4qvYhkT
5uTWC0P0G98jZLoL1WWZgv4EAK3xr1Awu8TIZ2c5Jd+j+9reT7AdkYfijJpsKEcuc0OIna6VuWKS
7AbNPYJOvKUVzVsfHJUzMcvHFGs5hMhEezd0iu2WWFYwyx6pXa+c0UpM2HntSEuGuZ7ytfeknsQn
YU7r/+rVF/xlozVFGrA6TDB9bwp+rXfroCL5PSLiBicYGJOKySdhOMbqjJH+b2aj8GzChEWskw06
cYFk2hyKRuAwJQOTErGa26VwZgrsMjV0c0UXr2pceiUohSsUpFyfjGg/IC4ZTlbjalQxLeMHD+mc
fW3V8FviadP9MOxKgXpnHADm3uEfvzl03MkJ1acBPjoTVXPEpVwSh4BSiwsrGtuOoWjmZSL92T0T
jOaNNhp3q66lcSdrfiS1vl470zbsfLt/0Dit0f25hFJgq5hsTQF8OddIZMfL8OlWphu1eFJtEc2t
adS8Zaal7hRkAMKbb/Trb/XoIceHl1O0v6oeu8XqYZ4xkWnigpG/dqSiRyevtXTfnRGEW+G0K/l7
JEiu77CZ0f5YX946tt1GBVbD8KqK8DA2EyAU9LHc9Yykr9P4g9VQe8hhHRx1hIwTUwDTFrBgek1H
a+ZO/s4Iqk04EOTb30JBKVavKbJE3esXmmhk5Dhnfx3PrIFkbvitVH+kkeHx32phBSS6bry/tROz
7Fzsl/bN8JjVf9qWnr2vOfooZ91S7ERAVCCZW5qSmD06rwQHzvrBwP4aXQFbSS/RAkL2WmwH+lgb
UbKoj+YIOxrwNCVFAl8BTPRIJKZlE+h1OPlHKIkHELJ8wncGH/ube3ScBtnapT6GDENITn5zrp9B
T3EOvoAGrd7F3PkyR5RsaDQRt0kMjaBI4QHYquDsDzXhY11I5A4V2zsh/eQGT5PyaLiV99sotG9d
iN9lFvqTczBwRI9hlGiAn4ypQbIdn+EkRV7sVuScTC9ag7ZSHY0esyQgn/63XawrP3aJ1jD7YM6C
Byiy9e0oAkTkpNj+Bn0XJFTFdP0awSsS8z9EKLiZfN32/0AIbJ7s1vI6pUa8lTxvQU8v7Fse7Eyf
SeS0F+wYFj1B0UfAdF9C+yehcOzPJAfBHF3iH0+ir7MG0DBPujObDO08Q52Wdqizi9cm1J0qqe1h
tBtDjGVeREWyLBNfMzlDKQ0ynH3HkGgb4ypXJjdBNMlJV+memJzyNVdyCKwZmERiax5HFtLM2aX3
7DhmwYhOBqNI6bW/ApuolXNDDItEcqekDHaRC7+ve8N/RMALx9hI907Yz4N7H3Bh+sKxNtl9C1g0
SGaeB7eXsgC8eztTKO6UZHYK3xjy9Lu6hcNkzVIRfrPi5sz0xAdDBAixQPg01ESM6H7CWL+xDY4h
f1Dqwejpd7dNR78gk21EEg4J4Unmuo6Agj7kM7RsTz9r1nEvwQXf3NZVTNtE/y8oftDQyZ0y9JIK
tU+HGsdDvxcec2rLClP6Qp43NUXGXXn+qrHvftzxRtYT+z5MGJkXcUe0Eh32ZpyQJ94UswJSu3sR
SZB36M4xrOxkQsPgWF7TyetQXytygl0iKi+7PXfJTOdxGIZGe1I6woVhJrLXxPVepGHAaPQCAC61
B3K6AuaG2Y/LpgW2W+6i6GW450Q7yW4cbpv8vTFWlnj1JIyVDeil0WjhdqwxBUNdObFSIL1lljn9
uvOli3MAgdbKHL+lZC8hXLXG6uGDQmR394Youh4gJTUffWq0Q80IDrg6RDhbcs37qJwOClxbfbdh
6rrG6tiNrA06spWFvcYjfWvKpoAwFHBEKLoXqJTjoVJmEU9Ghba4uRnabsSM8Y9lIwaz5y/UNDaP
AZjLxwMoo/jeua14y9vY3Otsavi1HVWBMMf2Cpxh5g5CJK83znIm6/Ghvr6V88W2hg9Gworo8hrL
nialvhaC69USA9zU+AvBurEkmwY2jebTXzS6vZNXaIWZ7Wy3CI1NBpibgUvhiHT4nPnFNbHnmf8f
/KCjzZnkbs5AJYk+KIn33bJoBXL3kIsX180HK8OaFIHRXVRN3X+aLeIsgL1zN2yR3nMd+UEhrpVH
vAgCGL6dMphiG/wmTKIwnILsJk0Lbq72zuzVIAN8dT0VYN15o82NIvVNeNDDuovaNb0nEGxytDJi
r63W2t/DjPIgmRoMygx9JqIQyxrdwqeBt+9ZkqgLAPSC2UhQ2+yeA4rU1dX5vWxuLDxskL/mqf7d
sBo/HwOVXAtZiibMH7Hyq8LkJxLcGpzfl78nr+csLD375XkEpg6pp/CqtV76Ds7ljdSh5cgi58H7
C6VEXeWmBFFOqXTGbi7ApKKJ5Vdraf8JEMUSgO49B1PkAn79QN+IyanGR5nT6lRuEIRdiFHwrQnm
pVmAtQj2ec8tj5cc5qDvB/RqSXT2tGxxcoHS5MgU6d61TzK/06TnVysNoO5NjzP1AsylZ+eXl56c
7A+irfOFyvBKGb8Ax+nLJasr+cABO1mGOKt4f3a3YeM9SZkN8O+E1ZtFcVSUMdqZ88l8H8FS2s79
+FJ4YOtdmb77mNPQT6PAZaXg+O4Fh0RKpYBr0GBJf0vZxd8g6XCJoV357A5awwVAEV/DvYqZueTQ
8ii1plGTZ9FZzyJEy/oYNafo0Jv8mpHSA4jc+nyUYBUT1QkeGPTyJQAkMRt5NYmojR1jIaH1m7qp
16NctF8jVlEyYVPCVeIyI3SAyzesC8mtnNbw5iy2bFuV5S50/B6S0vodPD9uCWJBd0pYUYwRKtPJ
dv96PwzixKvtsitfQ9kdtdM1mlzKeXL9zkEehTPM4eCXpVtCiyR9Yd1Cw6043KQpzfT6qpr3/Y2g
uiRcJD0COsY2iLhNmz3IINHZGeaMcoT3v3/vcg3BWSVByH3zMxH3BJ4E0CmddyjBYJuMH3vTmrQW
y2B8yOcyYcQbd1jC4fCREDllgMxhMLaVcd2SdnSkupyAGkkgL7ANTRno9PGNLLcx3FhgkJXrY9kR
nf3WXnuZySWjFNydHt7Bs+HTjLTnUH3O4nDJDlBAxGTFpuDrkhJsC13WM+DIslGy9dwctLEAKiuz
AZxgL1Qxjgp0nCk3x3TL0g+k3DaYA5YBDK7BsoddJut12V7i2a2LnpvfFllBg46iO28UFObjRkjB
E7V5twu9Xib+3XFyBJQqiP9fXlnM3aqsPvLFr4VUY51NIEU22s/DelVq+t9ZHEs5iDDniVK5Ez9q
TM95Vk9URfe9EmnEerHbUPoZLz+cKUGXa1xe3x7eggBVV2P1a2flS9ycZkP7lzNqo7gDKGkYR8iF
wwhcXppSAUKwKKMudBsnk6YaSv3jpP+O8RtS2+RZW8i2mdawZW4TgGnudYV1NRsdBqK+W79XNIew
1aqqFGWPIlNTIkek62UjbI9MreK2A0+mGu8g5Mo7HTI52PzpTQaGzXW7YFdfU3uHYeRoD+wYm1Zd
Lr9tFIn3GvgR1XBnvl3P4kEmbc5I2MvhW3kC5dDBvC1l+tID8sn4yh0L7Q1kAAGrLlT22mpmNbAK
8jWlj4ccuuU3o2EptAl8iRI5w14sy4U1/1qKqLOMUHSqIb1kSzzB9NG+1qe9EN8lRxUSAbMXqZQP
sBCj4QDz3HuyhtZdqXSHU6szitIFsbBf9vLLAeZK4hz/XeDgOYe53btAeYVLr3YkQoiQTFfUhDIh
mW3GUD7gIBahEbBc0usJIc+HiauEWukhBbNCXN7njqGD/lmM+NH5IvKiG/ZqcA/TURBfk6g7BDEn
UHSmTOxdGgQ0HgOqgK3CWxtDilPCZoFeWrHfijGeXQwsSvEELOS/1Gee3PNAJv0JZIiTguDnHcYI
BmsEc4et35K4y4gHHy3jiS42B96LTeccF+V2zz/X6dYSPv0mpmLGmyPxiiG6frBEiWw+m6VgXfTH
cjDWJr/CqCRfGBzJjO5hsJJM65+0hn6mNvsZGzARlz+52vbZF4vW6bwnbEVh4wd43FkgxaToNDNr
4eb1SoYho9LfOVANH3DrzwxZJA+AIS8XmQD3BToDi5DPaCJlfY8ZVpGbPBjY7+L84br2qI39BkRz
0YQu6ejJ+2EIJxIg23P7OX7xwZwLOvpYV1EbCA3OlA3npiVvoJLKbOTZU0HgQnPDvZT9cSlfTQPt
1/1yWY06twjlVpR9/9gJe1RVbuIM3z0gO6FZcW7RM8bCFvSUMZ5YPE4f4B+hu93w0EtFUZ5TEyMG
dnYyVE83ObU2ZiL03D+uyEoTDI7sm7QZXCmheasVlrxS455ZT1KrAeXd7D4VpcDHe0NQNBagsrI8
yn5Y553uYEgFqqXEimrcJDnYrYepxUrdacHet/OrDVPIrvcXKvog5PgzBHNjME2v3GAExlgaCi7a
Q8/acDD/TpoiaZNt5zI5pJWYaBIdxTLevNp9T2NFzVr3ays/F63DnRtrcF7wAW4os418lKklpfXc
dFln7dkAuZ0NnrMexEwyRqlbtEXCSsPXjCsmYC6SNXUcUKicw5IIS680KQYGvgijlIpzvi6wO0+s
YAM27ALPMuv50vgObG+DEqR34ET8KXroJXVZleSZJFCn4HOSw/GeMOPmi3gWCNPA5OMzD1WvvmHE
HGPFY4Nn7l7DbwVv6/LccJtX9XL/iUQt5pp0OOs6DjLNiFbZkW4s2KRtqw2espKQsNGxkGL5wkxP
3orP1ZmxI/y0rPvWGXtT1sxHfNRfZuxt3Sww2YzfqnrVFLT+9HlPgqDUsJNpXhU+gIta2YKysVUA
V2gSHwnE3elmGbIkJuEyJEh8od5sQdV9yVIKbgibsb7G9UbRgNyczWhmvAzJiYG6TTEGL9bffPfA
zh0qC3fMmh285PVYUw2QRgZql9O1zDpysmXZX1VXMLJqMCDgLNbai3tO9dxvhVrSIMwVqoXCDxMR
GllO2+ydqy7wxNcSdrjICZVMxGgoBYKyuMl/rn8ne8kg15w2weViz4Z6ylEzYGfW5tvfq8DcM7n8
eZH25s84lZUe4vn1D0Qx7PZQxApFb9jYTnMzeXLLs5KIoLjZ2mUI2ra3acYPjOYQgSbKxEvzHbgz
Y49Et68AHu5qDXoiWy2KGHmEAImbwHtLrC9MT5oZ+HtAa8W6qKhVkfGJB7xYNbTdxo/XDlLpWGNS
BYSYauAOXZvxfouCqHoJf7UYQXmBb2cXEL9ZAcVh4oJ0GNsWLd4nEyIwb/hWyqfarCCwl4cuNH8B
Cg+TjhEKu5AOt8jelLm8dNc7I1z104mum9ZOn7knOzo+o6b6HVV3LKHYR5igPYI7Mp7VrOtuThZG
jBS7XaIn9oO1pdDk0mauSDlIzr/e+bRDv71hCNBYWr1UJFRk9ADhldbIjas/G1qQXCmeFVWYc4E3
twu2kNLl2YbNUzxkRaq4eS7y25ZmluVglErMFkQxUs+1WY/el3gMAstgC/t2dvMoHZ9Jatno4wdc
/xntDJzjckJFsomTgFQBSvJ4RPz1P3G5kaq5OcZD97d5tmVEe6I0Rp2GB6wjyfTj7rmVLO5e828+
VJjnSst/lb5wBMuswfV1I0p9ejDY45TkkLIET9lN49CGrEP6lr+fZ2QSqHQEVL8zvXMYdvx8AgHb
rKaqmB3tl2Q1KhpZvMv8PJHAz8NsmJqfDuQ35EiorrsJ3d0TrCapRIHur0R7aKZ8/ifiOx3kHCjl
90sHSemwVz9VKcAXWffuKTOtKeBzMS8r1hvvUOs5+AH+j8co8IRpSmMb8sIUD4rbPovjWsD2Ndf9
wyos97LHFYVUaqcC/wz/sVyk2rkQtFC7Aj/Tf0GuC7TViQeJQrwS368ALAvNeqgS924H11FtjVuh
JAizSBawiHk8DJYa0ySiL+/eftAECApDn85U9nOvHWIkrpNN3/qNTEeKXDnbP1WhQqptuKnMD58+
oK10+l5XlhyqAX5ILyaS0Y/DZ8RYTkYSh3Q3E+2NF78Xsh7NBrhqvstZGoKuzJO2swJ+v99ycONg
V92fXFl3Z0XbylG5Dm8E81JvYmGdXkDiVB0ZzQ/Qz5NWuVFIdMfZ81rz53HLhric/8HmSbEp01ii
7vBJNv2cdZOJ7c6e+7idUDsAdQrPzYKUv3aP5aDTVp3K3PAznSOSszcmg9sgWftWiKLHe+sOYP53
mbvOXe1RZn7FRWz81PduyhB9cE1v9R+mM6pHVU2Gq/sB/ZIwTQVQ8W1HBGjDoQSKv/FnUlOeui01
sPdkmsx4qv4vbEfSWgtOOvs6yGtCERaQQvIi0oNlTOlAqSE28LpiOI3knYPrQCol3S3EIqA5XHqh
S6ckg8Fho82X3Ny7+Q7dBrEmC1PDFcSQz1TnfjCUGU21Uea92r/v082Nkg1QKkhsE6NSt8vWT1yg
2F2N8L2FxIOp2xI1868A7k5JGkfcb1hJQUCJyOfOYrHuIjz3xB8CiPQ4MGVWwHSJqM/16ZZcY1ii
R3XCKRiB2MFFF6YOZ6WRpBPcN021A8mi2ugTH4gPlcnX0C+CtiR1Hxl6gOUZgK/5i+eXXwcHrCxW
0besz0EJi3a4erkmCVKi74crbMztM3tdp+fcnEUNiaF+A+0H6foDGhzxMEWasqShkfbt6aI2Z1Mo
zolhbo4naHmNay4U/vYgk3J5/6QmkPwLh9LJvhm0YdK2Y0twA7okoaFV1LPoonA3viQ1GsoRaElt
QR5IkRpKnMLc9hlGSjDZYNLPvyHn1I/b8tj8K6BZuocg+SMi7kE7FQpTqgilPnxdPZwAvMnOan0p
YebTyP5sGX7UZ7sOf1aYsj6di39TdItdrgKnG2ODuMAcKU4btvQvO5NP0Q0n5aqSVv9J6sA+17tD
yQ1rcstBzXnUWP0IWtaQid6fJ3lg4P4+TdYAkCgYsDackRsheINiSZbXbgRviJZ2SuGcFUF4guJL
SXBX3ss4G5ozZSuYOsXoQ6RP4N0oj/8t4K9JE4SahZCFvenjE6Bm3OLIE8ACTJhJ78n2YB3PEY2r
NbwNMOJ/QiWtcjMeBhR0dInxZwAf/QFmMrEe8bnga5WdPIw+akftYY6DeN3hcxVNbiuQlC1WD5uH
H/PTKUsDyYHDVCBibre7J+wyoqI/cStl0nYVw0cEjcQj0XqD92GQpluwp5Kbfr/tQGhIyBtJe+HX
1rBDzDnoaKTiEEDemstoPgPVb2uuyaATXgMXXZE5XxjA7ElnoEUjrhxqZ63ZOJrzvgLotmm2uiH6
pv25B+9rbpS3HiZAxVnZtbol10FLb/BGtwA5yyzgkNQO50s8TKVPUg19B2jq6zf6zD3LD0JBb+Kv
5oolJlKDwiHZpzJOlk8F9YOlyQDfiWvQHrAEKQuYUC6awEnKLbwpRPEe102l8WZJhaot9Q7FLCA+
Ao43R6QdcKLC4l9LQj84Z+hKp88c95l7tfCjqj+pgQctU20ChKn2QK8fGFmXHld6zQsOIFixqKU+
6FfxEwEKFi++qNuXYvQT9/Qpw1j39fK76nXoy9C8RwuZoQsmvMKocw6N71STCWescDG1PE2qWYSi
4YnFA2xHQlcLheUWa26S1SNlbCZ0VCbS0PAdFbI6w3jhCUJPpX99UhL4zcOyaceetBPShMj4/ApA
fFt7kecClMc+ZBWrpnNLvrf02CqFS1HdhWdHYuziM5ZQqgA6ymNd82/NiBx1xH9HFTSkfZwUdZUm
RJNbYGLRrjONoEHVslNmuKimZqUGwe32LsdLJtOR6FjxXsBlGmZWbR5PcCy90VXt92OZP/Bmpk21
/MOdq+UDMfdRNAB1FjL/EHJfRxFGBF0xHXQ9f0bzjO+i6zsGW7Uq3jRBNA/CBYeyXIQ3BZl76YqK
O1bPKfD+eC420zCJ4X9HVDa1az6wX5MY5wWq/ll26aftVUglfv8tyAcXk6qlNhnA3/ss4uhddLpq
RYYHxc+NAy8BBHkVqpveho1ngovxVcJJzEDhxaMYjrq13ynbEXe6qiKgBmRwf7LUHRaXVA3ogL/Z
4I+RYx05u8BoSkR7pa3dzGVB7UVhTWTnt3hVmWIPgn78zgobLk8VnAt0eJepKToZLhszqus/TN5k
MAYRcXz5d3ZIJoTBNgj0nkawTcYl5oOODuP0dFCyST4H2eLmd3Rwbk6heFyI0/58hYBQieDLKVPT
5WXznNigJViG5Z/lWVTCxbsPLMbeyep3GRFI3i/mg1OBA0J+BLYsRgGHjw3VVGGTU3bKvECkUbMy
rXTU0eBA+N0sLW+HHceRDPd3nu5vwAoAg41ZGFBVXLmnOAiWuTqmx2svChdiR9F3QnIXYlVC2KZ5
diaL5j9ZnOVqISWQGQt+z976U9d2NFPJsOQJXYW6IIscL0z0RWh/5G220Bus9jFRYikPDq42yYmn
fNBL2qRrxixaajr6u3h91hhWBkrHVikzfbF466R67wGejL2U0n7HkP5gxOcEsp1ELAG49LURl3pd
lNav7jqS4PyeqPYKW8IBjOZO3yo/gMNpLQlxqTqNfj7Sctdb5o8V14zEbx1bFYg8UZHNESdlVpDv
XfYQ2TFUvpdo88l+J5oAh09AVz2WGLq8Qn2NYhwNh/4hCHUcpfu+HEjWOij3nEZA9GM4wVEkyRh8
Ag5ZjrFG3BMmM3rAn1UhSfrL7k+XDmAPltErKfDG5hFNheGdOWPR84uo6oZFSqYHoP+WDIy6kEHa
FvyMy+hflbFkskcLGvHk+MzcqEODMP5LCPeUsYiN8P2ARC4P/bCSD3PFBJRrINM1ZaPVT/2GjBBH
/m9yMB7JI/nlV4JaiFmpu1EsTSMsjzHPsXtwa3wUlgUx9kQha71dnpk/myAErIasKbGNy3zwE3Mp
EfIbWgWRdK5dRPmxwkO9FmLiY8UeownUHiDzU0b8WfuXD2goOdZStxmjrXBHCvV38SMZosAgpF4/
UgiBBSdIVYr4yJzECIPV4vrYgO7uMccj8ywPNHVxKCJ4Et2xV05siLIAHYA7KW2JCeTe6GWiwCel
vEVb94IIa7BAmwQmNz21IcPsOxUyWnqMWl1AdKEDPjGCyhr6ybEJsb0OPMRLhygbDNWJcRE5t4l2
IgSUOoH/yWL5r5UYaHSEAP/rXeKgn25mZmixUUtSNwH5JrSuz4V8Ae5CM9HE+gBHcH/drNrhSHYH
0n51oAvFU4+p6Yn04kPZ8XX59PxzgP/b1vYUH0dO9ScDbmrtsmgQQVsyqm94ofSAbu/j44xoRhqh
GVKyUv1uubWbNg1zPISExQFBPwJ3ct1ATMygPrXPasGioyGZrSa7DOl0/WR6b2vdfDBnwsoF2S70
TdcVe5s5kEusHAcxcoT8PD9pgXENS/2bw/l1Xh2WurrRs/+WBqciUyrFYWpgnzrDXFazG5PGsXue
8Zxn/SZozUlXhTrG1IoFfTIkH1Yw7kmwNML5hSWonWWzx0QN63M3eff5wpNLkH9NhqgQIO3csaPK
V7FPamLcjY0Wvjl6JjF9HC2UnZ4BtWkd5APrmQX+tDmhPpNuae11LeTH4Ss3htJMAgMeaAPkVsPH
KWDTe/QxahxQFPqpt9DySugMQ1FlMydnUOoFYyw6zI+sExFOZGxaO9ewPjjRNyI/F6jlMkl+97sR
zpOeR+mP8M88zg/pJcfbdPrCmdZ0QZcgkASP990a7etDMfNNz4StPfmjCpXDENmj+ZyyIZcnNSIn
bJKl3oYW+BMT8/YISClR2DStUblXAA/kMKsdUdRlI7Zm3A9/qyKzaiMQjAcw/rYS/qUUFxwPZlXp
UL5eiRZoA9uqIYs3pkAcUOjWDTSSKYETkTktSXUz6KyVFx3vpqo0D1KMTlN7afmgnU2i3ScD1tHL
pZXbvmB4Gq4hl1zfEfMbn4CXIMJP95rWiAaotiUTUgPZ+J0eLGiTIQmEtBBpefiWEloPLBDSTaTs
V/pxxFB555fhgjFqxCTS0uuWQEJoBWgpw6vO3VirNBPJj4C1kmw+LWT/Vo5WpD7DILu3AVYFZ69/
7qkPB7BlLZQ9+Nd5YyQNdxbdYsJyce0fgcxaKnYRw8QySK2bFNKAynCn07VLn9IfqU95GMsw6FNr
O6GRTRoRiu6gsEZwrXI7FkO6myHIYxeVFUJoCcUxjsZrGPM02pBuuMaVUnK3d+P5fCyOlnhZeFM+
YHh6ayg2pPDkajC8vLAWrqi6VL+ks2GcQhvXihwGultIkKuOXoxrUl+BdZMxfg9E2On2/igAq7Eq
LQpBnwMWQ+vURg0zfqHEs/wnnTnnIt/7aadouSimkpqXyAhe2EjRAKUq0mO2tc9m2zy4gksCGCzz
AY9z5dhQkknFYIMGtxcpb3Ce8iUJbZW0jj+uYZ9EKDZCblBDlJs+LMIeZy1OlAk1y7F2C9ijN8gm
7hKnEnLmjBAVTumS/Wb10Rg2jqqYCwOZWQX8y8sFOMaIAjhskHqyVGcMj93B/e2KGh7dJaqe82l3
UM5zyNtULK5wTnWda8yVEMQ3oq6OELe/CwP5ChY+nqfccYuPHNF9O4+azQbQyCB6BIFy+nxzSgqX
rx8dNzhBs8einuGDLycriJg+lRBnds+b2QIg8lQXOBqYsvRGj2QzV6LS+hIGoBAWt1KWPYhDvnQP
h6EiioKbq66AU4OO38bC5LUzYggxn/7umNX5nogRvnJIMRIxYljz6yaIcC0NCcenRMVR4Lw2vbhY
/LE8jM4Dq1NpLXZawtNE3E7BZyQpoOl87V2HIVcW4ZRHW41qJ9g5BfjhoFjSTfsvgzQx+r3dHLDP
h8O1LxRSNRIRHJgpjYxzbkVpf/5T7B8G1oXcO7K+CBJIbvNlJSdJXslOztkJiTY8s1cU1VPCzFcu
Lp6G0p7z1Kv7sibIWHN3qvJ8xblMVmLeE2bjq/W6JvuOs5Hnhj4BNPVkjYknOFJwoL8rmuvjjYwU
QQmOKyl6qpjvhJJ+dHfp8Z5DnAj8C25o7Zsfp6nnJpph+oRLXfQHFKMCdpKEhKDkBk+pOrospCHi
o7jaZTXUQKL002wpoJRijyCWCHn/Uzp06PRGrVMpryHE1Jzp9fM0xSSK4gSmgjOx49BsaHwUrHZf
pL/RTZOSr1hxcwwXAVL9p7f4up6kEuUokAhZ9UrbD3zIuvCBiiyUantsQXQ9bKA1aCh//9J5riRK
+/5pHWeBTSlBsPcWcuCJk8KU2gQvu41rDL0b9xPwJOTo9QSqD8qwvc2k8Uwt1uH4hgNqJwSIayTl
okviuVxuegIqQiOAsYF5AZCGyxnQXRCbXClYp+VQq+VLUAhaENQuFgjL7Juu0hZSB39XlV2+ZPqQ
xE4fn4M3mKQYtPTmfp0VWbOiS8qB2exhv0IeUXcB+YTto39Vyg0jM17KzH22pPE3EgqaIn23b8Vd
t1sahvcbd+biMR6FdiIxSwDY7UtF49x8fr357ATyM4XwEwp82YiVO5IzkSGhex6HlJNdBTbKowAo
o6ZkT3s19uF3OMMsqykmx97+OlVZb4pGnLXgt68uiWIkT0jIbz/sxwz46USh7Y1QiyLLMMyBlq1Q
8mtZloPO/PTXiCgxLCm2OqdiIDI4RRt/4NIc36Uz/3q+7I97vs+QO10WCfp9Hau8z389r850qfD+
StpjXbak3aN2rN4Fu9zYHrsHqR12Ag+uRJXY9rQLyXY/6mxcxr3nAQslN66mt4I+lNdKOi/SKzvA
c56pyQ1UPTpgSqlISJBGFuct0ND8eHY9GuRolstpTdNeCM+NepkJzTJaglgIA5rjYb0gnLP5HQPi
R/gXlt415kCQ6n9+LHKAd0X7eEYa21hnGECuDnRDEelbmhBvXajY3CDQZXpqu2+X5LDesOdCo9GI
Lt63ub64SyTmFP/PuPehhH3bhKMWEOpDJ28xQPMD9H2UKnLiDdxxgYwqCboT10fLswO390g8BSn/
D6q4NUik0UIzddENj5P9CbAw2YosSoFdAFf/nvEg4KzXJpiohvVJ9Ei1d8mPd/SXXhI70wfKA1Y7
xZK+hNju2H3XRVHr/Yd6z6zKioMls1R3w7DM3QS0lT08LDC7tWwPCWVujKdD53AGmFZlidqLLnc8
CFGxmn/dF6gVhqGtzCMn0A1IhEojBtUurOVxI+uDnaELsbFizztbtPiYnKfP7vvICWkNYBCTMo1R
w//BnH9Y47QZ+bJHcBqsHliSPdTR82r1EW/sDjt5uSkpjxZKqQLzfMOUE4W4PT9sBrGfDfFfV5L0
INhDXbrmN0skBxHXZXQLTCu5B+97ffkEQw8lvgH9nfFNeVAT7g2SObRLypUSVaLKSwwNK5XsaV4z
zCeNxxHxbLne5w0yyhdfZ1paC3jOPCkq5Ic/IXh47Wmbbr3+iILw+jcMGoMTykBb7taIk7d+T0fZ
dYPy860gr+RCafqW0rGFlL+FgIVuXCgAfmU/0aDt37hBpGl6C9EPeUhGiE4RMrcuKzw5oIxTrx2g
3GDYro6TF7kMHjq4wQ66tlywTcR6BohnulF6YwYAi/w7x0av/poXgm+HPGLoiK387KzqvONiGFJf
op9dE1arcXK28g1mbZj5Qtd1rYaOYFk9bxMqOZIAvrNKl8exiLJbTvcVbuYCd/AmpKkCRrxlb2Y6
jb4D0n9sy0ItOEiQ7Vua+NlBfvD2whThtNRuArw18M9NAVitQiw0yDK5UBv4JSd15v/ShUWxQc5p
E90fdyoEaEezNOjPlYdab0Key6+75InseXf6zzBMcp8Ga410qzl8cAHnkQpj7TZdExnl38voITz0
lZJC2pFhIbftaWFx55bKgyAlnIh5LwFCtuOIBQuwBGbw/HrhWhqb3EwCFtXIArPVae6qNMadKJxA
kKj6ey0sc2OVW3YNW8z5yQvbNwAgTf/WODmOtvovQtxs1mmQcTQS11Phh1HTDdTrB2ySiD7WCsU9
trhcyLE3quUosHGt6wVXFqqM8ae/PG/MFmKKGOMXZtFuttLVzOWK6XitygFxumJYUkkR0xYLV9J0
nw598XguSg5XkYBkn9NkvWPFosPk6kQws0PYwdh5Kz0+RW3/4u3QC6/l6zBfTXNGTYTZEEZmtatH
xO+Qz/Su5ZNcb7ih/mxhieyH/Kx6Vp3SX9pxYFQCO+j/vvOIQv3dgZjEchMmYbzrKdTNeD7loDad
byUhbAtv7UwBNGaA/aHf6S2RjKhW7xghH+w3RoDC1Nzdl8ygYOxP+4X+d6xAbrhW3IeCMm7tHgct
mtwNLBW/5MNrLENNt3a4OhqHNfxiuPFVUs8JSsRfI42sUVHJnJkCZxMCEQQUYXWsu6Wn/39IA7iG
Nj6mXDXlbi91MKALXJbbulG4iDiNk5COR8FbYn+0kUxoyh+bbvs+ZCB/Q/1YCz9tguprRgRIfXNM
9mdFNg2jgJpQA0cS5gqYhKbHVZhQ+zRtcooAmSEFcSTT+rU4N+LMySDYNZHR7yrKTxz+H5EHaS9m
5iBJi7b9R74N9cLAPlx/b4QH11rp6PS4uqlJQo4FyK9fEr3Y5iRYJRL0TFOfCt0caTs0dxC0+fre
czNiDOS2xpL8qwWZrVsNSFf5CqKD1upQRz3lZdhP7UgBuk5oheW/6L29xx4X+2+29XtgiAEu34Z6
7ponKLbaVetX+1n00qQ6ECNKvpJ0pQ1bo1wGmHGnsbt7x+LaztBOTrVw2Hl3gVJrWMqY+OaTjdtS
RH23TssNArZowyK1WGNS+UHoEiSY7BwunI4VJx0iBHEdWVbxSPG5ylR/s6PdadptzWh8H9Gmi9Yk
ezAHZCw87aOhy8R3S0R5OXyeIJw4XZzhTmoPQ3X3I34pmVNTtTCA9y/1dXYLjWPoKqsCB4SIr4cE
7cydvmO6oXQkyCi/svPf5C3AH4pn6EiSHp5AkiVKNOQBU2ThNWlbwnw4SEqnn4SeBqaNKhNJ9oSx
/gQIi/13MiHrI9bJu1jtkqiti5YM4I2KScQ3ah6b2DG+E7p3Zs6PJkvYIzF4p0c4AgYjaRmyKVJp
srSROxCfWbUY9e4+lexrzoPvwQsDPxmjZWMna/iS8TNcC3pVUwnz7LM5W8kB3urwkx9tXIv3rlQT
i/WiYGLI2LTGDjqwuoZC/T7BbOkGbMcMw8xmINHyWMq8kiOtVygMyV/VbgjFJi36RanzTWuKtd/h
OGELEQ6UiMRM2Kk6aNaujxljabEe/kmvCMVkY+oUPvgB/010mdZhQM9dyBkzLsHUVkorWDvEB/WG
Z0DUN16eVzptEC98AUSgasAnh7CDgWKwbDznk7QKHGR9N926/itGT2wSrygsfI6aOaSYexBzkPMn
U07gU6CMsUlqZxbXWVOLwiXnUCDAIoNzx/ge59L8VS2SF2yvce5C2ZmRbxR56RHfwxoFYPx8zDB4
DmP3Fx5qN8yqiTKpQ4bSP59CyTbwOyrlUjxH3PEac6IcsOfCagmJMYUpEKO9r0WshfIgSRhkFbyH
x3FK/Ga/PSs+AzmsN/lE+evNAedKnDQyN1LLBmdhgVYvPtu37VG5AkmPjzzteYe9zy0M03uQ0kHK
+sxIiqeGY5Kka/PfgbLw9ljFVf7d873nwB3/0GQJwAjVD1FSLf5vX8vykcAtAbXgpARHSIBoJ0fQ
VQDOkWkXg/z1AgzFfoinngzneeG22KjWhYlSbUKW+uQVxqUJVge5smmqTEnv2GztmizmKChqgR9V
87aEXAdmQkY7wTC+7grlXQSKrxoDbbwarHHYn4i9XYhBjCvNUJ1FEXZF5irrfifIlDrckO8h4rcb
n29MkjIQ6D9mSHAlm1ROOrNCOijDrxw/b/bZA8zSYETAxn/Lh1FUf4Qur86HqjYq074EDx2qAdRi
vgQPXl8wV2RBWERAMy9rYoqF1WB6NTPG44M7rpQ8o2/beVHX0HJvoTo+RDgHkfhFm8F+0BeUdsmL
SZDAI6DW8s/L89dZehs1k2H57R1v0Iek5kK8rA9PY0LiLQyiNrkRTBsMXXW6FY+S/0he5pZoha3p
K6OHZy6Unh9Mx2VzrTM2AiqfEPK73dywNsVrumYoWsRi+NeHbgYpillrfb2tJZIcovQsUBWQ5Shg
DwcQMa7r2auGqYVgPMe4+GNpaSFB+6m5lVCTVeQ0VcI8STIoOFaR7m/NwcckjcCS6Cz6e35raea/
2W6vhV6n2y9rrHAhEaEQgieRj+wpR+hBR2aX45gXqIbL/Jit/uJASNGwR8EWrBkwJ6zT+VKMrAFX
pvo486YlKZROLjLNp90urhr2muKx3oFFSyJM5DCSHw44usJVmo5qoeBmSdPJ84Lzi2aYL2ZB+zWE
47LlJJvlt4TpRycZH2A9one8Ug1nJroFwcfypnB3raA0VlZHxB71SEsd2oAKA81XjZFVFNUcErzp
pslHGcp9+RAlSH3q1hicP//OsYUmHtzuep5OvXFOyw19PSTxWQYCi+2dpAdm8xzi1dsaAZrdGgoG
U4UO58wKSifPAmbO/uEKMXh7B+7EBUOrv5v2eFVkVbfLZ1jDF54mW6AnyJ8HurERDfs5Ngcx9DtT
59+gQ4gs8DSDVR2T7Goa7q3zRZzMuU0q9uESveio8SdQJ8QxB12B/62r4rj7WOiVIblOrbQ4XVs3
48w/9pmT9Tapu9G3p3tXJEkIrnQphK/BbEZAwxD8lKwU+Of7mBk8gUQwVALKiFeIYqCzDwEX9weq
ua9YqlhAvSsM3w8v+0ibL/dG6255FGyJOa0qP077l9WOvPjNpvvI6hTcVs/zoloUETJ58ixNvfxe
2sn258x0XqnX6uPYFH1ZfRVDzSuvqoLisPXLds/57iiGm+LqGwlByDhWzzXL50nT8Hv7lBpkahM8
T/DBxHQ1HNtWjuhb5Z3CGGTdqx6XgIUcckiBoukMbBrkAr2AXrHdt6GuXWkwMGaZXbLbuTX9JsSf
9/DVAgYMaN1u053lMWZkufBZcPoc8mHTCvJBHv/D7H2/ne+CEYZo1AKaM2iiOq/5yXEqK8YBdv4f
k7wMFwzokgOs7bxkMQXThB688rMVuZE6bBCtFSwtRaC/BH7mvrparzx7uDdtRxUfAqjbyGOv3Rdf
jzQuuHfjvY/0I+mgAyDZVFcqLhOmf2juvXp9Jt5e0XSK5XywSDUVHj8i4OjVJY5eno6Az9Fxubeh
HPkn/ghgW8xaY93mZrJuy5TH9bmagfQVgZB0zUMNh//0WOn49HQC3SeJUygIWHLsC2R9YlJBi6Ft
BLKUDqUAK1d8Hq4AvK/NET0fbgr4myYQSc5AU/Ru7HfgVkJPx9A5xnGyGDVU0yPFcH/vUgMyzrlM
2+858BNtekcaNXlJziqAI+Sz+dvc6j6mkp5TzSJHk0heILVo6obEQ9rW1kaGbIeGdwtGaoLts1SQ
Nz1z3X0GIANc7yKOqa2rl+QLPNthO6uBzH4QK3AoBFUcEGRneLE9MkrpdOVldCqC4PY6kr5eUkD/
t6pYUFBM1+mjPfT1Da+17q1Oa/cwzziqDIeuRKCSib4jz+dXAdmFgVZF1mkKo8YaldaA4A1NU18B
HF0DeYRLlv9gZ8bR9zZKsStX+Wr0LjqE820e32v8hxqWQxOQEjCQBHnmhtt80z7g5Y6QqIBtkysx
H3Af/ZpWW36aeSGAppkYqb+/TRnJYYQaiZxwLt/ION248VEHce9GsZOQE4koWsci1ZoIZWBftnA5
0Z6Y9Aq6pHlDBlpgTOW+s8sNseWxj9jQgiAP+ZB/HQvnwYUXE3LCfRYB4rRAN4a3vaeFkLdtZWeL
qiUGYv1lbCGakFUrezewtO4/lvz2U93cjgAEZZ9adroDlGLaNkJetyjcO8YHkynKXFEjYcTwLIfn
3WGSC6sK0RgXTE/+etIe5Tl7AX3yRkk8BwN6xlgA32i8W7xGbz5H7zguNOC2h+RrvHjsl+w9R9h/
zTqUtJNCogajnoRg3snGUcBF21VYW2NVUeGNATeCcomSMLsp2rVJSY/hXCTB9BcmjTNSr9dBrnMx
rlRt0u1V+5YIW5KUlFBm0K+Myw9I8AujbQUEEN+xE2dBtFp+FMfDSIlCRkN5874xK5nHzcc0ySnw
BQ5GIx5+9zWrQCwxGr0ffcGUU9Nr2hkPoj2cAAP8oSZJmA4Ng2IfFsF1Y5DapCQyBwE3sJtEhjs6
2Uj+W5LJEaHB7udACiApe3855Ox/V18DnUiWBwovl5eXvWyK2WHJX+X9fD9LsGOIZPkYFRPwghHI
MvNUGybODor+Ywj7KisyBnfhla4dO3mspruTguq3wgORoqy+fdqnGZp7EuvHL6tTqHW66+gNXwmM
ypK7Xj590xLT1rTDvFtSYWxdKy3wLwXBUsDrcsEnNsoV3n28yNd4U0/+rrs2KfdlCmw71UrnR1ZC
laiOlQPfrFIiwqJN+h7qy6Nh6PP09pgnhttCfPegpZ1PszM0nQfhGh/Do5+Mw6dfokyakER3+wmb
1iH+6I3ZA+h5GoNjCcenINRVcfVHm/VWvJpllIm9UCPVn2qncS797mf11g+xodA/ltLstJBTwcZX
U53VuYZkn5JTsl/Vv2EQJB2nLauN/xef/C5WbS6hwTdZaIZc78nyYxfcEoVco69hM2n7ysiNXqDX
1B7l2p9pk3aFVFzvROVV0AT19EGtSDBnGsNqvdmNIlVX/L48pNUbNxpeQvYDy/QkTLbxmcy0M9wy
8hn+vUHd6N4Sd5iOCIXehIyf8BeG2sC3oYOqfqr94WMVY8z7sVZXGybBNlCII+HqShonRen0BFHI
Q+XcF9/BLark4NTDpCR7s0mCjrEwch5tSYkdYS/jiJ6ascjAif38t97H38EIjKtRi6bg6bpyI5Pa
ZoObrESD1aSSJclASO1w0hgEFRvVo5wdMYnk1rTeheNPjkmYbz3xXIAxV0n8E/6FinV3YJmpxLq0
uXLTkaP5+3PKj2oZrj4VjW57Y+f2yY3zepF5wpJOY9vKupmoM2klvMiD9o0BCd6NEAYWydMQRlaR
clG+Ee7Nj4te5SbzJN4uh+/yEvfdk1lajFv4oAfHiIxU2ZlP8wsdU7v7+Eb6/VXHo9kVNJhqd+MS
nRrgLnJysCPCPghF5xv/NaN9+n8mJJeKDociVzLikQh9vcIKfMqLnU0/RXCbhMu0787zryxjG4t4
4e8E+efKTScFoQxrGRsbGMuI0/sAFE2CmgESTSITG+0o9lXtrzWdxc2Y+twiDYbCq58me/zoZ4rD
lS2zEQcg8nxgF29qFAxOGDt5A7y+MLY5SgSFVqWJqpi1GLeB2xVRvz79uzhaunQlEWZV/z/mJ1Tg
JO/bo7zziijOAHbYcAt4oVDvNCyZ6SE3Sz0RFExT1Hyy7KS8cVFsmZZhVkmIV67afwz7l6R/RVAY
sLZUUPatzz18EkIV5ZQwGw344GJWvUribX/JWCuY7QZiuCtDaODD+BHIQQ0K0TX+3prZqc44BLr4
HLVOR4cKuLZxDhQfi28MzpTLBXZq/ckaSU1lraHShcoRkmzDqS7F4+jEXWP33WJeDNiZL4M6Umwj
rdK9d5rF7LpXoGavkiX2oukIgvPWytWMOZlJzkevzmg9i/vpitwyu+BKeAaOFdVgKrh5DiQxtDaC
eMgmYOPTMS3nQsrlGb+xAhZlCH3Da/OGskRxCe47EaFjbKYkwHMZm8caMsyFJlQcT2udz6dAvSVo
HncRYoZA3TT8J5E4MhvNdi83czPpOOm6KI2U5rwa/X2ewuRkBgmn6gFABDYYRNpng5rotlN3Z7LS
AirS/TpMSeNcxCKHY3bsspMRovQ9+p0IzAeCFYZht7eCWCGvORywiW+/xxMC5kJWZ72dmddpKHfH
hQ/8+dq0eEGlSvBSQpHAAPOEuq66ZzDo7hH9V90hBdCy62pHnvFU0PS4Nj2sLQO0nJiNt/4Tai0y
Pw+9izNnFAx91YACRTtbUnVFI0Taq0mKoifwCcRZz4S9avRKBhStHGSDA/4cY9D/7r6908aTfnSo
8LT+FK1yJwHqvA77UXclFAzOMtUOysLb6DfTCZIkyiRxWcsJ01db1Mysx51R2WIhQZuDHZHa3z/J
lNhLe4e9WEhUP6ZcGXC102DnEVIzdMlKCXjS6z2FdE/ZcCWRBOLM4+QKxVzJVvHegheQAZ1nLQkq
UOFviP3fh2bS+jKw127ty6m0Yy5H8hq+eJh62N+QXi5xSNYUkW77oNw0tiZuAw+ejCU0wLkl2JER
RBL+J77YvOTDXGM1fI/EPtQVGvmZ772KaL+rslGlrblOWYnT93R1mSLaYnaxD8aiV/iNkQBUxabp
IG1XDCZ0HBhhhI6MHubeEYZQE+Fp8uEa5Ez2hfM31i8fV4zngtILRtYCYXhZDVFNY2J3deHUX+Cg
y0knu0buE+N2Q7SepoHpbCc4eNJn+bxMby5+DuQtYbZMrPyarpFsO8Nltp/pDPEUpw/lJrMtphzr
C72e4FqsW6cHYhX+l4TVx3iRiUOKIy/6N6crf1gfcsl5AC3FLuGVR7k3sFcPgakwOP9umZbFpozp
2EB1vmEHrl9xHXSIs0CotU+AYweCaKADxLfbX3F2KY8OEmvPLQMchbcJ2pdSzilmWfhbgUShBXzz
lSwlSPdmTEgm8tfdIRhg0G4lp0N8nipjN/Jjlv2gqypXFKEQSSS8CAs3liP6fC5CBwrN7WtGn8mo
PUdpZ53OQpX81vc4PWQQmKFBrM3BbSnJIQD4LDVT/BrxgOOWHRP0Jr3KQaXgxW3pr/Eor727jFjg
+/zfG3WspQz9mEPekv4rvzqefaZRds5ld0pSlRHRHmTgqHw5yg1gKzcnVmmhpwmXgSy9jjplOLfc
FGsD5/kxWZPhxp9jnc0zS2KJPFLHkz3j48rqtToVUAzVp0syF3Z/MiZp9YZTEZZK936QAh8pp7Mp
SahVty8V2rLfaHM1kNaXw23Df7OlrVYG1OcVSle24Lja2oL2K8Wl5EcIW5YVNsDES3tpjrc5t4zi
kW/nFZjeXY0adNqTRlXyx7F4aUy5xhHnVb+FS0N/ig8l4WPVHTbIvkyLbLMa6iQ8jv/j52roVeMW
OpEbzBY7e5LWXdrlcrP2vNcwq3ruaStwMfyopLsBGhfDy8WBhIkTO6HnPnifzyc3kBpWWI74eSa3
YqGCBcsAgOhTjXdczvNk8zz6tSEFkAuyJo5Qb9ZEYnQZMiLdXwS/teVsdRMmzHSGgEEu2JeO6y4e
5vf+4TBvdp2fUel98zRuwjRzmi22TqA04Wo/MyoIDiV/EnH2Ns2Fmt6zLGLphvMHEuLYSBV+HRSm
xXfvD88sQSsKILAEBCKVizdSL3kssFBKQQmSFz1GpPi1gKdy7Nnlm659iewaBsVpLxn9hM9jqfWH
sMJsx9+0BJ1pQsfRCwjs8kZnOlfUikvCnSrP9Q/kRssQvSWD8HipX2sUSx0hoZpYh/OGh/WuloR6
E6/ITRXi1dQadjTXK4EquxZBNMg0siOa1ZkbJi3mXmx/X4sk6cIzmsYzM96nVerfnXFp4FZw3Jw9
z3yRN/PgvYw7mm86Sk1qyTAongyuzwfMdl1R6kZLVdrlLCAjG+50QzHtSRqZ7z1Oi53FKd685L92
eVeRzasSIcCOiqGxT2YBfVIkWMEPzcQgOShYYwzZeiJRz3sfQx2fHOBYszn4zLHDSrgjQMn1ZkJ8
CTIGvmUicz6/Wgpc/V3W4tA4ZEhVolmKikXpVRawErM7B04aZXz5RJaTDhaj0uwo/bnq398v1Uqm
nxOKbdqYlHjl1Llg4WoEB5WQiYtk3KUuMjrLMZSHXSkz4RYFl/iER2dmrAs5ImrSD8+qbJZwZDGl
VRaqUchoRT5Oc55Stn2tGZEiiJAvTHGXduU4MW3d2sWjoaSugNUvYhd36kU+i9Zm88bB3d4H/4kh
BF3s0w1m+jXpJaml5iZYGNyiMU9zHEWo90xtMvm1Rk0mI72Ef320QxqZuVsgpi49pq5SjZlGn6jk
on75tTAM2jcMTYDZfgJ4T8nm1qU2BxrsKINPFm5dYZhZgNQc8p8SEM78BSBO8SO9S6xgzyJpWZ+v
oQVk0pDfUhdiwYmUJQ1Bz0+SIGuV2FcUoCcMw7PmiKxqezwQypVjuWbK+7wkbQwySmjYLZD3mSZZ
1PcyqYwC2YN6L9kRGMAXZ3tKfyQxumm9FMjhuR730zvpOsYk4aPY7Ed6I6a4/HPIWw/sFUwINRh4
TlyDe9t5uiqhicoUPH19li1Gom3y9R711eBmd0yIHA+S1nwQLkrSX4Ay3TtzvpRQmohfPAxSc/FV
9aZtj9XBDsNwMRZPweqNLR3MAxcHn350ow8nYDn6AgIHApif3SbEnna2ZXc4Q8NZ6Gw5A0JclZzC
sGhUyrhtPWSeDRNnxyuN+7BuDkfmjAVo2T6vY8N6q/jU9IhUmXlz+wJ8ukLom/kfUT+uMlZkIu/X
Eze09nOxykpZaFi/hk/iGiFy3eyDtP9R3UnC/JBDY2XlrLeWQ8ghO31O22Jpv9d8OFHR7CeyQT3T
Ap7Bs9C76sTfTv0nOv9KehPh82mj726pMCM2bOlz1a34gJDby7/V74Q+mmysdKKFehu/fsnHMdSh
JXtK75lhl0pLHlHb/lX+5Mb16/bXKvf4iKpGgBSHwJ9VrpDwleMLHvf/nXRy2HpY/Bx/73+ZpBFG
uhrLSctFFtEV34IHFG4rZbkioKCUyr2fNCva1lbgO+0Ic3BlP1hOu0lYAkKTHx1Lu8nYVQpOWTzX
MV2LpWHrElT1hHHyz6YaH20l3whDYJdZRcoL4sRlBEA8tZfpn7q0LG6G35PGtW+gU1OXhO7AJ+Yl
FZEeNAd35SmhQdfRTzC5eHMmna3bK/pmw0Pn6p2k7EBHUkBjvqouH1g0KunPtYm9/sy/Uw46Vjte
roEtj3zHyUTuYsilKMRdS6BDxorjSvl/p24cyO4sHVizF1+sIYv2NyWSsaEyIb2eB/3fVTToQ71M
i6OpN6FKuk1m9cT8WPLTviu4hvri/+mazLA7H6qqkI+3Kr2V/qCjCCCgMEuCCYGtjLgaNtcW5o7C
4Fdjk/3m1CRpvL0GVE/GkFE0NvyCdAy6mU2dGM8EhjGS0Ddlkqv4uDBUgy9NNzvzeDeN97NnQ0xJ
N4tZjVe6PWs7EoklxiSWS7jMqERtsWUugfWIhN+Abm1AmbRKaf0fIYrddNuyGFYo4oncnl3E8+4k
dTl3/mvgIUh7vGgmq1crfvOQ0AtFpYCIebMa5F761vx2fGng7VSjl8caeHi024eX3Bm+toXa9Q/f
j5VB9h37KsjRhBkyRpdoiE6L3WQ7ksz1tvFWWUTL3/g3lGkrnS8IJO4Ub6P7VXs+JMHDxFnsk7oV
cf0DIkhwPSuBdiisErWbFRM7/vroxVl9HzvqhQVwCP4HLk4TgMzTF0+Fddur0d1Yn2FQ+ctdtlXP
WG1A+wR8BGc1WtGhtlnqvDbLvJOvlRcDwMdl+OgcWmM8IvBu+uwlDv5lJWDHW2ToDKlgegvcQa6m
eqzg7yQmd0gdpt5n7xVB8rsIYbCncJNPMlTUVGJ8xkl+fnooEhQFpEtXpjh7a7zWUKv4sg3kh3pl
j/zVVc/0n7M11Wv4s3HDHC8aQLe4Y7qZnPJS9kv4YYyIEKQvEkY5SLJM3LWpdUxo2MC+kz5XrrOK
VTT2JT7plP4X/VcOUfSbdDbCEQeZcVdEnZu9yVDYd3cgUHDGUBd7Uw0ad+RO/RSNmiDKR9P3/Dj/
T4MyxeYTvqhp/Mu6Kd38Wow4FK82hqLI6QXqokKBlKY0JOjS1H35KG2t/ZrfClwkTTq1+vZnxHan
Xm9AWRhuhXyac4NOgUT/yHmz5lNnxJS+Uraj3PITvPLujsOk1vss/bVWoT0C/o0AisnCOPEzbvxd
1PAYeRnvS2wB2MiLI2ZN5oGH7fnqpCGfTYrcqBvg+wDpHWWSGv0wpIrf/vGG0oK5/BLzmYf/YudR
DQ3BufrraB0+sRdx6I/x8HLB0nhHBCRIUQYYfgIYBQTJZjeloQddDPLGCGfI53XjlRqmftzfZaAR
Fj+StXcFN+/gvxfO7T92Fse0m0y57+VUaZPnYgmwu4IYC8kfQ1+csMdZR5gPodsO4rVZfF7Uhp3v
YIt3TRhbyoJ+oxuDMZywDI95GXYtErs7xxvBajSzyx9Pmi7ghxsB55crv8YiU6zL0+srXVtjs4WY
klzX38nGRnIgWDuTJIFApU8pix+D03y7mfTQdjRp0Eoyio/G+VcJf9STiHGGlPu5+Q3FrlQveR3B
Xb0++PrHh3WQpjWzWoNEh6Xp6Y//FQ4Q4zqsLYJHxZ7tDPmwiyCaDkC92xuXRxzRGGr9edjZTezH
Xc94GvKzdyfe9UK+PrTCMBXFp5fjAXJNd4ixSup+NmV0gN/ORmvUsIn/MZt8QfWffHnyskAIiRUn
9TGNL5yn4PyTuCQq02WEGuD6FMe8Di46LtYA71D+84Mhv19C7S9p98Lll/Gspg+AB/y0IGxBHhbU
kB1begx8RuI0JWAkOgC3NQMtko8u3SjgtgW0zMFeb7MKSwiUvg6KKb4Vdu0bLibhnN+ScFlOct3S
mPwbnHK3xBmSLoz1WwL2cxxOtaDEz3hZ/TbxyCvGN/XaCYpsUKynYBjMmHp4GN5R4qO7Q2xIo0hu
cOKTKqPTEkhHSt1uBS7AC4hCBPonHn4FSngSTUX7/IoWXO0C3/P3e8b2e0Vtc9t0HgM8Z1i2ypUQ
MTSpi+CPqSNHJkM6Q/+/mnzlujw9n3zTE8ScOvpLdNstRW8st7MLejTaLOQWOMNpVGPcIROjH2+L
byIzhOogVdCr1K5dtkmjyqGu0rpk01weTEmVxgk3spu6T8VZefHKXyhw4YUk13YkO9uJwNy/PyH+
unKwEqP19r/qfJuP2Zz5twtzHeUCuPL8XWPz0tYrNsDY6g1lNgpSorQ4cI932Wo5z1InnPzTPiQb
kCu88w32N9BDt+Ewqb3BtD5yIIMyc64tD3KsTlzinLV9Cirrfsn5arh53Mfnt/Q3E4gvTb0rcb2H
xbp7bCHyb5Tfh2iRB2ja0iipupotDQTEhabkuhMqznUX7RTh94Qn1cSl8awdCj2EujLlNEcUZfiv
yZkSm5V2lSfKRMUctrtIJB+6F7Vc72HbTvx9vgPq8U8SnXSDeASrk6SE2RUD6lcyABSfjMdIRcfX
tAiPv/i/tyHiC2yLpCzU41W5v4BIMd48ZRM5S4EQUKjhWvEFIouSI684gHkz1JqpFT/5kbAN90BB
3TO3wEAwyVCQuuxI3hLoyl6Ncy7m+mRQeOyETtS1Cb44DsLXe2bp593nU0dwBYg33jf3lhT9liud
gYESVUElHZVAYUMOKz6+JwKX5/m8ppJBaiyx34Ywm+xEZxqcyo1qGKxss+wU04AtmHQ0m+Ql2BT1
ZWDg68NKdOjeHWEnfDBbrOPo+rAEHoLnYAsVaI7H6PgkiT8itlDv1z2e1sOaY3rFiHQcxtX8VE5t
9QAl3n6vzUzDSyPJKePCSYd3ynTg77tRmNup8of8WLuAvBxiyGGDJ2Pr+xn/i4vYUZd//NB/yl49
l76ZkeCm5xA7LBAjZsLDWx5hkl/v2e+aB6mSOmL5CcDjUCelyAQHp0+9hSaIMwykMi2WsnANJyta
oFuMFrT02jtXhONh4Gjsm/woQhJ+2B9JJWOWjSHwW1Tx14minI32G9a/gJSOhKP2aDFJ6e/xf3Vu
8sUFxbW7Scu5qIlkGdGRzpSWyExEbTzf7EuKBkCY64nLK86qJkVEE3SjxReA3KjZshrjcRhJxvBQ
jMiC5Xm/4kCIfvQTM+Bu7Da7fi2CA8eMWZHQj1Hd4f1cX6EKreb4ZMdPpie9IOlEvw1J5BV4oE1L
HCB0jvyAvQTrjSqylTkeI9s8s5KS9VhWsnrdw2OAGxecK+e/DSd7Ta2jhe4WmoPFwaGiQ+odWpKF
WBjBgXhr77d3dHQWfst78AUzTwy4pSbbneqYqJ4DeYfmd9i6pU54NSlBTgt8cZXLVmZJYwhPHQEN
y048RxuzUXVbashaXvTcdQtradGUXQU5E/NgA4jRlQt5NaMXZ0q5Gl/eLdlrWH6Vt3Kdi6BgJkcT
zsQB06i461RZben7WodksDsS2QmF7r6vgfRXwDT8bx7ZmIBKrtrXC365CImeI+WbJDjx990HYA92
5/mslBdOiw6fYnerM4z7+Iher/NMEsVd+jNDCBR0quy9nbI8hYBH6lrgjQMYAjx1jxkAyTy/whyH
xJEJXljAGJ5w+ihVatGDVrdPBWZy4d2aG+aUnhJmma4W8ghyIq66QTGj5bCDNijKHp4rqGPp/no2
/+yTTamEx7sHSNEdwn1bx48UJBjoz8UPWCStukyJskcXa8fQqLe/jgmxuzVvaJaoyT3peg6xS+Gt
q1EMXC4+iAHxmEBInof5yVeOuJlJDLopCyi3k1esGfcxGF3pBNbLSwmuiJUltiIhwW14VyrHnZIQ
KAJlFzIOKvdEIHfLtgqFLKBFBV/0jaHBRzKqkIKDmwCa2VYxsWVi+nAhILflVBGCn4N1+ry6NDY1
JnnRZEaAKBxxbdW+kG2xTL1hVpWNzSCt1C6PvbiaLHKDpb06CbAT0Aj0h049RJml9Fgw+aUK3GQN
4QcLvfrirkuo1VvGvHtuwj97G1aUgxMiLYdXFpG+5oKMCOqoOPPGfIRoIL0RCXyqqzVhVLHFUq9h
yrxHHSURDaF54tlywHPErExk5S3FOzFgjy1WpEOA5amzWXTH+zoV5zO7iVXiQQvy95pSE5cc8WfX
fUFRFbnHqUcV5x66dTeeZZzW41QHPAaRylM64DMDZ1sAHHyBMsMlCVaTROP+QG9/goWND352EdqW
XAKY4ZJ6fNwf0/pnUCs8Zyle8NGWUVECFvmxLzZae/rfUJ3NhGWWBhl3A3MyzxpyOvK/+iBl6WvH
5NgmHamwfBUy3m53ee/vVi3I2eXjA/4CyrZHdWDx33jDQ/xBvM5KHBNghcTQx2JTrS4NwFC68Xrz
63Wwtbit+6IoqESvfJCPdh6rS5JgWX+ilEKWiygnzcQaY2l8JYGKhAqW5AYjY33aUZed0zQmu1DG
5ZohogFBSRoEePkSunLkRcyhGpBi/qxwMks3K2xajru6raqozq79mHlcffv8lnjxufJFvd8f5+xV
0G4WZlE/3pOKcUADPjzHeeWlaVPhIyXSS0vdX40f06DFE4NGQdCzHKkO5mpBcNKN9BQmFdE9bTEP
c5cw4yYhOb29r2kCqrJe4V76aF4pMOEyUM1zFhxAlfMDlJIFgPBN8H0yApALERLeP5Pw6UfEMAg4
QVw1b18tDSyOWksT/x1Q02wS4XUtVpDiKFQcr78JDurwdui/w1OAvtpuj6A+pu6Vj4V9PlwpkQWK
qirxshEJ7k0CVMM6fyd1BBbOaFj8Vn3gbgq+YH2I4PPzVDZTuGKGeiSGWKFytINmaIq+zpsqnlZ5
KD6IFePEIbyUiBguxsKr10+PHNwthCUqN5KaTgJQPSrTFInClxXyXf3GJ7v5FAZH1Yx9Wj25ad+b
XmfDgiMMArYA9eBijwrO2f187wa8IxUM2IWsAMs3fOvlO7ACpNdxhrij5hFK05oGQaezaze36J9b
GT4Wf/G2g/uVEONpmhOL5STcnIqPOrdr8rOh/bFslKDX83yml+pAshF71SIqSC6TUoEqCiNoSX2M
icW3hAyJM0e7ZVJCJjIU07p7SSpedbRTDZaaIjLJ87jNpp8Ytmor7K0iBv7VBeYhoHJGyWvUS1UM
McquRNLHwWnBVDF+0iMK40uQxlDmRTUQDcvOBt/hD1lFkFyJFA0on0Q/Af5hgSOJX5lyUrHvnXI0
F3FslFPgrJe/KPqlpNc/Kpw0ybHc8XmJI1PMntnPbiNh/xrvpXzxxC6rFJwX3UomDjGwZfuhdAox
WPGhQSUoTCSmLqA+xUEwNFWuzHHUKZhHtnNlILzKKzTZCdkkDCTCgpwbbsmNRZs13w4E4weYip7S
mvCZ7G398pgVmNxrjAplWKuL5yGDYTVVVoD1NRRVefAbKoLZ27cEP/rhncFToVqEaIpxw6Z+Vj59
6psv2lPgaBJGTeYjuaNYnNkCkHV6efM+yRFv5NifH0PsxDsSQWcq8poSIv+r/eInYCnTcf18XKC3
MKXFDUijswudH4u0sAAh442G4pngiDTAYgDknTaWMaJQ2hLcSgBqL7CGp4rhnvNt13+vct1bNa0K
qpJ29dTPjlCMa4AR9JuFBHnsHusfP8lQ9ujostZo4gY+2si/YB1I+nBHIAPTXFpQsg5nm+MIypOD
ja4XHl5wVYrQbmUnCDuwgJIpYDxyjcK8NMcFfBKiHjaCXB/A1khNiTriT7FIXyVYqiqxdF3KtSUI
qFrIXCWy3iBD3AxOuBOLadmurbzu7IKq2gMsXl0EfJ5Yt/25F+KHqIiSExOtC2my916a4ry/7Na/
PMvUo1xEWhzi3g4myafKNmajQ9PwObQ1+lPhezxLvhlJEeklgoRolzHzEWIliEqznnFo+3Q8iaT6
Ko5A9ai8T8ybhIR5lSldC3EHHoF4XKFtu6XcO7eG39ZXfgE3sqHvopbHiqc2sHGB/4clMd2vagt9
3E7KMz8MYUx4y77JLUEcjQTOX9MQA8psJn352M0eJv6yRGVAgHwDb/DFoyEPhJly0qiN/eALQuMT
PJQ9QJBpkuP8FzQVqG5YdpUXPYQqYh5LdD5hHXQE520wpbrsoKurRXzoMsQ65oq9ETFzI77mPviT
7SmONMCs14CdAtq+dNLUweOzeBjP6U8IsY3TI1NFF73ril2I6dMjRealFMqnz4H9HoYwNHOiIB4n
8AtJB2Lzw69bXOJeFxgkjQvm53h2pedeK2KYOAccSvPhERQUcO0R6fhzWsx2uvx8IfrLpyoRyCb9
bhM9ZpCtclKPd7QK2ss4doM+RQhAuWnPETl6MMdWp5RfdrzImnpOopPvssGnzxejA21ml5KEZ+MC
Idb0hV+J/6tq7q40hlrK8i/X0q8D08+iHdLWo/0BFhSoil4F88L0vLXxQWizArRVWpX8S3hGe0Ey
vldUPn24GZidEXMdFavy98NaYRPs+QtVi0OIz4Qa6Eh7pUhQOAEZ4Hrdp+1m7zN/vz/7LyvfeOvG
THkV/zJJs5qbow3BxRBqCrE/5Yt5f1VPRHE4TM2ftYm0QeJ4dV9ktnb07kLM9pIkq/vZIFbEFPEd
Ysm37/ZNs0z1052zla22k0v5fwq+KqYmqSkKEJo1RXQ7M6OhzULAIFE//faP+KwUOzz0Rc604sjM
xTCtojdJWQvCoO1g9yUQk+CoBQXbl4NItcKLceitfZHWd575A25rGZCQGACEKUBdVH1XuyS44M4K
Lm4qgLsneR7Mo31u0enO17dpXtwyM7HMQJAgWJBFr95yxGr7yq/4HrTBWBZJ5ZTiF6oPzFwDhidh
ifFN3Cn55dehraf3WAillzLEKBFXQJUfB2rR3huf1hNodfnFVSZxlONpFwCkejwkKm4RzB/WWVq9
gZfiYi3c1JAXEMUugU6YUw7B7/otKS+xQskUVrz9T2YGg9Urpe2l6YwFL3d8ns0eTfjjTOZCY1jw
k2ltpnVbZjpA6Lcfmbsge+sJn3he5eG3N3L3epaTgaAM7xig4E6302b0XquBOaBF8NA+42I8RSUu
8osmq/l9Hs+UC7aJM7HG656Vr9usWVPvqT9n4mej5TA6i92igHeWjYldrhdfyoeNIeKpm6Mgi2r2
kzKBvWH84W3D5cuiYRV658TC7K2g6UCqGNyrLAddfahLQV5xIuRVjchF5nvuv4+lGatCV9CvrYdJ
8MuQbnutN4rMAYSYHC9okiH+z+R7lGYMqU/OB8YaMok43z498py7Oxd6ER+99B/UM3a2P+fnmfEn
5KKlg0oXo2DTFZ0XiKTFkYiFFMHus1+pUhCdVZ1rUXFD89wJoey2o7TtfgUCKOxd1Cy8vSVpU4rg
R77BVV8cwXAe4hLnDQ6s3EZuGQUrvZ1XbA6GdjRQxOJcjMQUlUzNW9Avy4LJhAuBoavx7uJS3Oj/
F6fZCtYmdSwqpVsUgqLyXelD+TPxvV/48J+Vlqk7P2yyQgcS/u4R0ZPzwVnLJ5aEK6gvc6loIlUS
bHUpQHhH/n6dls3tfumqWOftOOAInFuz8RIooYIlqwB30qoh+PShgsU5lDdBeb+n/a22y+YfmLAn
0YjV0JhgmmictuwblU+Brtj7SYJBA29f9p5tx/AJaS9ksnjnl5FXKyiZCrv7ENS9itDvsARTn+AZ
bGrKkOIyOnXVKsQQLoaTjSvHZMQyw3BmrYdKVoNBit0lhc3LWiIr72fMckxPSxhX2su6F/U+DmMb
SevbPJewIxNZNKbVKDLCker4hAIaLagCsbwZjgz/kuzTxiHyy2+PPVCRqyly66gM/B2gII6aosM8
jApcM3H+jnKBkBPECPBhCJQE0MbcLQt8qWkK7M6gAx9pMe3WKw2jg+hfyRVp7IAo95aN3j5Byrmb
njXwhRyn9DoYb+tqAtL7oqoo3DUDnnLkhOOsFWeuGFwttEQWO8a/8qgF3ZXvvRnNyAbxCjsF4QUf
kwdVYdW2tLF98SFMzgLAvOXTPhzATMdCDkZlybe+dmJMfkplJCALY7Boo2vTDRqaRSnzp7t+Qntz
mS71VOZR7jM/cqlJ+uRHG8+/kQt4GVpmb3CgsCVLp/d7blRFwVeNgjcOacgKCkMCtLVw8hnzVgUo
l9jsNoFUXNSMPWvYCitQ0/Gi4GSUL3z+2olXFV6OVa0FDGW1XMAYmT9/d+zcdz/2uDTU80qLK2nW
12ylQjr/5l/50j88Wdf+gglEPcstPajlPgeKqR7ybeIQ8sAIWaLT7l7cykeF/mwmbmW8tmK0Yodu
92oHxgejCBJig4tJNfANDJRfc7izTzHnEyS1ZLu3bF28itfXzO41/p5lMsuIdFyIsPdT7rNcjCUo
RFVoYN9gU+p3WkK8TV4XlNTAesI4MHWeJJen6U0pxdK3/7sggy9uLS5typIQLMX6tA0sV5RZKPkG
M3Mn/JNxD7wkAQSTbdYJSHYZK3dfMk+qODAS0xPKad5T1NlDmDStfWrpBWMhNIvj/lsGND0GyvcO
llOPGe9Ojl5lejSNPdMYZU6YrlWjEm3wieuE86MSmo6OaEoBdavP459eS5fBA2/cp4sCmTnmLv0/
5Cq/B/W7Q9rzZA8D+UzF7kzdbynhuLy6l20cf08yP6BEjbwOZE74s7cvoreC5LwjjNMLH7pOohDG
gxtY9+qLcWAERz1+wHYshJBPC0yg2St31jPtaW9BwUiw9ya4fHWHCHOSLfCEvl/FvV4Skz/PTyus
GEPr9agZLhge430QpLCvoYsYaQNQIke3hynkkSGuSJRUTWBef4m4RcZYguev5k7S7N8Aoa9A1tAt
Nv/siLgxBA6DYNbOckBi5MWreCgJF8DY8goQFxxGuOPzYImlD2HV4RPVlz9Y5+3GGekoOxP/W+m+
Cwp9oASIvL0RiMGTzn92JQWuzsH/tWX36rMjSUzaCjtq5TVcC6cM+3nd2OwG++HHOOxpTemAeT77
ieq76i4Qqh3ZbfPpXMNjjtmyy9kbnGQDJ4hqRLhbYEb1zZ4cOBjJAnFkDTHpnoy7/ge1r6yOJZC4
zCegG/cLpyQp2UbMsGZCL1RRFzdGR1p9UZ3Dnso2te4PPd8ruYQ4MU/9bMccNwgrv4ttjnjPItPb
1VVF/sUbnVGjQ9qFrGU5vMLmg91A1LNsndnsqwwcebtVFi4plobgPzQ1tAdb6iZ2b+ve3c5Zins9
Y9cpGzNTnuAqSJ4fKhDCn6WTiHQe5jxrr/kFE6LZ0xahH1paNFuSeNeabjz1iM4e3OLJvYKOZxF8
+StE+TmA0vf0KGYnTFbw7yPyLgoD8f9k/0J79u9wF2GQlrruOvGLAbLsO4iD2krzX2OnDzN4Db68
73njXT1ngwG7Lh2/uiP/XDbB8ocNOfwUGNDBgNslPf/nKoHBe4gKtLIyqGhzKGqAmugyqYUrnL+V
d20Hc7uIbN713JzVURMZ1GBfSozEd8MhMlAUNuP9F1g+t2+AjaPUhXtvasJngWHIBdofFzOCk8R7
e0qhOYJM+Eoxi8gQAR+9/sWewE15TZP+MUAJp7PsK2sL6fhOOSiNZauCgYE22qtvdf6LzgGldZUc
wCwZapOWGnslP3GaZK9glduH7INptmlFOl+qZAeIKDN5GEcYm8hU0+j/iKelBdQRifXJNGzaAL1k
m3/voVcOdqxjSB49OE3qmqIUIuG1iWxdCLlJKmLpNI1p+ABYGHLKMotM+PfO2nx5fcU+rykt9RgV
UKwUkMUI9KZz2v83m/dnABCCiCbXsxFdtZ8c38rymDl5wdQsPfdJBCk0i8TmzuKLeSnC+wHhJOmJ
jtNX8dHah7aPNqGCr6MCgx308X6gXQEW6ICC+bwlDBdbLly+3HE77r+5oxRmA2N6y0nPUjFz+mEv
Jqdev+WkcnN0OsRhwpGDOwBecpIY9SZXhA76ojinbHmUnsS9sCvb/EbmhEE0EjZHSudblmYHoJBk
6HQzLjr2/3cwSMvp4l7sEmtIDLfUtJEYDsiq+/EBmubsdkV4sKT+WDlsiElON5S0qdPbS0heiF6k
9v0Ymep/lB1mTQdvFm692UmAUZHc+sGLg5k6RBOwJxC6aaBmYGwe1EfDHcNNrgqcNt0ZO1wG5f5Y
3PFcwdfMdvltk5X7bT4b+bTaQuxzz4/VI9wu7nl7KFmHcin6hQLbJiInUu2iT6w6sLVUoi34QtEy
4HXZPFrwAtgwQPNT0pESMA9ZM0dJgk3OQ1wDHt03c/Qe0lPym0iK5bnKFsV103IuHUZwzp8MxlKi
RD9/AJ3ofvc/t9YBeGj0vmcFf/tuKt40lKHKUYZ05I9Va5lQPdj50qdslqZL/v8vP4b5woETp7kC
QTdj4i3vv6nQriU6XD45TLYa3HeAgG5jY1oGNLTtagKUM49N3iMMoHlRmutZe2s0KRxfskVwdWds
Ohwj0JxaRma7IXWSy2sCdQyszNXnBpHYLzDIiWHOP6e9Uyv4pzGVUFQGvLNDlaV7nLrLIRqShO44
uiwzIMy1mYeiKijE/DFYAev9o+adE9ILXi5hoIWW5i6+VjdH9QqSVC0Nm7pKxNvG6AXwxEJtbNf5
S1VP9ZjV99B3ZC4+f8nJvTWaeqU77KzIcoI1NcFUUgCHltg/f89G9KiOmnH4MW3N2HVbaip756Op
YiQJ2OtXM0W0ILI14y2mrTv13DhSgRxvyINUyBRs22LpPw5Vh3jRck2AZR3hEc1sL9Bm4voXAuCd
WTQuCB/nn/rRrElX0hSSc26Bg5ZH87eg+dD9fiYczxLPPttbYw2LVHrlbYh7wQBUDkubWudp4I33
DqEQRmptZ4jB97EAjrS07ZYklAwJwfKBggW1V/sWxzHT0++RNhHfpJIdT01nQRAx/yRa/vw77kil
dLO72xWx5omlMZ+9yosZPkhz7XUyrPABMV9wFbW9PZHRl8zIzHYaH+wtN2hKDXr0myqOXmKpVjT1
T4cxYCe41Pa6y54iYNyPfd9A1s6bJrq05FdF/xf56S8oh18fYJ+t/jlI/AprnRf449LFKesUAQOO
J1mJZULwU32BI3htvS8Zn9nxnu39W9uDNLmRmbxVHHyaN9Ch25/iunuyw4mFvGOrhI/gB57+lRm6
5wukciykh48mxGUxL9QzKzZqgkypklaUp5YKOPZzW8JJNbTuUkoY9aLkdCChnXKzvlQ7vvu/LCBw
+EqamtxC88Pi1DlCM9BnuWr5NaYR3VIo/oIgXhxyePnpFipjQM3o7xqSxopluNNr3wL6UgKMq22J
MjG39RtAA1Klz+hJlupadZSDObasXG4vM/FflAN5zHbZfcwCJnyA8O8BvS1IunUJmaTy23jXYKSy
f40VMI0hc2EI4XQZ5TqAy0QD3NJgjMbZVVaNRh9qvZzFa1UxaJiaZrH/6VscvR7XnIe+hISE+1cl
Sr8qIbIXjPW/6Lo2o5cLNJXCJWTUTmchgyc9N4fKb9PRIch/EGYG+x6jF5XrbhgXqRbTblSYvJ+w
qdg4QlMR3QTASxJJUghEVIwOftAqg3+FT4J5ZGx5EwUhml28ywldeH0N00DVMdaVlePwLTM1z8Q9
l33UwACHye7mXP7vmkhQLrvHwWIGMWfKJic+BkvrggmT0axfCPlaC0kFJjD379E5mbwVr9JvwA5U
v8wOQLSHSUj2bInKWloLrQjYeYqYIV5UC1LPg8SCoCXMxL0Zy9AlXXUQL7vq3o2PaJtIbXCKhZ7A
3Xd0hCih6fJRtpIRmx0+NHTZGySgN2G7Z9v0wLoXunyDF7WB5JLHMetJJ9UoQMITx7RT4KuBynIb
10KzGBaLOo07HumI0hbNitRT0EcwugDbFgjCD8TtNLW4gqC4Ak713C03ZtV0XejjxU+KDG63hjlw
cLts2wyGTu91bi/tcES2rN/OglgfXHrx3E2TeltRim1+d+MUPG7sFzrYadoG1dkaTnYWcay5dNoJ
VcRLibBMsoTtcwGJx05iNN9eVRXc8viuK6tMyUxObq7yI0qrwxAcFGGPlNvpjA3XDvgeWkOgrMoW
IadrzUmdLsMEQeNf0TTfESaWM2KP7dgbXyfFIjZ/CW2DClqnydieLc1G5Bhv8NFrwEQG1tWnxyTw
uOSzWbebJ6UTDRtsCu4QUf+4EjI5GTNRyXCl7x+grar2FeWIVXBCeNb0rQ8qCGuOvO0uZuqCzDm7
jnEpcHSMqHnTfoIDpcdPG1B3e1dPKNxcyBY1OO1UZA0DWt4Q/cgUoohdyEsfA3PenZDXpdyj3vku
M7KegS9V6Z1shwpXikf4I9oS7ztbXUtHoOayr0M8y2PPSEhn1FZgdKS+8XQmCYFg3iOajWcLylI5
dVWDUNfxRFBdw42M8G+wMxoombXRlev3Pqr1rBPc9CkK2T77LY7LijulflOnOnuIBaAcQYvk8RlL
bOc/gUHJEpulaR/H9QMYAND3RJy3lpLBFbzMXOLZaURICqlLSk8SkeTpqaAxKQhqynY2VX5rDrFV
rx29UGQ5t2GBx5st67z5QFC3hM3x3p6eF0k/3Eojlqk+fFD/tuDHMbD7h57QNA9CTtYsjCiodQWz
xzakmfXtKtPydm07cpQnTfjfv81um2tFpSLDS801kxEXn0ugyWZeN7bHwTdL2LQ1nuTp8vVZOo9Q
yUQ702arvraZOedW7fLRPbPDKOHExcjketkdrgLfa9d62DiugZa75OsSV70MLVS1v42xQc6LZqcx
zQd1ruCFpbcX6nsC/gtiXl9MyptuzeM7RLeDvmOaBFdrAUGH3yhj3yFzSvbtRs9fJOFAwB1BXZ+R
YtbH4LCwdXADPC6qhLdXXWDSlexdSgKH81gQlQ9EmRQiqMmzQZf8TK6VNghZ19YLCx9SLLaJo8+h
9n6GOzH27I1ZClTKGkacQ0OrCrPHy9UsCitZSs5ciruPBS9UeGDbSd0hFg0iLbjueW3VBewu0xEC
CepEU2rdv/Pq7/r5hv2QCq55JSGQ1QaKqnWWkBuyFBRQSmEH/wbgsH/cB/lXuyy7AHxwhIzBTawf
67ylYZZz0hTERb6TZkmTdTD8Nr2ONLXLSvWN7PIovd+cLudAj4QhJ4Ek54mvLgXgtLpgzt4F9+QP
h8eG0bH3B5iw5ZZ6CjEB4TqwfYkdq0XXB797afNwho4bxmygd/REs1TFU9qGYwX4GKCrpUhNryJA
tsal9VZOOwh188uwb51xKlEKtgCXVjb3l+anf2gHMRFYFCB7KWPkwD+Nmdkc9euaXks3seT/bWSc
kD5Q9iBY0Tvhj9D09ReJvIz+b6zy/9tc/81uI3dAgDoHdGG9xW/E1sZMN+Fnfpn3ito/nR82+xDY
XaY/guyNohPZFUHDjDcbQOiFvmJA37zY1lC8cIGNLDIAA+apMKw+/4nmEeVtN1n5yqkww/dQ5imp
JPSpIckbFbRkNlCR1IeIqr6WFRGL0/+6kmBEGOoAPI0BAmxSThNygRi2n4wXdFNF/WQIl8DrEetv
8xb8HArLDgKDwzoUpI0PtA+iaA2CVaaP+vbKTM24DIprZHAp2NCeOX7km/ILUVXLXwctzqVEpHCE
qx7omPqYjoXc7ESrBszrYK77GuKfCOaSwwqpKIAKx6b+i648CBjylTJKt0Ygy1AGCcZ8ZspZRPg5
hIMjQxI/fmfJIa0DlRjuRMgFMXyXY306rxppgN58C+rEqxwiTIrkSQmRIkvBZtrBIIB47kbznYKf
1Bma6YTlzKz+F7Urivk+bcQ/goFYZSUlTcV/WJfm6xcZ7KO2geb5CEBkVEo0JDNAw/mhXCF8uUzJ
08I++L8Nes+qBU5gFI4VXNbGK4VQp61wOk0gBhegq73ocPO9wUwWtw72SeFguaZb9Qgj1ENwXI+y
JDsrhDmCRK+Sp0MuSYAQoreO+kGm2zIZsllJfBeumWFxWHnXwVhrLWMCnO14Q0zpxynJlkgPthrz
WEvoP6jfI+SdhGG+t4GVY2XuhOM25/xgf43fe0jgDRTyG+TfLwC9lX/HC8ZzUn1f6G9itnWxETia
0nd6yTp+AKPeQZeYN5ju6QNTNikH0QbYFW7cKDlTX3bHdPkcU05G4LT/vthANCeqFAY8VHW5zqZO
3WxSFQBk2XCC7fpgJfLstE8IkNezcMFJeklRISZZIWgQbXd+48XVD7itZ+mKZkfejUG43cAHHG9O
v40qDOkiowwnoWPTgljH08WDBlJAjMlXAXaKJH0QexeePrpbetWOzKqbvzgZlpGVqP/BLl+hsbCO
/asCj+GjTLyR1mbbZw2kg8klZjdNIZK3UtKxFWuqi0e88yV0MO+LvKApjQg+laaLPBaDa+IzX6u8
5t7Z86QoKqrDBwfSuWzT0JTHmqcqW6ruuCklCnqrxdp6hcaXwJ+WfQ+cj876Kj7lOk3Tc1Auhajm
oE5wKVMC+GcOyPxO/mQp66qzplP56bPpptegKSVWmVdymLYSlHJqduCDBhK2ybk+cXcDRH5sN9yL
a8BsLen8MOdlQiUi/LTYf5uDC5OE0nFPR33P1Rr9IRuLotFiTRPc+vMsjwIuzSPWAhiCCYnH8Ac5
BHuK0cp0x8zFSXo6FuD3QWkc6PVzEhtiWVdG4KWezBKx8j9ntV+ZNdWgWBssqh1wZppiqdMSiaqQ
O/u7Ms4tGOtm/JbzjZ2YOhiinnWyG+eb8/d8EhzLLnGW1ada6w88D73MsgDVrS8dhhvIBbY0kEkK
TJSciqWQqiwEIZm1QEqplkb92CpnEbx8M5ka6sW5oS20IL7uBVFWmtc5xrTrtcg+IaY3mOjWLETG
N+LTlEwqbO/WJ/L91R0Sgb4fQKjDtdRdWiff3VpZX4+e6lJJ4Y0jxgn4kUacj5QXHC2jIXikUKuQ
e15mzwQdVn59xqAp54VULFC07KVovaypoUJZLNfras1ZlpU303B4L7rGolh8zCasbiUCs15E373G
dZ6Ihvh9OiwtLG6Pa8DZr7rcDIS+v/Z1tuzHvFmRBw8Ceqb5YayZj4CqE294TOwmT7kTe9C2e25w
UWBHVmyN3EmZyOtCA6UDXZWPEOzfJTT5g1Nh6xcp6KM5BaTiZ5IB9423Zftyp6pNN/jXWeuz7GSE
516VroJVu6H3gi4vLZPxVZQV3z0+J2E9y9zGOaCHirQYTGdv/Fc8sfE/QIzgjKro1hjXB2MDxT7y
d5WuzLbUH5eGi9OLC/XwD73KpIJZtxh9MHSGwQPgBO3iyUuhbLBGMIQi0NVjtZngW7S57tFj4JLs
qr3nmGfS7M9t7SyshrEmah4c32JLg94AqtZyh/b7IPGG53ijmDnrH4OIcG0gGv7NuzJRsacS+jdw
qJTEQ1WlBa0Ih655GlcwPF+Z6lElig61Vp0St9oDvcXvqmvpdSZITkCXFrE4c3dxg2qCAKs9b5Vv
HbmLQ64Q9SLnBRt8o837ib5ZsKpS03Q9LYSfQRGI8shaWw4jwfyFqpkepsr7tXYAjxivVDIawX8r
y4ypnLfOLTu63JsoQ+Z78eVxZnIYS/QVJc0DPQkVnTpjGoqHKGf/xoaICGOzN6qKb0GLrJnZhD8M
TCFTXcEpcH5vKRK9BY3ZC22X1sjl9N67myiMEnj3AOUyajomWVuNRyp9zVi/Nzu5QlG4vQ8vMo6G
VfeY9K45JvXeD6PmPO+lTxcyZ0RBdZd8GLrrW+W2wDkU0VNgDduiFvQKqgcKozNfGc8Tm5x6cb1K
5HQvo7ZC3gnQk33jp+eYUr2wfo0mV5Fl660lS7lCeOjJb68ZHV070MwiTy9k9n25A3mB63Sf6OYg
cvve5i9HC0O9IBVwGvEpOF04yYLtC9emjsWe67zGEeiI0Klxfl4WJ6/fpu06huGB0d5bx8EpBp+E
SDKkUB6z7EPevbghQf4bePhQ+NHfqhaRch7jQB9nAR9zermc4QXPYm4tLLh7IU+9xjTtlENP7CNk
SFje2uJuviJAqmbIKltjTrnpS1L8YM4xM+qHcFSFJEki28Cr6MpCQP617Xmojv04OPzy1we7GO32
bSOIl9kNgdpTQokfp9792/fF7zk7Ca1Wog2iDFP3TNOJfsbDdk2kuO/yi5anTCkNYwN59JJ8TR/S
3U3oVVgtWyiYpyhCJIipA/AU3JdCZ5eXx6vbpMuckAoppAYNUCvVZcphUz+UYZ3VeaxZsHY+YKio
GY1mxkFJbY/ArV1ajBEHaxKh/S65uSKAuzWg8od+M+0nluK3NuJq8sMAuEGudIwnwaQZ9+lV8z16
fO0KKPvTcNPg6Q+PwR5/zEKgUwwZ0mkTh/7bYu2KThePYPibZBolYF19SEBzNrdaOzqjZRZ2TjJV
Zc1BeCj0e6hRVIp/hMlgIdzdxIXM/rT3uqfu4YKhreJZxQ7aMSwPlQ54/iklexkS1F8voMsUn+0u
3ptunK7QEaDtU7ALiQheMJz9hwKxvqaNEnIbwBMRHi0gRqtgX8E7ZuCTiIuE71lStFknskhal4hS
hi3qCgBhRmShMWVKAedqBtHPeS2HoaNhb5adnkgqp4DDSwToDNOMjAXygk6/DvTIhDYocjg+tKUJ
WXWHTGKFIWDjrIXmgHM5gKE/IR5gKMdQueIhpiWtF7fnesXM7soLmirTqrlZW+U25F8sSfEpWIaa
bSai7UvsNkmWwrIXvwZGWhj75ETTJ2hFe0sYcU4K1nT7JRKYdgyswVMuaoyVefJ1vexXQ001WtF/
k14nnkDqGfFNwIWdnqGLT4carVSDGQmDBsw2+hAXj1oINjEsWkhjyrkD1mNW6N9iINCxjjz6wTme
D2JHDfY1wpo9/l4qumvhJRNre8idJmZzVSur08AQPcv7TlDpjxFM28zd8Ny3UPjvCnYkdH7bZqKA
qCa/36wD0r6MHjETDmVw6SCyMir4xmvTboxMg97xbwop8RMeNR0i03evscfIqN4HErvwkdrjETVz
Tno+eFu1tkSvtoVaxb+659xIkslVZVQFOzex/kZg3TTVgjgzayMDF5NbF1pSckdVibRcHJ24mT9v
aFIjK9nMpAD5UZt69LgndUpFF/qtTdDOiKKN13To5b6Hz+H7lBV4jTmUQ/Ld/DsMObtsPEzELnWf
uK23yqCebh7ufxWrCGjACoSAezqRoHolji1R/R5zvL2YlkpEb4uUKXhMGRuekFcR7TTqcJFKkIEL
jqdbWb+8uTijU7N3wIcSrdMlBSzQGbiJDnqLsmrLG+/SvD+G/eI3tD2LHY6dAzIi/UR8q1pGTyHU
2lv7Pk6C4C0noT/FSILDIi7uGJj/T1DwgOlLMYYOtv0L4NUe438T0BIVBP/ZB6cH5ijoFQ9h4nHA
CcGoSRSVT8V+c+8Ap7lUOLa8f5BXo6jHqbsAf34NSfQ5735INKyBRQbFrbMRWlhCxfkqOlKQuNZm
D0ET9418N4shNU1PpsbWDpoimQYDNUZdeq/YfZWFkDFc0RO2PBBgoVuUnSeg8x/PEp0wvTMaDBa0
9l+XDUDbj/qRl667XkLoZt0dE5Xw08qiXrFTHY9rJf8O0faf8W1fKPXxq6zGFLSjge7Hb909IA+h
49R3IrDSC98hnUvghd1A7fMsA3k14bZTx/cCfFC7mAt3dbsLrEO4lXpHEjdwSoL5fGfM/XveglXZ
n2zWqWB4V3kG+LNex0GshMInbCBbqRgyp9TzKS6aQnwkAlXMaJ3fIGojaGDPgvQIo0qSr1wM/9Ba
YgqXQdodlR4mrwlbyg8owtnYEwHkhx1RpeMkxgIQUslBQXt8ulI3wbrxCOj7f4B33a22jLeR+dzH
L8cINUkfvEPGxZyJZFkNp19OlX0P6Ag7byooBW2wnt0HkWm73VHO43bxga4ZsovcKcLwFgRBfXTd
Ab1QIk2P4ExkGWzL43rAhWucKdRAjx3s7dByA7Xo57Tf276VolRH6ipylejoRbw9xCPDixz5eBw4
lR2HbbR2XSu+8PKc9tB/6OxAVR0zVeczrnFkPaR8Qx0yX5ZBU46OIt3nn7rrlzQT9G4Sk8C6nGX7
68gTbMRgbOY0/Vfnv3dGWlSYamDy6BNE6IfJD+eZlHZIxcTE4NVjlOsHL4IHBnL0LA8ipjnPA1b7
Cw+utDpSGIzstiL6Mss6o/Eto9K1JVgdpPE+ZBX26ksYES696wGYByiJ5j0TAFSNjNU/9qN8AdYD
xx8CPFnxcXPNePJVGG6/EfGrkFq3T7uQfXlGN2JqYL2w+T+EiNqo9EAOxnImyGMO3neOYNKz6KtE
QFMNVVvBDr0rYztqk5v4Sp9G4BQ4RhtojGSv2pcunhHlIH/OEs+o5C0+Nk06mISmnYBPgmigF2Oj
yFpI789JcWVzJOP2sycf+kX/hphGvdziBwe5K3mzorL+yqeFOTFh3JurrhDjdAlPDXU/Ai179CZV
b1wwvjbpBlrMRa0bBWfMIflFVrUiadqqRpzL/oxk9j+QlVscMRLtxiWZx9KkOYKJyv37ecyEK7vO
XDv+GJmsuz5083FyOdgWNlPqVfpXoIcKagQ9q9tqV6B/Y7WRRUUHgKJPW0xUCCTv2bn3uTxDORlY
hGHoBWGD1/PwIUnIgFn8Wuq2BGQgz/mNyApPXzOru7F+JnqiIXu5NzWZVt87JuRpQLu5s7Pl5jJa
0WlOYWD9shCLEbcRXzapoBATM6JD45fELiDGMMNSGGv1DRInQKhJ5Z/YkjlPVDpGMT+2CV9IjbZo
R3hrnesaStkUHekHSQSakLtyp/oDs5KD270PQAyJ0/mjQpGirbqdCzXn6yDrjMuC8T1GS5ClowPd
Vl/UWOQipcQkw55Zx5oXYxVy5ak8UOFWXQ4A4IQ9pCzPRDInLK1fykHB+5RfDTjqwSpKon55Tnmg
ZduIe7rM1b2cj4oD00hw4X8vK/Q3gvY1lq1Td7V4GcoEW9ZwXOiS9JWk0XnqNj1pHDORRw99icc1
YQjX/IHeZEO9hbt+qLVB59v8tUr49MYhwf2x4spoOgbx9EwBe2rxj9pkg9Kw9zgWBc3r4fMtexen
GJIUtJcmlllELMXmDHch7Ytaz7kt6ZCqWELZiqn7eZTwpDMBl1otLF54ety55iTgv8bgmo4I5WMg
gaoOlnspm1UB7NQoxApO5/fZNHqSPBPGu59AWg5mOvBk90AxinJ4nPBcmQjvNcCKgW4B+qXFmaN4
/oN+ME79uU61WwITlY3Z5pHKjYL1E+cTSAG8rXwTsvkp1V7qdj+nozDuViKlBRs5bFkPup8bD1t4
lWOltKbhN4y5hKJQE8FbgibcXIVgGdyMeg3BuUHN4Z6qHDgixHfwe2LavORNm6/hTwUtYVcK//F5
g19LY6xZCRd3xVppucYPlIVbCMdg17YsLPeLRRx1kWL/f+7gIU6gbbVgbI5nU4hL3gjCOVVRp6ZG
Hztn+SZDRkGM4rRKQnNrkWHGDONdE3ZZ4Qmz5xYqrfacT/GsMTdo/YFtH7nQhWqHvbBIYwxIu9kc
ylYpi/d8abngiYvPWRn4LjSQH0/1MwAbG38FLi3dsIO+J06nkuWBz8PRZO3SyF12t7cfuy+thFV4
m9jFIH0C5C9Ubn/Jjo7yC3mFlixS3wCrkteStFmKr3oQXV+UE8Kz9kdD4t2+6PxshCt0iAc+5f/v
0FRE54DTf+HfNR0P849QARxjXedoIuxK3RhtnoNm8trmhQ9+BDWzo2gNBmDcCM1kuKyyotnwVtDX
3gKnBcGazgnH0m5xq9ryV2KrgxXFc8Uz/8tLqnnDNnoeHRGYehRi2TYy+XRyHBfxd4JLQKeMHDjg
zSUldBuVPo7NYGuJA3SMRG/AzvaC9fYl4DOSLlJH1Jndf0Ottudw9rXXuIkFob3kDQEhBukI4wB3
CHCB602FUdnwLDYy76dDjaWEXqsRRT8YOh1m7zuhpPHsytNreB0HVhmWyYR+ZapLvm4vgwfc8NJ1
kZYwVPZ4hlARmgME2YPMkgFGCAYvSFoc4oSWuhpQ3Qo5WNAgDHaFt8aYmGjmZIOvw3FiNRh+xDWT
aWXBwiN9+kFIVDuZ9CeiStjR+h1xDRI8xP5BIV2ZWmPqN5DBEcRmVad3YhNkJBHulbvHtXYO5i8O
XrKARIN9UyhY1tg6IIgNPgJ/7yUoss5sVQ1vYgztuLZgh+1I6FoAHeVfUiLr1nX9WErPBsAT69d+
cWgqdMiNvhkFN+iaeN5Rohq9EfVxoBkxAYUluSltHAEfHVFYPI4vzXcmmniMfCL5VcjEuZZqXl3H
+JqnihrM+ObmTwUjpkidZ+zVhshHidDgZMhso1lsqYChFqBwJZGlffArU9eKKaqKi8E66NazJS7q
fZBy8Zb6dY2Jq2Vdj6fo7h+PS3HGtfimYkTPk505p7tduPIAqGcyJJJQMke4BIqQREzYqxVRegkS
R4npUEjT+3oi41bXPws5nhFfnv3Pi64tXni5ttlhbOQTHlWw3DaFoqbvxDP25d1ilcnNFEFatPNR
3JBGEIneYtq3wSj8vSWMnrFsFimFa6YDnBUlG2C/8sPBZ76tOzl7ARQfL60ldrrcudQ5NhAodznq
aMcxgL38TLmVC878fYuw8QSUYaOeGrNfvFgX+OELtAqGHLheJIdwDs+OjRLrko5Jb7wj6BfDJLP1
KXzxy30jZ0RqggpBU6cwrBkIs0x0zRpElZP9rvdVPBXWo+5miQtab29I1f0rHKWw2XtlW8w3jPc2
nINFbKC4Pn0tw4KRke9gfoGHUIgwH/rQ3KA7VcwodxQ78Kb+kTJv4YohjEdzhni1MH7W27OGDhn5
76VIQVhuUUbnynXenMZvWqU9hAVdHjg78QPaSs1Od7dXphKJBlrBG8pe2HalGYM9fSANJtVBqiJA
fzQPhwRe9iOMdwW+QMe+0/XmxqvLbexs99Bs65ZU3+r6HkNurBjZYRbal/GaJcxsVr/aeLvfF/d8
bR/YDKMGQ3n6O0rrIk8CKZco0lIOLtYJBKzPAmv0VzMEiUg+Me7otjsZVT2WuHuiZHGOwdscSCVQ
Dbq7/403fFptTPZjXFswS3SCkcukFOdKNFYhjCNKPMNi6TrqSnU+mzAqQ0SICfsPXMKhqcPR2xew
gBmcCUpJiR7lat9lnUvN/WHDeWJe5cz2eDh1oGSqgkxs2QSs9wq4QjLkMY0DlYCW+NrWck66rG1B
UTIehY4mEunX+5NYpWdvrzvWuqAat1Ve7BKlqzXGRyPvq8DKTLqFRtQq3DK4Gu3Iarepv/P55MAd
KJLzKj0QZPBp2cTV6TFLqKG9rPTPVTzv++k5pp5UKnO4ywbKAyjOIHlcgtqogrPaoZJODYwZdnA5
XtWQloqpeiNztQi78Ha+lLgyesMW376JWo6jaWESaXVBujynoYIhafGmrcotWHmO9EeKBakaGl1s
M+44DSxrsnPtxywstM9tJBmFotk5JwXidRSa9QKIa34G3Z8MEp2c/XGWQXlf4iV7p/yf/+Uh5pjD
+eQlEkrhebk+VA1erQLLOXE8Um3E8wvdL94dSsPWaautE2P6vO5Gtbx295sbhG3ofaOS++huWbqe
ZmmVuuWtt8hOLkalKG9neUGPEPGDZpt9yr1maELYKeoTLNseglLb8Hwa67ANB99bl4NRsjcvezCF
GlF9qUUXqDqeM1J6FAvyzgsvSckRsNxsubl56pIdlBA+f3RmWJ9moKouvf52Ssz4QD84tI2kKpQs
tdQFN19mAHnPzas/fsqJsXAKlrcyZFHqb80x33Fucw8t9aAqa8NzAQWImL2wZyPc8G3R55j7uMkr
Q6ryrKtdNkWv84ARHPnE0d+wEOgi0JwJ82J7Fqaj+v5tcXoBQCphu7CMlQS+L0dNmhvxkMP7RwI6
GWQJQBpo0NqnpiwVL0tGdV+aAaoeiXI8TZHNU14uPr2p5Yjw2Fz2vObrx4kagWgw6IpssnTI2M4t
x8lIKa131IFn/deUniIohYj8OcODC2+JT8YTfno75Kz4LE4UwBe6XeWYCmfc8/8Ip9SOgEDxrYY/
vCJ8QtU5CfunXZu/U/9QTRnLOxx0qF9fdRINyvYnZGSiZrr1oWW7+tntcQeU036saXbx+tRCYk8u
LwYyRVnairP2TTpAnCtiPEfQEIMHV9uvhG1kUG704p+u8o0C1Wi4Qch+BDFWDg1qRflVBU/Z6zbA
NssZPvUEkPTU2lt7HHCdbgaZDymZCurn+H/EU8eP/EtSGhBYzyTWOBiL7oMAXdT0w3VOXDwPxnOp
zD8DV6c/tU0sqK/5pwoLXIiRMNrdr6NNUgaH2A1EeTWtUd4qpOV6RF1w+2hBKGsF8HP9un6ZS+SE
4hDn4MuMFsCFfMaOZnKY30vpyrEjweUJB8IIB6wqJC/B9TqQReVGjE7YpY/Mg85297WWCiQZrutj
72OAqfUu1pVe6AlGEV/M6OjofVZtkalIorgzOzSQuy8WOqBB6obDg4mpwe4sjrMZnD+25lH0d85T
C5vBcR214M2uoJjUEylu+U11/yzJHMN9CF5KxAf1+sctYQ26nQ8PBOye1IYuYedrQW7QGTe/geQL
CxjK+OLMlurKKUX3GwABxJMMPTrOgZHnryNuamWVC/pOIjkV/GqVAHIJ+gq1Nu5+qxIt/0V9N+b+
g/rRTt1SL7DAtUsXu+GOK0lNAmg568jyizfZcg5Qlj8yDDtwc5Ovaj6xfN+F7aT8fvOVAhBp3Eo2
uRFqRvEOAUZ2okdUBo8C8Y9rn5UaJyA6LG23sAB5W0PfwZxiYqug6oJj1KZYQu5qXiv67Ct/dvzi
nf4a6pz6R81rSGsDnMSSdmKMJakHFbWvzwZ3cInlItO4cTIZh8M2c9lG17mlcVuj9+8x56I81BCI
8H6b+HEcLZxTVleUcGk6oIgCfE5F9ZgQ0f5bhfDh39YP6SiNojYsuJ6/yXSFznMYflPtZK8C4u/9
4YTrO5vODu7tvH+vq7Ek1pebCd20vHebQlxRIlnwSmwPhi/esTyZ67L/ftq1mHYFrBatL0nn14vv
dNy76zP3hvhBk5HWFm27Qhk3FvK9ojFDN5ryTCKRE6jk1nrGEkDngR037ywZ2Xgmk6eTlryK2Ixr
tMFN203wHtWkDw7PYVnJCvYk9JllJ3bhxhmtMDQV1L3mxZQZrYraE27JW4CEd8We1sKG34ADLWPO
HV+Smqk5z49jyWr4wjfd38/2lp8zBk8ZjBBBb1vCyt5D7U6zG4xjSnaaLa3VHOUJelvDNFooYWme
mDNICQ0wwZAiI6uH90yE6YGhinVbX/d3IowE8DHQzjNpuE44JRtwHipVldf5KZXlKdT+ki1PT+0C
3Aw6sa2OKKkWwXr3+2ZJekjZDVGet3327LusiyDlG9kOwbNMX8hc9l6yeV9J9Gw742Nucw1EhV8Y
yaT9HdsPdOrRNOfCQXlzm0G5cBHDrTqa0uMmbcDiv42PodSSo2OdRxsiHDFfq24hO/NFBLpc/rxI
d8AuPBN93C7ZpU3J99uYnJkGMwLG/mgO99ojt/zWTkf+VaTbL6G4jX1FkDN/LrXAanLGN1cn4QdI
9afsqf65Lh3n5LLQp5TvZGpGH/uvcHnQXT9vNsX9DNdN/OMIC9oX5DBLe6JnoBcBvqGQ0HofBAja
g4NeVKr4jfpHxu8bMoqioF88251H1o/4ygVAZtTy351Da+21bIMgRFHkHgz8QYxpZ2v1yvyobtZS
hI8wHW5cdvc0eB9sOZB3CVEq4gZyFV7UzPbDc9S5GKY73Ya3QBUllrXgxvugUEaddvZ+yGfL9PI4
QGL4YVbOcU8HJLKRo8Zyffq6TwI+tuOGmofaIYUilccH8iLf89P5GwWmHlkusiDXko6q5e26q3Pe
Cyto8+Vkyg/kVgulNoXXrH/mtH9nvXyhf3KDX3yvFpPZOl3RMj/YV648RdmRMW81tqG5HtUnrnao
iTYNSxWnAwDAuB27hakgZMt1EP4Fq5je3ieiZFHTok76PdMsCiDU8CFanOceNZavmtu5Paf2HMhX
8u2WeUL59KIcnXlLXa6iN28cM3rJnMKyayQsowS+IzZnwSpm5i8FtXrOhWVCl3lItAPQXgH4Xubb
zpWHy+JaVACMPEYRNNUDC39CySmHdGpQlrlaJHQAwJtwyszM8N/EpvKolCgF8xkfI0K7ZrisVnZS
6Oi3Vt5DKTNO3c/DMO43IIDvr69cV+lsmyghaNrgq4lg1tjlXQqcnawvM+548pL2OgwJ8u4i2fKJ
COak3N9O0hfz/4I1kxF36OIr3drpS1i4hJnj/vKY0ok4lCe17nm0Ddmut5CoIhpTTLPUuyPPLDjm
cxjRJ1GSZf3vn0rmbmgpBG3LXClYbNlLI6vXkoGKGysP68cHX0v281OdB4aJN26/J5Y1Tl42YLuo
8cYCqg9BiTBqCvBR8ZhqNuGIFkm8cj+elG+RFtFvz90zbu5Chh30DuHy+1F23MPSBz5q7aLQwswp
ciiCjhM16B1Kkd9BD+qJYi3HeCLApQX7yjo6D9qoFFPy3dxomJlhzelCjAYojlc01CpDodM0cpoP
YsjFK/shu63IJpZPxempfrMDF9rCByF5gfuyVQWzkraainzx052s/P3kvw6iElzc6preT2E5cJQK
sZVrwZwwcJ8KcRF1cTFXb6FjrfBJ9nYxrOKuRZk3mUUKmNLkerpbBbf5ZSiI/socvj9ayHAbb+WQ
PhvZVD7g/NTm6jk3YXCtN4gLLaZ8mVeIoF5g02h/03pU7fc0h89YFSGE1NFxkvnI5g0l3n/sKKw4
vsbaecKenVB8xZnnHNfymUXq3TNp9hqv/mnrV4TU38ox3bZLvmf8h3nZEOXq0yIeRD0n9PI4iF1r
bsvn8HhUoQOhuh6UYQkEgODruiSFn7iuy0hbOTBkw8QqdKZFhbEd56iJy3FFGjMDMNeutYe3zM7f
8mfNpi8kkGUZ3UqDJSZx+oUnmtm4HNZtD4jllbW7GuTPOh+kbZsWxT/INw3hbDBuY86QT0NOqS2c
Vbb1o1DmhJvqKCz389VjPTPH4L+hKfZqa5wBxB38Nob41MRJ03YemDdro7iDTc1fPS9KJfH37jB/
lx0eK6Q1DOlr07mrZPr0ITkuMyItKfAKN34TAE7YyFZDOCEkga8MEGOcg+336FsxI/Rhmpdylrcw
YFihZh1lbjmJHxLYpBAW2NdfD+YHq1gT83FbXtAhjZQ0y8gVtNOh1nkerTh77DfkSk7tbqKjOtdN
UPv/i3Ul9c2b1zFq9fDPm7j1KkjwOttdmrqoUQ4llMiLBGrt8kZpAY5QNDeYdpOZbZdhARAdqx8/
p7ZHO3PRIbr6F3wtmYqHtLLWjdLejo7ccsszbt9i3TXo4X3mLfRIt0JSyb+f2lx382dP0tTBsRCV
YxlqaEl655IDPatc97JqWILfrzTuDonKkwRmcfjxX/jRcOlXWm0nlBhQinIdeL7j6e6QKWWSzlm6
K/R1jf07fL0IxYMrrY8o2+yYYODeugTIK8tIF8i6UUCGlullZ/Bqpaq4ilRTI8dA7pqzr+jV8wWE
YQ36oNdnVGD5yXtHo17TKnMDQaeSRHUv+wH22JmNQ0Z3qbVqu4smXiln4Y9Y8EGsfvtMyRjIsQw3
VOhs70KiTld4gvFzih2yp+2KpM+ugYWsTaGGzyiZB+0ScxNBtRfuI6XWIXJPA/1zzFFSkEYRJ6jd
4p98RQdrBktX1XFcykxnj892DtiFRqf/EciPDZpP1TZuyLfMTAax0UTPlDGYm2589DnfMImqX2bU
qndtIo6CKzinG/DYrtuHkG1AghNHWsxN+k5CicTF6T2qnN6We1QZooTWciQZ4eXqce0tD6zKUX1q
oLePkCf1Cn9roWTYajHQSqe/wkgGQ2e1ofBoEDbm3eZ4ezyCwNNZdY1nI/gO6GvnZ7gyYtMgGu1v
54aXMIS/qs/tjOJCFKmhq579r6Ov6CLvHQkYhWUnyLMfG9w8kbTSkomFvGNPNarBTAzKPvUDIq81
V3kgAkTdGwQb/+y1JxJ6ce820yrq39ystFIAI/r4Ih9RAxltAFWFzO2Rnj9VfY0/HvW40cv2GUww
fTrREMGuM1NfrRvbMNIA2p9Rg6DBUTspglwU6kRfA1JJK9VnBmO8zd2Wqs/rqI0bZYAgcbjrXZHQ
njZEwtzEaaxv1lUkw5QEcmFwUHe/fP7MlJJEYG8veH9Rb00WwC4z4dJLNvcaqx4BLfhjUDyMPYZp
2lEE48k6FWKvqEu5qphJ/PyRA4DE+z8T6A39nHwDjFZc+lmgFb4cYb6NnXwAAV49wOCHRGQiOQhy
VtXRu+VPmbYaGY/1eZiG5qSSEXWBcD6HYCvBbcoiDsiWFREMHBU7v7z50oycTtlu2W7PZ3augP02
zz95nB4Zn+BdX7lNfGUl+M37ZsAVNTFzr3wCnXbPaw1MPgBRCXoAHdlmLsshqg96/W5UaaLug5ob
4X8suvBaHqwhVdpV1/bhTQIj4tTtP05yuRDyKkRjF1nHk5DC2ntMOpY+lH941jj4l6WwZn01mSsq
nA8N65xi6a8ScfLMz4mDpWzelz0ijAXB1iJIJyE2gFs8W65Tfh/dU4kjUJy3vbnzaJ6HaZt2u8fl
khpR5fWPQn0K/MlM456TezHGYPzUFMUhHBw+7ylmRt3Nm/48dLMeZ7PW7Q0RhLBEWoG1HOHoDTnU
8ROGgioJ25tvYlri/melAgziy58WD/cx3emeESD4EUquQtHhgoj42BgwpJsP4MAM9K9Kzhje9kb0
DN8VCygrLsEShyKtRmhppZIYNuZ12uIK8nrE78MMdMGesuddkg4MfOs5RvDjW78NTzBpvDnsTRYQ
hVuKqupufZBfHk27TInMhLyKDRWDthytS6aYYffrCXGUCgyucZ95HF0Dp4ZoKWIdCXVF0qXG7pWL
Gm03NjY8Tyoa8tcf3+C2wwCMssLOZziYLC/HB/K5i94CrlO3UKOXW5QgONhHAuhfdntiQenm3Ipp
WF3byKvLTTXv+9BGYymP7qfMq3KiNehJGuDZsr6QB+3DBXReQIfZvI1WGDRuBC1b2sirKK1b8+vP
MR5pcKsDqBnrSrEPUxiT81hQAbv55yTmAGDTE/DDXcR84QO750gq29duHEb2UD99Gg7pnk51tay/
fYkF8EOMyYcUmBn/lM5kxBo6Rrv2fDUGX8Bs2UQbSPAF9Lo/MI/NNSLbmoGZXOjqa7tiW0IZxE0W
dWgF5K6KfdZBCx9Dq5+7xpPV1f11prSSbgDCVZY3a4kPTiP94OVyTHlnAqeozmXCCFvOU4kOZdqN
iyG8xlNIMW5sKZYoA8ntNdj5YEC3/19Go7gBFCLeMQsimT7iE+8+/OlpKn5hDubdiQLXEMZEIdGX
M++/iURVTsgN2BzWDSLczGYNvbcEH7hNl7xp/WD2WPanFFmLmES/GtObPJUkfnjMX7NTkGDcnpxs
sRh0qP2LDixgKqlb/jvm3/HKwCtp1KTFfN1hiWy5VU3XbUcg4as77ouIXeTRb3qEkqGe7wPVEOIG
2zUMx+xN5M37m2Md3ykjPqZzF+zxwERdiDZPcLusDNIQ0xCWWefONm7YENeTccQfJBgusxmbsiB7
FREb8O13bq8Klwvv5lyRMghrvX2jTI+QXGQ7bOBr5nYJVYtwpZSTZ11KQb3UaXrqble0HaXlxRtG
RjNzICV4H8SUZRDlfO0ovl+8ZucedsgFeYVSdJl3tpCffJToZvbKNV/0o/gLxiO2beTxfkaTqsus
UCIe86adaHKr9Z7Tc9DU9avsvmKfZSC7908ZEfAp33XMd6qlsvHICU523U3N6FESR1i3YhQxX2AR
YcpAE4AbWGF2bKBrRCcfozkKEuCIOzKnUlmBHNxFjQTbQxj95XwbmsXDbrSnj+kaAOoKsxuYAH9V
nO7VQwAMdeD/3yO6+1HoHpPzDwtShhMLrYN+Euf7qg8k3B69BCgXyX6/BxYe5pAAjPrKwrDHxgzS
AlMGe6DvOznrcP1oKZ76uMerIgO92+eRJGYuX4pMjjgEV81Aas++cKgzFkfnHFAP80RF6o2P3GZH
/Lxz1Kk6Ppjg9d7fmYY8KzQgoRXSfJk5A/gI2TPmd83ScmnH23OMM8HppAFlxP4gPVErXrAhUPp4
RHsIWGdegO303Pe6oG9tdaRxv6vXuAyxA7BDTE9ScNgnvEWCOzj2GRIBwYTJhACj7Bwts7pBgbcT
KjxgD3xxYU6cnbjDms/1IIBXasuOlz/RiCJ9G8J86UC/KCBKtDBM9NyVWLUKAYmsPBlgT9BOD6R4
B5KAvXhgyknhCPyUAiTZ8mWtruC00uPSrxNaRO+6x6I1yR3CSBuecuqeD4k9hYoDwK3m644xEdwD
fJzgWjgFe4XfNm50UTQV8FCpv/FUikCMkxual1iNkB2KFs2OJ+RJZuO5MGhhbjP9n65XQsYG+7Wk
mYkfqk0bsaoexjlB96q5dTI9hF9deLhWeK0b/zzZWDSCGI4CXlaDHee+1ae33U2Oc+jTquQCmQ1L
0q1Mi3quis6aSMTetijFydTJvaJP30LoIK/0jVO98JU1dyi68oXlWS7jAE63bGKulhHqUULEvOdM
VALxxgHxNZJj5Q86Oaec+x2ab8a/ahxP9Ezcuj2Hb3PLgsuab8EaJgHCa93NVmHhe4ceiky6N76Z
6jI5prFdDwi7lnwOS7Ei1En55UfEW/j/0MuEAG+FEnkKMrmTM3Op6N56m3hlxH0LNVlpGcyeZW5E
85j3aCt3dshD46BdUU6GHGiSKz18/Tg6VqI1yxYQiGDnn8nsh9tB9Bm7ZJaFkngTikHcWPfcDEyO
6A3eZ9qVRWbEKzeIaYJHnL+CdV88DSdbJ+O2zhJZqOebxdD5j3KVVPzcT5OVIzTp630xe/7FsA7s
qqAASeXP/hp7d9kWx26oV/F4UZi44D1ITyNr74rnJXGllIL+dq4VpRUyYsK04tJ9UEY+HyFmIZzg
2OxgPEyY2Q5oZxmQAOrbDU/SLzgX3+zmFC/PFiQ8dc9/oWsJE02D81xuKdGxG2Z5dROt5DX7KQYy
yiA8F8cnrcFMwaApDMP9RF9P+DpN6LePmwr4h+ui5tQXjstgZ3wshjRaQPQiEI0+ROzFZ2S4NT38
xraYNX9KMlR0x6azOVen5CEcRFct0xOzC8Wj1Qfub8lvN0glW4pQ4CMLr1g8cvSCcZk/sbJucwwX
ANKJemJRJMXPXM92gKIHI/33FqcxNWncUwhi0tVwbnvlyko6tJHJDwI9N/TyGNF1vVZbTesu3+bL
KNgZQYOlDBvzUaViKRfWfw9bLtG747yAfyjnEDA95KkkHhy83f3BgqtOBoEyT0MlDkq3YHx/UOZ1
XtwCgVy4MaldNJA28mteYUGEGs1dxKabdL6ECqsgnU+v5p2fiePekOuJ4jyJSKNswRcjPUvd40L7
pJd6RG8EZ5XianV98WkV3VJ7vHOQnlmnckGh6Cl/gIPbrahO+mE40AYOvT6wg47MOSajkgEBpThI
5NoVgzbNd6oMLOE0aBZyED7qi0XnkQjBoU2pLvmS7fZprpoBWHUUGhiFwieFEGNK/3kDY532mMWT
d5yC4L12P95KKeokon+rFWYdM5aMbyaKDhsTBix32kgXBvytEOA0OzyPbjmZamt7IA+lkZbFabRi
r4Um9VwMjFKEIQJo+3SdDNIAdHSmW7Ds4Q9I2C1+NrLnyeY2s71zYzCDFP2w41MSqrrTiJfeLpDS
7X34QUtb87RRyiFRQ4heEtpD1kgB94BQmUjdLFbN94UPXz0x/y+vicPMRJPFbV2x3P8tNelKsp8x
KM1kBnVFyUqRB2HhsIqeeHOijUUAu2QTNFJ82902YeO/jloDcgfdjgICGYxpK+rvemPTgkCPlMWz
3C9BQVswo42ZpSFZ1s23A34sHG1v0swv4z/rkcH6xjz4DQfex0WwhhS4C/FaYRLOQH0XStOTUBNj
FL4Ny1kkv9Mt3qIPzDSotjocNpUiGAyCpuXF1dSSwaNZFV7m2sbkpXgULXTHz57zW7qS2GPeATDP
S4vlOsPChOzi2pIjFhkqO3u5Dj4DR/Qa0h/hNu14lOVS7esEZbXGVT7mx39WIirr/UZGJqu6GW6l
MuKLVoYMJmgEa4AQWgUA1qjYVnywn9cQauMG1qFPNHI+Ss7bGI3mGhvs3/KclFGelA44GhLjCYvB
/ulX9fxtwXWiTESrdSZGn97az1R+ZigK1NasM4tpkzK9GQ2D2qcZHc+fpUyKjM9ph/4dgma++akx
ndStKo/pJcrQW7X5gLXnnnjWRl32nju1PKBU42fjlyljZuMIYvPJGSx7GS1SIQUMDdSEOcPKtaLi
aaR5dMPxvmS74jv2eIIHBAC5RRzK1hObaMtg0AJ8sa+s7o5hfzE33MS8TnhprzTGMEfwgG6+MTBi
/NdN9dXjnBNOgM9yJEzDki9ZUwK8e9PbiAiOjzYhs+HpFqKY4dH2wuYKQhf/V02OqA2sLKUFiTxQ
DiZqyItUrS1qxDusw+9moGYOFe6SdB4Ey9YMHNfDJ2rOfC46MuUG43Y9r5ihcN66UQVyctt60Oum
wWHHdIv/ZO10OV+9x6IDF164MydfOujXhsOnUycxp15B8QqVVcHVwZ53T6syl+rfQNzdHx2il+ln
mB+setcDbdgAQNrMBuu3r8OngpORhjUDZdI7VDYt5RTXvhP3TFfI6B7B0OCix6q7BSgcejhTiMBz
IMxQWhBp1MpR/AKxjzBVvPtNMk1JXC+7cMNXtVEueZp2M2bUXSemOMrK3znA7AzZigIdK5HUqhDt
p41nGpf4aGbavGew0iVU5EIS8slJwOa5U3vcMUlzhBgN8FE+mH7Y4uTybPqLY8Ddl5hjl0BefkYg
u0QQNvvWqiIS/Z1O/wS3H3aMnKNxe1395e/UVOAVE8gENF6PJpZ2Bh9hb4BvMvGU5u8WvviAwu4K
7shL6VQuM+ySqd6sWMtMguOipUtyXj4eZzPMmoxIGglvuwDKLeRXNPQh645bmhH5obhLngNsAG9y
UZF1YwVgn7+c8SdjCNZQWD4aA9O3wJC8YJSmGrCHnC4uv4jT1l0IFjBsg+IysXpN6E97no2VDFfD
kdmb1GP3A/xb1J4nRS0BP25d8DV53rrkbvDzpNhS/0/WntVcCtz3FL1+WgS/jM/vb6ylteSmLoBt
l/QguPZts78yeV//xIAa2rvFoBJwPGKBEWYn+nqouCvi9hE5OOMm528iG0s45Q1eDCRawLUETgFj
kZr4RnhdvwEwh6Xd97qkQAlvQWjq64xUKhuYSqNeH0tGmolC48YGsS0WaXAUSsZqi+wYovad5MQW
kDPclZNFIZyrO2DAoZ98hy6mK4vAhLUiTAya1g1hIeZuUTVuwwhWUA+upRZ+VQpPFYcl7lhLgvnF
NW8fDCIsPoDv2gMZ++t1hpKimmGJVyR3c9XR/dQJs+a/xy8qPSl0sU1eusW6+vp+3n1agsXClNAS
o3MWQl+aKTNtzG4WIon56gYFqnpvytbNu3Hy9bmdiJYO9Xj336RaGn0Qqc8P9Ul3odINmrr2CI3Y
v7/5LZv0C8kRSCN2NOzcnt0SL5QI0kop/j0cgYiSQ/m4H3DFTmb0HaOWybZyf3Z+5qcp/eWXJySI
NDTm0YK2xxKp4Cl3V2RKtGTdNmzcI4shdWsT/I86gt3AoXm4q6D+cx/wbfTlP1dJw5UYx2lNiJFC
HwgvIWq2SCnI9peVC68FGKwhivHRDdmso38E6PsnCz3GKySAalHg2cR/lziL7sJ+G63xBgn9WN1h
8g1RAw+ImPk5zzEk3TwzpP2GFO/wP17VqupNNTCV8DXdrrvIZL03B71ItMPNlXJURBviVFKTKNGd
ajAtOTDY389AlYne0MkZeixt9zKd2Yifw2ZO5gRjFLQfbNNF1oWmx+jDs8BIyYwx+VTchZPAU2fx
T4mONrLq/orl3T3d5WAvESl0Q/80jk/FvKPEIby/Lt3nkxulJ6gpcqByGDzxvUWdXc2+MBQeLV0t
bnAPxEZFi9kc/V2P3/d3uvYmOeR4EMl+sQ/Fui6MqJIRmXXYw2fMetapNwL2Jfakr3sKCqz8yByp
YWr0DN6HiGFVNtJylvf/2xX8QDqO6ttev3niIx1VElgJ1Mk8p+kubpoJo5ms/WpJmBFqG9lntVyQ
t/rE1Yfa7Z9QDddZ9Yrw7pdBx3+3wwj5gSDFG1k6BD5NDXCRhuImIKW11fk1BsHKq/zsZeW/+7eF
0+FhNYDLMNGpyYbwQUu3SsxkJZrtJX23n4YIciWQYB3jE2sKQ9T+F/qmaiXEOczQC/8FvQT/XlBE
i8bsz+JfERTgMeghfJupSfOFO6Vu8gzXfPqKeuByOWXEIHAuIWly9nqu7GRuux8eF+EmRbIgMSXv
UYZf6rbV/JdBqTgPaeIg6V1dkQAeh4ki8ah8z/L0F6EDXrpQzNgruERM2N2MO3Kv5NKhUkMPXTJI
kKyjLdjEFHDwPe/LIlxtlTUU5+SAXw8CPoJJJYVS4kG2f20EIhdvdbMSTe9JzQ4b3MraW6q2MPpr
2gEDImFkTg6JWjGk70xxU6Pf0yiAyyKrT8ZLuLnJ/MrIXRS85BzqMZJLz7h+ZU6P2RK5RIarx12N
I7dp8CYrFst+0NmjZW4sq1/VmU2bdJB1tfN4ORtO0QZ1N5xR6kPmoyDSAFMrczhe3L1pe6tSzJE6
2Q4ILOEIlihPg3Qco+1mCWS+zehVk2719ruUL2+Wax/QfPhAI2+AbpnfM3DAQoZKnai75K90nzmi
tBqjCmBVYtqYDHtPhCG4iduxL2sUFMsoH4ndnV3Gb4XZ02NG8lSJBXM0nXkIgp7mX7LeXB+2hjAO
kl7/z3Zpe2Q0CkIKws8D0qVQm+BB+CS6uiuI4SnQQBXoBdj1PubDRHOHCMuprbkhsr/oMJ3WeiJw
TQjPL1dSap8m4mJwXpMCjD0vGLNqEmSIPNK2NaBN+flh3XNkw08/wYjhL64yw87Tb44YQNRWzmxC
cYbTEWCYvZhpYUnCtp58zYeqIurfIRhbCkqriZzPnoMMNTZu9lZM/P/D4NbeBTF1mIzAW2kX9URC
747VyNMhW2b6M6ZZ9tMzjSabZ4GKQ6CO7yGtycrNtE2oNWOj/JQE3L4sNbZvcPdGLsHqX4DMcSJk
M6448bgWDUwsVC0YXY9XQ0Ukzd8hRzzV7x8JPVzG6iyyVXu1VkIqwRD/SSh5+5U7PTtcdpF4bCfq
TpZ91uMyiVzkJScv6HYrm/wU8aEke1U7ctIMW0NcGnAS56Z3y+Sz3aELbPSBwOr8N2tyPKCUz6QD
0mwiMpTlZg2+kDg7ToRNlZY7FECrcObG2ov1GIiMkr/Ly3hSNItF5dHL2d5C8oUYQzk1tFCVbNR6
DKJ9fN+9HY1A+9ryXfhDdtYAIPLPZbGlWGUGaCi6In2y2HBJqqdZD+zfIqpMjygKaLPCaHGvtp2w
bEeyjgcdCcHMNZf0iJKcy63fn8J1kFUbnewO4LXAyAo70SAfTL+bsZUaqRwe/k/h5EPLEu2mT8UW
aU6OCIuC/WmL/hlJwXbQCS0L4ws2fgCUJo8ek5vu30M1nJ3ubix7FlCuH0Bp54Z4ZAWJs8jYILuc
npKcBUleosWcTE24Ewmfym0a86KXl3enaLSUj0K5ue8qN5JduTmarVtOm/phnbt1gN/AoFjdlVtK
HlJX5ZGiA1b3n8xHy+18LaqBlgYnIhH8fKIe8sk/I+o7u13KWHovoDnrOFSEEds0tm75m6I2DpGa
4bOuFByUK6GcVZoHpf3L+IM2axMzzE4762EC+wj5WHRboCHqwzyXlhty+eYXzliUN8aHUxobXj4F
f4hZVIBJrFUH9LfQMmKOczdAuDC1+sH8ZXTwBm0CX5tTJEpXu5lKWujBDZo8+eZlJLPIy4aQ0qYS
mG9tF9zsAi3MiHv0SfywoZXVThyx8XjzV99FF4EsrTCkXrI6zE6uIrUhrXhbvq3e5D6s0g7a4s4C
mUHKWAzEYOuTSZ6Waj7oO0LNFznBLbSAFBDyJAiV5XF8cg//UIAgMQt+iY+VP253s2YbUCefmjlI
socIA38qC6WJh/yPdiGjxubBy3SDIcaoXOeqdY/EOtRaLF4un4jKtYAeKotyCmMXjneEjoDgk5nt
Zf6W54nqMLGg43BAE4BJzDEc871W8/0nLjtgXSZikEnEawnjO9tziMeQloxjJJE4X54AerLpdyPW
aL/JaQ+dsAchhBuI+KD+KbxOuB6DO083pAZ4Hw7X5TWYPkAIxBanavbjC4tgdsE8m0tF/j0oXPct
WDKUllj7IoNWLW01pgHr6AciCTBhoIyF+PjD6+aplSbGzH29TElvvS7l09PArb9aTcHOLS5QwV6m
ZG4OJaiAXomqK2qrpOBDg9jr4JMQ8lsUrC+cPvEAnfBr7ZOBgS0iQDhUm9/fMWHjIm38d8VkaYRh
Gm0BmPAvE0AlbrIJvaVa6mN+/kEf1GDugMrQ6WjTgqRcI5eTH5zD4ujEQ1K+RP/HFQTSrshlJSZD
+XTXAb0Lf0PaRWXky1G0beFWvwtldd4KjYYnZuETFDuErfMRDg7gbtYugSPPNCoRHWnavXRGG3iS
fvGAWnnu1mvzYgRiIj2wAHPKzNMDBwcyLE4tLJoQMRe/RhY/mx8bHtQ4lxRYc7qDuU3b5R14aCKh
0emX8H7C64x7WNEYL685LqA4ILeqZm7unSjCwiPP8odDom9Jzx71pAKS5IhQ7dzbkmyBQ86PRpS0
jcPMYfZlvU+jkH04ntWr3MsOkh2M1hpGRJkq8w0sGmmPolUyYcWO24groTz2Yqnm1g8PTM2TAMh8
irivhBalrZeW05AOqa7mu49OBPBF0fjIwb2g62C2ptYIcet/pl34ill0aySfGccQXhfp5AqJ0R7C
XOQLafLvpF6iSm4vkymMspzcrgwhkYO2AJDAkS4hhBSeXAIMSy+5mUtiN+NTOGwDKCy40JU8kgVz
Aqoe+uV8zVZnhOUbc9ue1KwWQ7W9FxbUMENkK8Jkgi33W0xCI6nOWCw+QVzdudc/8ZDgnPzSHPBm
C5beNUNXJrQtfURvmdP8LPBIki5nd+mNhiplqEswRzKDpaiQRWo1cz2yE44Tqmf/hoRkvsgDXUc4
gexkUXvAGErofu28AP4ZVuugPJSLDhIDexVBoIfkmSII6yrELI+sGhLd00LCj7IfLCIZkzPDi/AT
TTg6k+QEojzMWEw3SVoBKgIMm4A+A5k1T8z7Y5Cq6SKvdy8QP+McVdXkLqNwuqyfiCGJWM2pWjVj
IG7ZUQKc+aG7CH9AvjBIU0Diz2IoVBYVotbPmbOr7kMVZmMUA40Z3lUuFwyyz0KMhpCsi4j59ijv
bESaz8qEaJbUUwRIUQit90isJhBs3lKGeHkgAQo+UQb77Ib614Uah3qEUCbnizpgaY9TWt74Zpab
rRZEEQcWyWUNWI8DxuiH+YFC0Bcdf/hafMeuZ8bNmeucV8IA8JErrtj9LMyjVrsYm/KuPu7jy/DV
FkYRCub/0ctvSQfQSJfZrl0q2Y2E3FmJYUUo2Gb+T9OvVHnqEmrluBxcgAziyLfnOBEcllMJVzoD
tSsWKKdd0q7h9rHRRGylzr7GRctjbp70MhR+7UMhCnmGmCuGDmj7EHbbyoHQmHZ2ryhGpbs+yaml
b7ZgzdlvOqiPhr4TvBxnQEByCZsWYhSiyoC97ujPOL6f9QLOqH20ao5SBtZpz3aN3d3vx9GQkxOr
xSQek1xQXrKjVaE3RjpSoGF4HzCW4Ke44MDZgAHXPbkPe8hPj9w+1YmNOIoRZAFtW3qpGhCVV9Jp
OCuYgZ9PfDvm5iKnfDlBlNIPBdg3TZtQV6hW4eB2o3IyW921Fmsb0sXYJz/KhYBbgsaiFeJ9fEG1
O/6au+Td3l+XwgW5mUJK3bd1PrQMfKTkuCyGsv6uTSxlim1nRADdo//5XvXn8tylKAg3wsVx6x5C
MDnCJCyIkRclm3ZL0qydsJ2gWGQ/YPD47FdCyIMf7t3VGgXjYnmDAyKo1eQ9I8h9aSgWCd493SgZ
1H5KG5uHlU/++5BW2L/Y7Vi8zC1J4jQ+3YOzXBSl3s1vOl2z087lp/6FtHfYhN6z1BabTuGmOSwg
J5fOH77xpQCQJvoWLXHG0ls+/nHLiL0HWURm0O8XbhQ6EpxMZuJxGyB4SAK3ok4LzaTFPGG4lW6H
K/7hPrURJ/uJOnmA0Zk7alyuj1SrrpnkGTNhJWGC9HxWkn5HsbyGUNGYBTAWdEEtpDpDrmE3lEM2
mHw4sCtxGNTf60RtkIKXJVz7z0bx9gdDTkKyHPwWUT/6+20He7M+eSaOCbFcnpLIYLhLH6RkHvsB
EYtrEBWE89kYpA8ZmZWZwZj8HqpxFBC+77QQbnh5GcCGRFYK4Y5fEj+Er7m0TkPb6Uz4M0B/CvD3
azbSJdERr97BpwQ6P3ehIrIz0eOlCqxg86y5T49b5kIgA5v7ouu1irDny4H0Ex848fHBdHeRartG
WQcrJYrpboK/2Vy9W0R064iE9F/oR4f2zGx3aArotw5K40EOGbVbRRt+dW0OirhnoGHIql88z88F
kNCiS+Kj+cjNBOZOjHlPhJ6H99oAunqM5Brs8earwNYra6vj2g+r3NlqSQDY99QClXno1SHDYuOM
RSzMIb3T22GnMKz4qpjEf9Vp4UefaKOTr+D8u8VBcj8k6c311WgyPmhfdMCExcdeW4NDGmBG0+Y8
AOv2RqBtGLCJ8mDOXojRp7LxrqPGu6ReuJuOniCkBHaVbQDchrKzK3E5rtElPMEDsFqqlQGxAE2W
xqpT03nyzEqquFoTDoxHWJS56r3bIBDcWXrx7uNOiXKe78B6iyFgu7olSDXMS6aqZ57dNbE/O23X
Gn+RriSBZlNpnlYdXrmTDrwAYaSpMPgZpxWSE5cKuP+zovDQhH09RY6LOc0QoRO5H/fr3NMFLGW9
2ePGm/bS1Dpvl5oh/PpfhUUwHHqkjktgmg0SOckahVC9FAtI7fmhKalm76bzvWh9PXXfQ0lMAF8e
pN2QU975ACOfgt7jXF3iQKL8s26TtF9LjeLZviJ/04/P47B7M0Pu9WdJz3bfHfG7E//3j6F9QZqF
gs2QhjkGWne4Gr3WukWPlUBJf+Q9u3iLXWpwB3jKj4AAWfpnehAjy12X6kqY9WfzBBPb6Abo34Ct
71AlkLCt+itmxTq3u+azogReNIqYZYk379HLT1IJIq9t78rbIc/yB/WpKuFSexOdhhGwpn0pOGbr
7v1T75d8SkOQopYjmT2WMAVGuZOdRtoe6IrBkry/rBinW3ds87jtcnAw3Tu7G1l7bFDwfCRhh3xW
erpff76tHjGW3LJxtGFQuqOA/f3ee8GXMaXVahGqyrrUOYiV4u1gGPOnJKuR2rp31dhV20G59kom
/J561lMeVIOHha8Om5Tt3zn7IdE1h1BspE375x1V/uKi58xKtg/+NSrg9dOyL5o1ZKNchRwVEdY4
7DTU0y04IyCLtcWflvmdC87jdq66sixk0xELQ47eJRNcy3+Bv7KVeiDu0LRiQlpVJLiAmezfSAHo
yFCxzsP4sSTJ+5CMBWd+LSyg290fpBA3Go84ujqHen4oKuoQ1tcLDbKqul+VbJrYX9YMMZDgCuto
j+33QmA1F5FF7qXAlOPb+HizXoabq1bp7B56l9dExdKllpqIbIozVHzqg3ZJXgZratl0id+piDmx
hFpiixn97HA9bsnEHDQixRf0hHhWEkMbOn+N//XdQJKAlF/t2OfNh2nEi96lnaJXvE7sapoZa4Og
qN1aiLL0lwABf7HoFBA+4HHlqzBwcpS9kw/KNMLoFZgzGBCEvzLhcl1zJeIqLwUBnix82WjF6czv
p+9ALxxXHo2INBfQ5wTsu7it60GtnQUp43kjn/nBo/A3bj/3iZWFmjqVQumY3xHK1dGBL9MEF0TP
eKd7HeSnQB8bsQfoohE4j1SwtAM79WH0Ka3gcLsLrHge9vs5Mi3FtkLk95+4VK+ls/W5IWL9ppxg
pEQVWd/wXBwe3r7UimaF6qXtPAIOxqbEIHby0LeDqfFBqmq2laSjgeV20FvXDjdiMBDms+nS5/qK
G3J/bfAaf0Q71Ko8W9neFjR+ty2o5cy07hkvYl+J/i78surPNA3inS+tbIdnanc2DWjjs8scVTRK
XJYNFH8rSrulYRJS6OpH745CpnxS1tMrbrv8ROaN1luqs/l6mqbyJgEGUQqZ+xD+VctvVTsk2JZs
d8p+XoBQgiZI5+sUr2IP4T0n6ATk4tHJappkZVNZum4fUbEW3NNphmUYavGNfMyZE1cN9gQshVV6
UajdiJvrhUBKNB89vnP2OfmbUsj1kRrlNPpNlcX13XgTc0bUo2+tWnjNQaFh5rAH0qoNEdj3D+d8
AsXghcf1GiZXSCUobwyYU87kEFNo+4mg8vH4+3Z/CbNtSmMFxclvZB67hJrTUgo5WOyj1nvGGDFJ
WAanwVKAy4ToUqElQG+f8uHtT448bSqFrJoV3m7z2cRf02jo6Lo6JHAzLhPG8gSArH61cduIvL9h
xROv16BCH/eHpzu+UHJ0J1TNUIcLqJplbE5C0JtJoa9OVccIuSOG4lStoA7sE/B+4xtcvMsSr7Py
HlJQ/dtsFpHGfSHLt8Xj66TrG51lRE/SMj5vruvY9jgQWAemHRHhRr6i5T5OCEOy3DUV/0ofktRE
9XI0tcuKJ7cmk13Tzoi/d2wVGkjrn27BDGeF/hN17tigGadmDwyvDYlBk8UBQLewLICPBR9SfGBQ
y0vJRmoP19XIKub8Tn/wVMbHv6PmOtbjq1P3WlOPiaOnfwaEzV78Au3VNz218fLE6QFMeAG14sL1
9xVq2S16Z5RO3PNB4Rob9n4/UPQxefVYvvgHSzL2XBi0oNfm57WDgWszovEzVKcSmIR5tv6stCgJ
w8uZgqLyAixCyRAZQenzwmFQm23noRY+44yEJegx15JfJIWsvePeqMQqbRgTWemoQjBBbPIx/+gR
zNLrQ1yngFE0d3LBa4HlNX01GQLdUmbp+4TtAlnEwpqpoGOL/4bapvQMXWmi8sdLhNPtmZ/9vpyr
8FvIWwhI0Hn+ftf9iK+uRP/QxNh46nRplUKESd04BB+ohsdygHNEEP3jBC+fFr47y/dBomaoLIXR
bMTvCw+yYZZpEJd4eUeVEpjtnFXGHEGeqvH16CBA9lklRP1NFh1+UU0lQ+LcPc7kXR8KjP7MLyaB
m/ipLNzhpEIektXADeMv0GVphN9wEMIYpkLuIExEu2dgKxPvPaZTcLJJFykUEQOZQFxfdsa8KcIT
VfS/AxWR0i1XTx82BCqWohvx6tsMDGo971wA8/HAzvXhonzI73jESQVjP+lBrUqCLG2UblyaUVdd
D9KejUs/dtK8ICEmXGh0XDyBq/rM8LB8nvPkmQBzLbmLzLfFPWl2B5ArB7kVPmfvIpTmal0Kmk0M
YkJ+kXIGoj+85VNz8yWuZrM8yAtNSWXcOvL+eKCvH7wKLcXxInkYnZxDPKXw1kcd4SHlTf10Dsf4
Ty3ck/W1uPl2HRTDxgTszEmiVZJ6H0dJlcH0wYrXWMx5op4VUr6bkQwqbqJNlgZ++9aB3rzUq2Bl
wThA+64wGD0awuTjRCXFgVwIYozQ+D0x+H03EJZRUqya66dDKa6mY2Ripo5Tt0Oud/G9FY3aF9Z1
r6+YcGJdlDhQUcLsA4nFwfTRa0818gqJ4icZAtPU3O9TVS6ifAVOtMtZ7HJhvw8rSlE/PhHYjotu
USfM1Uncjxtw0BKCz5OrkBjO0suXLiYO3mEzC14WD+fEN+1RbbSO0nyYJWkflIkmWKGb0MQHq8QX
/DAxmKX//WlViOSsKKn5Ek82xfdfJ/nlVk2+kP/yJHlOIlLBMU+enfY3lnGyAc7iAgHyfxqzDKp2
2umsCrUqiYc6Xy53O4WPvPuslsQGx8w/OUI5BenNg4BkUSRXAMjS9ctsmgw2NNoTucOQkbF4DGh9
20AVYdmJfbKZBuA22pX487hMfpHn6TyOEw91Ny1IAnMvNj1BvLXmyOLIr4fshwwRVUa8iy6Bg/8k
k8VO0xziyEFgFl8RHSk4veouZNaVGCsUf5N899T7u3Mrb1IcJKzJbifX6E6LgHyCkGYBM/t7ktu2
JIoKmuW0wzX1xN7OTsdDk56ykxzJFyylIEwaTNZ8383s+hwKRtq15CJxIayOJQTnqoiAuLGSh2ug
wCyraK1p2BnfR0nFX59z0TzQESXXt5ykBzRW3AE3iz7ISxaeZspma2yIksT3NdydKOZUVxjSLSRB
wgyO46eXMHIGvNaDKqICq6VcbFyHGL+Dhfj3ETJhgwt2OZyRG0ASMzZqD6kJqen2J0jJ0U/ayn6G
kB0MCFbJVa8Bffvqx3PQFNoUYpyfOMo4yvp3Z8hRTm0jUByjCp1QpjJrq/DrB9CUJgJWMglmyeTN
ClHt077FI9Plek4RFEO/SNkiChnJElqYw830Tx/FZe21jFZOK2bG64PyhFLVPaYHhhaGDCkJ7hib
cpTBMeUUpQBYd037W1oTTvJcZSExt3JHpV6qDfGigLo/L4rdQbpSb3czyLqWOkIJBgMCzDEua34B
/AdJC9bpVag3g8gPJoQInxaHUY8a8HzDlzIkFSJQnEI8lT+n1GEnu84UoF0/Dxa+S63B2Z5t+A3q
KgYxwmwSqOcwi0P5MS5IFPByVYxqXTERdKnEzWgxf6p927kbs9N9HZnaV6YMPBLLyJZ30Tw9jp/3
2LCKtOQ/CB+ape6VtRpZs0S7/GYLbpFdKdvKfVKaNfFagvRmI6UfQIPEghqKjyLfF8jbH+fyp/nT
gFQsqrgi0k3cs9RR+chqY3bSaNkjPAdY0SIGA/TFO3h0kGvHJydf6gBB+LzHuI7vET8fj7nHdhNQ
LAsNCQ3B5VFIgnp4/stLoofFp2kRO1upR6ZlSqDXAIx2ogRwPq4+eSa55W5FQYOnqoAtl4cM88CP
PhjdcVJrzth5mWHGtzGBi3G0ib9WtZodFO0WTFE2qZAl1ggBX2GTgNCuupfKi68kwTXGiXToxh7B
csAiu0SC7rgDm62ud8n2P5N4JFY+wrwjCZkXgjaBDhFILNb2FKloQ6jR1sp07VIDPJUpxCcO6f+0
pBSQdrKkQfnGOBYWCzuHkdxZWfW4frvyibzLOG43RTZIiANUoXcd7Me9tsnPfuMaVo2zPQNTjqcA
jDBGz2XqsndaSLGoaoPXmFmvsSHaYVbrZ8P1wtgh5oWuCVHmqgeGHzSMs7uLGS+l56cl6zQwgl8I
pAuMpvMHWqiMHPLSbrkxyg0DeqL0JOCJy2pVjwosWR3n5xihld5e2VhGAyrSuFA9d/0TCPi+zpzw
yg7UhOFJJ51zGl4gf4ZOM4oqLJTwUuPNkD8TIsyGgJ+FZHvjUID+KzvcRysUCJsDzJR2bUkl+EIS
8Oowf4z8IYuKGELSAlKR0z4kV26Zi6/fHidbdxB5MMaOlQCj0B8Qke3xYjeSy4kBfcOZIwqcwGPK
sXB8Th4DKWNzgO6wfDh1a/NHqpw1DRVAlqfYv8e5C2/TYDwuY14sPGu8DYdNFuHIj229IG6r1DlH
dNlWhjSY/0oUztH/m5CrRVR2QwSAvtIqyFSQ7e1fJcwbFYULmJTSRawgcc4BUeiRP0kvVC87WytF
AjuoFdF74YVadUKBwzE7fPp6M7/CrBgvA0MEMkoKzeMLooPXMM3TdlIOO7GC49qCXrzFS612ve0S
n93jEIDLsEi29yVPt9XRvbkdqwySH3IfbB6yd8DQ01S39l8h/wNsjEO6z5X84nxNrrG5rVbQfbqi
gdiJcNJ04xMdm/zEMBDfOV0jIIkB9Jd3csuESTfmBLWU4w2ecL61TnXgaU5HtjCoxRH9ZcBLoR15
wo+kbaOesZgKhxhrV/LLtVpdz1jF7SG6cpr0EmvDXhhcKwR735I4A262Vrd3EW8rk2D7kqSFwYGJ
1TJZ3Zu2C0WVKLXlC9vd7e2/rwQGnJBFvIiBAFHqdsKBOeL+6U3bdcHnqoRCXzvCrqX+wEY5bmke
tL1lUsV6AUMgbV3/uSvgxhvEuR1HYIKvKUH4Tn0TcugIjyFdSZjbKNPYo9KjwlxZA6ozdr/t5Pga
ucG6+A79Qx1LnZQDoouek77C0VoL4rdNmwaZtOOP4z0aN/rJwFah6WOyP7nqNP1zx7IzLLI7vTHh
o2KsTqzmHfBZrxC2R5mTaTMDbpK4TDhg5bXeg5emUW2um2Cfmb1lZWY6VzlJqBsipOrgZNgdgT0t
qOvrU8EKu/g9HJVoPwoccnywnTRxml1oy3QlUUIhfYiI8cUa1Uwl2iTAXkqZ45v4lxp1pJ5nDVPU
AnNC/ex0d2+tjLIkeC3FXoYIbhFB/H5QvB1UnGZGk95g5+qOV+YMjNzov0aor8pUxsI9HnEANAaq
yZ2+zpQay/PtH0fX4W6B8bhpspTGwU/Jnf7Ib3COPed4IDumavvC19Vf3nwNFWnm+JIIEFBAfamQ
Ehmu6NBhOQzDtJD0CgioH3raPpSoXqS9yNHyaQNj3L1oZRuOtOSOJC8tpoZ4FmSvCLhHKNsNBeai
coVdEP/GF/y3f9zKn+C0/yV9LJVG/g+XHvsVgfSf0pyUzJR8SW7bEaSvQUAbcF4EafoX46PwE11J
yoGbQP2ZKUlIw81Gle7yQhb/ulNmr7P+UwSeavvooEtnX0xYnNtkUTaA6LB2pCYa+FgeEaN7/mbj
hkCrqrjqfAggP+kA1EyZ118vGFCh+l2EsVtOx/uoU9PE0U9esbzgqd3JdSsGlX2uEWVlxxY1Hu8y
lz74IIAED7mtw5Sugxq579zEk/gdK8Q4EvnSTbLuUvgPR8mh8YNqC0zPzbsvPMDo3mu5ScwFU5bn
zdzGsHJ3NHp37FOlh+Kn6cohdrP71h/D/X3DSNO0P71qd6oF73dGWa/8JJNlbb1pIY/dJEhtpESV
TiwzA7NZS+vqwvd4e+GduT9iQDEjy4lFmotCGBipJHaQvQo72KSR5QHgSxZRcioB11rhaoBglfx6
ctDXjn7Msd+51bWokAfHE3IuE0xoLxpeDNq3JE6T3XZ492gg1bmS/dRQRyHk2RjE3s6wz5VctfEl
2CiEz7rm+b1HijF/4sQ9NJvenjoqkhYj2Sc2imRad1XN3sxRlXZUH3BXFhPXcAovKxKDlbGLW5CT
MjwKt0SsBfRwgBJSDuIpmt1S6woYqYMl7O+pmN4WBZEpzrl2XJ4/pIcxPNF1OFfa6vxE43BsQ4iz
daMwAy+oT9gZ9U21ScAzZ97hprnr7PiQPj4ScRJEg8wHoki4yMSmq7QpChXySpsgcg2UdrcaijRo
SRFYEuNuWpNBr0Xzx5C2mSUle7q4R8XODZjbHhx4uw0ihrPZ8ik4rCPCSysLWB+krWLLUg1Mlgmu
CBpWvLhCkqTpi130vpnd8AbPertv4j67ntJyiNEXSkQu+Myemf4pZMaSZ911RS0XEfV2NYWJoaYp
H48EwV0196hNYNHORwS3mcf4/HBJehMcAXBY8Gcx2Ygpj6gUiV7daWy+6PlLUbnwPlyST7m5rnfh
C7n0kuX/vwlMxOs9x5DsBv9mY4R2TbIfAqEOsapU8og0tMefjWuKbhiJekAq303ar5+ros6Sy3pj
Zyjvaz/olhm2Fl1WDIvF/uzhbHSZNQ1lS1m7u6T+bbBuB9hddcmkpp8UtUDHG6DPisVFjG8o7y2Z
KWdUZNQKRXKZAg7EwC5IF5wi5GaSVBThKTEEuKGIjp3UEuNHYe7MFx4wL9sTMf/RXU/jqCaXRdh8
ujcbyokSls+G8c4ih0CMlH4DknBCFfo0/IFTiVmQ703fq1dReEszx2GwvgV0xO1+JlE7hgjbAHjG
XeNq4wM6ZTc9f7kWMdKu2Z/iBdy5efTY6I9jx/1fCEVfBBErybQJ3NtC0lszt6JNW9mkpVXmL02q
3X6DbFwlmAbdqoCaBqToOjdWraog9J3tGcjNBPRPJSxKovoTsaV9Mu+DO5dSDa62N4z0V3JCtugJ
XENuF7D9MYcqtemMqmwhDyGruYRUpOG6efdB2Rij2VKUUbVOv9smGNrbzZz4sksLgjGezXbdQdSV
ry5wMGm8ToBa3Nu7mAI1Vr3rX5WqLhJ2QlqXJtWiuCTO44aUPTPWZn1sN3XZm68IR94+JhqxQ8BE
6HInw/tenrCcXFdzkB01EP4S1a71GHca1N+4iN7+WCNHhPRNZEspr8/hpRJFhgIVlA1ZQinlGF4h
r2rP6StpIb17v8Uo6SUvYMEVJtN13MqMBeOGcAqXFxTl91jNnno6e2cijHVcQrF3QYNbF1tICARI
xUQi7lZ35c9zEdaLkZDsynf+v+H9gEzLT+yNWVoUzJcCJp4UduEUgxenWMGBlsyzVszitKX2ijPY
zzhqSWK5gmkYCmNkY9yBBnwe/rGsTCbnreir2hsEPhVgT6bNDfr6uaeHFdq194VjhEW9vdQE1u+O
S++2SHaersUA0SJN5y+alD4dmFUVPfei+aS+y7k5p/n3TQKTaRstkHyQktciyB1JgGe3mfT3NJwc
6yQaEnzkc3JkwaDFuaVlU4kM1BUMky3GUoXvvDH+WUh3HMCO0/Eubf9PaX+lZZD75guAPIADiUPy
MjTVmhsg6Y7zrXK8OlH7mYrM7xYVQ10EcHTeXIVnmI4YVRqy+d2RjlGlvrz8CAiLKNubPntcWL9a
WfWEG/xz0slnUahWSCko7eRm5WqWBPFqi/iRwWr3n0Jqd9yVXAzmlTa19PsysFCP2lbSc+0NbKSx
I9FXURhw03RzYtiFEQqV7VmdxjGhw2Iifpl8VGr2uwC6gn1tPyr7FQk2xiHZe3OSzZXxG4EtudJv
a9iYBaiwGDN8t6FfSk2J3Ji+68vIsKz8wo7N0S1pCDuYbHacaam+msqXCaChmuYmhfOZhEKnUuMi
JJ1oadkJG+qIskA9zIjmf57pZBSD0Dkbj5yGGLs6Thfc6RHf/WvxBjvrATbK5zwaWWNHe0cDr4AW
t4cy0jjkdxplR4n0lep+0shnGagH+ISNo2OSw84W+pBT+oK1EK9NAPet1uxH9DQt8F5r+yxDNBJM
j0UQD0PlFx4WNAxz21V0zdr3CUViJ9ZpswwkfFrmVjQoMcct1m4NNCOv27osOqbbyoiP18ptpBA1
RerkxP1GWw7rC/jnQTS+6013NFJez2lFdA44CRcTwSZmItHtX8nz4kqyY1lqbGfj+Av9YTsO4X2h
qmio5ohUufo1VllachruJkwSdsYLfgIVfzQ4jx1DWl8HCwG76Jc9R4mEShYY9+2DJfc0NAepF+9N
gesz0TD5vIpLdDfRaC6RAMRY9AG5JrKHx51OgXYydpEUfjzGcZGe8dhQjf4Re6bedr6ipwoYblTd
Lm+QnzAQUJjTTSxvVI46+wbY2P1bR1JVkyXaJqW1bBr/LkEk/D1+ffSDUKiUORXV4Gas70BRXECc
g8vwiB7a6s8wbvZlfvRsUWF5x4g6hEump1qzSYIlWlhwnJHDRYXzbN6OBG19iOQDLwXefZ9bxObI
Y4K3HX3wdd2juKgWoMIOfoEoICGPFC4I00garAljYIQ02QR6fZ0k1/Yv68eNJj8uxabDkH9ZYn86
0bBfVDLPp50eeEgFRpBbg3M8pif9ghuw9mpynE5StVFM/Y2CFTn9ZMnmjJ+Wmkry0FwoTwwyIlbH
832d5Xl9hw3IJiwGCI4gPmJ4kK0/s5WttNJhLfYj/Ovm+x3nyyk4j2Ey1bWSTRpMvXYslP/XV0aw
XmsveeMtVFqRsVPjOCmiL1kZrlAjt2Ds8ZJTkmw+Gq/4w1Mbs/vlmOw/N8OeODPbHoqRapL+KgTv
tM9Hlcv0mkrzrB302Rnw81+JK6brz6HFdqf6G3nqGYCwqQKyq2bBbDFBTArhw9CNFMDT0fasi5kJ
A9vT/VpkFCvsKcRgjffTDqSt/l1Yo2MjKxjQ9jaY0BFsktUQtKGzCxHEAfocbA+hptFb1bctS8p3
qvJOiVGM6O5g32Y16K2MT3z7bEP1NPf10VUiC+I08XUo/v72C5oUUd+0j3D4XdThz1voDpzl8TOm
W/qfURW1bleZPJh3rNOIyPR+1rW7nzI8tHBNzsuR9V/mLeY1VWyeS1XxWk0rkq7++PSMAbEqRY3F
/xCcdiOwMPAMznk7bG9uwZXpIrGIXmzEjW5SDrhxs8WbXeiEppvFQfh6pnWp9Morw0EiojoNE5mf
+1efAOn1IhB8Y8BTHL28jDdR1TlEkSHrYC55QiCc3MsgsnwEx9C+ERnHFF20V7aOEizk5nbDhTOy
kZnxvD51KET0SqyfYcjDURq6mJ71mFPi2+09+VoN6pvIZ32A8XuhJaqsdvB9HfQFSDxUlCVOtfn0
aReCwWRN8bXbdHWFWfQtnqJvDAFEWotJ7Yr/8h+yqg9tsUVUHx1aFnOZ9MWCYyeQ6MQadY54R166
V5l2LoYB4bGiDU+GXD+KrzXpqG2v6Czf79n+tCfcP2Fr+d/0t8JgJ/luTwcMcL1TQdZv8ZyLMwlz
LJoGCz9MjwIWohZGhx7IM6eFj7W84RjK7j5p62ozF21lzjo1aBPL+NigJRNo7YUO1+98/CRHkq34
LSnWD4JJ+R79jvkrGNuOAuurHtRJ7fAgmToiIh2dmml2mBes8hMGPWoJMY7BN2vVKlLgxA6OD7i+
E4JbXZs90mqEjJ0cMmJOozeYTM7Ia79XjkjNpcSIH1HUDBQZ6CD14yAGuNI76XU5D9K3pEV8upaX
MSNoJ3gBEJnMRUpxMh6SqtEL9WkE6s049pI6otZwek6+tJUzJMGqAw87wUCmH2q6vOP8i3OgxeOB
moh1xwjWJthdYbB81fMXrwnWBXcDeMkt8dkpUzfPXuTUBSz7MeK4UkanhpqlqcIVVRg5g0H55EVj
3LdKssXQIr4NrYR5RDNlSqORl3L60Ogyz/riDRFw5C3ELmtNxuGemtZfPYzdhnejHAaFUPapnpcV
7sBOkdY5mxGRUkZr/O4LCQWu7uGSM1TwQ5MroJR0l+rmvGCY115KaPoOhT35P/kd2UY5qpfzQKtP
5sxzARyHBRAymTDwsNxOkvVrw8+i7yJmG9I99MhFqmc7Ich+N9bZ7xRJF/JicuHQvMfBmBPdcJ7R
+BmParILzfY2PtyV/dXmR2ilLxaum3bVrWOLY8weES9tf6Orj+pRMslMucDxTPeuIoRVgxstsbws
ljNFkguHs5GVKRaq+nL5BfbMXe7+iWjhieBw18raM61UFtyowRmlbXhjvbpdJ83s6CuGvcOvK+ar
mRuwZU39Ba6kZxDSsJuqJLZw0s1Xwk7xO90pEPzZqP/4Wtkv/JhsO5LguEOHBdv/H4nJpjNEMNhB
37qfcMEMjz9MZlQvad2dr3XCzxmNbERmF7q1ZkoqWKWlWHVgRY49rnaZM8Jgbxf6qR63nQy214yu
MDnA43EpjzZIYBwjQSjNDx/fqC17XrT58ljs3nJmikaukI6MzoLDDbslaODyKwqIih4IE3RNrWkT
MNDGrSFHEMlv0kzy78rXUjIoWb3WBPvHkqkXrLI6WkZGLGhFtSSiDdsdoOuc3TPpTiN1XC0m/+6M
OAwjn/3cfjqWym9CDYro3+eQg8H4VOaVcnbn6waWpFZO60LSfhzemVgW1hyvO9WLdVL5PMMVCo5F
aF10qB6ziHHV+qUQqY480tyikHBTDj1/tn3qwnILhjni9idehs4YeBoxW0lsLX4ZjCIeNWqfYqyw
cY1jMcHNHeHsUbKh1uSRDndxS/+FboSIwtNHm+IBc/TYS/DuI9O/oDftq1OkJw8PwUNCA9CiyC4Y
QK4Y2WtAQhfOccs1mCTLQ93lpaIcOOFfXQ6darM4hyZDFmAglIEVkcoHmQOUFxz5d4Cf02Mm4w2+
M8QRzpdey2RjtAN/vjBVwATH+nGHHBYK5zGIaIO/rZq9nvmYroAzf7/pcksoi+rWfReOe9kFMc00
3B2Ve8NGbt4WpRnRk6n96D/Zhd8i1RUv2JJoYuhlgGPyBnZWd87Zk3TAetGtpfltHSVi7mzQnWuT
pEhVKUsFrVuDscuh82+4bxOQLv8tSO6Yqh6+twXBr+Q8gkWpiFxGj5Ads+nMxudOoYo3Zyzh/Jtg
MG4ckxW1sKSYOD1Z1E6MkEqAo5pnW2aU8SCyycHvVUAQvM414pexxdb4aTBUjcyx+i2fcLo/5F2S
W0Il/D1yFdBS21mVuldduJ1oD0emYmu97MbCDVAqlehGaCt7AVBgb7U6/cRQZSbs8Xhv1WFX/Mry
yjWqL2Sd+/ulAPAtr53SKLsSnBlKYcZiBdwCPH52qwwqkpGsw0eX8I5KflVzRXywuXuMR0lPwbA6
DDfTWHuhwaYjxIGKIWgka99oOqch7fGFQ2TJSibsCoHmJXRqA2Q4qNtnfxdph3TnJhLdvbxBuuNs
cHnAyNB0H6qT3r/QvDOa/msybEwSphDhpJqy14nAGG9FKIpjEsVYdWInH0eV7jc5KNudvujeMn9T
aNiVxjdlHgwgSUUYaPI+fRMc7Df3WtEad0Q6Bl8weSknIPZj/lr2cVGz5UAZPbkmDIKsDHKcOZf9
45MC7f0dwrRATIAhFI1TJzNF2bApAbOtFYb9zEJ2JNQ4qMjXApZtYuuqrOCTRmbHe8L/knVAkyue
ELNcmBpt2LvBh5rkmH0r5ZMU/14CLepRGogPoZ4v/m9bE0wNQ/ItjGfknUogEucI2/HP+hqwO/NT
wu0CvizxGwVJEpdsr4+UaThGziRQsI0cPdBSYnDi37t3SyisMi7abjNaSniSNj94LUCiPmuhQwVj
lmU2bhrQUSFTfIAgTItFhalUSIvXzOf07JHnVkgs9N1ecf8n3nWTdBFcHzG/6yp0F6YWmnagK4l1
d7LJhKUuwEWr7dKyM8/7FAGw0T5h+vergHQLywsVJHk46ef7+jCYQvt58xy5i+PA5pcWKBpHMt5m
UJoZXjn+l7IImgkls+lE+EGnCqFiYdS9mhh1RnzgCvHFZHqjQiMsM0ED624MFQwOVWcV9YCzocxM
sKQ7xFIvPJjaKkriCd19Ws5OpUzFNp5J/sxG92LP5b8oSQcYBwGxbU4RwPjdx6TgyKs6qD2UVs0r
sgtnNrApYJkeN43THvovx6VBxfrB8bIHAmCPxej/OJhKwaYCCEigKES0Epa96aic/bqym2KsRwSW
1w+41v0L8BFAF/cVg3XxvlaS/3PyF8UTphy7hehqoZ5SOsoppovZhB7E3cGkr6ohULjkSsVTGplv
SVYumya+SshtVgsJoNl9IWt9X9ScOpZWMQ8IFhBm1DWGf4An3JIpu241sy3amI2LQNDY7COCiBx5
QkG69gZn+Rf9Ud94mXF3da7hNzPt7vR42w43AzPHVCBWH1e3bqFm/8sM0Jn4/rl/nYVkZS5d+Ece
CkSk5GT9bnARribxK4FLui1ewGzRR596v1u55knlmbhHquhs9gOUzOGnopvJYW3vZi8WyO3autzB
Q46QmMItl81Aw2kSdjtWnbwgbbCbCOa/cauexLhAV4mpHkhFFwmW5I/zS3HCIkT0+n0vfZhF9211
8ur3+129dQG14s/m8ts2PlvkXGAQ2DCKiREVDcedWRzDG8bkmttnCsjcZNTqqRC2VFN2PNY17LzX
Z2xymZGnCeo7Eea3IdyQ1r/xs+ncKJVZbHqMK3crGHSsrYoYBGtcKMX9jOfZfqLDHFU/i4ffq4Ef
yAIRB+c2S8ljWIWHCLVDYteSpZKpfwSC9i2AkbocUVMeLrgf3sYzBXpiZrcvVUdwnUUTonoSKK13
7KOX1kU29jeRplUig+uK8lOuX3D+tmIW8UcqeBhBsfrngzWMEQzWihO/anA43UCJXI1B4YSeE8Vw
+FO3UknhPWSzEcB6mSPWfbeXDkhNLAFnrsXe2nTxTSJuQHiMnPAymLtVJxX6XkRsLdFjhCNfcJL+
QLMvwiOHI3EfT0/dY4AhlccVx+U0jjEnkKLJdpDHIyOwlrjUcNvwS02LR8OJodBVn9Udv5gDEHHP
FfbQotnb5ynEME8zJ5vBVqXZSmGpic6Qe4iKOMpt7pLGny3SfdGCMjyPuzuPlKiewBB6iXIxD/D8
dwLmJWw1O2gl7SVQ4b3TO9n9m/u9Tq1vjyIUIiKvliIitQALuNcvZ9jX9gYHgJ8CteXQFLVI+V1A
M2A9M5hhT8eYtSkt5AUniyar+D1tT1U1ZlYc+qk5x3SR2EQctJCfHyqFj7rBBus87lnBSgRWC0/n
n/lpzihSqboh0i0e0zQK+uS2Yi3TqKy3pb1kTG04D/dYSI6q0GN0GJUyZnYb6OLb3aXtVP0Jbowu
CjVUR5FZpSo4U08BFieOE+VN58iD+eHuHNshrCsTEyEYqEPIcbjFOtcRGxRBgzWZGOBJZX/07/1D
MJ36eIpBqaBgh/6GcMWsDH0xatDJFzrBgrtK6nBlsY/szTduaVNwMsMlheLcVVPmulmP+kqdU/sI
bILkuO+rRcC+x9jpO4YiY1qYbePoFFzEm3dlE2oFVXenF2Je+I7Ft+bGvReQQRcLVEZ/C1pzTgCh
72Azwzm1GknoDatUXb5RIGwm59WvD5DtAf1LltJIrMZ0vygJSjJFvVZ2zzTYwDF/jVfvnqlvOD8l
HPGWsv5bCWk6ANZgygsyF2B6adaitZk7WUcqZS36cnj13b8Ey0wvaeGrcWbaEDDSyvErU3M+SLc3
Jd8D4rcEh2Go5bGgNo+mMyq0H4ZvnzzPLxR3RyY5logpxb/vQp05A3zNJIGwze755RCRPOYyNye4
3pC0e8O0BjuDZEWfDzDB4eQIuhEK3ClnSWLN1rx3C/tpjzbTVHdTwq1SqBnKcUDBG0xcGHd4ykYp
dLtJjjdufdhIeJUq0l/HB7jMxSA1G11baqE3Ytw4AWHnpAIxwXzuo0I+ub1GR+byx1nGh0n7UXYL
ap06NbQR+ypkb4tMOoosh5LZlq4tRUXzarRt1Wmlm3DtMDpdNtd+7bHkvRnVTfUl6zCgewftdZfU
xF0YOgAt9UZIjbciYuwCgn9Q0bWWZH4fsyQ6++q4HtmhI5rm9JwHZbtr6LV0U4BoZu2gKiDBL5So
z5msaLiFchH5CCZKzx16emy5Zx89GrL2HeuiYT1ha9kEmQ8D/cwTWC3xPegZFfIJzlDJc/hrh2ef
cJzF+TCKi640tH42SpbasJao26vrEvoVwt9vyP8sQdLRKmZHut122VSAiYD15TP5Ex93m9bupZ+Q
XY5V2Mh31Yl3fFKA2NPm5xRYl2GRnV4DzaVDPBPM6VvM5eRj0IWjH8TPhwwwd5c3LrrQLFUul5Nl
ltG4Rt3+TjFd1JmzkQFxh5azp1YiwJCTngzaOAgkVD1yAmUkjmrbqxiMTwVZzY5Uy7VZzd6fQcIh
0o5OSQU7AosaRRYYCSh8+jDEatALdA1pAjU+pR4QLUWwzLwk+iglb+FQvjlhJBw3gczj57IF9qQO
Mrbkid6jurqTn7Q7FAKdYxp4Xo8ls1ZeJbuMoLUm8mILU/iuGc6MyZX8Xk6xLhYMucd04O71d3Nq
GffB9Hv5rss12QZrI2oQp25ssYYjjW9ADe7nKjsgW9st227QNDhN/y+JiGF/+4wMcADri4RB/FJm
9wY/kKe4m1lsUyLS5QhfvgId9zFa7V7+i46Y5e7SRYWXv+eOMSg+l0AjaYRLSa172tSsSTn1DgSN
qI8OoppE2nfG45f4xfRf0DeH9njsONQgbuejZA/p7FPIGRmEFIbQ1LYiUPeehs9T40J5K87YZ+sp
Z9JVdzlg6Agdg03/wvK830AYigLWC9pRv+8imqLeJQUWmj9Qmn2A1WCZJ0IwbOHTAfLYYswoui0x
yAgeItO0OU5fMytwMXjIepl9Yy+EcYPzOGB5vYflo23Oz1uFLunpBJ3NPjoAnEFOlOGthkB/TmGc
CvHGWMXPxIPAqKhzCfTnDingrNJ2C2UiyDbEWu6hWFbIhLkP0+QGyLmLsSujx7v7Cokuu4xMp6DJ
H7uZXN8GYYm7zCWVINo5s25x8OzzoikkYbQ5/3UP8eg4qfUajQ8mPTdz5RAFdfxgMnB7lfYnkyFV
5o/ZPuC9iDuLde+kVeP/HnOaGp1+MerIbBshidoaaH1OwG9wnYxu2JuAgU3l1ekl4SuEX7JzQLkw
rKfWtlZ5c6QuCgGMNT4zYQnfDunQjik1jiJyGwNQO8JjZSU1n3POHonVF0soNxdl/LHoXCzzTV/D
5vQlyGGxE7f4h240DvpJL6FOTjlsE7xg2iO20j/xdLLdlCvYVxumRwUWCDbHGdarCR+XnjH381aQ
1lvodfHjt1FtzX+6vzFp7bEbb/oIpArmYJp3GLW2FZ8OkcjDPoxrrt+1ixR9q9wF/5tXEaWNQsOT
tWkqsGp62nsmJKcGLKxg1C6yuqKAE3w/Qn80BiOSxk36uqjxQcuKfZkMI9VB0JKYHc8AZi0GqiGM
hHBdEin55wfwDV/NIR9vntXyjLgrCLJlmnoPfHzibiG8Ye5pJ+GUv52isfDnH2ZO0J5LVmjXHs0/
ueQFaHkx3M6TmdXefDUJ7Fnb9Zsh2LG9ZMFHqDtPABSFSuk4OlJNbZcYVj5/H4GiDkhFsl5XL547
QI9BifLTymcbYWjV/wQn3ZfO5t0Af4wqDyspVw95t2xIn8oV/t5mG1hSJ98g48mWnaUvyG5MFlf2
EUCN+5V+lW5H++Zwqjukhl0vms/DcsZ24UWfTsd6/5YY6sOoofJrFE7/NyInxOw5Jb+2LTY8pbzp
qZJjPEJBqML5phuO+DwsKWXkcVdlCPZ/05tKezCxDNbhpkN0s8BqudTNFpXh9EgWPNapB+4G8ySL
sUA8LbyXZjF+8nQS7ur8UNpMb2yFykrIfQrank/zQ8GTXJ7a8V+OlSArRgWFYYMRounzbrQrJqbI
skdTQb/nkKb/Oe6TSeV2yBpq3lsrHIAsCdQ7CCOUR8ySqL8THqFzfydzpZz4OSzlcB7t7mr+Xj8H
AWhhh9VHGeEuUmqSltSnAWSBosWRsUniZpsxaI+EzE35Z7ngjKII2zlBgzdU7q5ujH2zv0UJZKEB
I3GReF3L0DNai/R7jeBg0TuZzOlqkVxBKu3kmcPKi2ugE7Bi56JpsU32Ijcw376aZ92rqn1jtVV+
luYNMPJ2zI79qTSxhzXiKOORCxfZgk35ZV0T+a4Mw47aFi14gTwIQq9WGUay50xKZO3YjlLWZT9m
6gxQW8s6/77+rpiAbi6FcO1F3E/K4Ivqp9Be3DRFlJ6rH1A79tQuS1Wud2tuOMI3kER1yufzAb1d
7v63/5B2/jNEiiSsLW3bDbkdvF/hIN8TB2iLGI0myFX7Qpuvt3G2Mf5CNFUbOKaJFDkiwooTPFeh
Q5aevTbSxdqb/8L3o7sc5VaWwi7lnifgInJbHuSfeBJ7TSTGPujKWJxFaETf5mly2Q/LEteKo8Zw
y1wPFzOEp6DMXY2zsxRxO5OdORa54el1rureE5puHAZlwZ9U53QvT1oIn3IGnwC+/RLaN3qqJ2C8
5x4sYj/HrhnpGbJ0+EL53KmriLXnXu27jcH56LsLuUQdNt+ZrI2fRGY0b6tgd2IzTB3WRgfxSgGT
ZCnw1elBcQpQ+DNtLCos9JATmGM+lmGToR0bY71p1Mhqr6LLDrvdBFNltKiRrGOdiMllB+e7dsJV
8NlY6/fTwV0S5p6z5iZicgqnU+9SbFqg2i0byjBU+tW/Pn0y3MJUhSxw/8bejqt03EAy55PVbKh7
7YQNnq8xQARoYKO43jpUbNcDXu3WwZssCkAaZWCUxlU9NXEkGL648FcN6LcQW1HDf8TWJ7Ytsyb3
6bjv2nE6m6N/1btxJtoYwkh71gOUZ0fxhLW63+NyucdDOoVkuPBUk4suCOOg4Uu4e8PfmaDGA5uY
15tWannazhVgMoHo5Xp1/wRcOjGtCFIeZu2dgUekqfFS/QUiRyndrCAWiKlXjPsB8SAiT5/by4kq
RHXBF5l3bATOMv87XahoD+S6h7ic/zHvE3yPH4lslhe8HM1X7RP8hrfFuFklgxbwIAQnA004H4dJ
o94iKO6uNKtRLvaPEUxvtotFnYDSP7wdVtCHS4pBTRnB1HsDFk6WCAMkMeRFrrHfhkArws4Vg3Qr
gypy1EhsP4EgTuX0PyxJvwC/IGKowb41jbvb9yRJqqQYi26FaCs+VNx+lNUd9u+YCL6W/mNtSHSR
0OXXDYIfjT4IdVuXA+cNjBIMbGxGXR37jlzxyYHMb6L7Qab4sq9y54toKDXE770PAulQFqUAV61z
HOh/l819gpN35zjAJIvV2XGwaRK0oaylBI9EUIUdkWS9tKiGdiGbDfLVywwpL5lWH354IBXZsmyS
Z2xgnF0M1OUEv8qNCt2brXtb5O9Y2LLlYbf4CZxipB/jjX3WyjlePgYTUY9EX1cOGe7NFRpweXyj
1U2KQvLKdguzG89lta3Duix8WQu4wGjMBPTyaoa9Ydso8xLpc00rVZnRPxhnWbUSC0QQqRLFORFW
PJUm4dd2ajRAqjAb7124Gv2/EERKw7lU79asI34bVyy/snorxodMSlZLiWUlmB0ArgiXow+jhHHR
Leicudb1DyiZPITB5zV/8wzgy5tAercl898pytPYfb2X/itazDnEpYHXIBCsrNi2sPenIFvpUem9
nuL3ryoT/MbXozODgko/pC2mO3s+3nsBk1hDqDbIE0MdUe16H9ABZe72nH8Owrk/7fSynElijo/5
vAoPtuDPV4hx2jhkfH4P1bbl5yb9XS6jvH9KS779IR6261fDHRhSyInsAVUIFXYtTwFnVl8ECyky
VZrmnBBoxd5fxyJncWCxI6lImriRmFw5L1i0frfPM5Lx6xD296rKtPKrWBbotYcEdzcjNF8Evv+C
ytRhsUCyRlWKrhX47CTKwGnJF4wiapaTbIP8QCwkMurkWV/29dEcs158PSQ4RrUNU9ELd9ZUIl57
UNdCfK5I1M4ifoiQS8JAHc8Fx1wDP9DEKit8kdNIWN3qPzRxfN0nPK7cdeze3qmOZw0EXXdydDcQ
4Jh4cr0GB+bKEtJ4EqArTVL3Lv94SUNtpLd+ZIHRhHl+gbokUP1xvbEhWDuG6cvqoakaDIcq0tjb
+P+AFH300RrdhNsFeURECtxSkILlmY5huuMMLsi0ZHrG5HLBuAS4asCRQwIww/HaenMzSd4se2KN
kkAsMyK50L3HQWQYHcClta8ylwttupxah2xVH9b68AN+ExauQSFRcfa78hTRpFbVKZq0V06QCCle
USVwxJUbZ6M8ezipO+VywLaYDdmMSM2+OeFXIbfLMFv4huMGxyBb4SInQcihN0zOz+5oK/ibhOyj
WGmPn6sswDkA/JTeYzo1jd8PqkAxccxGwyM1jMVoc+1XnAnyJlmFPcB3PjltPd0qjz83KaK4EplS
Ea5Gpg3aFHJKcSZoPTkKinVubSld3sGMgaaD7Aqp+bRl8tGn9dnmWsFzU3Zkr7/82syojlPwySkW
npi0jKo4xHEwi+Rb5q+3NFuuvbQnEZKQKwB6fLOnQ11pK62eMhFvjwprDbJmNluHJ8dFF8hBZqRU
wLXxFueIPqSjRAeXzmMA7MH+v9ByiPNR8MDpJnhGj2PKHGwJNnniFTZtGhzmbE7Uo0jUKCTjtiCn
tfEqpccNVz7QPBnR0nySQ+2UPsTTy3RpZszGm9+b1v3+UHvxzuPXITGWF/roPLk+ffuhI+467RmF
deonXaWzAwpknFAYd83tM9GGXgYQqvK/GM/6k6byhW8iWCXKMjMeckXayigoLDZwGHlaV0Ew+tKQ
/OkfEzUpzZJo7U3Z1wCOYDZNZeeXpdawm5cl9GiWGkvxknov5i6PZ+igbX/XNPzv3NE+5lryWg1m
gXDZmpuZ0T5h6u/fPCj1h1qsyNzORC9a43F8VddkL7l/Juene8ICfAICjicfSqjp/Q1/e/BH0NVG
o4pNJRMPW6MoFGWLVSXBRIHadAxis4kqzFZbUFb/bOFTS0dSPf3I+rkCDt5G1InWwB+JhsMmsfTQ
omJJJ1AH0o2sf9k3YEycQuSZkixgt7m/4Mj+dQJlx988EBZEUDfCXeGXIDK6uuIQIl5gIJGGN9zN
ahy7P+HJKqWsR8B4xlgoW3uLEYI8i7lYejAl8xL6njCD750rJco+P2FlxIu89n7ZMb5qL44h2bHI
brbKQIC/4ENWctrUhSpA1souv9J37M5fquk8Gq0Tfd1ZZWNgAn+KYPHGrcK/7pW75XPN6HJCrLfo
FWd5+oKQ2Ft/4gwH+PlyKZ61ugj0oaBzEOE0VAl0cuJYrGWKx5KDhAEH/UnZfCttmQk8ZzKDLWFk
N50pCP2h4NXedtd6AgEjjy0JmC/SW/gUYDXPume7rig3GQzpXOhELADmVN8ErxqaUELV0kHhIXXa
AojAwpY1RDR0yPNzx5rDglz/eBjrjb8l0GGRLT9hq9CdoTIer6+qjsgA9L78PtXu2sK5Qnr/1E0U
RBNs9h9qyZt2Eqy05FFQ5O2uvER1HmURgAq2KX+4MVBlrO43ZqMhG5x4Kz3H2lgOwVYkHB4g9Yug
jTIUpPfc/xKhEjQ/0RN8V/q9G4Xh9Xo7OGLFuO9yasOkcmnCqkOC01lkTmZCtF/eQy0z6doQTpk0
3YtqksK7Vt6RzCGTfDDR/1dZSrhKwUMcCAvlNd1XwmbQMxmie0Wrsmtzbm09+MVODYeC/mx67nKz
gvvxe95HX9dhTymgLB3ThjwqDIKJdvsiTIR0u77LtSY6R10+XLIOcmE37cXkF/FYw9PnP0UVLlEc
qt6wuul26QTOnbwXCXIFd7Pe/aDKPuvbarG90xgCZ0v57gRMbPCIUxD6XfmV8ZccwA0RahkzNCEI
JwCqqYRc80dNRLZR21hLhFVReH4ZiVZtNZOsOZVzc7JxCGpgofCxrUNQEfCgSVn5xDzmLT+wvMO5
Gn5yIvNGfYbJcdmce75nafoN7xLb/u2/P1uMq72wArFfaWldXj06RPhe7Eps//r00+QXWtst5V3V
35wtqBBKtT0ACrXHCp/4FerA0ydsGccYcpCXOO2xdr4pJtwyCAbywIukHNKPzDOaXF9+pQx5AApV
4rTlfJK+dBqYRWaGfzvHRZ5MwZRASF2wWlQXht2pHZEu+7WBbX+CXfJzZaHDN5TY4gaeORM/bVme
8O2FIqWA54nOr3TQ/2LhM3If9rI+2M4pbkE0hsVh3awC1r6K2w1TlEmZnrcz9tbNPUJJV5csJEgK
WJnhXWm94xWq14KHtk3ilMC9LCXOr1UDhJ9LxU8BGochVVJCIYGKHTxoLyki/I+wmiisUJATY3o/
JB0N9ONkYLbKWmHXUHzPdGB5MyM2Fl7VAviEJkI/Iun+YGGy8T731BTUYgYatludTRgwwHS2PDLr
ADWNLokYtST7fZ5KUPFdsfVD9qRkuYJqXWI/xG8uuNeDA35qpBDrlHD+4VJlIMWAsAj1TwR+K42R
D/TmgEy9hnq0t+MsH+YySN5BgDo0NPkrBIfj7sLlh6umGpmoyKrSjvJts7XlFp4cp6XCqgwoITNo
P6Zx2LkUbiV328UKfF+gEFbewpMqiLi7TqkeodW7IrIGdOmXhzFO0Oh4C4jYsvqDngIOxzxWzh5o
eEYsCPsxkTxLg8avs4Tg9D8JJJCCT3xjidoyTp8Ms3XX/+QmmqQYjpoj5N2PnkqVC7YccV2BBTa4
FdhxTWSTs5EPtgYOQ+xeVF79gwalOQa7AaN5U7uzz/vcicHBLtZPre0kuXe2leJJCPLHN+dV1wIr
EudXFmJq/GE4PSIonF/mEPGgVPfUn4L9w25+KAkajhBUpgVb7PCNVmQ8JFvu5ptO+a83Z9ty0RRZ
oEuxemn0IbGEp5g4KE4kpjUxAQ0qM3Izk+zKeh/7O6Yfrb8SIolpAdXgyKg0l2wtAzyJftmCEtg3
XBWerWX4S9MyRrZjBsxpIdJxI5yx4GiquYp0bQ3LLdtvocCkoVmw9njFXf619+1iKvhBftuMJTB1
An3sRqBHfCqhhIdRzcPaUAiPdtfEeIjFaSnb86+0dVMfjIE5D02LwqU/UbeSSyKONC/cIZAPv6g6
4AhWVM9Q6yFTuKKFBFvqXQx85Mn2ZsBvEik32ZophD11MI6VP/TNZVzP5JpQQlfJ/5+E3jeSpvFj
PRsQq246hTAOKWcZnez469v100GJsFP4H9vsu/cHtNDxp0f3q10mV+FM5FamjhgYrK0CrRNPdud7
EIE23aoOPvKh9zoHrL1QQajRWT1OeTNTVXm5kavsq5vQPO9Rz4ksjSUfZAEAUqWAFRl8oAqlaci1
a/ipTGF4ii6a9q8MmtNw2ZOEZ5kUg6viXlIcLYiVIRUKve/QsD9nr6K3Y3snz8BBa0o+PdYx1iud
5BmRrAeGVJ9wyQvJ3ENH4WHwuiQ+0w59x/fMNB5pwqPr4RVIHTtBiVcuOWOHOb1RDLKG3BsPIb47
fx8d9bLcDe8PGrIy9pY34mIXR9CnkYad4a3UZMDAmBxj9gDv2cx/77WFQSsaH/gnAO0V3Nsk9LQD
G+7o5ksfAO4hBTwhusP56lLl1DmjYNrmEkoVL5brzd/6SUk2+a5XnQzkKBW4pvEYiDWLrp9Xkx67
iUhX0eAvNHCSIYPuepefYUP2A1wWKgWNR/fNcQcRJlNBfU6crA7RkEekFtKF2XrNWBBUqYZyrMod
v7/Ha5EGqLYoCagkPqDXbIjZvj9NV63CNd3RbeuBqB99Y5Ne3rJqd/CT2t4cuANleK+lXg/Zd53u
MbTb5744NUpV9vfF3aQUL0udT6dKmaHe88p2TAB24YHbUpZZhd4OkuyHOq9j4siRrWZ+tuIntL/m
gKqYmLJmcMmczkO9hZM5RlutHXY8Pboe0xwYGMQo2BgSIrcuj+n1yXMyIaPF+zxAdAuVSCYpR/eP
xu/81ReA20RYiWMCZ58rCN6RZZpLfMsEx1ZAspMXaNSJHOXktr3eoSyhmgYxb23yE1E3jItePf6B
KsY+LUlOZb8pRgp0zToX/gY6vhl26uk9XglyEA3cVaG8qv1uZhfnoXJU0jkOgBYow0GSYAeSt7qI
9qEviLiQr7cTJAs7bvd4K7d/Iy2CFwailxG2iNhvFuvzPGk9dVCEbqpVNvb1WTT97A87jRUYJ2hA
IAr8pRw6Vzb+jYYlagJoXCyQcUe/ay9wHvkxZ6bbjh5O3llTt5Nt443uT68rOrx3yciaJ39io1E2
uL2gukH6nldCfPMdZS7wLC2aL9iA7hPtoF1obZ/olla5PcCGBfNcVSZtjbrKqnkJsmVRdauhLAkC
LLMi7QAitdEge6rw8SWv6JE57Yy6E2dDHNAUvNNlL2dbRjhZlM26a3H9OZxxJ9JG6cV17C2OmMbO
1zlsO4ONmoO3O97uhQv0Vq2DRscqCaPX+c8+TLtmmGn76jlI7qKUz/R3IXhp0D5iYqhYkt54YWiS
AQFJnbdswgy4gl5dI4+gwXbjduUpif7oG3lOBDvZ3HzbP0oM6Z5brGTMIQ14S9BCWnImIYpH11Il
MiEtRwnkBPJ3K8URYwy+xSa7p7S6gxI12TFbBpGzpFrsjyQwOoRN4JTg1TdSYEsK+BmBoCjMRbhs
mAOTt7JEBtDbKOwUX195x3ii1oZHBLPLTJq9yTJo7pgvfnbnCfWde6w8Vg8C8/npha1x886JIiEt
cNS0DexPpxUGeDt4dXBKus2rG4UZGCgXL0fPHzpQvHG33SVyDpX3KgGSM8K0EBobLPpoIeGijL04
j0yxVa6lGTPLBpnFY9SDSuIfNbnNAsq0XRTSF9yZZB80BmyQjVXQdZpHCzYVe6MbGYqOQTXRA1qt
WGtZMx8wwqmayBnVJxWIyXJMkFXIkjV1RW7opm8mf8XWsGdwXEwya6GvaS+JZpW6trngumKI38/I
peFeReIyTUSZdfJzv4WrhVIgaZ+EZ6/IWOfb1Ml8sTvdp0PMi31WkM5mRUZySJYzLqrT9Fju6vCM
f+eyPg/qbTHuEXfdCqm117v5bfax4C7Ehwy+FixHqVXkqJDsEc95dGrPQ/2YnCAHriNXd1NyjA5q
C8cK364qVCQRNK4fsiZZ4MDgyvAvqf/osD0Q/rvWXfyROAdP/jvvdvvKVpFMc1wQMilNHVeMX8+c
dhEsU7EmEnIy9jp4IS3Yj1IHXh5k/NFUNnfYdfjuGyATflzQNA0gITaWRCratcOuOSWQ8ROOhGIs
K7JtljX7fUfNV4q/ot7z46/RLehLrtRfOhFX0BJ7//iulhRg9/eqwWPx2SYpO9MYIOhnOfrWl06K
Cy9pjSuh4BTSVXrIEEbKwXuYEexPu9fSSFBdR3oVJOrihusyg8S8ef/OPIfr5/s4DIEq8xMFX6pp
basjFEB5Wsz+jmIAQFyWLUPz06uWxJTm4FjAVQwVN5MjD0f82RGB7UVC0lE6cw3pNLsUxo86Vp3i
JAYaz7aKhxIZIlVQ2vI9q1Ns8MUAra2zBMUwe6IbQmbWQFlmWauD7pH5EAxxdoqE5AOeY2nRcR4+
HtllsGEadXRjU1ZWsv/0xOe1QugkslhAJHtoPSe47SAevUBkEI94nWvdj2x1rgp4NRgJZzPKACJP
rgJuR2qavz2rC2/GZBdIwOWlbUpJMIxKyATguvZu4p9e9fj7B3AUp69dnj3DyBtpLj9gCenKt2sM
0fEVUjYyK8DsFQOul1eiCgMP7JWVu+iF9KDJbGbg83L9UJvXfRHFySPThK8WnYT2sfYdDItr28i8
cI5IzMbxmmtHcMgtcz1nYeWNGb7ukm2A6NtvMK/oOzVz7t5P3BkQcj7n0ZMrZhDfl5okqrjTra9o
zEJtTwvlhfJvRim16JP6KpyffN6lXUjsOT8HO0eY1nKY74UzAeedtH4cXSQzCw+zdYW1BKrDQ1GG
QYWZRta0XkMlbwD9P1yYHW1TnSju+9djHX0JHwesC1huCA7BHNI9O0C0xORMR40Alp0tOxnJeZij
lUBfzqjhsrsEaK0aprK/PzPXrfuMkplf/V3Umq0doz5DjDCiLzKyTZr+esv7fOEv799iLIhGK+Tm
glG95Hu5mLWRpaHDlKwCsDdIBwwzvih+04tHPKjUQA2fyPDKPb1K79WnR1jgUVqM6X9pexM0Rhep
oXFjPuzMgnocH9592iSxSmdKjylkC/Emv4CbijHN7KOvk+Ms7kD8tsODnDqLDHaBixkuNlXMA6fk
w6F5bXY8lL+rPg+Sjr0kjzT6tN8cH4FJyM0TmForKNjLu4MXkaVpaXMxM5eiLwnKFUXXXJ0fOzdK
fbIBOkJUMt43i50mxfTf66vPkI0yQJaMsUmRdYDDC8m9ML6a0NPZpGX7zyD6bQc5xO6JrmOEdlwa
uuOXe16Mij56cW0T3EJD0W9sXeF/D8FuADa2PB0XSuVD02xs3/7pQRBQl+UV36yhimjm7Do+XDjc
NBKaSCSr7aJP/wJykEeoBCnVm0BCjDvxgKDWmin6Dni7w5W/A9at4gntVGrb630zeQYM+rIXi4zm
dKEXv7qj5Ou/q1UNOPfUXeld2GoQL5BkVAOszzUHDsnieYhxz8NhVSnlIbHkjTOs2xM67rxP87Fb
OAdcmkoo3dfS0Ulu0VXHyxWwF+VyxYdcn/NtlPCrCAf9zbt9eex45p+bkhNrtjwmplRe4npEJnMS
/m926FWTcHhRbJ7ILMg8mOtDoQrgEtxDC9Ie9o9IG2JUeTCGFaihE5QtkKfEbBHNKM6f4sjkbmxL
D80gXyDB3wZUmYPNvaQY5dZf9afIp8zFeKBlwX7IjG+VSalDs/Z16ClcyrZRC6XGETRZGNnPr3W3
dJMUWmCaXkgQfrzElyKc6ALTsE5YUdulvyS66xqN/YTl7M1iJkTqbblhvTPBeaknrVp54MYhkJKe
ECuSeiN0kS6kGPrpoWHTOKdkwRaYUjETJtW8Uf5vpQ2aGpzq0rdi/QM+UK2RbYr5VCGbg5ZhVwLK
2kBICiuLkWkF9tTWJ3xT4fv91L0xeSFjUnk6aOb86kJAi5yMKTsoUcAeg6vhLcUw1hCs4w8f0DYh
mkP+zZxOZkE62s+2VcxQDWT7KhizpXbil2T+FQWT7xCxRG34v8fK6prjMtD3dfJua5PX2x7FEop8
4W7/JgDj0m2iLZENz+RgHOYjWnRL0LLcvBzaCKLcs4Y9WzgmMRTsZ+LW9tfCgiIy9vuCyf/wxW32
iVdCgJfg/drpT23wEDnMkRAwgf7f3iHvgpSkLh7e8IBcYYOEQhQeR+j5fYnQ/5U7h0cyG2KBW65z
xEbukydWCRABRKOKyA68sTwcsY72jQe7jynwS0RNGHb5ua+xMGiZXzExYOddbIp1m9apOlgAOQRc
ObpaPurJZyx0dwB19P3VhURzk7sBjENJ/FLqhLJwPs17VA1zLdprA+Nk4t8Mf1U9kEHsUU8mQ6cC
Fg5qaIR/MVeaKYS23fZD+zGC01p1g7K88obVDkHbFpCfBFEtbjOqvzlTljiEKG50Om7xf11MsSrI
Yd46r+fj8kbLxQYYrCWOpUnxgrLLV3yW4NVpL+Z1sychzHKI7h7Jji5LOD6Z8adjhZ8murq9P87X
XM9T6sFxUHTeWmP22UZpopzmddy1i7USDN5qxCbyGgpdyxrR0ijS6DAKHkEl8TMoban3hkVK9Vob
tWemvwR0siBGyXng7oW0Y37N7w6eqf1TzxMMCeculKMBPsWJxSA7tQcCyphgJvOFXQ6beNz9gKoI
EeyVG4PcjYy0jQQG11pCGWwwXOm88+VvdyV1NcM9qkvqyUkNDYF/teamNbXoVJONTYd3q/LEovlg
SSm7yOAtS4352W+L9RiOaZqq30guqBgI8v2jyQ6S6XFZhNhkLod+5Ae3uCoxa8jKnMIcGl8jADSS
5dE5f6w0aEfcIebAyQd9c7eg0ZaEiiVE80uZpQv+JnzdsQFb9H81OoaEhbTEf251AvE1PoqkkNZd
Fd4n6XQCEVEfTNbv6LtKx1BnPYjzc067gg42z/7BRvRwwNr0MYP+1OvMKouc3t8UBFSKqMWoxm+P
ATTGT7gcKjclETKDAKA0v8yAJXAzDtGQqITPXGS59HKnqx+gjexoJBJMB/5oRTe4b1Tji3E34qwD
jBM/trHvYxcu7ZzR6RXS652JRjgisxea/Q83Xf+LwT9VfWo3zz32NPofPn4pPRj5eAww1L6qTovJ
pgENQx6j3OCzBd3xlpJ2LGtzM1cVV0W3vy70/vAaEUI0XApPV+vf9BGyT1okeR96zP7gcVhytgf2
zofdz+g/nSvmMbSlcwFoiO7cdJyCTTrTNW9HBLfLiGOvENDZO6T8mcMzvoCM7+KBY+OkZzQptGd8
C2V7ZXVFsiQmoLd32Sg3P8dkefgFUKV4gNA24nBBpxToW2Kx1jmbKxknwUJ6bB1yrbltDTnKovpt
OF9bQ13pPD7RSJ/k5kfy+kpvaz7GjUKVFgBTFw9vfAft3h0wPITQLwmyXtZMewwABC8/HyoFCAza
gULm7lBvc6cDI6pOmt9y+mXS7tMuKbn8sXgoWw7CBpwl1hL5ey7iy7frSDSEYUbmC+9eOXesALJm
WEzTXnRZ2KyaS8qDUzbSaKN0orb6MRldsVtl++ouhnotwrv41fogYgQqAr7m6Uemlep1GDPXX8cN
r1huPO7G03xpLmpthpcoPs/IY248aVis6YVRULNwO2c6pziSIWc2B7j4Sw5e268BIHLYAj0Wo6CQ
hBpsrjqQtZZrI8nBruJinSX1D+7r/syhQ3YizQvfQSolYrBQLu5vafxYVTvnELxa+vA9u9tzHKqq
X7f2AK4unDVMt3qNje95GVdVb/U+mfxCxmr2EcEe3kSa6Q1lD+jnss3zpo3Fjs7yXTE+fIuH9Joz
miWCDz9zyPYIEnMHdvnktrUbIO1lb9AshjiF0MvR+030MuxsiNjMmCPhwmfYv1C7qiZdsOwF2e6Z
vGEeecB4yK37FauAygqSkQ5PXPIrrgtA6vSB0sMqHvx3iEgeVfX6TwhqfrOksZ6UAz19IOHm78Md
epf+0je4G/2Qu9lHtH3/ieYiLk7rQAyQ6BmGyDSOOxhxacQpZo60csZaU+Usyr1Dtk4QqUFqty84
xGpcR/TwzBnSuoQvV2CnlqCOc+cFwkp2lY3MGvb/4y2Qiue3HKviDVEZBLTj8/7I4BzF5gGWU92e
IYpUB5C2144bFLqgtY10KfegRk6d8oRMSpjmg29MoSogqUnGhixrCjJD7HEuC4bMz37wZ12i4iyU
+dwbfaH6fpAJg9HgZNGd+/A0ykjI5QyYt79Y+0dgHt+D5CkPpx+/sktrayZGH8SfMycJcgL4IJw/
dFfyDAfODvoYClbC6a6SrXBqT2rxWBWQz4+UHncQXYTXvFwDCOVoooN58bkkuqfwFHsitpT0+mpv
/5dncNGNe0ksdBZDAVCsTFts9LHG9yocYt42/Qw9Thyxmj0syY/DejZUdRjcDyLLPOYc61VRNske
Brz6PDgdVI1IWFaehJWKka2inck14YvQoMMaZFZ2LxxLoDsXdHoijwb8jV9XTd4bYWbOza+0obMF
ykMOIioAv+67kvsD07ltsI7ehksxclRyV1MqGYDcnBEPcLE4gwJfRmOafhlVVQFeaKGeov4KU5TM
59WzH0t2PLItiMf7lrRk/98UmnOsI/0z/vpDMLhR4c1GNwSiwCsahx5micEz0C5jQ78YaJUfgZo9
ql2bYN1bFHPaOcU2csnulc/cO0xoyV2isIFB4FpmkBs2c5gdcLwogetBMJXwlIpKYp6en1jF3Abx
sMEEr5TUJYkFaC9zdif0aOBqtJ9oHSdij9wY8BXmoPwkJiMtIkMOF5spotFjtWpv/IS/N5Im4H2R
P67wMiP2LLfi0czffnsti0Z3lQQLD8UTXR3i6LHSfKebTjWx7UhFZV3gt8Lj/jEJ9d66n6cXpC4s
lFJ4KBVXsRwPfXnC+7KEcJWDjXG0WRDu8qr2LISgtGlk6MnyUjHKJbMGV4v514tDwwalFEGidymz
JN5FV8WwNEIXmCfWyP5NCQ9akRAOujlnFgv8qppqNAg//E3SU80FuMOJp+di0HGM63e3p3WCnAoV
DqH0lwnxUhrBeKdbsHFCNV6U+O03bJk5tbrvSm5OFqj/eCHU1DQ7NF0L70ERlR96SpTfPSbz5K2i
Gsexf3Ikhx+YP7F667oxMCzRv3L/dj+istRgc1c5L60zVsGCwW2VEHHtFU8n4CDcWVMQutAq0hoi
AvnJofq2Bvg8vZQHTq2/FViKLTiHGllIwC+iQlK8D6npMOACiLfQl/KeZ6veAmWGXxV/SU6kDWTj
1S9ehoKLbAHp3SP6ZPBQ/loCP4QsCfCeKSqYuPve7GL9pbvwIqRYe/TFL5bVqc/jkQ65tfxLT9Ay
HKjWtSUbprj3lRF9xWzI97jVgEulG440pOlU3VijhI1LhWaTsGZ+Mhj9uSsUFyDDIsvxcyvdlJUl
SkkebTRQZXaS7VwiIopbyYenQLgydLXY3c9vMdpvDukejS74ac3OBHkDL5yl3ekAUaiXtl9i78s4
hDSLjfOlgH8RBjPiTrUy3kBlz8YRS1OdQPVU9cehtE+5YX4zqUUdEt7sIEoQexteluaPbdiruM7f
cX+grsXL5/FHQnH4ykFlV8fdqxyGFZ6ebzxb7NBZpTQdO1rLQC0uE895zOOBpJFvN5L/LTuKDxTp
PEqsJ5LtvWHeq+Oa4+JDs9tE5lhuFFT/kfkn8MrAsVh4eeLsrU2HDFUdWcDfyu9JDEwWTGQ3df+E
eRJ2xRlZrdk4FjR0YNguJ1mm7UWilNwvL7mKVzwlpQsBBEleP7QgSXXLu9g1+TGafNizLLuppzCP
6WBCOlA6xD3rLDBdTsOUKJu4Tc3p1csRMLp8rLwqUKyiQqeO5pOXtiRVyR0TRJF9YSKtvs5yPZU8
ZcKnR75AQ/wGSGU0OZhHMznhKhES08ImneIiUH2P449C9YVgb8o3srTxBEP01bVhNii+CoYDEBoE
WpEkyIwwd9NvkM61QBVzwa1aLk+rDupizv683uJWbYa1cHADkx8fzuP0FNL+8WUK/0C7Vx8zfm54
TqxEVVdUdSoIA1kVZGtCF+3/29vJV0tFKhkt0NLpIrNr4LPsDTJkAmO0zcYIvjQMp2wnRMdNlrPw
mzbu5364TudxJVJK+Fkm8ZTw4ug8nm8zVsWomoGyJaBYlg04M8xvfx20mqIiiGWt/g/tlb163W8o
piwifKsj0PCEzQ7SjPYQXIroYrJN9RJx1b9NSwC4oWUWNKulreAj/ILGXXfIBrlp1soX1CGHYdct
20lVW4o2OBLWekQ2LNt+qblCXMSpXzRmkzvOoGiigCYBLMA6s1TOPDtZQ/FKc31UMeWA+j7hN6Va
SYG/Eu9IgzesR3A5wcb/vBMg+0zaBKHPAsFNnaDlIbvJm47IrBMPBDhch//Hs0ITQ6wF48yGHRHK
t1ZwqWMA6dZG5EkerUNkRhqsQ8AqpLR2R9NY4yZ3EQJltYRdDbhaK8MikL2GkHZRmgkZQWyD5sve
qu9M6YqdotaQnNZaHcW3rDK4QVdJy3RHjn5vixxr7+f6Tp/saDfzuYy9dmpTDLMm9n28TD/OC6Ca
emHqJpwDVA/bhKHdRi0awETr5cL8uakW1LnAak8hGzag1a02ashjXu5T9srCQCK2T65akgLGkXj6
5fFOQ6gAfr5FtfgNNlIghi7bOFoSDoBNDs/oTvCDOYhtROvLaYeFR2lF6B4m6T7sNQF++3la3BFz
2C65E7LglABu4NGsFj0dJtCPSdyDNGiIXb74OogkAkzCQk6FEHoHumbxhsi9nmNWZkU/vzBgsTZ0
HG16Ac5HBZXStUmLQH5qXDmIxrLk2X6h7IZBH1vjuAQ5tCYEqs4eCRahs0AnA8zgxjiqTjFLhWtw
2CruH/ZkOVnMCKgE8+tMSjqxNDpS/yLal/HKRagJLqa2Zae+d1fW1pJSDyxZz0TtOK7DAVdvJ1W7
UCWvmpu9XdJdhSDpUNRmcVXRGkgylhPiQlnXRAqi3R3Bxk9XpnAEWgO6AEAIBnoG8JModCJ/Po6G
zyq4Bls51bnm3KDgioeIb+Np7a5bDI61WSezcPqClof9/H2bSbTkPgDh4Des69k08trEeJXif++s
7TzD8h+gRyIjbG3I5jTXhAP5eHVsnfWO+Duo1GzEKWD0yjaLmULJZRszvt9eHHpLsMBQlUbsbT7I
0Mo+xQPY1EEcd5zBEWzTy0JTJXCJcEPxAwur/gmcKjVuWptwPd4k8EaaavhsfPYoz+To+VcraEaR
QzV1Q2aZ0oUlcy98VdWoHUC5EQuyxzE3ooRMMklFAWI5Zeasd/w3J912wicTG6Cc61UHwPmKAD+0
r2/nw2sflH4g1gVxmQVwmfnByx+rKPf7PebTso8J8P/qsxny6qE/yoKjqu8azvllh9f2Ne1/ig1h
ZCSNFpjD5L7jiugiQG0Lp3pH6i9CKF1LycskbmiKIrhF8cuudOJ90eiYSVTAKyngM0siQVhOHejE
FskY2v/P7Sqtgo7ELGYR7PY0eHQsMmwlO4IrAwrgzspGiT6fQFnBh2yb31ifIkv6WOQ7Kd6Iglwl
eOhYNEUb0TPCjuPtGr1UwoPa89AdBJxFBQcdr3gacg2pSwylYKAJxlQmOpzagT13Q3Eal9PYtrWM
dU82xBZ497aTsDo71S0OGVVpf61WR1QwquUNgcmTQnJSYx6Op57DMqaYP5d1HV0Tveo4MsUMLCwM
EbbNsXWfFXBVyTP+He1/4Aa29YQtJr+sL1bEx2P1+ptJWYDSY0LiHTbqhFkoKlYNSdg/qVZe4pF0
Y1akVOXNbvJnFVpU62JfXR6sVZRCg/JOCIuLHFr0DO8PnlmJI4+3xJbTPNHwiuSZ0OGwj3BgRCzP
SaNooETfC7ghYJPKIy0/JI/QiOZm5OjT1m3vOhEbg5/GYpQcvAQ3J6c7eqRjCkmaVVIytXLxBjvv
ORx77eRzINtO7GHeV6keuKsxMvGoJmv4TliXyURx7wm3p/hDtFxLM8xtgi+KDj3ZJp8h+6VIWTNv
+wPOiiTFLsfKkEruCZC2QmEMFP2Iuazu8aJ8w3a/mqVAoyjgn+M136QKIho1owMBzvmzx/38A7/Q
qOrtnvssaySSFvmQ60I+cKMufzo+WglFUjq+/K8d0YrqRoizb+jaqclk9dzQnwf1CXjpBw0uu8XB
7FVmlwzlTAnYnznzxf8Pc5nnhRjx9d+k/1xwXXX7lTaS4DCeyrHqpp8ruRTV6VJ8QQR+NVfDT/Po
YPPuNNoUQcX9SdBjfGx2Jy+Oegeaes806DfjpYOfcUBKkm/dT/K7bzbCRagPcD+ORdCUqz1D4wDV
UatiisN8wVReluj1VdtMbRqgxUpX6x1+6PwXj9Ci25mqZF4FR+oTRL+LqG9wSDN7quCdglIicWbB
DhriRvrgYqDReokR2xchDc6HFXjmD18O3JE1cYf5WdYgkfz1OcZKrNVe6hml0n9I/v+qOgbloUCS
AkJYp6862KJLq6b5CdqhDdCatrJRPi4M7b7G/HkKFN01TsVtRcofDtTlV0qtmbpCJtVTJMCavHrA
kEEuWNPeAMexbP0iAbRLSYOrF2l/cATBsJ0ZosYOVy7+Bdggs1w8z0LFSOC2L7N8xFQdEkR6N14M
EQIrGeVpAQtzf8JHGpBhuptdR7wIbjJeA6trLnmL7r9CCdHVs/k2g7iHIP/zQJMT4iCI09q6tr3M
aq+/xTLA2rF2Az3kV2/vfPY2uNJ8xxtDUVCRDH2k/AR4cIR6OwEtHP8OmcGQEBuQ05ZMwlxM1GEV
GehKqlEn+jAwE7dJRN87AWlWaTTkRiEZc/J/1+xmowzbZf0UhTaIMUJmgPa7iqP3TcHfUDLEKis/
SVdM0aRNfqSA2Yrtn0KhWx22S3Z0AJ1dhPN6urZsttkvkh9D6T9f2cLjTRYn5o0sHswcG1alIQN6
k7pBQsJMaSAHoutUCRCeTRR90LAV8n7JUhYjoINqL5OGW4WV5NZKG/Op5Z5s8Gvpr490pnkpCifG
vyxLI4bNh4FL0dPqHh0vmnYvfxT7tj+leY9SKhJU3G//8SQw/5DT+Oh40Zth6LdHArLgrmlzdoBK
IHO6A6NY8AXCdnFvVpaBbjTZ73ykQaknX8TcIJbWb+GOgTk8AgAO6SbYmMXCSuBWZrUtznracqT6
09Yuw76wxyQZJQNhSmm5KLcLiwU/Cv2SiYKPq+l7c770u6p1k+2vRgO8EpRTDlg4gjffvJQZ0zqF
QR/+BdQqOlW6SMFaW/0l2/HClobjAayT5ChYxl3vdUnId+uIBsb8BAJygfx0aK2N915B4QmmNOar
THhf719vtM3k57cA+UUPOenv6dBSm2068KZ1DnMu7oANC3C5Z89lkICSkFFGllvgk4dD/ZE6qrH3
P5RYx3MDMwYRR05VXUtT8uXzKFyh5h57iILYZrxumvybpcM4+fbhNARyt83ZBjl4bSSQVVhYIZys
mfDLqmqAsAbTDuMnulLkbQW/qzSdZqJASvMNeHXZFwC6qcLftrTFZgkhk5xUP2B+iz3fN8/WaRsP
vrxrb55LDn0fkGM9hwth31mS+pvAEBn9bqB3DY39x0iDCBWLXOBJeC45OtiIBgpKqOlYl3K5EXYk
Kp6oWY1exl/Ol6bSf9piJ5UCE4wLZCbMDUKY4RqXK7mDYW2TC40Md9jLoQhZU4PrpvZRDl9h2lne
l2lAEWiWcoi7Zocnf023UhcsioGoTmg73MFTmgLWONppA/s4os8jJJR8I8twjnFq29GxCgodWrSU
b+bh2l31m1P9SpIai7fNC38xyrEVrpKyoxcQJoObKWBIWpJbjaasYsNInRWzUo30dvI+wFL91q/V
bcoK6VroHQmVQHn86NU8NQYvCuuUO/BpTP+9Qu36fP2Rjq0V+utlhrWlFm/9I7wMdNHtKHL5ZgOH
KIrifuBB8gC3pHVald/kFiUJ4nT6ziL1fIdlekFrwTCYo9U4Xmc0D0qeQKSCEs09t8FTZh8WZYVs
d8SY3AeW+84eIxBJfDeFPW5rkMRl7Hr5fHv8vi/F0LTmOmJxBMYQUgm++Tcza6I5KNCQmBc7ccHf
sQJ923yGphlxg+5HSqNs4UkFOPQTa1Kt9DxR4yrsvGOYZCPwhNvzT6KnJ4+kCkXt4Zptc7Iqw4M/
cc5C3umFXPvhN3khvGc02H9Bev/OBNsyT3Ab3GkKVPTB9KaqJn0J4K8Cxng0I09klBHHXCV1aMwA
+j48wIpQtW1YHG5GXjV1jJvRcM9RBUvquBVA2o77vAhqVTp/gTrWBFga4nRSMVRSQ8bcHXgrGK4v
ePkcmtyb/xeh4BggFdDiZ7lxDB96GtaXy27fIg0ilzuSDu1d8d4OZl4jVuhNjJPG1s6ig+RSYT1v
+OpR3Wy1SCWmxaJS1/KxIdf1HmrbqSmvuwqPhKzkhjbP8pG8vl1unDiN1q9L7sPbLDcZBXtdVkeD
6zqZRITsla+1WrpS18ywuhKl+hNXETJZzjkHk6nyHu9Nmyi0dn/mTSLY96KIYqm8jElYzjlrnyno
UMcq8DuLEhUAm0j4iJUTAXW/T8lNdMq/3TliSBKr6LX5r0j95B3w3FxYKzWjP+ScBNnIZMJo0GAN
/5u9r9OcPg1bDTibqbP4XvXkAp4J7NAAnCPWi3KI7JiXJ8+vVIikIgvYqaFUW8n/C1wCFFNvDlYs
sENseDfsQi7ERMEqJme/zcr6UYmarXe+TBdLXjBmwmC/Rj4+EGNu/V6a4L/BLypMiARxkmp2DSAt
sjcJUqJrmim5Xne8eqULGcmX6y4EfUqoiabcs0cM72sZtuvG9tsO0tK9WVaOlrMOG6sPVlr556Ld
JV2ft1F0ip0fB522PvGmfyin5iFacmG0j3YKG0MH9PJh7iJI9NQj9uUh/p0Rb1LOEGWKKpKigbDm
TxSmPFuI8ia2WGwkCKuRFBodoNXKWkbe0/AJ1tow/AxGeNTmX8CqCsrW1uSVLxoyOm6rHUtlL9GK
xAT07sMklP8y04TYiBPbSG0vhFCiBPjXLcUld+M1ni7w/eJks9xKQzCjBBeUcFESyP3o850YE5rT
Oel8yM3dexvPwiacr2Q8+re7FHn7efNjcMo+QBhtMXdfZKQ8LTSGWXKVuUNdGLemNavmslk2WJJy
Sv+0zQ2vCy4pFM3PdCbR7jjxpWTTyceACiLem7U1T6gVY8HnjcggKf3I4RxPBrBqYgNxPA88KyiA
KULxF3sExpH+1pWQjeuN9OAN9+mpoqeF4D6f9zO5k+HkH5NcAhfxslvnr22tyzXOKNqKS3PO9M++
LF6jaZFmO/WZi9gl6zH71aqBtLXdAxihlYHXe2TSTPd20UqSblXzM26Cl16QvtiBynvM8Cv2hSBd
BJ7KmwumMHGO9RgAZdKd9LpMXNvAfjHa3OzJ4adewBEdnvuDa+U5rM3RNWF92cMXKuKWQOh0eJiy
AoZTPwlfmMTyuPCrkOpjWhufBeF4AI369HMZvAa1EzMwBrwXiKa+fNHzVSsUMORPU4AD0KqbAgPg
Y7O8O6MwyJJbraFprtmopluQYMIOszIDzeN7hyxWetmgWljnAEn7mkmQUr3tXhOT1dsXIgp+nqiU
0ztIgiYAQOS1s7IyT31bj6ZEz7XmoN54Np4eb67Zc7T+Hgs+85QcqwwRzUMcBtSJr+2D63o49Rlu
fbiuZB5U0GpgTac1iIvIZlFurLCEsZCuTwH+lj6uINjw1wOPq7gxvVujPdxiu57TYo4+2FiJCio5
qwFHmzLaM7kAnZu8XAO6QFtFmForm5GJfI/e8Mw/AhVFjduLP/AN9nCdQujJlXN44k2myPqfl+w4
a5e7yATgrjEALE3tS6lhLU5oCCH3hXBubvxzIeOe2sJ2p0br3LPOsZB7jDIRSJw115hfHt3+31wJ
XhcCqe7D9T44Qc47fEQCc8vqh/ULOy6TQldkvcL+KmMYz1YLx/jQ2qDZ7JKEOZbuoNCTalbHz1Ek
W98R4F07mpmEK/yf1JgwG+Y/HJIbJ6GUVeHrpxqS3F+mutd8icjbqLQvn4C4/WMjj2TOYJ/RBct/
S+TYaTmiT4r9zWwRvnmkP+/Lca4XOySYaE84KrOWH+jYNO5r+kZjGDKTJ4ZIgq2tDeZ5/dujE5aI
hC6nxfrZLMUiOk/yb7kQwlbTkg9+oMttB2JxU1w6ov1FjTm6RIWcfK1Jf9YNU+LgJhgAGDz14gtK
xKzs2bi2ogvpc9cNZlT7gVu2Fmwm84vyb87NoFiQHl6F+UYGEzVDO4fcqL5+S0b6Ftn+Ne6GFBNh
ulLpE7jST9cYrruGVLRq3xYDmvvHas1fDIY/7WGxm1FN+Wt8SMdkAS0dQXE3aoEyrHg699rXG93B
HuVI6DW/eRe49QhogYFl3gN+fwiI9WVRErXhGlyDy7wQ7NO+vB+zVh6lCWtLns5sMqX51F9UZ3pr
/UL4vCXLDJbg+1mq6/3PAsZCSPeBJe7pfV2ewSjtUn51Pj2leDI1b/xLOHWg1P10klc8n0vFN1Dy
dugD275a6qqwUxniIvwll6tsISWbgMbKEi82vI55uUtIBSfVK4PqJmzRKPZvrN1Ff447Mu5/69D1
+nlcuzInLk7+LMZ8YMy/CvJ3jrE6XT95kcnLxvFjV6ttdDlAH9St4DMIz/Ee5IM+ZxkCJLI8nrW+
8QcUA1tOFYgoiIjneR9NzT3UrKr8p8gRy7FNrOKo5u1OebwfhIGfxSQOemD+Rv9cYkteS4AnYh99
6r/FUvPmNJTEOdJ6mdcQBL7fUnBIGNvy+5SzoYR8j5DQs+yZKwq09YrOjvvVkDyFR6Jm0bibjua6
PogeczaEUnkpNg1W3RNYBMIEkmqizw9QH1faxUwjaLGvne1/U3F3KnLL+By+tc5aSn+VWg9d7OQL
QgOnuK9STHEy2RKIYqO74qZWpBBocEE2nLD6oY/UZ1X+EMiRRZeoZFOqO5ilEUVff2Ipd9bB13W4
9uvfGLhLPcUxlrGjQlzW9CFJmjU1wgLGm04pVx8LDu/RH4fkmhuKoLjBOPrcR1mu6ikPXxVAeQFN
Q4vx1rKB+if1VXPE90CpDmdcfW3Y1kWJlnDyPoikW2pzGMXEPwY1Tftcmr19Ooo6s6l1LwMZR3ax
Y+b9Flal0CxhbuWy6j1r2iLJxauQKTGd8fAGgkznOJbj8tHOrgTDTEHkV6XcoPs1FBDYoVcngRNp
MukM3TGwvM6TovesEvNGvyymBD3jIKXAlwwnjiXA7rrwgWpWZIvUN/r5gMXmp9lDRqmvs35Q4JmY
KU6vPqyGrZcvT7XoFpxsX/nDLH0y6rQnvMoK0gKTbBfROKlvQq6DKGOGzFGkj0KeJdi2BuToooVq
8J/Ria+L6HlpmJGAqcPvPj1EaI2OU05D9o7fMkhOS5i2SA/+D3GZ1iaTWdYbov64CrUKigqLQmXE
G8hmJ1YAIMkC8FJFAU41xXnVot5hWQPLmf+SZwhd9apAMY8zX3/O8nBE58AOtFuoAzkDMj+K0uhP
g57JAvojcfphS64qW07Bck697ZgseTCS5jprwYtXWM8+x9jNrE6wVl0HDEHa9Te9gLVBsSH4RApw
aY1s2quWIg2JTye9e9xhWMYGeFk8DqYbbbBhzkkzf9Fgy7XvaevrxlY2z+BkzVXzU/gmLKmyvhsv
Wpt9UwfNyCYlhaISJ/kZE+SAB6FdzlKC7SKfsWBTiSp6jlMgrGEqmYFgh3FWoSwnoL717rcthgyM
B7bhunnMs1jkPneqRc0hTvZJhOm1tjbD9lO7NQka7pY9O9np9Aevh0WfrRlRtnLVpOl1eFjrblec
5EmFzyY+ryQvoNTjhGGcCeUwLnAXbW3xsfd0Jtn1sT1iXhHicgPQafZnMuilfTtTT30lKotSk+U7
f39+broqkv2UDyo1tShfqSI/16od4kZnL6YspLEuU0o352OqJU+J3eeN2xSpH6WR7jjiZdRkgvWU
a0hDwlZ+souvRZrZtQjqqXjHNV4//kfpfZqaJjPzl/WvET1cqX8dqcnNAhyoEI83RS97dspR97Ko
0mOaVZVHQMnp+31osQNfM+dAxP+dzqA+HN7q8SzkLJY5sjz+4Be3KIO5oa9A2EEMuZJU4ets+IPH
1fU7dtC7LcFyZWj5FMaYd+tDMDpwcW9pvmDGGmqznASu6cop7DTfM7NNJ6OHxLAl4jkYasWSCRpa
esRkyXTtw/yLz/2cpBrOATeTfPNqbrJcCvShdFiv3Hipch5tADjsNhvmctkUftRhLEOaIPfS0HIF
TcI3XR5XSWlqxLWHgWgkwXfOAggNvy5s5YlGiYzRcSczKNrT8yZ7GAsDrNHO2DLCsoDwOqxpWeLv
11YgKa67FQHOTjtz3GUyzV+JJm2+nfuQ8fbsjdr53Go4l3FTFGyaI9pYc9OumTIK73Jp1kgfmr3p
RLkaEyYj9uyWdvETKGBmtKFPAEfNvpVO4xNBr8E4EK3hYfSLAbTqlySE4/uBrLwCnFJAxw93SdJK
6U6Uf3YSjV5hRy1uaODe8u9YxSPtZLygkk5GbR6wV9bDOILmF3t7syvyldWXK8zma6r+K5MLH1PJ
QscfcMLu8Gq2URFpnaoFBCZIeG2XbkD9siLEAiNFqHmu0lpOe9xD93CB+E5N9/FLHnZksjBBNMPL
Unxt+J0iZB7+NwaozKHjkXsW+NwUORZyXTgs/r2tZYtL01iXlg9JM20iXe02UxWRqCLCIkhlzDO6
WQfDrZNzvUO0kSMLlcbxSHKRnZTZ9RQht1RP1jVT4ZD+ouX5+6nCEN5aMpO/PzdQm269lfJqDwkv
W5pUtG+KkLKD3Nhzkbn/PTUdP1hn0wQS0s1pf6zmhs6OGTXeE4+7ovDfivqpD564It/2uUn+Bkjn
c9S5KkmwfG5DwozzFi/IB9bNhlSr8uFGlKWz+aMgVoK+Qu7jtFI6Sh2HIYrXyhsHN73nmVSjdLkP
QIpO+4EDa9jsZJwoVsloPOGYxOaWzD/l5PYV47K4hEZQE6MffcSVTTjQUQwIDuNbp4lOT5/akuds
xeqWK1zdohzqNJFWia+YxI+xRaqJtaz5pSeMKjr9sw7Fh5yIuxAd5W9QGGvADU63WWwuJFsbH9bk
TgX/36aObFXEoL17+XBzi27hCHi4JovC5usr7/eu7v6hyn552+ALDu48dvJKBbjLYbuIuRQ4bq7o
qvc4kD6jD3iYqaZVX5ldSOIXMoCVuAiRAJbfhh1r/nAubo1x0E3FytGWMOZup2erPDI1EfHZUhBC
AGW4azy3ooUOZu4raQDKXANgcdv7Gre0Jd5sU+9n6uCeQAsEAT0Foa7ymkN+E11gnJbKWfrlIVk8
Jk2LObtXLxDFrfeLWXklMsYRvHZHtH061sYX96uU48u7lt/cwmDIlv2W0vnlhuW7Eg5B8+bLs1jk
VOCaNtuoqkw2KEAuq5kNxKnbf+L8EKlhAV2dP82m+7pl71X2JqSn44aIgCtUUtFCcW/YsSXSrnr4
06fNHZH6v6E6x6dGoIuRyV503SCCRZpj1Ip/apeSDPru5ClEcFt6rsZnlfUVUbyvgwPfN3UrePzL
Vs7/VJIqKnJYylVFzFsbpMbdQSXJDNIbBhoE+6bFYAbcpmop/wbTZlCRG4t7E+56PCLPe2rL0eSG
vu32DAdN9f+82lWrjjN2JDsImGBedjBA5iHRIUK9YE7R+Vt1IAOkebvvdKQx3fYe2bes/NOICvEd
qjo/bt8a7zLgJbhi9jeiwZ5u56aSF1Y7d8b0psT62cw1ZJ1V02K/7GxY0g2kyLUDp/xFbw6f0wfD
zEKLk26hJXVrFl9hWnc6fkoJfm9QSdEpwRrDR5c0shIVpf1C51WhQ8AMlZFZIABxbxaiUts26Skz
gWR4If27trLLHAZBbwjpqjJVheydHQsUzxP2FgypT68X/zVz9DDmXuxarA3b4HZtSkeqeskUL+t6
dC0tPkBy+FEuREy+nYugg1sxLDPMymbn2NexcUdqH7omntEIEE6yvPI16J2geVK/Fwj+cCF3GQk9
t1MK7LSvvaxym52NzjtNhISDv1EK/Hch1GOfmh385Ze4rGXji9S6rmG1Xppm3RdaFGW7UMBU0hKB
f0JFTCTA98Whxs2+45mF4chWG389gd6YJqXNjEN6nE1y0pkBSWAxXOZixOTSjfvcw6tY2lf0ZIhK
47wMrQo1M5mWvquSKdQXJfp/1smhdQ2KQUjYYCo8eUqXC40+RbX4hKhK89l8WcSdUUw3/FyR58PW
GffzK+p7SDfK7ZgCCxth2647fOC2eIlK2EvIU+KVlRl71sUNWdhGV4hrW6uiwG29xTzMCbthOowN
0shrWRvNA2D2waOuBS3nI+PUUyYRI6siW/vO1emH6ZLdPHkydyguWXRK94Og/OuNit8L8C90PdQc
m6uFwOBGtj1UZsx3e2F2k3t7Pg5U/K5kVwb/UqljBy/e8dwdOmuC/Uiaukh4MMYwZnvS5kYaZy+Z
4FN05UZrFO004xvGzw8dNpqkva3a8yYiwPeCxnobEyE43R9v5liyzEod65z9S8LTbrcfreo6t3h8
lGJWtBcqFms76NMl4kYXNIIy/KjD2DFR3FOaxSnBV8L0HnDrRc5SlzsSDmqltHtRPjsy1zmplgl7
HweZ3Kr3BV1kBE4gSpzGY9JbFNiztV7XlTe3UPfDi/Phy3jPIPhBPYKf+ZE0nDkFQfEKpjVoUHrH
F4kQ47K9rjJzM3nuU7wZhcVsdZu/N1PEdZTX3/iePBBc6WUsUwVh5Y4A1dWzS/k3yWdqs8dtqljI
YJjEZpJ297QTVpUF6ySJ+lrHrCametJGgLTJYwIAUnahKW+QjRBLkig3fFPe5vfTu6MjU7q8HBJS
YoXnXYSHvnUBZjTft5entaFH5giBpYsiA3kQKDOTpR9ODBqaRFfy3t9MoHnZnHACkkPIERevMssa
ASe4ozR7F074OtyqyJXzGrym7k3hM0d09VDE0K1balVjBSy/X2FTNJMmfvK48/IgR6lMmyWYgZqP
ZOhisKAB6KnulL68MIJo+oXrcFANmLbI9i8j7/ftrb4dMxjpB/RPxe4BjC1Itg01QQhR3MC+KH2R
ryOabbXfrVJGuKd1eqQ15V5zvBnZfjkb0ItNY3I7dLvQ0AVCDyIYAL7dJ8Miw5mg+c60seUdJc72
3JGlzLm4BA/RP3sI7JDzdNZQWlPBCmVWAdznk5b3wF2hTLqBivcnfPEMHtwX76lszfP7DTbtNm3k
5VBxLTgwLiXvFjoY72fuqt9T4NyFg6zYcQt5t787j6/hOTq8CMh5MgjBqpDVPv6fiBKlyWt/QxK5
TSnslq4edrb1vSIoCDDEYTdXO/P3lv8ijGx4DRiwOjzry5zEVyVx9OCpjsD5qGM5hm/F1yvQf8v/
LtYCe/j6o+fDciiWNbTZgqb8oIN41qLI/b/h1vM71W/WJ1x+NSv7jGouO+rM4W9/ZkSaTW5wOrkM
uBWqGBLxdXmKPUEX+nCWoIIPoWv7ScbmswzhfQ5Ssh+1jo5++Ii+1lZFCP8Eq9HbUL5Qov6SOKhm
EdxgDRwOGxFcdkqiI22gU1so4Qar/yzkOuFa3w7J6qW4SlU7N6IxftK6qGdEKS6APsdoXqtrA33T
0/R7k5rk6pynxa6l/obsQp7k6/MlWpGf4cAg9QMSvow5/6wc5kt0jV/eYOILc7rxUkmIQPgfTkwy
+zvkgCSwAhItXTDDZ1RCzvjyHOP/acCz4siRyqA06JaZFdyIYPv5Fk0rBRZVhRIbNTLWvlWG62uX
nw4g3fNohncxESzpXkCjO5oCV6rlGaI7g9fFBdjMZ9wVH7iWQSFKUzkigCwyHm0Ebdk9m1Ly4dnP
8gkig0AY4R5UpSsGgpEXMnTRy287kqz4H+dHcTGolRo6+/O1OZc7ABUjiYj/KEA01D8RWRY9PmV4
9DanYZk7rMoHWYz6rIZ3vO0Lf6vYd/QnJ/9la+g9ZFuBpmrrJudggz8s7FFIOB6JzAOjGNGU+DpV
+zzBwTMFAWcuJuj8sZx3JQMdhvHnFcRHClO7XeX7s9iqkXgRhogMjjd8Kfvk82+zwg+D95wX7jPe
2VcfaMET3Qnm09tRjPgCKtG53yBf7XaWW8lJ93omZBItxL2oUQt7M7QIqSsVHkCS0sox9zL38Vbv
G0qpO3uyDQhVKaMDKcW4nyu3PK1gCya6RjQq0g33Iyrhq+iLecVDf4mIHjf4fioSjYTCuSdZh9oT
z4hDXvcJdw65nTP6sLxt+6tAIO75SN8gwxRng8FFUhM+0AcsFwhzJVEexWSCtFYiSfXnNpzmR1yC
wkxjZ72KnoeaRRssEZSJKSG2wB02za+Gk4TOMbiDrFa82bcGiIo7O4ph1oeQOt/B1g+vK/QoitS7
rF4Jx56zWlgL/r+SIXhS/fxBWmMSwmIamqoD7EndOmE/KGEAL4sFr1HlkNDjfPK2hJr9mQch066Y
sotK5iWAarXQ43x8UzEWVcRJhg0fS5u6lt1TVsR4itUC2+FW98WNn0anywcGmWmou1iszaI35KRE
P5m8ppM/7anAm+P5ZU/kCBOkriNni20o4tqdUgCQEcc2qZJ67JJZoor2szsFSgoNRCcYPXxA5BXy
9SbwvG8UgqY2Jpp5uIoCjQd7i5c0fkaJL5VzgaEzQnysMwcnqfKczSDhbN+TyYOSNzENFR/c7YJT
VU/x7NOIzNAS1nwN0O9O4B7Q8J4VVGaCCob7lo63lDOnCzMUaqqfVzt0GpllkQz6nNNzMeCSs6de
mNpPCetRcEFdgu50d3SBvF2NA0y2zZdgD3mFJZ3SGp/yH+S63MketQEZaKUgLBMyONAnR32q4pBW
r01zo49B0B2v8ik9qAu+KPbGunXH3+eOHHfvJeU7Yjh+SYF/kTiQCLl+iMTtYEVb+3Qb66o2TP0z
R9XYVnDqk2IEkds8XMZ2C7bMNYQ4ty67hBOtg6Q1rZv2yYUp8mz2kjUNcmnk3bDiYoNVYUcBi8dL
Zmu+KS68DUg6Bq290YQALzbcCripFGc1yl6z6Bj1GzwrNOiwENxVHvvBaJ8bDcgAa+PBwK4xReZp
1gNLUaQUr8g8lymzmA7hbB7ien9UgJ9w+S6ITrCKqEkEbydmhXKPOm4OqbAFb13uzGYbSNkqckgS
w6sd3b4bECh4h+0HYfB8qwf8ujsXzUr0OwpFfk9/qLx5BQ5+2nuNJ91zB0+YaltMZiJIeIkKhCX2
yC0ZB1xw/q9Sof8hdOkVQTIECflmm5JRWyTfGC+BR4dg6FRuPsavmXWm0/w0DTcGB0mgBj+FSJHp
qqhtwC13Ar0PVVBxoFNbdRkHQst0MFavvT1q/ENuMFHvIvKKmj9Nfy6vY+Ax8gGtBrWWsSXcklN+
qtrC+LJJ3yoXfDnN2IWUtj8iC0H4QqHtDarGobCilPf3U7/Iwhgoz3wijvD8zQB/Yogg0w0SWDEC
V4RXTMSX7vn+ix4/URKYqsF33ctdKJiUK2WG/KHgbsauSp2Y52iILhmqkzKn7YHZKFYuqWgn0Gv8
snVSa/hdQhKAzLz/Byey+xHp+nqw1U11NpmqlcjVHR5FYa4JDIzJnrzVPc2Ri+w3PbKX6HKoL5fz
20O4q9I6xtWxPOvjPdsiJGgsj8xq+G5VMcf+Ches07c47ESrwboRq093kD2UsbtEcUHXjnPqbRz7
2fSU7ef27nqdDR+UYqEo2g86GWL/EOo4ZNpYIwS+VBSD56phsDbg2alpAwvtocNQex94miXeZrhv
C3PXnaNyYRmBgXIrjlFU8bilUf5kMOftVUz/usBeBW4oHe8WTOvvxRyU0+Ds/eB95Wvb1wreAp8n
K2U8Pqlk78P2/TkbRXtBI6ClUB8FNjP5FM2/R4f+M+0G8dlEsbaBcyRHzIIDE44T1sadnPEk/iUP
dxK4Ced2thD0m3lXF/cOZqJSIA1SER6Pn4DnrmW7YUpDfIWrcr44siQVKQFxtFIJmHnayK5Ck5yB
1MiEiOz8+F1e7A1vRzEhSVX8FWHzzHZwztHWiJA+b0mN6GZzpwhd0JAfoesTsHN41Zh4gLEb6+j2
DBox4SQwD4Q8IIz2mlyeFzvz8E1Ivtt88w0BeRerXkxqG1pCfZ6iCYlKooQsmPBkn37zRYOqqqTd
4TZLNFjEQ0wPlCrZmsFX+8224mRdUDbjnDiVYpW9g1oedjg1HGcFs3gg01m/Zt11lQcgkg8uAbGs
b/eXX/D2/jO2HdIj365rP1xAMfGMMPomyVO6vI9X3bEVlcKoaaD9XBJI8FhgRw4t1LRWwErr9FG+
Wzplxh50Nt0HPPEEqLOcE64e5OROpBmrFVh169UKX9y16zXxLAv9KK7SsGG7yfMFYgMWivBS34sP
V457V/jZcsx+jQKVzqq6yL3C48YIKYu3P5EeG+Jpcw0UPkS9oDye8e5Oq8sBCnubBeHblJuzCwnM
pFpp/Q+xet6aDSZVnobbESFOnkICuPf8lg7KkXAIcQ5imHvTNPq6xaqHk5+ZWKAP6BIY9x75bl1t
TLPADrgo2Yk/wpCKd+1DCJaKdFu5184+aMpxysd1npBP9HnsaIkNMcjasBFeanavj3vvvodet1Lk
mmLZVDHuxPScgUxhilRrhn7CNCQsQ3d+QHNGYLDwdjF8bpZLBlPOV9HnuAK670gAoF085jwJdCvY
yiL1OiixdOsntuz3IvaSKCyt8qdyuLc9VtHSB+2dNe2doHhEV2+wsxQvOWYHVxLC/9yXO3XojUwC
OZKfasYG0y6F9Rjj+hcI1eE4fCL5oSL22Dm7y/CajQWs7A91zCUZdgHHhEJP7LkBKGhW+gIhj6DJ
0CauHXyxufpCg1LxIigRLRiYazsAndrg960oKU12f7+SSAxYVieNQPcqXkUT4btCwmAJKsd5PkE5
xEUXF2cIeooJG8SCGWtVyNBNT4l+wrMagCUzF0kU7zjGkj7yxaLU7hZ2Tl0uqCLbjbnH6m+Cq8dz
lLY2IogQee5x//U/fzsqI1tLbhq1clJ/bI3/4/kTcyNoR6jVDF40Bb2KK5e2M/TSYBt+UccaR89I
3sGP4DuLFdP+xap6dacdKb3p79y4TGBd1RcrLYyIptUTFJARFOKwb/QwqUWtnZ07AapmkijPmbYP
mIJ2xNUzKtfzAEC52UgcysqZMsNbWOmGFkN3FNL1+vyXDrZz6Z/FCpq2tYMFOBCSENXohau0S6x9
sYwn6ZHzhp/2VQYUl/rLcxhqEsUQzM5Lx7CYzYXT5yllR417bumjnDRFTOELyrNo9mdnJPeg0GiY
5BPZ0ayytXUJ4prm7ixAexebJjoAE7jqIlBWaVWfzh/+1E3qE/DChPKFktSMC17G4Qnhf0Uo9/vd
86zliawG6Fgn8XsF+qxqEUCjbAD7TbTOkwYTt5V6LSJZ1vJiKwEMs/i7cxtX58pDw4HvN4rsdz90
N24HDFv1Dy4PEMAoVd0LhqozPh+HFUpqHRbvaVksSD/ycWx11vF7w+4pHszfrJsjTtbcckOQUGSX
0uNwsZ6z3AWfNBMAv2pq43J2SDcNe46+MTCvTiDXo+rudbl6m9arleIOoN9do1K3MQqDzDVyEKKi
gTqTsYI12FoGGnjO406AKNiMzpqsJLKYsOZBSF9FND/CsgCm2MQ3hTx1CmrDvAz7A2K3BLKzdk28
Wo7I4ZUuGtFLlnLvzYfHZE5E9t1Mi15Ta72Ku5HEw0NS3O44VkwMWdooV0jguh0DbetR4jK4rQ/w
5aYWyOBvUH2fi/rJbN6GunEQaCiKhEUXzh24U3+ekGDKBHPeOL2/HC3rz9KdGeJVE0WFJO+7Os82
TNtKxLy9x6VX5OQfRCuTiXlhzAd1vrdPaj9M8soig/JpHZVpZYpKDVnK40ZfYIEVu8eJS/2Sgsjw
9BouTvEJAUd3Tv64LxRcnOdWb1zRF3lQcJSkWpVO6vlqFoqOBEx1IT9mGW1Rz4nCfxWWQ/qJq02E
z3BMPnKeEtXG8I52QOLwh78S7+jzgIe0nG0HcZbJa7p1qlcpdgxkDA1B6m4NZZJoKHDeB9vLdVNz
uyMdUerYoDxE5sBGl2giduSPWw2jzjTXsATHSINxf3Qjw9fhhLUBdJI+HXVbkMDL3jaBA6jdygQd
+NmiHOIGoO14mCyx2nu07QtDNKBe1SNjmH7ZxUgE3o/lPZ6WL5mtif8tFcf4++xtBkQg7KPUmV7A
ueEqyl5sWBMwJ5kYCX6f0fNqPSeCsEPnPlJeYN7ziSjSsMqe3yiIExb5eIum+CxWUNXnHUxzpcQz
crHiW32Ue8GDgPTeGcE1agilHsUY64/4hBTTEQ+M37S1lSLNm5T02Fls5vt+g72PjxffKaZLOEIT
iE/hv+Kfwl/3s9DChiulXdS67tHTKScTTv/QvU5BQNKoa1efBoUxLm2abB/2USirtZTMAdNC3D9y
lwfbPbUhjQfCIPy/9m48Hf2dEy261qVpftuEz8j4o7Or21C8B8ibVCPyStmjBQ5GIBcDQJL+kAqE
/5+s56L+b1jOpiFAHyueomm3cD+/GyribFIjDtHBeKjDGexGiv/ZjWwjQ0O6JtCG4iVwZOdzVpIi
Zx1zUk4WGr/zftJnbpf/hlmUYlyF8n+3+7pvrZti82uPxRDHeLFm8It2qvBuiQuw2YALS/GDf+AZ
ksvLC2w+9eCBrIJEC9vj/iVRyyU9+9MpjQYnu53TdagAyOexOts6Un6gVLnGCOwdgAYFfbx79ufB
coxr5Q3BX/KUv2loLVibLIy5anTiZg2u4h+DHAOtC9IopC+ggEnn6ywq3pm0B0TaMTfurcYIBLtG
yc7CAwEO5UyxGe1SfxJnPqp8mMjB6WCQx7MJiQhSisPvfU2zEFPgsgBMhF9tqPvpuXCL2woJB1TY
jGuBef3xiM5CIWLokoqbfb1MAwB5+9+ZCHPELCa/9oPMrI5BfJro1TjvWs/bt5h3FPTYG9nSPbk6
Wtjq8X2uNJOXcfOikr703GyWbb3vT8lzh8o0XXDg56Xi+RT8oO9afFJBQtsB5nmdF8Nc/VGDtSFE
WMweMB7LmyQ8SxOg7j4E+hg9qTEz93DQ8c7OJVMwr3Irfhemb2Ol3i/MkDRtwCiACtwd8ZwgUgB4
vZFaDCJIpLvPC1YXs33+T5blrxEKKbLmvUT6/j4SWfgopWV9F5k9jz2URFGUcJ4qHNEnD4lO9a49
LNu7Drbf4QoGrElheJjVFr/mTI5FvyK+upX7CrjaCoWs7qxxDw8w1ep8BjGx7lhHeOSh7BHQT9jv
gVREkX6AB39jsLxoCy/zPSCv+IeOZuptJ/5Gj6kxp+xJINYS33BVrJG5gkyhLNjslpiOvnxv5mTz
/2GIMx1TUoNC4NoBxjX8t5ruFGklA6nRv/Z03YwW4MYcvzK2ZGO7HRjU6LOCN6sMkBXrYRP97G2Q
+OqezN6B3puql4Hk957O5DNXG+7e+VaFAPQRsGq6MAFKzOaw0lR0hXhSEel6441Xc3F7kKhxPBzX
AzoE3XRs/P/vHqTsYxTTIPslbi1J/jj8wbUV+RNR/3x/eH1qWzYzVuNWlWg6PHLOX90b7ULXzgkL
eG2CHZYH+XDTkskFcuaKgf+mSwmv2EL0MqF/kRTg8wcVveOCcTLS2NrOcOiCueEw7T8K+dMyhBzV
9xfxD52x2s0idbTiSX6Y49OzqTaU8xlZP4QsGNkmwhWTAr4bEAP4MB3ycUpMk3TI1PyohUB1/Yux
V1pNEmScGgdv5z/PUVLARzyLNApTYXCF6DBcQVvkLnzCsrw49DxyEBidB2ULo9zVMmrOMzg8/q/q
1rlcB2xiS9+jMnwxSsQahAI+vFbQE/yY6mgCuomCkywoBPHS2aCRUOaXPMu0s6J1p6Q62Cx0di1n
lwBgowyOWIaHxgBpykCEpHDxukPu9LjmVc0i+Lkzhry0IgJiafPYfPwFqBz3rWzlsLhDPt3gCJ9h
oxb1jMHHxiYzmAYSvBt2xEkIbkNacw0yP9OWnOkdrdcuDDp3RDE0q673UPg6RsbVWALEqFLI8sQy
x2nPUREvdX+j3iW5Ld+1cWVh5Owh/d8rvRfNrfMVJ9CXvbyq/bBvvQIWNFrfrMzLEPMnXRGR4HDV
V5hFJr3hUEHZAWJuXfURyYcTCbd2swDYtwEV/FcsQjfWcwIE/yHt4Uc84mUJ9yoo+nLU4Ag2KGwe
lkAm99SmKtTxF8BJMyayeMkmR34cukxKxplV/weyFhY0RA3e0MQ11vkFNKOP0z++V10CifU3k3gO
e9GgnZ8QO4KLhkDyySPJ8WirdWE+jVJoQoM9tTiMvC5HnpEDY2Z7fDIIzmn26SZC02SnlCwUjeMF
WR6F96M9oCNnroRSx39i29kGtN5DvUv4fSxf1EJfd5nADqG2/TLe+JBjLpO9aS2Th6oa7ZBobgaY
M3fxyqi8vikMgtkmMGLvyn7PKymXv3hpz5f0gV9I4xlXOQYlSoriHL4ZWiTG+9G0ZrsuFcTWRrRz
6XaGMKLo8F55U8jAG5cMAaknyq0Awn/PYglefpRK/DB89Q8ltrjiJKLVb0B3/NMUIawFbZAhXtEc
vQzOVjCSYAyo+wugJjl4tVhoe1yOJiGPbkVBk0lN58ztHzdaycZj5nrdjAArdrb/i89gWJgk7c/q
Xpqc9E/VGHRJsK5bzvK4r9xFCziduhKSB0oqP/kay3CYkfx3npEOewYvfBFcYvrsYKz0SNMom+fv
BJjLiFMDEQD/xbw1glHiF1nuMrBvj2aFqob7B7GE66blgT2NFkfe7/u1kkJDdmH6POaw5Bc28fIN
+TLH6iF5YLEG8GJlemKutmf015EC/iDcmOLj1BtSQ7pFifDQ+3DvTqbRR8Fkj+IGCyJ4G0qG/qDw
Ell2gl5mHJIHUdWRXlylKjA321N3k3fKux5KqzuCH+RsjMT0/aKOeSJ/34Ofc7xbfSHFjN/ZmVf+
pyf0fHAaWsk1GE23vsbIMJULhDXjxOo28HlH7XOjFyxy+I4XyxitMDJm9o25Thtdq6ZCrvFSKJoZ
YUT/gywIWPCsJHsgy3iqJDHJ50IY5vXBDnRWZPaeCMMUPvQu1v47AD6a53qNZg/3yNGjIOPwMvaS
MEqVnT5lRZ+J4v1h5WY86M5GbWFFCCHw+RXbTg+4vLW0OvUO9Bj/MRB/6lkSomxm3KPheLHWCUNn
WNCNClJu5ERwq5OJhr2j5P8A8bQ+DtGF9w/F6w/ZDt0stt41ZmrHr3NBQAaLL7Ps95nuNr19fa0b
cAsPlsFjIiuMhqEgHOsS9OhkE94hnLFpB9T/Xq9R9tCoYUV1VKk0+qV27bjxC3IMcpgXMlAQnkzX
pGU3vKBlbwui/MUv6Rd+25viYx98mNbxBjFbohR6za60jNL+D91/VBSv6mpQuAnOSkvO0AF28Pk3
YBSx1vwCY6mzGUCnqQizT0G7sGEiQD/xUdvWlzV51a5iEL/S8mlOwfQpeTWPn4a+0vEHFiws/rty
VDfKm/TlYSOgu4k0VHDoNx7BCOzovw4kg5OUMYdOv8KEBK5ZwCLWsODwQsCH+DvnZV+zAiZmj60s
4ieuCNK5d+GVkOFzIIRTAYbmZVTQy31no8KQqA2/JO0sMsTl6oD+64z24ImY6DqkSHQE1RW14kCX
pUhO7E4kK3XDJw8fQrt/pKn+kXBAJKwbEZJIfKoRXa6fneagl4Rg8NgTaaI1j/7/42nYUdzYsjVl
TKFU2oeB+Q9Z/6woZknzT9oNJbEeBy8iJqoZRftXwJd+6szcegYO6pvkHcX2UPEKG5pyUsF0WEYr
6CEyZskcxR2BB2KaXS17CsPvA9shG777Nq3hqX9zt5vK2eFb8x9uzSz3w9HY2he0obLxz01Ti3SF
slXTq9sDzQVNAeiaJq+Re3Dkd5JZqrc2XJkDceuJ4Rn93AvxG81/B6IBYN5IW1KXRsab/fj8CRHa
Bt/It1510d5LRvjuwp1rhjPaGAmZQ0APEEw6LfRZpRKA06lHK6LIBnmSc5QC3YpkWp3ozYPRIDz3
6fcPY2XxX2GIKynzVLUo0WJ2xTG6nOeuogDJS/vRUG0fnBpANW+Rx/EeQKDjlLKMYbIbf/wxp+B5
3Hjd+CMC7suSX+RtjiI3/HJS/SnQ5kbFBUKrSXQs8kVr3ZvHAauqvKQNNvNXHM3EsJntHpzYtCYm
EeMEx5Ff16CHTnX5vWf7Tq1tkaDo1vPwRxwMvsQPfXX27rQhW/yS4T8nw3nMraGn8Nk+o4biIAJq
tgI7JS0ZtdxHiCX7PK8T/4myz74ZDvuJxNNBZo2fph46/4k6IAf1p4UhMh4NnxfuDFQnjwACfTlI
08pVzT5+gr9yH/dN/AjgoKKeqfbEMGMyQPGf/6iWIbLBnPzyWuZ9d12C8+SubewTxbvnhBjHdeev
C3amvdobvm82ITvbdiyS7QjtT1ZTpyg4UJ/r3fYl6vkddCserRucWJUeu60/kzKyx0AWgmcKhjB6
touMitjxjATJ/0SEBiJGr4ISdu8C+qa/g7vElIoD+GACDwNB5yssWBTC5NkDBNJYqRwj6u9wW0H3
iUinb4KCRa3E4SN4O9com061j5Fz+k5kgZRFaTvzPrye/ktWV4CR+EpOcA2N8kxxvQM3VMLDFfLH
Oq52jvL+oeijpVWTJQNZgNBcLbXpVaJ9Z6SWsLdintnx9U0X9tG7AbCFum6vjnky8vr/so8Zti8E
m5khCRlFkPADRF+3DwoHb4AdfteNw2Sz7Tw+kcCfEF/PA5P+85l5mJ5VG3q3eBVRsgA049sxm3/A
e06sa9mLlfBWeKI2B0TiOVocVlmrwSCtIDSm36NltmpjQcDTu+PtrdlpaEgeUh1ykWmCN7kLWwab
Y+4LnjXMmd9tTQF1L4GKBTCGrAaiQ8dFcvrVuHBIPxIwj+JuBAeCHdxc4ArcB4+rKilgwOG/MBO0
V6MTlg/povA17kpIhdXqfr1gFLn/g9PCcLOxrLQ30a4Lz46ugcyKHzTarSVXmTaqI5717nSqXJoX
447EtqlPk3ZoMqCG3JuLeuslMm4IR+wt2E8rD5Xu0Am4uXoyr8MVPu1uv++KBYA/r+fYASa1nhRj
PrtKWswDMeWIe/2t6hPC2yCQyX+KzqiYwCbn/Js/k+2++3jEGbZwfHruLOSmF41Yj71KPYpWK9Jt
J7shnq0On9gV8DPqzNVyWgd69WVmt06i86AZHqwiUYdnCDtJkz6l/dUBZhEv/mpp4wS/jKTM98dp
lJAsOYVsm+jL4Ldux7w6hTGVd/kZC/DNHMsxWGXBFOhVCA2SpCREygOKn+JtFj4EYvUz5Xhm/ELM
blkFvnc21RCwCCpiOsC4i6a51Om5DfpR07T5/mSE2V1xmX7/ejLue/PvXm8/jHt62m7zx1qlEqg9
oCGXGlhXmQGTtdjoGZNYTziJsB/rU4ftfkb01aYK6vSYXgdJgNxvpeGI4YSzXCp8UrLNcBmUy/LO
LsXaKOImzLxDxOixF7HbjOwf+n7ZZbJGMXxoJ2gMtdbtxYVx3q+ubuiPX859dlfJkwh8hsbKGDlX
E3JAIrou46vDfWFUJ5KJS2gADDjWAzB8kKqWhhNBty3LR4Df6DGQXvll9iifcgk/+mkfqkIpUPA2
LJgCxuxtebA3Nkk1XU5jjLlQqkaen8VLyqYF/NUuviMdIeXa0qKe8ki49syKAkdXkkEsBMuFf4W5
y7B2exHI4AFW6nqcskyu1OD9+oFNeUfEZd+oLk84oTSpxaKoRbWnldDR70aOISAc1oxBG299TIwp
+AcRgcJfFLwVszYxoIVGkf8Fp1wNttIXkGbzcTfw0W6A5vKx4j3Uu0FJCazrXxxwB+QoH1sTVAb3
OeKB49tgTJznNrpFsY1jghViwLkhY4NT9VuDv7sn4u0zOR/2P1A5Y7NwKXJYdXEGPwPmwPSunJM/
x6Q7hfzSKLezIFre5uM019LeXY8jU3zIwfnZcOM9FaDmlHar+xi/HWusuYxRQFWAmklAuMowhlio
GDmhPJZQq5K6gEW4x0L1cx0P8D6hSvl9rT7FvGjkYX2B3LK+4nQF0ic5rHXJIpXpAvqWKm8VCLEg
iECaqHh40O5zJxeFXFNw72l4whNKQuqQvgDAFgBNZIG3NtMRwjCc10AluIXJuCyrrvDZyKpAZPIx
dEUnArsoQEX6te6QEH/vnz7wcdHgH+PhawS6+xvnD5So+l7X/NtjLSVLZ2p0wpnN29IVE5Granhf
6piihTdFJ99OiyrUz5jcLHAkc5CC9uReMQ9WPw308JOgofyNokXyyIwX6zWBDIVnFxgW2n/TbNKH
BNHSwCMYwOLGPlpuoatddQbvog13l3/QOoY9k3wbESsBOGHinLoRaFU4gH1J29cxpVuiQMflLj0S
lpLxhJu0vzcT7k8sfZwijRVjbwuUfYsJjAnNFXKwtkIUOKMjiuYoCy1Rf/GnRvTALemzwS29W52I
AwNTVHy8RcQGQ2+SmSGr2zQRtU7syxtQgcmjKw/Jez7Up4UYtQMbOaKvVnwoaB9F3cqIGRYzgw0x
uKgezr/vRPWY0fk6mh0yfXwz6seQxG3CNvxauChYgyEFAoLWGZXX2YJVKWPJUzDVg5W4tcZFPfEJ
KGr/gTUbKjWoJ5v+7IMnP6jbastwsaT237nmRjCDDRFSuXC0wEOIHjDJrMqUjJuT+ZPdhMQwOhl0
6TV9SKNKBpgqx4+tOnbnhhcAjmcYfIbhrBp8C6Kp9cN/R+fOSLff9YtpYApV/P+PJ9cWLkJuOd9X
NSvKAdUCQMhoDzo0xQ3TfCrHPCWbHJ1Uh/QhzrYcNp4LUGZ/W98xq/N/2ex8ViZTe1IZrcvk4adZ
cfaDxGuTlMjIy20hbKbxuXl3UTDvexTDqlk3oGtaoCEiKf0mNopFQlnNb6xHNOZWU08QYk0oGk/Z
1bphFDSlrA5/3hqCI4Yuoi54hfhsvEN2cDtpJX87G75LFihmnyM8Z9YgAunxjen9hVI1vqDUCOuN
+Qj0BmGurYrsTB4qkySsJlKyyGFrvCg6QChoH2hdeos6cREP8NwJy0AInE/CqMdw9Lopv8jofR0l
cgT5Sq5k8XNNSic0JqXa5frkAg44dctfvgO8G3wj5T475BzVFXzMN6Bsnt2Npnu6DqvcKzeUtvKi
K/6Y942uxZ5OODSaXN4GLfgzroL4QMe33mUhvz+Ex0f1un38Slh/y5scA//H9kB1s/gdDxI2bIlT
si2GSwcn0LOV/AaSLMSf2guWckAi65FtzdCYnLGTYmNY3fW1P/z/S9aLs6BzOTpVoF5Q0Og+hXWt
Xz2hkx/seHGtSfF7jzTHI2hDgBXnpfvAZSCjuq1nHlmyHabgKk6HDubEEPC3r8EMwvan1WXTGdtL
JxeMGQMILFtLMW+QWy2Au55gBkJwsmAaUNUJOwC5AYk/knTL4+nE+CLu96EM4HdQV2kJinbA3PqW
s7pVdNb0PsICRj+C4C7Nai9ijS1yNx7rmExqZBR3ubxRkYmGcgVeud2GXYwSC3jR4EK3n+jryVaJ
98MO9dEXjZGsqvy9SOecrnIqQ3FQBpWedjuIaG+C6qx7LydRAjcfOR4vyUFwIeHNRhxSfMHikLZk
EcriEcp/dGslSlhSU/Kq4uTfwD4TRt2RmwacBJ/ZdC2soZOo2nTkjZuoMN9eNEqpzCIqPBExkNmc
ht3+vypvnO5tDDmIx1soHR2KfaQ9gXgMkQ5u2a5PllT/3hlma2k5zTUEeebw3yPEvyHc9npThiB8
+kiO1Lnh8/PbS+4ESBuZtQipLJhYqYHkBI5oMp6DBxYwa917dtK8AagpjQaL/5O/YE6h9SEhZQx4
Ky+IjNcfppk+JBZ3by4R+kCUCQu9SlEsOOA5tAqoRvUobEQDVLqpA84ymOWshJrsgKdxfWmPuQBy
oTLdaAESbkQXHAVCogbXAq47eDmwcFd6CC0AoYjaVe3N+Ucz2605zzNk+mome7eBBY5pDAe/zZ4Z
NZhcix5XyAJaFTVmAzHERjyqsa82ZAU/IlFQBV0JASZtMVPPwwXBb4o/EmnMpr2lrC1ACLQUGDAw
ct2Lis/p13B+TsKT3pCrtxy1DXmBvWWkRFZc6RW3iROnBcVi4kQCXPTAcqGC6c6nkfm5zk7kp9Ym
ezc5Tc6RHCydCRJh76jtmXOdPmC7e6+YytFPCDy6Cn4X6c+Ec/cCFtiWErax9vxe8D/Wc9ejI7iI
8e0pYhp8OsPgMcKaN/YzlXbJu3HL8DpKqUeqGjqityelMihZMtxaVww3JLhj6BQQfdKodhBnOMT1
WEqmWey6uceaxNMp5bZ7fAm43LTh3/ObSWeByfl7Y6SbdNEATEvj8w451x/Uj1EGH0jLe/OiQwkj
Tq75Dt5gUjsCi73H2BQzHco/A3Lcj6XVhBmO/cGlFuBDz3hz2fgcHFLLW4MyU40AHKXRnNPFaTtk
ozl89YdHIjjo4/1mAp6mNCs8owVrJNztaHntaUXN0hNnCMqe8Y4b5Em0j8cZk5kObKknC2qxMEUK
pWHtj4TDabb547sDvq7kaTXzAAvCIKsPjsrmwurT+Ck2PKapsEHWoRyOnOnzUx352GlT+tay2vbi
zPadcPN+f5st/KCjg1H9mHpnekOkUx8A/olphwdywVw9jXkBpUxhqSTfb9DRKeAOEPkImmGLVNTo
+dEvKaFyaqe5BQeSR1VZRqWo6kay0N+f/JzgJp6nJrKrbLuStEoe4iMlH9e5r8qzUqv5K+tmTVz3
YSksfm7RQpYb0hG+ABmpi/Qot/dJWqVZenjEe+YEoJWBWck4NJzRH8t2zDmThl9Kt5ZomCQelP3d
gN3LtSwIbtsyEmgHJCTdvUlFHmQ6ZjEIYnU62AZr86uGIdLY6jMpoM8bbaG2GhAclrwTx+XUAjyE
KCoZzp4MoXK1d02HGmDbNl4Dg4Xt/fb+TcQrQuNRSxf/wvroksLgf0dHp1rfaaek0DDjlDRKPSX5
gKcJctWh2Wr5hXkEtHbw1vKUqVl8Kqdjcrz9Roc0A7hfXhwrzkNGLf2yvq1HqD1Hc/N8Ovl1Pf6B
uJ4NCfJuXE9m5Le5VWPvke8ETOBvx7pI2bkvTd2aPIQrOyu0DDz4mts/TJiiYi3uD8Mf+4Eu3pH2
T1A+Fvwk2ORhJO8X3yaBblnQDmOu0sRP72t1NIjgU42oqozVjcHpWn5ymqTXhniktSYpWldzcxb1
KWy84UfQRiOdvfx6TyM0JwcKeoo1pMZw4DUSneDS+fATp4Hg0ch+g5uJK3lLHG0PAcy05vwcPPCj
OwenY8+2sq+1LEi6gY+qGTVQn2HxwZ3a9I0kWgy+VAZ1adqUJFKHmjLS37OFPq7Vj9tOCiYynQ2H
ufx80XNrjOB1vLs97wWM0Rm180rLgYDFtPjpPKOhGeAQBkttqIsZHmZ42/8WFoYsf3drsQL6xVEF
Cm9/Vto6RPNYBj/yXQI8ZPInepo93bPQ+MvbSc7d+7i01nfIrFkyCSD2jzqAm8TWrWg034M5E+vo
avMKhKTUr6g6ajPzTDZRc/UgYhRkbetAjRt7TDs0VFjfT12nxv3KCa/MyZ5hF/vkzJPUflocTZVJ
pSiRYpRd+fkXSMe1Yix7AGjpSKJ2Y68Eq0ALg9iOfXYV3JpcStht1LuEEbllmfz8eqk8dFXqjXJV
DfX2obXrT7HmSQLJVuwTypWxPNQz/DNMdQOhOFiWe5B1hXqWHBLPux75/eSERm78o3/avPZtRFUE
KPEIQICOuOX9gi05XTpgV7tryWgYoOviQTZCWyp6MbwJfGAOBYSbRJlkMAFTgWXneqYt5ucI2VFK
eVo0FgTmrvm+vwZFn/jkNJbx/pHLntdN06oNwhDp+D/G+ommAfoUtspcB/MoZkT2aVo3zAb05a+F
joviF7zMGLd7zVA8ant7/FPJOfsLnM8xoFH4McRg+129NY2geIHUjRWbYFKr6H/sscz9dXBBpc7f
fqtPzecIH+hG7EbFqW2N1bukZQGQaMqGIyTSVifxVC5yLb68tkiJRGG/+BjfwzDELW4aEN/qqAA6
LAVSGuwQUXlqHOd2w49+bmFBV52m5rEIUQPlx5TdFfuTN2snTS0y+OHmObuE6AK/XkiGUVObMx4o
bMSxvKXmbxErAz8CK/y/47NTl3CT5a07Abc+MgXlN/KdJrXA4/g30YIWftVoXHLhLtDDhVJ7DKvm
QwAC0fpsciZuO4ICe5YwYp8vJW8DVYiGCnIoqrq8IjD35jz95ZNtb1h07AQbBl2f6yEOjJ3o9QBJ
CTsDN7DJTiwWbJcdJU81Wpy4Sg35Cjv8kZCg2KMka6VWK+Fbh+WejJDhduGHw7xdXpN7IDF4e2k2
0Vpbgy4sTMi/U64l7xqpLV+duOpfMHD5OFkj6NEBaFc2dWt+pxVvTMVcAxMllhGhPZeyTvWix6b5
hYTOvOBn1YmashPw/qp+baHcPkimzeQRwDEdlyThzqDOu1oIPFlTH74x0A+jwrO/1YXLc+GtZUOJ
YkQNyo8IO0qd+8xjtZkPl38dpbMnN2yPCoKTJ66Vr4Am2D1trfomOYTh7ZQwulvW+xow7uhMTVoy
6tUYkoZBX18rd/ltPFmQ7bAxbOOoa6DsQ4tDCOu00G4BmYea22eRwWxf8URnFgw57KkZWutEyE+P
YP/Vw204Y6UpSfo6jKcEJoFmFusVJE/6ObFVIFZAmrhbMa+r3Re6oEKQZIBL9cQsjdIGmB8CRBkY
vaqB0uoqp95JvDcYgsBExbF2WPF849xD36urB+ndLZ4yoI7leUFPTc/EOpX+XnIzqpOeJwicqbeC
RFgELuBnui0qAWkZv0UtShoC4q7FM/G0y3jKkVhUalWqNItA6wOvJUJY27dA04QAisFEtxybo5x4
t1NoPFx0XgIFdh5kBgIfWiHWG7kPD4NEqy+4UKgYaOspUkmgnxGmLK2VkcFPpp4aSqcH8/Z2ewwJ
Q1cUdmtMvngMqpDD3HsC8mMmKZHiZ2QepZvggOglQcqdEaulhqqdb4PmxTNeeJou7OAMPmv6Qznr
/eZ0sGnKPCjnag+sq7DcCs6nM9tWHYwm3ka/Vy0ZyOTP0pVxNKeA1/BekeQCamF7M0AmBf5rmcYx
pQgucWn4ZrvBR4MChdKtxfkNSKfe0/MgcOkwihaDpUHr1K4hh4NOvxvKtaPa22+Dr1VyF1KxI2rS
w587DN/kzXl396yl/NiG1wRIU8IXjJ4kXNfeiUlAwg2z4qn95LrvzSNmLlSy2AvXVSGRv1T9+ljf
30rQWGJ1c0sDP5bMTf60ozs3GLlnR1F8wFlfjGZOB2+ceNc59oxEKAcbPCOd5/6jmBsBYGZHnI84
QHR1LWTbmZoBmZacZ3/aGjxq2U15hGx+VWAqC7ktkD8xIJfVLC9ZL5cou2JjxjTBvLoK9OnhB85Z
XYywAZjESUCa9E0BmTv0KYp5xKFUBnvVQ/+r/y9zDfU/N5L004QkarJJ0ZdRoVtTvOMrgSYUHf4l
8d0+DXcm7gfggZmRriFKzeU8eBQru91/+EGCrCck6jkrJA2neCI4G9SSAld0B5U56iXhJdi3Blkv
bJUJefoBE099YtA07rtGHszHYygdoLd+Am2s1Ib/RQzlr+4PiCpWwq+kcAyGPdwI/veVOZ10PBwl
K07nc+1rV8Vyt9S+yhNP2dx4c5PlaeiSiU4xKWAs0hcqn+d9srtYdkS/dLV+w1BoUEwwMk2GnYkJ
+DdMFsgA1Wo2++yItLQs831+isDnKzlzAjojtC3WlnDDAXb0YkXyYAXIiczXWmDmDcNl3Rr75rVz
QDmUJPEvCn+NS+Z7HAryrobXyjblSpBwHOjlMTq4+gZrE1V8UAGLpAsDeQnVuDwg0CAVjh1HIPDF
P106ltkAK9eYjIHjRCimedGO7VGLjLVZMWnOfB6w7u66Jry23/f/e0sGVY8uQof/H32GAdUmEjcn
TCuRIP3l97sjsrDDrL+qdVbweTcMOn2mRDwTLQzAxz9H9NeqN1zufFsi0fT7AveJjTlgdG9RoDZj
ZGR2r7tr4lguc+tpmWXDAhn15d/yWGoJpnTmMCY+NEshQGNLlJa9aiKyUPldQrCh/JnT39Odoicq
VGM0yB3ktcecQvsHs8To585KG2HzdfW+Xo8gQIOhziwqwF1oDPII6fRaFbGg1eDGL1sb/VQ2XPbK
G1cht41Z3b7cb04udZ9Ylxfl/z22LsgMK2mbIAldeHt1TKuePTGvMwQy2xAoU5KxMNvsvXvrGyDA
MtjHFFr8CiZIWGCJ7xe2i8hP4L5mcuaY4YlOrsu2Ldcc81ZsOmiOnGFDNoEYR92MhLevVNE/6rnR
dq8Rzd+MgHLPoHO7lZF+ogxmHOfqV/0b/KFu/rW6A+FFE6ru6cCALAzOlccdPyiveXUmwzBFITtJ
Oufe2SWQOTtAkXFv8VnJ+H4iIwgiqiFHEP79vJrDX+9yXavgcYFz9T9HjRgZJHG0c3Jhsr+mW+cU
33yLUyzLgHHSa052FMMLe8J4WM62iuPsRxWbjKl52idEinUM+w6RqyG1dOHtDC8VYjTbBgf0nTXF
ygvOJIZs52YWh7B2YMMIwG1CkwvjxmwVmDeewAQJLXbAdo5BBEbjIGN1lkVpX8YGkbRavQn0slIG
8UcyNpQgrABoAsJR+N929Nlis7O5OPlJk9/oI7LubecrPmXIkfBd0gwnL8PUnyKy1zEMHOKasiaa
6JDeADcUzVKjTfmNSK6vHNXOIA1NJq5l58IIMeDAxGRR+Qod0Fnz9M9zSQq2mcPc+3UnULk8a07J
xVUvZEHCvsEYUADnrPz6RI9O0dYT3xhnWnOgD/3iqdzD8YDs5f0p4k9NpLotyh8ad/8jvIK0oB6a
ciso+3I/LYgGvLPtfOEwTDx6Zstrou9LRwYciCXWQ3fUICm2bajhYa1eqOROW7sIE8f7NGDu2zeU
j0pVaPjs3P1KOsXhICaYAF2HpGX8lE+of1MJtvb5TOjUQtvdGJphisFCftdBNFk2eVUaxxQmaNVr
DnuHU/q7DdYG7+EDwAta4ZVycABQuduh5yoIEUA/0Jw5fZYaQoRB0NxxUn6hNEjhXLgH3dxzIQds
2sbJA3v2aci7RUm2ye0eBkfh3KUBpNFZf2tsFbHmEczs/jjzTAigok6lClVaW9DhSzdCXKLcOQ1x
7oj+hmjhhiu7zmF9a/mTVRT8On8XHSZqge63pA44gduDxYfbGt/t3j3Q8NW5VP77o6B17L+HDOm0
EzlL2yfg6XZ3aAzec9kce+AluSezAHOXR10j0vU5XkzZ9ALkrYCq5Luy/b/5yKQl0L58H7/+jWqV
R0id+getJMnNBdknZoDsjV4iTozVnYKPfdKSoj3EWyQ19ab3FXtd4KqdtRrjUzrNI4ijKexwSCAA
uXuiAw3ac15Fk+x0obNHS+hZLZmFvRebpuyw3qy2gN13EMxa2nxBd4VMpdmdAPJd0P61sxMFjV3Z
Z3vr2vbr3fpx91FhnGMh6kvb2uWjl+gnIzaOCCFk4zACh6MZS2aO+Ndnsl5nuiuMYvk6PuvmH/So
/Upp+v7vhtw5+S/Y7Yqnz6d9RhbkoP088qR3If9Xn5cCnoMNLAgSuvXU+3QofQkHSViyj3zdGLLa
QwmECPiGbGFIZft3w25EXqAZS0ne/mY/u7crMZs3ADwYeU7poj/QqyyyfSN6d5OEzzFUD5hbvUdU
6ArcX05oOpW1dxORZOhaSRpGMkRTDD/CrVbXHBZx6R56lxItrAki85FEd6prpl81DIIU9vAlHk5p
HML/3oHDs8Exh8dYeio5gadLEly6zbJmYIdEP+dLPwgAJXUPCfWZwLkAaCst7O0ERcw1MFfjB00O
aDCLDgHtayU6JWRfNfBVy1B5Lc7ods9w+fM7mmEV6dcg1na84OvDHgfXSXlYCFs1mbNeVSC+8H3v
w4NOtA50548zbbI10eXxiXVmSxcuRHo16VR+mE+V3T4CvhLNshgFYzlpm0+9mG3syRkKMD70UTfx
AorlzRdUp89p/C9HUvm1C6f2Ptb8iRqOG/4fZk7klCISkYRPFUXzLZE4q3uDkehi9THzdlqm2CtQ
SjDc6WZpUKke3MAhb8jtFY4nEK2ftZjDj2morKByB6SgOslQfzbhOXzExlEsXgeMT3FzYugeoxe8
eng6qGGydfu8nnItz9WJ0E1FiYu7nJ12qXK5gfNs73LRj9PTGdmZGI3bXyercEcB9C9uPH+OG6z8
laDtKqIYkjaJjF8us56kFbJ0Pl1NGzSDG3guEnu+XLFDh5HvrtbLN5mukxWgmA2awbUGOoYMfEGJ
fDWE5nWY5VtgTCbIct42GRzgE/nM3o8/y+16C8Cy3qNOB8BMAgBiIz6VOI3cb/ol8AP9ai37V0Kp
1LRhLv89MAmRIR5dk/vI1YP4yfIDhoIgizb6CybGYYy5STJCJS+BPs1E2LH3PrkKNPowBQiounOq
+PRr56GJ4ujOFYU5Encg5Z4P9N2V8r7jMr6MKPlJF6IRdpGDy3MbJG9A9hiDo/+tByRxUkRJTU5x
0ILHCtLEzsyIeF2Mv+DEAVaWtIkhLgEh4sBE6a3JgZlsh3+l7QI5o/JbQq8mMMHH/tDwXedzfrxs
VGRNj+KjHPvcspV3zi+1AH34kYd7vRdF4GJWR10ofbl7u6GveP7eUXz/NP46TQh28edND5HJYihu
1vJmKxHgiS05cF0EGsOwxujCVmOgI+soDh8oo2vUx48LLiQdjvjiLMI5C4RZ7A1Vz9pPLyXpAjcm
0vCpT0n7LbN/arflf2lQnrLvvsnf9BRRWlc4TaO6RBFUfp8qgfGXXzbuTA8mp/KG1k2ANPCJl8kl
OPgn0xPL/LUWw3gognjETtqU7HRj2ki7dIUpBF4usUq/pFg9dF5ykyG+pfodh5hIHZOQfh5LM60P
m7Fff+it2ncFRDQc9+Ui7UDM15Ipu9Mrfl/7rxNHnUq3reCVUsHO0dUYeya27OEVovJ7mVYSPfFU
DNiJyHyRT8Hz2TZz4t4KmBFkJ8FMzCKx8u9D/EqXQ1t0S6GLtCw+O0YFplFXJdfWI8Es45SG4xq3
aE3KkPOmRerCkq8/4/CDmPTFKpFy76K8GUgxHsehmx3EA0X/rWaPLojhi3ZkICPtMnLMqWHBVpyu
okOho15ZMW0Um129rAv74U4g6vS4RzG5vnUc2RcKGBkIKRCm4XckvujVQYIsEGnuJaYC6PAfXgYx
xCkL7lBvuAHAE62NxaBiZqf5GJn8pGIysURfbRbmW/AqUOoeTVKSrgi/87bWdogIysKpG9kANgaL
6cLhHjuCrMy8xScgPefGbR9gOb4eZMfVNEvHmEvMeIoDdZ+YRD2pOHiEJo1jPi0CLSWALsyBPIT9
fZ3VRRGafccSZPNU1eQI66RnVbzDfavdt4B00OMNtX46DdBVdoRiNMubf0jhJ71H2rEn5UeCFOuR
1KFnilFmQijwaMi/9kmbwy4YZdCKIu/cdWA2QHGXfwcoULJfK/SAvmTAh2r9wsvRPCRFH/iLvuMl
fwsu85Yql7kiroWhVPiG/TZQTIMm+eZIECDE39GaPIkCMR3ZpEm9Yh9zbsSzr8iIIbGqLAf6ybYi
Fr1IA2Xi2ygDZJlViB6Aoau2m7/CP9iNQQ1d+Przr+LNvQsi5mzh6/QH0f9L4ob35NuQlNangO1d
gTX/oyPUNW7pPfHvsmOUO1Z5TDvswl1aab1FukhfSBz/FFyXXQ+2xWlyifxZIDYGNvmWnE9w4LKv
zVi9HsnJEKTUQmv+QMJjlRGgsIAfFdzcjmb1QT09ZP4SDiIVAv9Y2viBQRtQ0b7wfTt2LA4o/hdr
68ZQKzYkWvnBOcZ8ZjrbJE4xJ26O0/ma+WRR3B1TsB2n5Y2FxAMChAaWZ4mER1jDc7cbU0iagvaO
GeouZIIZGteY/HYnD8ymyiyo0nVVqWSl9GA2iuieVTS3u9lCqGSkAy4n6tl8aD65Tnc1VV/k/cgk
qFN4rapAroj116qDg4F0hY+58DEJL++BkdXAi2gDuhJOSNBreo/G4+vJy31Ah3/+is/bTLJS4zsQ
WBYOVI+BjjQ9T2ZQQKkJF61LV+HHitC6nQWMoTzZJJuB6sqAxO2x1o4lXr8jUPXjYM3iA6JTlDOF
N8emxnUavurbpdd9zgyzNbFpi6waJrAegZwevFO7w/2YeEBqNBGhmf035Kjz5L5MEdsuxLkDjvyX
8pqr8BrN7NIVVhAR3DZt5JgGBn9Sd1UhmuXnU1amSGmQVnPimqGa+TlAUl9XK/353bOPEj2MQfrc
t8Xkds5B7JQejOtljJxpAX2CjWkf5rOBCS3hAHNNy/zRIcVDE+BCvNOMm3paRtR7/Ck0bKhh04Fx
081/dPQOloSsBB27yQgBis8H12PU1uIiJGZp4qYP696nmE6iEIGkI3ftWYT9gVcFRlSoZAkULVz3
oOybxW4cbCKNXBJnZKEzWx4uoCunySTYLfTb4GBupuID+0SfjaZx3NnE/gjd1yCpZZ/ccDaDOXOz
ypTAI6Ebl24UsTH617I0EK1ivnL5gkkYu7iTTDzco8wiXChwbMUVO1cZLvewPbIrVgZJbNzPzLLK
dj8D0SoPilXwWY2ftez4KSrwLMQnJzXFxdiOUI760cnjxw9qAeE4AZDBrPCAt0tRS+mD6IeoinCl
+OJZjG0sZT/NFfe1OcJStXt6tJgBrlbYcjWPrsx8Felc572KFkmRPStFaJkfP6wMA5SrCrPDDG4U
UMjO9dnmaki5fJ9P7qSftOcdjlrkYojO3IlHxc8VGC4nsUoeaNn156riQNIC6Xrestxn5Q+DhC2i
s44W9fxfzTyti7r7QL0wfqSkpszp6bmkbFio0F4hsE5Q9OvKTty7mg0/6q1X39J2XOZi441fp2Eb
9+DPLFzDSbZBRjJfJGy8ch0j46F+GUByC5lHCeP9NSzdk0yUY3S4PX0Xw9SHAmrKCLDzWheLHpFc
ZqNn4jJqXERbMRJAFeRacIxBSMIe/jkuvY9/Od33tgkxbxDvTNyf/kkM5zLPeCFHQ7BFv6KFfKvg
zWP5UhrpGkknZhL/13NGPg3It/hlpKQR9JoUEMeW3YnQnTTsPOrT8V+VoLpv4wKn6AvsKjGxhntM
tT3EK3+Gl16FJWvSUjxksehiOLtq9+WSzIslqDuH0PagvyztG7xX0rSKTKj2r0CT5hpEyImTKdYI
8CcKWAQhSwp+id3283UxDWlPIX7BBnabE2wbk0SPVGZxxSlvUEHoexC87LIZHi9taso24j6tNjcV
ZgKO+niUcnV9kXoIseHmKbAWKU7yralJy0aSO+Ofxb/cf0vMvNb1uCsA/al0TbnpkbU613raB0I8
/R5ykuX+7zVhfwri7I+q3TD0AXKS5AslxKhOthdy0cjWXzlQlShLZc6YFATJX2j0leo2KDhTp4G+
P9aCL1y4mzbFOL1iU24iJKrW+jLe30TrTY0rF8HBNm6ChCNkjubT/5PxO8b13reWrM4Gd5yfoVsG
FsxWXaig189ybvRDsO1KmEnEUXIRcHqq2v9I6k7H/VTdLEWu1RxBdM28yLryHuOj5Dt1DFaN3w9p
KPwB0Lmbp8s5kHJTPsLcndeRUgY53cN5PII1VDdLcgsghMMevqfvFQWHFw3A5GlqvXITZDhBTO5k
wx7jXxbu7V8ETCrTIfqbTNsK0wlRVGZazmbbsEKr+k42QSefR3zyym81KcHGsghqm2Vkd83T6c49
89S9+mlnia/+yiOn0DSfes04pRNXQyc07gLCrMEWgZpqM4YT0wf1BxUPY8h93FIdj830a98xjbHH
/A5CnwTzyoBgtdmusNEHxNSqjoGa9toWCHejlepVnu5Wi4jJaWb8Sz8ZHZeFIvZKuq96PsY7ApIa
yv/qjYRGqYjg9q6sqU1JfpqY9G0dHFIEQjyjS5q+xJNkWpwvXtAk0FEVvq2tR2jAqSgCxYbLEAYF
dpi/O8hfhVUFfgw5Jx5Jta/uf3wJd9/cwkp2qbrusXHOR60Nv6PelLFWs8xiKLf2NMEwWGUA0dWz
mF2TCJ9x33jag/01k7tLH2/ogg2dZOWmC4Tzvbw7C8xZMxKJYo2YU7GqRCaNLyLC3NrCUhXca5Nd
j+y9M0Mw70Qbhn4WjOwgnqCWPc8gizEqP4JSgmTuNhGRJhGT6KHidJl2sZ0gJLQPCKuXvNLSDAjS
uaaUWbupEP/SeXbU8ioRIFyh47bBFnLoNRt7kW8j+MqaQLWClMuyz9fSoUGMWwzAHbL9RhxkXMtF
+SFfxVsFmdeekOKUXNfCGhYxTrxhjdzPE2PbvRaGg2Porl3XxMJdoOWuckKBUGW5CphtC2yN6boA
XJ3kvihnON56MNvOalL2uub449mFdmrDrvhVNG69TrxP+XiRKWxX/7A+WF/Jsjn8IBLx6PxayEtj
fq4UlPFuiMLNNy4840x9Pan5wBL1uP8ddCz4jYaouCfmg7jFD2Gjbf6LsQFY6mwO/YZPINGoTVw+
4TFhMzJeRygGIvSDk+ygWy6FWWEfKdUta8AyPC4vJl5oKd09k2ZIEgFtZnvi2BurSqwqfXg6nEH7
czYdezR/GkAuULfO5AzN3zDIU0j3gu97QnVlanvDnp098/pfXlHhEbJryEVlV0hPC9qXPNX+pLym
li6gt4VihskLJESZFVHwsA2bRObbqbWCoTg4hucfNdFehoXQ6aja2EIMzL755Ix7/srWhan5YS83
yg4pqHOmfGCpbBHGIhV7UZY7zC0WcQLrfYmS9zyNeHsrerd1HpZpIZ5AgsK4oyqELPj1aYYO7wV1
0SKMgHx4D2AcUshHZrE7n/Lh5+ioJF7ppwTCMepdeFwq//4i9OdtHWcitYYIYuWeg+jTjuyhGjKP
UNOUbdwI8jtO4AFsVmV8v/B9t3Qw8jFEosoaYpgVg55M3XpjmNczZheeRlupynNqsfP7vQG1ALSb
1cVFzo/q2ozI8d9Ffv3v7kv1EIcr6dg2hShoYUFgDoGs4MkIV+qvqR+RazIxOlp9YnU9/k/uCRdy
gCmY1Y7OCCtV+uxIvMeRq04cc+dqqPgbMz6OmvI+/num64KhDdqjy7PQJsEWh2BjEztP3oYoc3X3
SzjnB2g2BpYDpGY1l0n2TcP5vXB/9Bud/IdBNIcXrpbsxW2FQv7ZwdCorm3+Lua0MQSVhSfFmXS0
+4OOuEKfCcT/U8SqiBIFhPwE05er7rTHmh5YFSFjcnfUZAFsuKqL7rgBfmj1ZV77e72/dWZukni2
fgAQ/DxomIyl19tof4t2vUITOeOd2FeexShoEW34wyRVPVS4Trd+l35/SO6PobxW6LA/KHNqp5QJ
QlYq6AjcH9x1T8dd8rWb+9oU4Ds2akcwjbaIZ6rDdYn4OZQ8yXJ0p5f1mVsA9xXrTe/feBxOeE7z
eisbKBo1aZMj03U/Gj5M18phs8iMXDcyYTJSaxdVaSWyHNYdyCWisBTnxeaTEhwKHAoGovNHE6aB
tUauqsyHlArWW5saBciaicKFBOAU3ocXULtvjm7U0N28x4it4jP9CTf5nD118WPjcXMIPGfqcue4
mz1ocprIKK4Ob4PPFseaokrvmsXpExOSgVl2XwLykBSIN8ZdYKHpF24Il6EPMZs3D4um5J3oxEk/
sK0A6su7l1KIAXA+hfQ5i0ReaO0GnIZj0bGxv9VjcSczQ3oKJ8kGvvicNo/VsPhR6tNfrO2wRkjK
G/8ZCeZnm775HnOxfDDQ0XuM0IhEDVQHzS7Zlwi3DVZmt+h4hDuYb73wOqd66EQZ026EkcouiKHo
sImzWXFSgLAouY+3UnpiCjgNGTY0x8HNipUHN0MwPc+Mbbj0MF+cl5hYx+KpfYN3yiv590dA0l66
ZUimEILWc+NjXGVtuS+TXRPfjTlginJ9UUQC+n6nIpdg3hkHk4jTDOhsS02A3FBY5MXbORq3hDL+
KlNbrJ43sCpA/48ER0YeaxPgnAGaY8QMF8DmVv7LZHBUe6f+BU/cy3PCjwiETTUmjXp0KV3c1VkK
4a12MzaRdWgN8MLxBYRPvQSUDLf2xRoikF/VD/3woJkjy2V1GkLrU23grxKTP6shfFJK+ZBmV2x4
8oe+0/Ruep6b92HfAa3XqCzxzZV3N3JCQ4IiMnvbda2g9W6R5nn/xiOLECx7YEcZ0+lN8p0FdEvO
OBRwMMuw0QHnczAxows5QJ8r5mToOBWCkPPh+D/zZLuLUqwo+JDQVaBolnH83vEd95wb3/wtInHX
J5XdCqiVOcRu3dSszpSZvGFDdBUfsxJlMC76gjvayGhb23yFvYawRLofCqI31uvVcLVI22FkW1g/
v6knPLMk9DdMz7ZSzDAYQJtITsZhyYI5JPF15dXQkoimmSbAwgUsj3srI4zGMeKKYOI0gd8Yj+7F
Ga/CNlYno0BYxOwtYctff9LGG3F5pUc4CTvyLqb8ROvxEbocvXMtSfiXePFSQZz9YB29ZBWpSV3l
npl0kfN9tKh+7I/ZoB8awuYirSZv47fg8qR3meMrbxa7ESzWpdLgd28vU33Qwme2BBTKRa5mG276
HuVqgQ4nYlw7bTWde4M8sMex210HEF7czIey9kSsUhn6Dr53VgdU9HbRKNsdcOMdLk5Ze6lG2BC/
SKUB5xPfpHGY7iOA9fX9WZ3TWrE0kq6gSvlzCqRrEcBatuwNpn3gPGYvG/sXGzeM7i3H5XxNjgof
0oPpuEU6c1pWUOO7t5q76dlvpXjMiARoyLUs1B+wykSfw8JXVXEQa+FVG6ZT/TZLhIxR/NdGAQEO
D1uY6mOwEZfQ0MXjJsCWCko/vv8tDfj8gp2MEM6b7ASc1nzuRFC8N0My8RQoFGaWMP1LRih+Q1tG
yxY3MeQKvyVV/ZXmrdDdeweJWYWUaZ6DKD4hxKj5N0PTE70zJSe2VcRsoJLL1lm483DVH8l+QtSR
tx1b12hJGsnBgVAofvDr73EtfgtWMGW1ZF/2qPZfw+HGB12/wqJQALk5jyKn/Z07OcxQSaMeoFuJ
pZPrJOXaXlM9lUPpQa+3k6I9yoztKwTrAsSa1I+9ozWzCv7sqtuglFhqvgKEtsbu+dilKxzvNCf6
KgKON7IhM0aSMnn3WWkUSkMKF3DF4RUOH6A0UieGSDB4/vpTTORllDaVfOHYPb9KCUXSgQ4swBNS
C9qgFara4MNKZpH/r5iAUvseIvDTuFYCRREM7xVxUBLJ5T49tujC4DOGSIQEvC0hxQUIVdH41YPc
tugZaExu164qpREbP4hozJO68KFRBduXKDjCYVWC3IKj/Kcr6fXHB944HUr91NIZD76R2KO/WqB8
Rz+/s6muyA9dNB5y8wgUeXWj9FfhzlvjIqadsn0+jVBFFqTEg1sIFayNthUkarQ4lr6ODJ/LppPL
dJUCEhV19P4+/7o095ZJtcDcI8IjCkrrA5DI3M7kBAOT5p3WmCTV8P2XYlDvCwdIeGq0zbfIA6EL
dKMHneeyWD2W/ruA5atHRi0LwFg0XIuXjMnt/ssRNvwe1Xgf6RwbeEFPcQb+hEbjfGsCWmo9W9nu
GMhEU8BQJ1Bt8o/hVB2vsA1G8A8JZJAngPSPZkWqgkYahMIdvI/W6O/OnxcR78mlyWMlKrhjic8U
IjljLHWtiwPjweHYZ+H8hYKfsMNBZqlIfN4GStsrAJFPSk9FLlh4pvWY1NgyC8hm6JUe6OHkSP8v
CtN08rISiDwS7XJYZcMJ/Y/H1klQx3POfqYOHxUNIewSkH92tzG1jnGYIE/1DCrpxY4em/rO64Hr
145QJtiicBk/y1+A5JYv287DDDLKCgfEN3FQfrtNqlZtENYQ/OuW1DjX72NDWAq7bK+CokNygoMZ
1QdzmIPLQnBADIbMDdtiepsxNq6PrJtiKSZrGHU8IcNZ7F4sbhlZ9XSeidF7lKNtIGlPSuraPpiO
heujX2Tg64/RMlORt6KEsBZhO8MduKhIXWjBGT+At9v6RWzAuk3JDJLlKezSmoaKVBpHIyTs1r+C
PVgUrunQf7QTFL5Iypu4kNce6bgusctj8terUYofh4SoNAzKF4aJheszlq7u4sFq80lwSc96wi2o
jhSemByqZIHXnxYaIeT9PjnTnQ1RTInbka8W4FFC9oFzmLAua1ihr4m7+RTueLphqII15gNgZSB7
1fhz1DSRUVvakLkJBphLgLEez8nhhRSPOsC88bahYrSCL1yvDlII9ZrOb81BISFw+VD2+PDTkfu6
77E38yYe6OyPdU+bNpY/u7JoRMAxznxsxNkmVbbn+uQRwuKvN38E47yTil7OcF9IvqC8vtSwbbYq
2A8jcT8BkDqLrRu/SZLQH2jqKWMTU9iPwBuNQTJAyiU91xOZ+of+j5Lmdgea4LrMu6dHeA0zVJFC
f+Rm1CnCaZVPmcGjN/BYs+/NEzxh+znwSrpB9FtD68uHrPcf26arTMGNjL1Rd5XzotkM2UU1RALf
M9HuDQ95C6K43+BBM0VZhsYiRXrsm8j2l8qqgJ/x3KJJz7Thz2r6xmLm4fsfxOknRReUKYbfv6Y2
dOesWXVPd1tx8Q/fiEq3d6rRVwrkhPFJuJT0r5axNXvCi5H6Q+vRr9hlOQVBIyFRJu2rnmuAdDhw
uOk4dSW9L1x2E3Q4Gc3nQg8ZrkCp78VQzrA4Hb7xqVB7SpWQDtNLzC4N5k+cJVBdB6+gdUMeFnCs
ci0Eo45a+3HFeL9uZ27X+owH5+CAvsh/CRJdt2kVGeCU2FTf8NAJ/qiEHX39/pFOYtMTXLGI09Q/
B4sKeRU16Kp78H3LZlkCWRBu3ypXXBr7XJ/RdPPF0HdlDbZ8Iaxp4Ze18AyPcRSl59KGtbV0ZatO
VrlQD3aQVBKWq8shOWVVupzQ8z0dZI8QncDwtlXz0++PvxOTaj/w1w6cGl7K6uzWK7Dw4CFuTDWB
IGEybuJ8d7OqUPx5zJXW8AxuZMv5a5DStKaVZwK/JARvSwhViO2pdsK2LJAmbZzPxk5KD31djUDE
HCgebrvaf+sKt/iMwfYtwJCQT7MBwzvTo9FnNZHjB6jEzvN0tDbaBYm4lgIASqqJBWV1cFeZpx3R
zhjpbnWTvwZKZv82QVbAMBRGv8YXlnYPx7G/gu3THDU9zQmyFEIKWH/te2nz/wi9LbP7vosX/Wdw
8IgOA2f4/0JOj406sgj1f//qAoGkxT/mvjBMdAyR0UQsEbHSrYlo0bK5S18U3J+bunWmIyC+28h6
KhlK6uyZDY8hJIBNw2Wz+279nG9gIhnP+XapQ4mLXUvt3hSNXjb3SPAw+68qQFhzKftZuY4SrrEJ
c6Cad451MA6Yt63adixfDEZGW77ayUN9pSpBOqG6ufTPzhgQ5u0Rr5cxzA/jxabVOm2URslCpesf
l4To2pIUr8RQ0CdrQX/b/kt5K7rTP9mlL+MCsAEy/eama4IuAWxrykOLd0cns7CbhF7+cFMTUWVx
BW49xegA1W8PPc8QoTd3Ycg9g4lpzLTEZ6mVYA/XJCdFF6xdvLMR59XO9PnR9xpHHWJaf2vb/OlL
7Vf68gRvKaRz/1yuNcdbxC3Kc0bGA5WVYCIHg7PWSF8UrvnWIxlzm8JXxz84LUIOPiJ5bsgzMx1X
yojBAi/isqZnv95oyMB01fqWXiVwF3h12zs3wp4kkGSW+0s8mhTg4neMtGHEL1ayLakilocgQT0S
VDp092CKeacJlMDZOXnEy+vw669RPHwtkgeu33c+iq72qM3J8TzSzX0wixrX4XW40Jv2GgpKJqyD
NWez1XWG0PV+4dhMj4J3kJ0n3mnON2+vrWzfMIywHRLC8HylR2tSnzXOqtLixi3Zo5xS6KKK1hms
uT4bq42Z1mt/FiTxkXedcPfB/xfboORzX4O7eRPGohYwDJJuVfwpRnjxuWUA64SXX16S2YYsxFW7
iPEVFtNiMgO54EpGXAF5ZMMoKxeaed9qCTgoj2Mks5S1jOWSH+SkOwHgloNg++rbZjKNxi/BUZDk
E4tuCv2k3X6EWfYtpqZL48CpN+4MLGCZOxZ6RxGuxYjXvh7hENBSYytgoJgxqbSCF/nDIECc++7i
vpt7A27St4+K0D6xWhYWVsjBwNPyl9ENFpUe/HxtsgQCT65FC4x/F9KzXpG7JYiwjaedr1BI68HM
xygfH01MjlmnTR/v2oG/Fafg9XHGSzPO1ejPZSmy64Thbd+m+K5v0JfuruWmTxWN0p5hCFOEv5PX
bsvIUJjrNrFhGU5UQxUbVW+wb0vnO2Cea1K9TeZiAQgyFgzVbCR+U/cqYhTCQxxfrQZliR6lOTao
B2HEcdd2um131T6jxHNkk6P1or+l5wANtsnRE2VM5tMZP2ZyHZ9ga0Z6XuuCWxnIQ/P+PrglNofu
YayVTpUnjz3TvaC1ryiquGOrx2OuwlYRm/n/my8N+bxawgQzm/bYYoa8wmZPL1dt66hq6o1WpG9d
2zTIs926IM6V8T3D904omAlv0d0PKL8b2mxfGdRUen3rXqStYoyxfd2MLU2yp3PsQ+U/JanpghJW
8NGiJEqlm0yVmjmIL94v7NBr3nHmv4pfvMFAo3hVEfw/3AbbmzxF7va+KqV17qt4jfEyJ+OzoSDq
MsUEEGbDRo9VqUCSibl32ZLBbp/L5hwcxEWtMGAjHnGZYXII3xngk+0kuszadI9MdIMy7iNVSejT
nOtAlqbTXHm/bHoHN78msBCgHb5/PaC2HT8VtGREDNsX7YQ0raY86NBU3ynO5k3mQa+3pCQbRZJA
37IuOu6z/qZlaAjJj3eMpGFjtfcbnqwX0EMO+r5vp8l62d9ZyBFWuS0vUaaFwDjKmmj195bYBq6R
5vKVDknDgzkEWPzusT1IRQHG9fopYkfEkMF1UfwWMTU5m+NEXsLssXtb0ndca+kCty/9d9lYpnkm
a2B5vLCXAylH3PLvDSzLRON2vBA8qvFs59e/jvXpN5V4PnTbR9jsRPGmHtepL91OILAbsbpTotnZ
d3w2uQDK3l/G+gILQyucw6sVnv5Fl/SaAbEu4qrE2OWLzL7MEzwGriXruvYiU6NIFgN37N6slnYa
bwFCIDmIYKJ1rbY5EkF43FqIyHoSP3cf4+vHbQZXJxqCu/C2Gf855+jR3MYWq6j97w+CjfIrakKT
uhZXXARcQARrgGUUus7RJdpGCLUzAWDzum9QMy/3OmO/gL/77uR1cyL3Cnq4pUNl/I0KBZaEBkqn
8HE8LksTmigGI23JBDODGnaAQcWNJha8t8Gps8crfiRyISqzK3fwGwwrOmKM/2aYPOm2EUxavFOJ
sIVxJCx/gzqz3HirVkk2kxbVJS3GN7CSZG0uKDPOeBgUucv3YfFijMcNuMtp/oIBlIncqTRTkgnl
vub1f69fI3yaMsgDfVRSvK6Mt/j8X0uCyIHvix82TIgkGwjAc/zCY9N57SF7cZCJ1S/vw5UCvbol
iIKVgs6/X4olTSZZJse2gTfPQAtu7RMV4O+PVlJLMNR5FnmfC728GgeRQo+m8qVg87s+Jvp74J/x
RHLDXE0vTCAv/RoiNzhFaXElm0ANopTzhpVCxZgyx2qPwTluUnUtetmmCAKphgdETDUKi2C5235h
MZ59w+wvmbGoZKh7xhjMWfl+eCCeu4g/0CCdLpenmDIxDuFi6yqOXWt8LaQ+vzae/q+NzJ5CoDFG
m6oo8nLPeIirpIzmTUowEeSv8pFjgLxq84JJ17cKqhZAHRkZ3+GyOZn4LBwTam5y2mCiq/G+qUw0
mIB/0A5tCpkMCO9gl/nrE2zjnNEHV/eKLg+k3huhyn5o15R6S4Mc5VMtQGUXPMNIYFhTX8kVCV12
BY2W8/JAOnTcxPtxWBhdKicf80hIJhuZfrSEwY8KcshBm0WKQVN3Bap1HTfoGA4w2HdK5ytDLkpP
qSHxEZv/eeQcFir1r3Yj+0nOyUCpG0fJi+hEpUfpcOAiBmC+v6B9ceala9ZoYecuclfupU8pUJJW
LmQjgbUWTiKVO8BMnqaf2/9rkDqLItvEyDCQjKiMCUMpg2xtQfw/QxWWxjbl9aDLdMUvg8seop9U
/zZSOFJzTEI5U004RjpzRzKjZtuIpqxQQ7yKVYD0M8i9Rx0Hp+ukanXHslJ2TwzTD2OTZiVL9PN/
LsE6iFu0CCkXT5rO/Smm+c50KIkVeEnibrTvrsNEMunligK+C1BRJ2k1ZhxKDp/VrXI+rer10/ym
3lhwAVcdbaqIoXSAzcp4ne8bJA46KakmJmzOPtRoiih3vEmlILdtjDQWcPc8LSh7XbDsn4pxcSmC
D1YVcxPxtUDqa+cdeOV89BwYNdj1h4hcaLCnirSpOfGb1vhAKjijcXnpTOjgGucKe1jbTJHk5zIU
kSO2UpS2yYXT6PhXx1MYf2/iOnSnNfGiiS3qw3OFlzzTWR51jInnkM86TwgSTu1/kZV1cBPDbdBK
OZ7SZg6pUvT++39zsvdwMsBYpgkJXe+fNtWvjk3falVpsETV3gxq6+9M4KGp/+Ue0FSY7EG8nymX
b/Q7/I8vTVF5CmS0k7kGjs/TUsVIW/YLXg8Ylb3UKr/6s/FImFy4E/zPiErX5p3aJAc/vTYtAQP5
3OdfikSQDsHZ4TxBAmhoadOZ8vP2KiFNYZCn5Z34G3ysqNyWbSrun8vaySYW2M90Emstc4rRYIFE
YqjIAwu8nOZbsRO64NlBvwHtgOScByDkUX/RsZL/BJiWjYpf2hH3XGV1/U8+WBfYbfPGzxB5g1Gu
Of1kX2xzrDNAKh6CvQKTJxVjsm4sKNerzXKtPw3NIZKN009vlentdmHiW05RQ58ad9ByeT9suyTY
LY9MEeYdmeWRI+xnUgr5EAkMIL9BtqV3kTnAqElYGLMTd7tzo1uy+yNCnma+htaeYWZfTd3JJ5oS
QyCx92W0ShgmyxyT7FlghPcwurt8LD6yaN2ayQeRbDK/SRu3I6G4Lke9xHJuhLZx0/iZ49TVsWPg
CSrT3MIloJmC/41HxEJCNGahy8KLtMZAXZpm4rtAO8MmDuwX5PV0xv6Vd5zebnueRrz2hySjbCx/
BT7FBY5cLRVnFWz5vFWs2aWeKl44VZaIGUg0OQfX4mnPBMpOsh72XXq93Y8aENQsjgiEp7kf4lXq
ZWP/ZcXHHIvFknee8qQndVJ3qkn1OqTXjgCLvMKfva6mBTB543bT0IbCITS/xNpkjgN+etsDpeP4
Du8KyZk2LUdt/LfGx1B1ry2TXaN/ZgbON93GhWw5CYErPbrZenimYtpAiROQssj1pR6RiHmmWScS
1EaDPeVye+aMQDzE7uBLJIi1ohGPIbr+rQkBLQMLAQhJmvleltJbD54tYOSc4R3ih3FrMIJAJzKF
HnC7IsOpACrYdfjzWYHIKN/EMGFiPIiZiWTdEU9cxqTZYM6+KPcR3IbZDCkjAIxRkrhJ8FoErW0Y
7YD/ZwGl9hpqpCoetYLM2xIndFPeSwQiTJL2wwIE32hlpX2ySTfjLYR6wM/KK67loWu4zGm+1zMl
bsTP7MWRA+H4Q47au0j+1lVggLJSaV/CsmW9luTMVq5r1n+pdc7GLdzEW6q6pxGusI9Diy9aCYl/
gwQINHAK4ScXbP1DW9VdEDSBLI21litbW3oprca+zOCI1PBbqcrt0218aZXN1VMdvgWmYVpNjKwl
itvvBkgbrcjri49RjJn/yMgU9jOTXW3QDcWwgBH2FFk0sW/zkFpi6hXq+VLqnAXDUcbV4HDGQRZa
braK+PyKNbdUAHv8DC8TxELzko2QDTsWNMqeSxaw8zCbV4/mIPHecWayvMhguV8XaYehG5zvDdNx
a9KKJIRqk1pQgBhpQwmiDLaceBuySIeMTKzDsBilKV9ZmeWDgYPB7mL6mnY9Nb+lJB41AqxQy2iT
eghIgUwCBk8EXhvfu8m0xXl0dMeizc8AvLS4apG3vSMKeF8AQ157U3y4Y1XYsHNUmZ/nfQ3Z6GL6
Da+bv8Zu1Zzyy2ucBYgkWHtZFUpEtdROa7xS4PUpbDW2ZSop5N4526idW1Uu5uHtFX4345Cwt/DH
002VoTn6vqMAwml1f/JYkmiqq2nWmrOd02KB0vaevU7o6dCcnyMqUQgJYcUpmoYjD5KMFX/nw3Qq
Cna870y4nrzNUa4MBDcxqrA75zddDdsBuKcvbM7aLIxlxX/ALonAOVE2/951aOIZHBg4pBJCILYF
QfA6pezswBCQb6RYqoMsmd8ry/LWsiccWfzG1jspE1ao4qA9yniSL7yX99auJDzqBWXilN5byuM1
1tbhlMeHopqWis1oi9Ykh59OlgjafJGo7t7EsL3IuX4vbTV1E1P7G219OfcZnUZtqDWDLjFPcXbB
B/onlcCyat/EGVL6tPY8robMUA5+XVKf+oG34aK0RH5qDy7291vCkCLhhMOeHW1YCn9HFbf6w3dB
sZse/o/aOHbRFwf1w2VYcVBMch3iBLLcSSJUndqQ9oqWqtptxBIMgy/Gi1WjHMfXTSrN3fhahTyh
TrJ5s3uIlbLlhiRjNyuADTdSO9B9QVszLW+i955kWtag1yJJLf5lItEQyucfYqt8s5Sa/PNw6Qfv
wsURviDq7s24PGv1a0kK06PmEpkL9upVjSfEqQZ2Fnr3zmkmwCvfZUPF1wCdtmesRwsQFOWqHJzd
Sec03YSvju0Lpc6dSKQ/7N8g9MVkgReccpQ1qG1/FJakrRucfcswlZu2WFkAyq5kVFn5SJ2Hu7KF
zYzFMHQ3qJSge7Xn+RMoSduvTuVp2e2663Q41ic4Fyz9lZ8Hd97eK7IgDuU2IQKv1gV0ch8cxDVb
VQoHQcTkyKsDIsShCWK+z46mpKWJ4RcRfZTqLxoXi0bP0rGYk9m8F3AwdktT4675HenQI+yqCNlP
lWk8fbZyF7POg+xhedcFfg2K8OcRTkLGspKjkUUqGfV0qHewO0lREeJf2sx71J3G1J8P+tyPzilx
QF8H6P1BDBc3rV3dWMyF5l0sg499XZw0Bq6/KgaXUqVyVuGpSdTCK6rVA6RdCc25K2Uj01u7w37v
w3wbI0aO5qzGVBH9iOUom+ZNaIhcY+tlA3vHqV4TI2PlgPiDI+IbPT4zvPYmEyaWBPYhX0u8stog
KW5iX3MsKnSG2/V540c1fWzObX9HTE9aZqzk24qBcBPTXSZTLIakVKMVXvxgeQPOHgktUQDaEd1m
QzD6NaYgPT25xi2arj/ZIePx36KloTpn5YOor1Mw96P8BX+9ftlJW7+K3777fsdTLVhdXWLQiRog
bPyjTUnb2iF7ADopIRSJ3xELwwxm2V1x1MgnzhU3wozhHimMHqlMolPPYXwWCFGmSTitkMct6l5T
WHuy4/6tn6YuprcfM3DImTz4Pke1pY891ezQChQP70rYqU6A7ZbVGx5wNJHg+7K4Lxe0Xy5Dtzig
B0ATTHwEWtphL2kdv4vJ2fwMeA9nedEhfaQWTmWYHiOcqUvmeKslpT7edffI4PhgtWYXq6dqOgsM
6PlfGeOndgjBovknQdiQQG/ten9uBCjacrAo6KmGNVx6A41w/I5atCqBY5b3Zx2UxaIWhq431XST
Es46m3DSNnbcEfL5ncRsCfG0l6men1R26kpNp8vQCiJu2P2WrvjonazOY+CjYl4qhYymqV22fzI8
7DwWldTyzZ/GuRpR1wJcQ41zoxFowQ86XPGEXqkM26+P5wENgiqQvcDyhFV5aWmDmtWch6ecqf7J
49SjbWH141eUZPXdZ57rjzXjpWh6NsFdJbAIX2F1l0hCYVT4+ftJzradNiZzGX08i72x8unxRPVE
gYHodqze/MnV4zksOYRG9vRp3W99ZmIY5FCzhBp0wJZCucFxpF3MDd0VUegyr5wo0ZhHAeeO0HlO
DcWoDZWFRfYUUOJeMr4uaTdks8GfhNpLUVC7irGgWnV6G5I46aMx/tyj/AeaihPtfVaSyZRiH+uN
YuWto6d+IhV3PLmGNwa7av4RsPzfIIL9f7gvAe3V5fBWzkXR+38jpbOgYxQISuimbF4/RpA9EO/N
pMJM8u8ao9oGSZH1+n/yD6u6j0dQ2SymLNG3XhqTHREN+XJ6R2bQQPD5cGicO9jugelLD793SqH/
brUtnWT0QgvUJtMyyCPw5ksy/bD3VLf7QsoJiplLF67X/a+N4I/JvmUz4qIc73AiXK7UEfY6Afa4
otqw/0RjvKlaiquzvfoCiWNafVkeSZXHjOrLaFldkKTqeefDy6CBc8tueMIXG/LzMCdylU3NabYE
7B0pO1Gxwuf14M9ZM5csLOsafVSojGE1lEY8e4qJIIWft/qmvRSsQPHNAC6rMP4zVh+rltMKYbHM
/5emPMqKH0tnMoo6t3P67NwxLlwrQz6/4WI0nhaNl+5xngantWnQcfXoAKWLR8mz6OAu0+n5tlLZ
405EPoakWovDk3rsl2NMSs5vfxnm3VfSSLUF+bIRMug4iYI2WKuuH/o/ZnEzNBgDUqWdMPlKseyj
Lx/TtjYS8P5Bcxc2817tePStGXqDbUrf8bn2XmiBUoPM9xNfADYqPlPBFMU19mByRzssSoEvkXli
6DQiNTCGicrjHGjEAGGeQvbUIRQjUBcqP78HJUKgDaRWH+JXPN6qT+5XuDcLxZiIwZOfiAUhIubu
afdYm68I/g7mEO7059U44fKSFBb8bXGKu55EEiFuDURzva1Fdk8aKcYh8plOaJ/nyEiuBQyE5222
W72JqUVrN8HXyfzTpWhMAGGWZKofcm/o1yYiVC4J0M3yVOKGvzr4CjdFLiHLCoCZxYt9qFY88AIu
RtdUjiNZrx8u1Vs6yFBqtD+j8r3VDTtQiHd/D0rLNi9b8WaQQLSI4QiC+iHkZsZiscKyqDgbLGXt
MJv3+vQfmWpuKTggG4PJaXlOSnI432YHogLzJ3/0aYvhu88+ZwqEUbPwQYWkMBRCdbXvtUhvyU7l
CmNjfAwrVNkfr6At856UHsLuOPQcV2C+jxuowVurnntIEbFfJAGNGqGzV2N7ViDkDl0IvlnT8Xev
F/Fb+IXr47SlOQM75SQsXgJ/pQYCUfDFLEh6hrk1UqoklHtqm7uIITUL1tS9ydxZmYFlq5qDu2W2
W5goFtQuZlykqSWGx/yL+HZMZpUea/J0nooaGYPKzdgRSFhn/RMDUszV/Kc6ifPNKWkJKeHDpSWv
orZeLUHDcjR5jQRXMwA4P/q+nsvnNFNj/E/GKEluPJPAuM+MPAhysTYcPPq99YMrr64bP74+/lQa
HNYOcOhFa6kXMldJ0x/2GXtrbTzhVS6LMbGY8OJihJJTLXzozKgIDFgxTrTuyxc1dT6U3ONmRzcC
uk4IZtl+SqtlXjAJ3B73o6dXjL8sP7ZdhG0wYWElm7BisSAxpEF57bUhXSDNGaFic+EzqXoS9uwt
hbmH+e083gsxtrjk7hCHHSiZ2bAZ4lggoqr7U/NKjgT+vs9x1zSyfQuxfdTcytWKHt21IjdWCF64
nvJnPEXZ5wX59ChGJimXM5oGvYYLHsnOhDNQfoFb7x07NyDvQNgj14C77UuvsN6B4y0EUNMigQrM
2iiIjyVd0KfIEPBVqMq1wbOYAZ7FRmF6tbIGjbvUccScMImLlyy+RjQavtesYElWuj+/PhtbwcdX
YEPMvonWsBA+c6BFLYgeihpuK2I0sVfMuFNbU/r0s65CCtanyT1bOyWQnDaEIld10UwzNovkAkxL
8JYR6nE0rIGiw5iY4tKFLS40t83giBlg6cF504FUiA3eyjb0EK00eT4LFOt1/ydDzS1QQmVFjclo
k5RL5xlykx1s29tuixF3iuQgvKsUM+ZDMEqasxg7Op9yrq7PxLBl9+cB9maBklp3jzKS0cAmznd4
ABKYs2P5/K+inNwoS7ANK00LrTpVuiqIipE+9WpM2qh1UZzobHQ6F7+Ncv7+jV6ZbGuUiRMF4EV0
cs1Pdp9SO6ctL7TG7Y38A6aGNMHtvaPvMfJomoRHGEZAFE2YbST+RB4Kr+rnv90zwwzDFpa6Hqkm
C6fPVPRQvrJUqMmCmUO7CMT0oXhfb6sl+NmWBsAvOZnlcxgsZN/Fkh9R9Q8Do5l5/PDgVzW+Ksbs
gjZxoTSQPNiqKBSa0ec1URRoB6+USAMKO7vMeFwAlhenw2mb7XYLuo4C1p77N4h220Iy0ieE76zU
B6N2kriv9x1W4N3EaEoUj4/78C7lVOs6bB13EGjiLZ25d6k3jCFMuda6wo3Re4hjxYLGYOn1Jq6b
C6LVeWJKSb06ALCuaREbDPLQ+VF+lxTTaZGJkcRZ5ctfO+48i/VwWVmbn/YoTCQesoWrugrmACgw
VSLIs2g+c3gmMJjT3LzJPiMnrPN15p4r3M4P3SOcYpAmsU4izbGpAv+MFAm/Ks1TjDr1vx/RV71E
8eXRNyXqvs6MAZ7W3r1rFPIODdJ7LtTBRMk0U/67ZcxXpFdIxzsQEm1k/9haGv1QQIPK8zJO4lEq
7vFB95MoQ4YfywGGWUooCw1TyDjSZ/EJBY8A35dL+zELdcgT+uTyQ1IwhHV3lmH/nVVLFJ+NeGtK
uRR1R1rSdO7dmprmBTwlfX+LJp7T4PTXVw0uc9Tldg/MjR/zAyJfQSdlWLMBOuGvd3UeJu6p/aJS
wwhJlyj3Vxad8LBMUFr8IqcNOT9Q1lh56uNzc59juj6s3hKrKtzMenZlmNnZhaXlTXTcynTqqYA6
7J6tSzZBneOdNvUOX+1XiaWaE31GdSuukKqH8NjAnyafHsNMHq7mrpvTvAdqSRzqNftD7QYuk/BG
B8nwv42ekxyJFpMUe6jKZSmiIvrYsSVua5Bli2vYfEwO+kL3QU++mYSL6WiFhy5cTZEXZg76W9Ut
cH/nR33vyqbqAjk4PYUAHQSckH04t5KbvSJXd4b1boodaJSrex529+D3oaB8NwAIvKwRO4tUWxoH
kCbgECcUNRE1pNXBwEUcXDYvaKap3MtRTSXSi/0kQE/HRQ0I0Sr4dgtMe51C65p39ADObiJADztT
liIDAI9mEP3TIQVigmIPw1o606FYBgTwqHvlNznfHqTPhp81ZXqyGP9zx9ki4DV76HQkEJsNGS8m
IMvyPSpG9d+8R/0FxmPM83rz7Et8BOBILFStZfiSO/NOXqsoL98htSUrioskZEp2eLY22m4z3tq0
IUzHPDvsSobeXkKbu7nU/ta8Y9QBFUV21FDTsDFNaI/54ot5HgEuK+UOGTwLNEyMeMqncMesVBWV
8vZU1Elc7+8NciA50ubVOck5oy1hdNZfV7nv8snWJbH/9rZhoKM1oPheMctbM2gYE+DKXMRVLkVj
Yoz1C+l4D0dA7bK52JXs+hDrxJ3Obfa4FKC17Levy/jPAQLDGUF7QjwlJQ6YdguVvLrRv93AFPKR
am8quqJj5LRnw7PauVjAnbbaVHS40I8/EBHhLc/3+6zJYpBa78nVO9fMgiccbwSsxP02P5QSg/Wq
jRW+vdU8gt19Zlicdcwd9QHefvW3b0zex/5Ku+qL9m5VcMPEd521MK8rrAApaw4v74ancfmLzLYw
RA+JtIlzEaUP86U9l0tJzkJ0IbHZv0MM09q42Sa/YyKjYGvGjV/gFRhEkzFn5oQqQygPMZJc5hpY
iAAQc4+9gmR78Fty6PAUsZOOl0c8/1F2lgtMIdXeTyR9diKG2AShkP4usZ8/4gB3C/xxoEVKHUQV
x5IwkePiQSmgmBVNuCKeLPOAB+u93uSzhx+UHX31rcW+oR41o6GAb+g9jnIlaACTmQE9MJjSs3Kt
LM0JpuIZ0ULAILmXubTf0HEUCfWspjCuwEL5eYmsyhBpPzC9a82NTbDkAWqxjuzGvEiUmyPgr/2z
/rrIlBCv1YUJuEW60MhakgPMxKpa0KxV1Ii7EVT04WCrwmEurfba1fSwmVOihLjgR2ymwv3nALcw
+PNwdOM6pPKU7pjx96BrKBA3djT68cOtUXjJPKnvMC2OmkblZKHwCwuI6zrrBHqYxIM0DgKx/Zhi
wMH7mKRNxT5P330Ls3V+WVxJMxeIiKf9xe4p7vpNd7n2ZSG/RGkn6lyOXidPVhTbcwIkjmsa3FC3
iFwilXc3L3DJa8uTXxOeMTnZ6XVgO8o1/WN7Q/aHhXWUXjDkIwJ67ckWKTiRMv/CS4Y4JdbKo9h/
wDvpQV/ecsUzrNY1wxFtnrYVdLZw7c6ENxrVw/cbw+Xfcb7OYRTJ4LHWru9j441X1b2z1mBkPFff
vYjmPUJHVBU6oL86JtlTNCdspbv/XMB1QlloqYo7V3IPNrqoVub62Gc2GuHPZIUYWuM3Sp1+CK4v
Gepl9JmaTK3BqimXjkch0UyCjZqOQYd4w0q4RUr2iXlem4PAlHylbzoTIi8TmkP9IDsW+k6B2knq
brrbMkAuoMtoUeiqG1i1DhOQ1bpCwSjO1JSXIbQAtWtgI9CbbGGczvhDpcU3PIXNqKWxbuAuSOQP
2FZVg1n3C6bcr+cYYR5NBPqUZJDYK3gF1emt8acVcI5JBVaE8ttHM8PVEAmvV55FFya3dVApIbGA
qCJZecv7HKY5n//Zd0/YCCT+WGSVOUzt1wMJtbX31dxcWK0+DLuBF0/V7cJyYkkMaWcNa14ZHiQZ
xuzUp1wYwbUZohvsjIt8zdKHeomjRVi5USmzKcF/v7kPRp558Kpc9buHr2vut4Qw4HylqltbSKwY
DMrF6+yq/LwWalI1pfaJJ9uppZq906kULhJSm5dyCcgJ6arFoXGdG9/t4+S4XUbF2ecIxVVnHdC5
IVTVZRbhSAcbgOeqIozkP5SnzDlyx5o49eceQnMjJUK7uCn8HFRH5oxiAbAWcO4VkLgKz2E0wR/z
F/3WZGCRJjdU77Sll+tElG1fxYv3kh02SZR7QNJUwMF9YmXCfCAeduwnfpCqvl6n/lRw2AXgx2Vj
ATfRffnS1V4/t6DZWP62krDGhRcgBbyk/ONx63xK5LKI351A7ydijxlHYV+waYQ7RLUXAsHtzeKR
mdH6hEc+HDnXKWZQArazwCpfFC08li9FCpzaOVvdV6PTXBV6rlH4IWPPJq4o9SiKExDzkasGfHwC
rHOOsRCpTJ9YnVYkJwW8D7Wf0AofqzSHS6QDMnKCAtRUdMFWwflnIXzsbxXfnHWoBE8qS3mK05KA
DofeyGZoRu/wI/rbC5rDf3kP+3jbafOrHoWqMJRNUuvCgZ3Fzlwwyrc5sX2rHHdK4flxDFyIrXjH
xysXt1DKb5dncTOl1i8dlB3irN+JeUu43kZAuVmDgfSEnWQQUpRgbhzA2MAIVYsgVGraslhSjtiH
RwHwCyCi7HTi535CeKjaGq6iTgTxpniy9M+HCtk+rBrJ7BgHyar0FR+2GB5kHX+1T32Fs5KNlvTs
eEUfZfpUcoOtEgyDP+sfLYFuTrgbjZRAGKOLNxYNDiTcqEr6M/lX3mwbfwEcz1A+LjIpfepzcVii
nyQC7qIzEmOsJq3hGtn/qAPf2XDLj93t0Q/hp1Ui67an1+4zSOxmVJdZ+WmJF+9BvZ176bBJisdc
ORVYONqmruTVcr4aStF2tvMNdMf8xDaOivrg30UvA5Ck6zdMlkBEKnX8eQY47sF5qIFbVGT0ZFUF
iD5qnQPH94WEA1G5IcuoqIdSkOeRmRIxCXoEdXcxfgcYGMomFKYHKc9Jj73ewQ5QrNcI/pzYkN14
VX27zP5pCOskb3gMZl36W1x3mK+jXuMNNZc512HzDFAUHHUs3J3PzK6Rv2yD8LY06aIyb5ZhYXDM
pYZP+me+TLLXyZOEJ3I+gBTuMtSgMThE9vADBzyvmoEhzvCq0SGk31BP9aUMLzmV9pexnURjj/hD
flKOABpAb2QAA16kQY6BLnh13rIrnYcN1nBy/sdHZRqaultnGelevzrx2LvpgdT03QQblDhRv0Yu
Mq4ERGb7WXuDHxkC8vdnDH5n20SkpMhMpeHx1DF7f9c4NIvgDgqOGzKUOQ/UEc0eIoE5C+6ZSisy
u3tfJhBqq/I7f/y4qJ15dFZ4crZD6KtOVkgeSbJZdEGZG3QT+KTdIpHEjd/zTmzOkWRzbFT+HEoV
KCNP3azOcZbhMLL89hbYMOz0fVJ3B7tiWZCZBE/i8hLOOawmNNcWhCkXvflmWdFu4AYuB6vgzdzT
8kzMAMfmtwdsU9V7HJEAlGp/5QXMiD8XtTmrqmPZl0RNEa7R8JnAIeoYbRnZuFnSh9s9Ha4UVTJd
AdLaTiQt8BIFKsIt5fa5cd2m4E79aRVYlX6CRjYglfo4hRas8fLgIuKTqMjiL++v/o9akyI/32OQ
j4nZmFQq/h/SO/0gL1e3LPNYK/XB7hFI3QoGgBlK/xbmcEH8BvJ5UqyaskJjo+I3t0Yz1isj6+4/
iaPuvs0CaLdeMH4UCf8FwKgXjnZ1lWTK1svheIOE/eUujg+wjvkdk41PTL18pLvI2E65NR7jFDcT
KEthG/NdSkJmKEqk7grVKAKMC4OcsLdhxgilMYuY68528McP3pIxIU7bhMDiHQItzGGMr+vA9omC
P1rPMWMFcl+jSP6R251pruJUZEqYbgYTXSdzukaVjv9o3nzqq7SZYd4c+2D5OnGywB8+H+h4uJ/g
oTLk+PsJmAtbkhrrY10ncvahg0IJSD4pkOSx0F1Fkw0cB2IxIfmO1RX39defmEvPpkxlOpgQxr/Z
RKhpUMAh+yRMQ5027qz/4jT9542OFpUCRzkjMZemq1sXG8gjGOvK7HasrTy5kOLws5t/Vs69l1pv
0zOTQE7iiey0J3mumnjwXSWrdHwoU9mgeckn+6hrpxXm6taJzcYf2Q5mr2pzv1jg47mVPO+F/zbf
NeXLFijxrv3ER6L/rFyoFbk5WCPdiVy7C7a8spNwGVJFVQHYPX4b7NmXsrxKELBCvXw2yRXgktId
qVSPqz9MscoGogLTxKa0eQb8/gK/ITfJklY6OBUBeHvV10iIsOV/hiEx+2WIJA96kC8zSUHV59TP
QDpVVNwYqDySZ9Njif76gwY1LrB0Wpq0X+2CpmZyoBgXDxGiNxT5vl24MuFgZ/CjGJeVkEJ3N/tR
jLZoaKhjYQ1sT4Le9FTjiTmGbs+me8qlkoacTPOf8areuxzg8Z+RHEAC4pwGlqWWFMZT/dL7shU7
cuuid0V3HgtVZ6HDQWx2FAcZWNNSzwLqkf5Pm/QTqXElC6eYgxkrFd97H6YwihQqMnKV9r27GuY9
sYpOT051tTX7LsciaTYetoERpupbp6HNpe2sbImQmbGyTRO/xriZu7th9L1rwtF07dUqKwg/YHVs
7lWvTwMhtHZeD0mRsdoaBJV0ngbtod+1NN4pW5nxstudvk7rOLISLBrNxPwjQZYRFISK48S7DAuN
nMsgp34VEWKG7MTUVUfLBswg8ywcKnLU3P3Kv19nGiVlDN3v/ppuGSITDHUfX90xryHg19VfUks+
3/drypVk8kDp7QdQav1kUctOmfh0mIkrkj+EswJHnIcDGJ1TNcoNL5onz8UD8NZSQI5WbcbMXFbH
5rdMmZEJX5FbLAOPWcgvZ5dCbFs1XD8ikWe4K2ivvIdBJmCDkRle7JN9YS7XeEapZdgQJZa0/2Wu
/kPXmbKiuI8Vpn+yOws3DBRZMUBVAxMPkoDFR3bWHl9gvRkE6iFZcXyL6TKVNXZLQjbURRc7yN+w
YETUhVZ8+Allmo70IRtNW7beItzJbRq8LgP8o4dr7B+W8konp6UIBNKe01KUOr1xQjwXvcQW2H9c
J613iwvB/8sjI1sOn0ajbHnC8dvBudfl7JGa3eCgatT1eOt8WobArardIwAN/YpwYOVBBhTmBEqX
+5jX/obYtk5Cu0WaRfFnkclYnqusdNcuxCQbs955uo0m4yBnDJtN7MurzFEnASytav0r+GZ2iqsS
A8GsZa13u17+IByXhKgUejbNN2o0PeFh7NSS0BUnM7UozoPNxTCBZ6LilRYuL55egjLs2WMNeFm9
4LRHVQHmBV3KEG1yGLP1nkhy4APyBpTpalLjAZiCkMrk0wZupbL8WTINoOS00bfZKCb7mDM6CWYM
HyVlOfCmnWuaNpAWfoEt7D3HT+aN6uMlKkYwbR2MTrUSRt1QSlxNY673x6cG6YSKlojpn9D5rtl9
nLmupS8lcJUIvhPpNDaRF2Tcv0GvENky5xx/Oij/+pB0Oy5YqwI/E7uga2GFpuYHbZEC8jqpCgGX
aFtc8bmG+1kk+ti7kKQg3oYs30+jofxg3QkqVJVS0TZgWrHD4jnOCqYs97EhP4E5wv8XFzC+ASNd
LIkPxQEeKAve0yf7Erj+AKF2XBxXDfCRFd3IpjHu21cdYRcHeRkeqqtuzCjKaF2sIWpPCNvN5RYB
ssKSiHJq0OApTRklr3wc/uKixAqwtZ2S0vEtwh7CMrCiOsdgq0Vi4jBEgkAI7ZlYK/acM7dMgWDR
V2GuqEEPVB7ahCansCOzdOSoAMJ/a2P2jz0Pz9QNLoYQZx6ioDiHoYQs7FEBseJVR6ymatXSdnDx
rUD2krxPNEiRU9UweyQp/xf8iCCcz3eUIv3o6sVqbvte/kl5r7lob5fCs9ipjJYpxH2vVzKb7CLx
DJetqAmkMXrB9S48JmbWCDWdM9hpmQJDBvCwLc4z6o4p/eDIAoOobSWc29SuLk/FzIftDo7eT0S2
XwO+j1/w9CTm1nURFhm9OFBL9PzpVJcY9avgYPPoSlDfABhldFmCTJ1gFGtiLsO28Y+uePgP7JJw
gxdN3ndvIXDpYqtUTxtDSQZuvqKZJqR0X+lQmsDMQzD/xCTsUViGMt56HSRu7jRDHLh5nmBVnGYm
Ncs89sv1CkXFKpPsP8f04XJKLmYZm8ho9fb66934MQ3gK8rjWF1PpzZub/X4SpK8o5gxckDP0gwI
zuO2iE3pG/Rq0UJbvqQlpGEtPREK2Mr6Oib7Nzc+ToFQfOmVuQc+6n12oNhue1fideUkn8sABn46
V8WMqm7kjty4TXwmwmWyg0+ytcKvwN4qRtAXGpkJyYZe51SXQJ5duiggUYo8yv1Q7/jZFscNPoi0
xpX0XLXXYLfY7l6wRn6xkoSfqqwYOSAjg3xCHYBPU8oSH1Fwvu8TWiNrNYEycDB77cWQYrR79BLw
po6Xe7fEjFMmnlfZe9vYG7z8TAy1rgMCqXyL5EyKVOM6tnKVwvaIkgCf/SvloHcOqa7vFlXwTm1q
7PtndYg6U4poTKfFOFPpVSQUuY5FsqLS173M4cdLqZWhuiqN32pwHRSuNWlDSSSo4vtyixlK7nxG
ie6U61trhp+yYZbnavZzr46t60gDgYELQHKciygJHX+oUPivfHFwgVhF0dNRF2KKY8+nCa1mftsk
61PLToKjXO0BbdwLgVfxv8bT7KO4loLr43WQCFox7O87T1UbT+DCA1NC3NtsX/qXbFXoFj2ZBMa4
m1EfdH0+hvGHqsd4LPdX2Dkx+ATpOVNhncomZipGs4i36jVAbxVXu3By4H87qHeh8WTQ/cZfM/Cl
3Hbkvw4N+W8prh9dVveidE3eisjs2JT6OPDzdVr5Yay9rKlQEYCRCuc20kizUmz/fBxGQjB4828q
R4UrdtrS2i8TBfqDVcrGil+EVGO6xHBa1TRCWIKPY8335SuTkjItGua66y90y3YcMsXGPx7HsevH
YiKRZkPWX4wCaQ5Ka5Ax1+ZdBMMUDdpFqJLj75ihRvnlp4Rhro/dAVhmc0bpTP4Z7oRSS2qowvEG
SfidZVYYcJXpOKfW3Z1BlndncNhChimPdJs47U0sUCbg+B9HoE3ZlgYULdZtqEHdjOMSPpRXoLN2
eOJp/q29eA5EIyo4lYRjR3QHlZe1Ade/BqVij0jBl0UukZX7MN4pvUK12bfN87rVGRxBN2SENglH
e1BAVGAnFHP5YS4qhAOn5RebpCii0gZ3sNOWS0f/+drq+HJdU2PCBn2OjqqSJGO2VG8QclSOCIEH
DRNG6y6pmHkXAfuhGovTQMK//MGBuqFJLZdaAR88qRmEenJt5g6wgV92k/pQOEkPKseRX7H9sjGW
rfvWPJy52YDiBfuJtLacFi7lirvoFS2CFN4bCMyvhtYMKn8ezYE4wDeh5acf5Z1ELJNV5Pi7c61m
qrSrx+/rV7chc2ByiPKpDZmjONaU7+MmffbvfDoRbZMfM1aCls4NboAWSOxWWSYQppiBIqrM6tgl
VzZxL4zWrd1p+rAfo7cOA9L5EdP1h1Nzq0tzX3VSekw4UCmn+T0+wpuRbPktD/pbjxE69y2MxE19
2XJlnu7Lk9ZGY87xJEdGUrifNS+/9zgC2uW9vUOk7R3zziiXzCwpMWNpaVubpl2UuC7JkXyVWZUt
jqRyoBz4dAOiLXV2XWscwzQne64+0amRtKBeJKZMjj9SgIv/LoKOGJRLV2GYZQndXKD8VxXfnc+o
VvkFhnUZWR+vkXms8EPK5sSlVSRcR9+e0B32zMy3MCBt7VqRYIyHCJLtl1fKhl5MJ7wS1LMNEKr/
Wm2qEdspa18kgkKI0CkQhWV+SsQs4T6QmZWZrhf2AB/quJmqdvx7WLi5WwSm7H9VfzsWg/FrAP0P
NL+NnvOAXD/Sb07fQdpTwSywaqpElye56xuMVeyyXuQdQnSNTeP2MH6RfQ/d414y7O9yEYlZmkuj
YIjMjg7ccDhqzki4/JSiIZoPLrxeLyCSl97BbpgPeXpQIEc0jNFsUuICwo/8CxnLESCwB1NV5ZdK
HmzMQGl2tMv5Wg8b1q8FPHuuzzkWqsey/nqmQ18W9pcVioqN2k3Kb0WDeEKsVwGcn48Uah8FBaoN
luUZGOO4PXjJpHqPnn90MkqaOWlidGOVIeODwn7N/4ZliRLUcgx7qH/vljUwIAY3tupnL1xe4cfB
HGMnR1OqR0j0Ndpg4gAeeItc5phjyyVsRIDwxzltWLt2PQXMTwzelKb8AT3YQjSW0P8dyCXcfj49
eeEZi+QkknGOvjdVDtSlaP/qDzqTe+/JVCrkOmyIIxtpg+abytfZiAhHHFjwSG+KR9JROnshRKlI
fH8qWDTFoV85KnAGLIY+zuLxhr70SiPNtb4fxXm657EqVQ7cG/WSAhwWZl8z5OPm/gmUXEcEAyVu
foUz1JPuXIeb4IMd47kn0p555XsOMe8UhVaVs41qODaUgHfh2XWRhaaFPlNZb+WbiRgKDpVNdYKU
rN6oO+SwZKS2GDAxLJLizP8AWVZ1ou76814Ym+ortGwzCHAKyMIl7NTCjjOOq2naWKoSEQHWw30l
ZwP/0qZVvMTRSqOW2pRH2AAP6Jx/4y6qd28qnnodzq0wD3ayPps/DSDXqO2zOBuMm88pS69t8a8N
Yp7g2uV6XoFlNgyr1bgZ/hYSLwwC+mJqdvYGt765iX9J8zhYrWlxAW6yjRnPmbYn96WVRyMRggb8
3hmCRmY7faKX1Vl8mnsKCD9nedoO4KPKM1U3WhI/krnjcKayzCZFC9MtlJqsWfX+96RES1wVqlfs
w4eQgoHpxNup4aax7JF2jwQtaq2Ya9NzlT4qnubYJGs9HkbDO7E81Ms7Ib2ngPYwQcNmYhtCHIKC
d5zkFvqhUoDuXrDBNn6ATeI308/xUyTPmF5kWf0Cs3MwTkEPujSQQRj9f6h7oH6IC8TRnBt53Edh
vEeCT1T3mnEch7NH/JlZd+IlYTRj+UT2xw5AFhrEClWlersy5ULzHOrkZHRpylSe3b/GJ4+aVa4F
4X1XeivNccXST87wiFPs8ZNOMrdj+RXBW3MuIvrJ9A8Gw7vuMsWYh9EkGqkBTg/dyr1CAK+sdC05
roeP/sDgrh4tXlH5AK+NipVv2UBmL1AEIiWSTlnJYoh/Hl6c2pauIiK0zmnQiWWm7mvDzLOEIbFV
1U9BEpZL2xVdqBZGLPXHGnXGlfUq+nT9O0HbuDapbEjP0mWgrQonnAZ89l9s1m+V1O77NRY5wBDg
zmcLXd6+59iSMFfI7l1WmwcJnD72yXxqicBRsXIvMOaattZ4Sva44kFs/uXTuvhCI9/K/QzFnvWV
NWxEzHvA0pbROaSjfQU86pu6OkLFq/ATgwDOWiRwVGnVYhsTaq+HSjjt1Am5jy/3RCgS7nfRFoEh
BoNZEBWrGyAPRxxk+Kv0sWBrXClKe+gYTiLNX0FWhQqAna3PVFMnr0TI2Hlsrf7ycYGHikbBOrXS
rt1cx7pPMbuSBQsm12gVUXegnp5Y0PkZ80jAZFrHY2WMyhOy5MGceGEeexjn2h4WIsQDoHiOwi54
IdNhpmDQuVpvzQBsLJY5ILW//Gy0wJJcm4/qK08y8XutwGbiCmj7v6oO8jwEPr9WvuOT/3SicREv
OH+L1iSz5mACLsel8IROArmwkksKQ7N6XeRoMbupuBlncPO4+0rDqEMNHetU3fcDc2WMb7EaDUV+
jRY/KVLuz02SBMLrsJ4BlMZExdXsCFmRotFQ1kYBoWB1UQJaDiFnpBbT2FSeJZtcUEatMry1DZiv
tS+uzIjgn1yodI9RDMbcobWi5T2NNoLh6xZsqkLfeoDggJp2GUzb4qFQ5wIMpOyXWrlvVrIUDkoC
6eD8Fw3B1oB4YcmSscxqbYWbEm0ISZPiiL8pqY0tb6mxhivDuIAOfFcCUAtP1jB1I+baYZv9mIE4
iw1iR4Z3MmW4mFWkVEF5rGlPagRy2eENvFUQEV2tWp2Z6iwhGrdq8gAlVAKVRNapyngsZYS2i8PZ
l4spmi7t7bmzYL5c/570Pvz53mDl/F9geitmtC7oDSGCUJgvGACCMs1iHz42MbLUrlOyRnMTxTJg
0IR63/KCIxh5a/n0byfqalWEy0P+OtlmkD46LvJ7anvT4bJvuPs73i0OvomrZm77X+4Coc9j+vYN
i6OVo55n+2Wlm43AP4Durab+qyCfTo9hJ7XvfFXkBvT7D10ctOyx7+2XnT5J6J0TnItLHxKB5jbH
ZXrZnES1FHh+79TnD96ofFjE9zMmSvg7kY672XZGnG61bk3FqNOpgXXgSSmfyleiZwiZLsKJpmOd
m39We1aSFkLmXSJS9txD1bnCBARJcgOsjbrtlsRydBz68IRvscAVFkLBW9qv5itF+wy+NESLilp1
Z9Zgpi18U68SY1MtybZgEzbDpKvYYr38xtWj4MqBCuY/pSD95sdmW/NviaX6CwFEWB104yvxIBQz
i+oNrDyB0aa2wNExpVbPjBaBXkd4rdl3/kM6pX42SZ15F7ln+s5bd3JCa0y7hjYVEZBKYEvhlTJX
bE1TOrzulTHcwHfFv0gsNDXtv2rRDKmWa+Nnyj36QgUjx8e/En85FOistQSkeSp0L63InhuoDLcp
QSQl6XUId3OtzYyUyXj4L1g1G3FcHI85ceSUZCzkxBIObofr808+Tn1T8WUFrhcWcdA/3qdnlMG5
1w2pl9jBpuJCV5aQ3nYTlImY2c9PByA12BBDLRIs/noRMlS8sECL0G7KrQr4zOtItTiYpmdxRa+e
Az5HFwi6vQQx65o/aOvJK89GsJm+nWircY2A2u6/CWTehz3XDW26kaL/hrm7O35vWnedBPczxqGL
Apv/yKQKZ47EDbJaSKiVAChKJtPIdkEoHR1To8Caw6Ylhkyc4eGdmXWFxYkbf1zFWqcWWB4IJqtA
RKQNfSTUsiCvO1R2hKKq4jDx/DygaaMX/YG1aVEeais3xAGXzMEnlESqTXQr8lPmcAIovK/SYXkP
jyg+eddOMxCFrFZj3RyR0W2l4mTQrrDD3A/27fUXZX+NIre96BJ9TWZX421CAp9xaqujZyYBMsdB
XmqotwjFPoFnmLILg/KoRtMmOJ01TxSHAPkhz+r/nF2CbL6cSWK5q1zrMLMaPjLXwci+DKSLKqXZ
r+h3AfQH1sO5g8QtKADtzECpdt5tnGB1gVmipakC9TEWMMqS83KdJAhr6mQUjj5ncwDS/lLVy9F4
Z7TBdUh/SQ/R1sdXO5RcjJ9QzzxCpB0If2xiyfZbxExjAniOIHlEBURB3vlvrXeQknKOU/XMMjZ4
33HVowGeo2dYQw+hZiNXR53ok1hYAtbY6IVnfTpbD4BUirY33806poFH8E/xH0j0BfSlGKLunmaN
G+ekO7VQ5jetIRC+BqIqZ1rInWSMCEdYtzopVoD+fxpZFL0zou5ppAz9wGY+iicz1FT7Yowmlb9S
JWwTGJVwNNCWUp8sQq3cPexAaIlDSpQS6l6pAFZxXNTTKacEcaled0taRmbZvrnoFqSWe70C/R78
shRp+RgukRwuRlK23sP3qAsyrfj1a48lEyrqK5II21/JEO4kY8egAcs3mK1wVaX9NAC65G0DowGq
h4Lre97A8M/DpC9Mycf6BUz9RlRT5yl2qQXXlYCYIKx0gRjvMycpr8xeL9genu5PEknjaYf47wuH
UULmgDG2bcTgEbJkUacWUmQhHOjN17IDqU3sLUXntE8XuZE5hOZ2TTj+OWA09nH4j8T1LtoatLgy
VmeXgr4HDIUfyLLKzWMBTrTVJttzhofwSpFvRWG78XXhOunkYmAsfue49G/l5abB05isWqushvVJ
zixSjB9nmGd/5OyoDj/isAEDlES+pb5ZDkQHtgZmOH1/DTi0r1GKRL9yO6n2RNkdi1OZPFED8/KL
oAAzyIFzryPE8rsHpwQC5uUdejkpg2ZueWs2lc+NA+ndKZMgQ3qL661ilJ2wMaiBW5FZa49sBxXw
ypxHi0cGV0W16ykMvZwWYQlKZ48Yz76Yi5JmHie/70sHwu+FVTVntOdHlPtZzc1x6s6DlM6TAM+B
K9eo+ppxfbgg3bCJpx9vImegslPNSjZi33OqYr5nddYBraFDkB82uE9uTZRnSnP14co3eJoT8vEm
qRge7eVl6VxEwqkiHr/jxuR/1FwICjsHdU/s2KTmPGt0tMA54y0RWQqmZsG54E4vFxSs4k99ptGh
vc4wMnm7MmSS0R+WRWLScqiey4uRtNcazQ7/I3AEPDt3+24p/xtLQaGz742E7w/TOvbUxEt/HUDa
TcqIP8RuV1JxJTlGDLNVKxackmi6rmWFvdNfE7H5U8CHR8Iz8dWP5ZwavoMUMB6ywr149mvd+4mB
IqgF+UqAlVyZzfvJZiPCJMQcKq0Z/7pJNib4UmZEm3S6B5PLZ2L5kLUfiUI/bB1PLpoMFOwcdRx/
udLQDlPT0Lr6ksIvQO64Weq+CJvOVzZRk401pSisG6vM9n8IXsvljqIPJUeicqexu8FYm7Pj7fRh
WIaNhCLdq632cOf4n8CUND/ieFv+SsZnIYexNu76LnjITjl95f2iLM4v8IL0L39t3QBg1/4pZh1x
7dzj+lTgf05sXeTHIm7jaJit05h48C/GiYtKWFT9gpIgCQ47vmdl0/PgHcqJL7cokAJShU8EmCX4
E4BsZJUgkoIRF+uMO+klA3G1b0KpTymF22uLpD+38nAQWvXDEG1ItvECxShJ0HOJrBnyO85cyJf1
uczbeMotO/nd2nFfRrFlb7SU1Q55gt9SR2CgQhJy0MmG182Ab3jw7bH+4W7HTXJFjoG2FiG0v9aY
XlSW5RIRUJQcplZgnuWTiq18vrVaxuQ+SdPvLqU5HwnydAMEz9BGugyoiuxQOGYaqlum0d1ovy4a
TV3H/GHDx0zcUn/yZndXzUMk0kmBXx0KLpYl1DVSltzi1eMIKcj8KJgWgGpyx56InIxpcME1kIFr
L5WSzVZDqDq7df33LjguVM8VKG5naf7ib1z12YpqCYtfB7X7vnxTETKLG1Zc0j5A6u4k1kuT4oSr
h0fLifKQ6AaP00flJMEQKfe30XISJZIQ6sEiKIXWCtDqpV6HfRWKXb4BWG3iL+C2wplHJta34vP8
nnGxcR9k+hVQVQBjjAaR0fH2seohweGwRG/Klj2yHxbjbT5Bz4yuGowjudl7wJsuocHossGFRwZr
YCWuFonASmxf12qF/EzHeDie/o39xIf2YxyqhJzI2mRjO2IyAv72WEGodAU7GZsDj/hZ9usrbTp4
ZsurIy1uEMIivZqkezEejx/RSM+LXhT7wFckMgKaguOfPPg6QxE/4kmKf40jJW1LkvTcGMuxbM3t
SJTQr8pdPa0sEWhinvEJN/O+92uppokVSK3K5SlSo8o1yKpadYIq9M9TaUbWYZwXQ2oXIGG0JRsl
OwDIR0nhcCock3XCvVfUESUP0lzNbrPhNupdnSNmSyrZ6eP1RkmSVOk8sevSnS1y+l/j3DXaZbMm
9RMKYE9yZ1RdOzaDQgxNg/L5/i99fHa4AqwAJEn4WJLKvm4wws057LixJmKJ1cASFGJnBU67riXV
y15nsEuMsmWqFu61YAcxA8zmjAJwAebh8LYs7fdFFpdmrcRSZ3zGI2ixjnObmwVw+MocEIXGEmGY
Jv6UlGXOyQgeJgQoj1wyJDvwfbRBn8cLh7USbmMY2tx3lqooTruw4FpiuEMx2D3ITJaYcdE5KguX
9fSVh8x6aqQMS2o3ivG91dyVXVq+K49NB8XGiM2lDalzaWaB5ylvT3JKhbnJR3KyFWXShMdIAnyr
KfKQcE8Rut0p1pkzEiFpacQWJ73Ea6Tl8yuU0z4JrF+9nb1TlBD2j5ZCTH2+z8qZP9JCTOjQVIps
KVT596ohEWfMyjIuX0TQzolsUwjFhOByBZAFdS9mwVAF21hpQbMj9r/LS11azwzvefRRDggH1sy7
RLBNCvUJX0QkHUeXsU0/kKx2f6jY+06NRibxtsNj0QjcMZEjTc9Xe9W6n8BewwPud69QwcIW8JdO
qQc+j7CFgAu2mR/nJxXWqJb7wpb/mCp6YKjecc46rGopJ0WDtqgo7IjQKDEaOD2TIeB9FSyk5RZl
FgK8w85Tjx0gvqkN7hvfDdIJ0MfaNzD0JXi/05gvqRqBO8IqrlH+dvf6GQdPHsIWx4cG4tTszOdb
t0ZNgTI0pWfhpj9mQNbtyLlnoZUDcrLVyzzGrTXL017CuCrauhGdWuq1UNElWoJ+hrlYjq2q4FI/
Gndu43PpjrHK0hE4j0DmAtw/AgzJM8QmHQzFs1LaVpEiFnXEMvPv6Dr6ZgiC0y3ZTqSmD8QzuGSW
mnaFzH9PaT9hpSO986XWP2V+ziJD0ngbGPEjEohUWOtXAxB/fTye51Ju4YZrBrwYOgqcEZnjV4th
SqrjZsQjQWuQCzSIJrvyblWESGFS+hviGNiFwzHPMD7+m+TSUbO0cJJmbNawV9y9NrO00dl5lNz4
pFHfdf6q6o0u+4xtyJAoX6AlPL+4VlIz4IXj7YMXkXXk6cQrNt80yXZTToFzHqjp+pnUW68l3Ftb
/Ne0GfozKWOrPdqQEkNBrhujFc6KywfwyM/77i74PrKWVU7xnbNyjlvYtv80NYPWXzeE9cC1Ek30
3wKW3JPVeoHdMOdLTDa2WmN8v1y5DkNrq5m9X1Cuq69b/0sT2ITaF2Y90NYo7wDb0c1X5u0qlQO9
f4JG1l41ENs6bjgm+cLYZAYO6xfhgIdh6/gJZBvdlhaNKmltuFKhfeJJa4dWEsLYfkcYNxJEVhy2
jTp1BHqG4xFPR5faFej3B4CoY3VZ8YIVJ7p47RvjOZF+ub2EYbI+r3Ro2lGtjNfOa8L20U7aEvn2
WZJxX+on5sWpA/vWDmuQKIekciJUB8Y/Ly8y4s/tfjkbyhmVa/bdNIyyhJqsEXHS1ZqLVSBjYkHm
ZQKKqY1JqJ2yWuEG9r6BVoRPgJ6kXGlhhKdSopsGJft9aS0MRFLB31X0WG9IQeI5uq1SRC9TyELW
/JzCJk4zsP7Kp71S+Ibso0AcX7RpFeFGkAjQxW1uZLzMLPF3K7EqQY7nG1O1g/Uioz1znGGLxAvB
5roETvga3AhUTAxJ9BNWXBiawonXW0DiTVSuOKiW508pmXZu0WkpxvUpLUnTE6/sOmibiBZqf6Me
cUe1p7uro+AVGY50egoxq06MZdl5kNIEbNygG40JYmBtNWgC9aBM7TDjSZUZstLtWq0l8pPTo/fw
f8/Q3SRu9XmiFsdk8w9w+nQnoSilJbzWDKYfoSsg9ExFWjF7CG6HSIdqUBzChRscVX7GgrWrfz4B
J7TvlCWjNRF1gc+ZXZUy6xwaBTr/IXR4Jx48dGK0+7YO1l84CbChD4l0t14lFOIP7yjUEQoj2KQ1
epVBd5IKWWDM6fStl8x5AalYjKKGE/LaHwmkaM4lANgNIVLEcneKDds7bqrwlvza3a0AAWlJjeM2
9E+Vxrd+QM3EvzmEYaSzfBYTiqX2v/FnPd4qfDm7UwqgFszyITL0MpRuAYp3MySofohY8UgRMNmF
lwIPZXGBgFq4pMemPWjiNG19y7R6yKjPXJKyBDhF52LiMVh84uRx5FmPOW80tRXF28sa5fZuM+EU
s95P8N6vpPT5JMJ+tnX1tANxzfZIAP9aWUVrcm7hNTUcRoenB94yPXbWONsNT9WQwRx+9ASQmGcv
/rGyd9jBZkgPvimXVJzgDptcq/ws55yBSiC3Xrx72xrdkdll9k9cKzhHZKeRgFinWKZTKGgfTPVp
CVqmTQesIUnt4CoDaPqTXk4cn6r3/pQVef6/s4ozSLT3c5uQ7RMPtVlYXiE+DtpCMd6fPTUhui66
dk49rEFGeuAcjXOO3Rz+IS115g3tXZkMN5hVqH3qvwzIofIoRj2E6cGCii1LKztzCs6dqCilFiDS
F2JadMlZPXxS/Si3cSF14hYSjGKaP1/c/VbNR0gqMO1bFLaC9rBv7U0YXrXhejm89lRP3A1mMbWU
LuH/nDq3fc50pgJUOk6TE2IoRsQopBZ2lwgl0gB/KBb96/AglJd7JsjL/b05dk4wbTsOmN926Og9
YDD3m7EmlDsm4QjzE2GyLMwvR6QrR97ZZoddsBJM7TN0CEEmJVohbnzhwgdFxDqKasbynZKYA+Wz
ceCakjI0H+zErwfWHxTM1S+naMjVoS07zErEanZQzB3h999hknb3DMiEYdJMCBDSwQBDPVRHTNNa
grNCDvH0l5adRHdhQp9yfx7eBKQsWbzFm9aQeHSTYB8sDIF2uabP8ywyDFOfOptp2OhAXDo2iWcU
i/iAstenWLiO768SGaWBHMxXesVn231TDnavPIOiexXv6P4XnKOtlk7S5pDCYemtBYjvixZmHEUf
p+hsrS5BQ3749YnmSN7xCFiVe/13r3bQmO1pL8eUJrNReug2Yj2Lz/wVu8kNkfBmqDdmTWSl2w15
/JMxsW1cSHBSpvJVrb/laq8vdDLRNjKaX3aw/iCqOHXTycVt+tVbvhe7zeUhxjVnrDDDNJ9KfHUN
/70fC6Z4kGYMr2bZl+Z/ZlChE2fgEEjN4qJHGnU7JuKvkusBK+jQ/tzDKvIIOdmRy1pvVYs/SJFC
RdwC6Hck46gZ0BrNaUSFsK8dY9rKKvxwW5H/9oBiMQrIQDsTqhMxqMyPPVeS06NcTrSC5ITxc9Ey
JE13Y5OUmXmIK+GyRf9QOf96EXQCivh8wKYXbsfrNI9P/z+/I18DDDaEn5wda+IIT8KTOLtBlehq
IpxNob6hOnRncCIctZpESgA45E0xmjE3kOQfUQ7qiEeIMPzdZZDRgvBQjqoie7HE6iMAZnu3Bndx
z5GPkdeR+oYcoeMmfDweP52mCn8DCQ1uEUVIrJKLzv49E1tMiF8P4ZFksF/nidjuhoVcNuTQHqWh
alefx65ptFhNUR1dIph28SbSqY1NIENZJ9O/cwfe/A7CqsT5BVh8xLoHtYp9HUp4VfLBchEY7uhk
4vFinu3Yxr9OLjicoEC6MftxvDNVOyZ6CiC9j4qlF38UOGDd1EhrkuzosBy/Hbx3L16dj3kv+5AR
pzjkjbUitw6+HYrV/qeV2ltSUTDCbv0fCUzpKMZvWLsOJ1oEi7OHic1LgXVffQ5wX9EDV/OiqL6X
PjYJ1rRsHP2lDCx74fhSbSv5A/Yr6GFsXRbRFZZsIWTvXeG6pnntFILF60smhj16Q0YH2YkdL2FG
ygPog86be7eCl96x8aSNFb/5R15K2GTeNXOKjigO7UTznUXRSoC/RQ2ze5H+x2d6gNwTG9E0pnEp
xU0X2hh1rW5HGsUshwO6iF8EcNuJGjQLJvKbCfPMdzP4pTdaaVxMgTrMpwBSnLXBKGD9utxsdxGa
Jjt8OXa+fnh93V3n5NCB70x5CT7cZUhA0v3IHuRlSxVYOpyIv1pDmge6mwFyk04KUvUy9YLTfQbH
/BMekIcklz82KzHPPCndAhIDCnn5lEbr+GDDt0JTkURmdLcE+pebXymhQE4F9kyH2PJSkqU30v0B
jtNDn96Pl+HhaIkNN14kH/Ovjjfhbsrjxv5YrmFSygT9A5aSPJaysOskgv7xr51tiZ/csiw5LHtj
10IhlC41P7raB4tLjUFEcz+HO1fSyhqOl3rE0mz9ET2sk6+FDGbrTWIcR95EB2NqXGOUHPngwllW
3t7e//MU0+VgOfWLq+FeV1xmhActtPDSl1x69ZoV4QdpLOpq+8N3RV+YTo3m2z2R88Xcub+ilcQ8
Iw3tSFoRh1/GBqpLJ164FtNgDZHi8TpOcQnYUsy1gydl6/QdrhaMgJkMVl/6bPoNotwKTW6DM+a0
Xrpl1l8G6Z0QBK3AoRNwxQUQhNG4UYfPBB7VFEHLhkfoQTeM7tQWy19x92lFa7Ov9e1Lk+m7oNNw
GyNPf1giYoC4MVCTNkUIU2cw6Cnrc4yak3UZ4ZZ6egvFe2y6BTmFhGOzHMnDKzDtu5Fb9DWdNCfD
gdgar3FrA1TXuvK+0xxS3nl5uxPUl3HSGbm+AEcEO4e4JvD5cKxwtUI8nANg8we4jQQqYntMfzmy
I14FUBZwiD5xb2Y4hQ2fWscVtU/GOIFcb9vR0zKCjpOQXhJXstYMV91NUHO9FjHZDx5rjAolVN+b
r17CHL9Cu3yVBWnHotEcpd+EyVazgjtulfjMcW9WrtTjylzqMjhqaxX3xn90TMLmHTnRQa/RWe0A
pqi3MOqywjBCGpxKHn5uWgVolUYoRhAaFCpQO9atvJOn51Dkcp8mYQj0rameXi9jtPm11nTMhTPY
ffuGjVUW4rhuL0ZkbqfQOwMKVFNRzmwJAext3RgoPczV/orkEq4Ayoxwn97CcDLWW3IY2/DjAxKS
9KylzqfvXQ+m05B2bKrZlW8ztf97o9eetkPmxeMH39PLhzybRteOVv0cb+JSAVzyHz86uY9qyjRF
ZgnLEBVwSyAGPOtHAquFZB0gfH/FB3446gYgDwvvqfhTVH8IdI2lZuQlBOjWAaDUif75X8JTRUuW
JnvP7zzZiwzF0FM6XSgJrERxiwqZiAVAgAl3Zsyntwn9kaldBZbyGDtlHn/4kVGO2ynOKfyB7UIr
tnf9NQxDhYRpRlLbtC9RdQ697bgiccU678nfWU18V4Wxlho7pJ3LPumhu8Bh7j+eMu5eRONhab0J
pjAKrP+RSu8Vy409o6J1fBKdBz/V3Zzz0vrngzwCFcX6P15ZzjMSDHe904L8vvwB+5oJq6T8O4Ew
XiOL9x2VDFUwa/NUVo1rM2SJ1figbPitqYFK/ZltTvjiQpMtxQaIsgj76yh4IPIUP72kBjjeLxye
m19etUUibbXRTLyngVzNW58R+S4uMCq6Im5Qyv1xdFmc9jkyzUCMxI/L0VT8wbR0X0PvXzQ6vN4n
aThhdBP+8CAIFh60fSUlQP1E4/mr7Cqd+Kd48wXUGZTWxhUuRHMDQm13ANs5pcXJ6sKahjA+QzjM
4GGK4cGIdRPPxd2cDvO3OF6TwwBiJiADIHIpA0+YwMh2dQvaC/CCwtlNnZYqwxK5SHLLw2y/tXKk
6/D6TkOOfxlhfm4/NIfqHVQW8hx/HycRHsNjTJ7lmvjoOHmU1zW3UOC2z+mOC9vWQHxVsgVbN9u3
LIk0i5ycplj3ZyRg+/OJD8arjhjLNLV0+xMQ+7ePAnFdTvsK9D8rbGMawveifLTzQHX2J6D7FkWq
c7027BmFALBI5HIdQY69tOkjPdP1VWuU8G6pvXibpHauuAW0pFjgRdP1tX2thxvShRNKXFOs1Uit
tl8lNeIrqpKwSpzrP98CfFAqt1y7JhXAyQc+KynJb4W9/xrm+Bnsa2I/o/DuOnsvKFu44zSkUX0i
O1EuRn9R2G024C2j1NkflVh8G4ZMOVukoZKS3jqlBaQHNOJGCgvxoKgTRgcQX1mkGoIad5P/FYtC
8Ig4hu/HdHuaAhkGh0WbJkGt7JJgrCX/ot7LD0aez6uxumvsLw8FoBSGCNAU11C9jrw+POIO9oYb
nSPCTythRwxGobuEJZFQnjltttRrD9RLJzDHIKT/vkiWjL+M0FxJkUOuuivNB3FopsksnhNKGGaH
Dmoxe0RvenPnPQj+oNfP8KXtAwlBTkCrJO5YYhgV1MX4tkmdEwdIQegwKQ5/idJaDFe1CRPNwFRK
GifFWs1e6UwA8Pz56nAwvDbJzWVkWFO04zCbDlDYAbEBevOdCr1IwR+Cu36p7uH5Qi4ttwa+qwF2
l5SS9RyBHBQ98sO64FzthSf6BRNI7l2VwFVZsGr8t82a2+JYMxUTG+rjIPQDfuIO4g5y9F3Lk9NP
1vVilzgC5NVEwWVNgQF3DQppzrwIzQ95kypgwpHtsWqFsvCnIXuJcmyNb5Se1iELrXr3d91CHGd/
vuqaZHa5z+jQPVNn+QOv5e3i9SqutBDHCR0m2NQcoYWQeTS+8iW54N+yd/I9aM7zILWm6oC78OpY
BpYsw8pZBTv2Z7Z7WNIDtdcBiCYsM1zXCtDgPFzUVLv+QHwF75sj3GFNbPO0ti9ehFeBDTEgLF31
yj4eEWPIhYVK3pWqkIvKt270fs3clK8e42ZzvuL1YOqcH4B3HU7dsHYgdjP4xRZ7v3BX9vqIBzEx
aoCD+4Mc8BAR4tRig/bDKQ8JhjG7FhaGIUFI2cAB2dTnzTgcxFnxQ0F1oHE73PWlWkESIrf5IE1K
7rRSiets3xpNZSGiPYLCpvu+UHWMMgbItYNLilmPilbTY5bqd9JqDKbNpwKB4HirtAUh5cYA0mdG
6lGo/hMYzmUO5vMzGmmkjuXlni00dxG09Xs2GZZP4elA5pzpvw7pndyIzn8dyX31Mn1miW2naIcr
quPFRDLvAOOQ/AzpMDwK0xPcJXfHd6zqVExFcWOTrPhQfoqLWYHT2XVihemcL5JTPXm0fzG6bwjL
o1k11PvgplaTVak5x9tBHlJ8HwvAItMUPDGx/OLpgCU5TXXriEfpnsgpx4fdB8BUvYZul7AoPf5J
xUA62V/F3ZOVaYIpsgWPatPwaRS/vG2xfTkYXX6EVJGLxxNDMdcMF9ThNNo3zj/3RBU2Rn9ED9M1
mT4NW4p/CX4uBNmaHHsqIylBQ5FHnxHqTN1kcLGeXB1qvYZHVQHq7JoTVSD1irKCP+L0c44l/JXE
U19dus0lBLT9AqFzhQKk/3fTolEKEhPxvRWytRp82fTPYF850pgGuyNtkiyZFXLXBR8TlI2VOlE3
FjcywWyilHZwKoRtN67azvUQi/UBfiUkGpBBP1uklhY76Le67krZfn1Hqa67kQVlDVzrhW+/kdoE
xJu8QyTa8iaeYdkgiEFwz30MIqSoUi5Kb0zaF9EwyjcniNncPDK82IErTRRmefM5HCU1PzleGo2I
7iTtUVFfbKlnbDfXIFQDt2+8oPtQauYgfM8bnYdUcsB1/1MTapuzAi8SEPxSlWT6IG6SNV+R3ycu
YHYHzAZrlpTNELbVhE2AX/vzyxudr8hrqqTIims/hSQDvbkibtFCVFYFbzNyLgy6d5tv88CJ3TxZ
MnnmFhKYORMPH1Si72cB1DI1BjuCYe/0YtyS1on1x2VAUGD4M7LANlJwGCGTLOZEGUQX1hjiVY7n
lOKD0SSF51unWeLzT6yPl352MbSNdicZtBzLqPb26PKeHcWnoqxoezOTybAQWoCxUl4WWkZL0CZx
8TD+UOTOxF/XcLs7X60fruhKCJ4XSc0f2nuoZE0AP4j8CqzRofXV/U0+sb4a5S4vuNd28Kr+b3/h
YByGdk42+J+U1QjQ8TKxGlLlnoYIzy5HUt7NURQcv3bNJfvGG1wqO/LU35toyyeKEp5v6R6q7ymc
/pQi9US6aITbAqf+ZWjHGh9yfhl1qKkS73K3ePzLUcBizfQx99yh8BP4SCDGT9+eMtnK1HBKQ0FH
LCVa3qhMUmJNQoS8MQXUm+qNTYO/e4+TKSJ+aW3ya1/Zqqrumq4Cj3wEJCvI5b97YxD+aoCFgg+S
tcaWKm3RX4yV6E3DtfcaiLXcoHKLb0m1fImwQgxtZydTqicdoNCTGT4nXYeg49qvb85EYz90guG8
dOUKwlaBGeKDVT4QblKz1QBAz/OWNye0OL+af81m7CT/3MNS0attR+Zb8m/hxlAZj6gej5HBvylH
roM3rXr1mxzf21JC6D1//JClwaxAKuRG/5XVrHiXmpcewt7B1wmzJPoIC1WiBn2nDdgCBtgC4/Nf
TcUKn8hhZvx0sgbmuiNxMtwd5AZSE5I9lyu9aIBcFGm9KCuDy3G2LGgR1JC3xDDolkpZM4fAiJrk
HGon4yO7kcNc2jgGyrMOOs3EL+UGqR70r+/vmGtrp3+I+oP8mBbc98bkHWKYhfOssD/xXFDwVdu7
799cgIHoATERBFWznX4KAsg0NllQk/3nLGXwFX1h9HaRBv/ov0iM4kCIhIxIOOR+6TVr9AqQaJhk
9wKyACnAzH2k0dmIyWic3lCWhr7QlKVBwF7hSCF+Cp2n4T5Qg1CudhXrvu8RLaLS5RD63osDqALW
fjElaUEuM9hOhxsp5tcWHUEQfiu9kBSHF6YZ7yMctQ4x+dNkmKUmT3YFOGRqUAtRi9542id999D7
qbI9iGlSbEj+RXq2mNo14SVG+syKi9OA133WRo2wraohPHrU5th2NT5ZbTVrbA3b/5JazHniybjO
8hao7UzTDLcAcgFUBTBevE40khocbQyZAgjqUBVzMO0t7WpcRP0Hx/cRnHgiYllvGV3vpeBHbV2B
bQAsj1SZR8ZtrKepbRTwqHupRL9ww67ZSbm95/a0npR35gAdoPjs04+QdbKPuyjdwBE/9zWuQegw
+HkASKtt4i1BiDEJB/HUIYfumOoHBpfA32L/3snTOyFSoKL2DS5foSQjDBYr3DIXpffhzdZq6+yx
HV7Gg5y0hvB2lOIP/hG+Jx4JqwhWEtAXevWVZQYQkBAlXWm6rWP/8TLdqZiQdUwNpzsfXrRKpEJr
ZHDdAu0eSs5QANUvPvS1XOsnzmZoQSg+Ybg3GEgpSntektheMe3ercPGE/bHvD6XDKfv7jLC7uu5
phQMx1SObnNm4CjUYD/5L9l8DAvCkZY5Yy1XWdwIoEXf33qZbNtJseB5vVWA+r7eoBGTFD5LPpZL
27748KL2AO4JUr5C8r56MBBNoYwKA42Lzkaaz9BB+H66LS/fiA0h0qjIqywUEtSLWh0YfTQEIjh+
qdvUossBeL+7HcLWKfY6yOz9jYbBr4FIfy7c6e/+Agq16QDLkLtdAmybdIDg2kZDYPy8xiyNQXMN
rbmHyXB2RjDRykSHEBYpp44x/VXW9GrtrxZfOZr8I41qUUNAF7G9W9h+tkLQNxj41dtYihk/l7fa
dXI15+0xD6mvN1I4BXXRN3dMHDob4jp4kMfH3CV5nscwRZptO5rv1vBAsbRf4bW1gsZMbecAxiyZ
PfKz5zZA/a1y66E0jUvTr5O49kv2AIQSexauKs4kua3s2LFRfwaxZ1RG/yftsWXE3FroDAwiJV5Y
K/0zre7Z8oLYMVudyhn74SReR64BlsbxJKVfwz55MY7kM8NbbIH4yplKopV1Og3lSmC3/lAJ1OGj
3gYQ1QYocW78spnkccXNcX5jZENTMnthVWRSLkENjRDyIGCBbVyIqRZiPypE0BAZX2avnEDdBpUi
simDI2BndTlgX3N17h1lqS5BYKC1ky8zsSOwNIt0yg2CDs3tzqvPAW18EQ5mgDFzCoCjaL1vUcdX
3K2XVYUBkM5nhzT5Ep32JZ3lhljfy4ls+0zuiBPo8Ea/gAEAxfguaBK+B+mAtJM8XMZFJsQnsrjE
Ny04SDYVETfFYX3/Zf1g1WEgrKCX/ixpfqgT3rWIBxDluhCBs0/oMKg1llApxYEgV2dAxmDaB8B2
+mDHXvNnYo+pPhnFPeQA8RD4eWNrTKte/QTHGr/bwtfQzDmzWP1NKDyRcYY8XkOvUVaMYCHp7Bor
u6ThY0GGvvCaYvxrc3Yb5+HjVcMwjuYItxxbsT7T4h/deSivA1/c2QVdH2jLuPDpt4LmbYw9PIQh
D6gtt2jp4JZ4KNeWBWxeJ3vQ4/a0Lz0e6UiUkQ13H8mRJDPaMYktsY9Jb9tdDcXGOFm7U0PMttCp
5JYhY3iSzQH09P5V1Ap423JXKezY/byf9ujQKRnMubAtOn4Y2djI0GG1DIWRvYbUbqjpfDIEwjHI
daSOsCRHw0MnPyZe9D7+NkXGO8MblU2C+Q5p3QmDPTzr8NzpTEyxDdaT4W7o+Et9+2kCgPrBno63
E4hoUHzl0vKhCAxzEqsfED5SspMx4ScycSXn1OiMef5Zp9DeWwv+FRU3pUzcvpAB3Nh6fYs2q6gL
49W8xCBVnAaXgSSeE2OOdBM3FCd6xiENkz9ZMVZ1p3dzCJu3bLZ7j1gGoOwQSmh6L4BCkN5/4uVy
880Itgo3xh58HzgYVHTenttyuatq83j1FgDD5S9F1Z2ulf1Okyu6LonKshKH9RNgUKbAJXR8t/dd
law0Q1HRvB36Hj/qL9thvSFvKQcjwwTvNL4IitVvz10DOe+BIAV3OjywsjVwTfG0cU+CT/g1kbPE
9wn6J5ZQunZ61+ucwWleG0w4vA8LZEOIa42Oz7s9MYPl7gkzLvEAXUb7KzMnWIKJC2Vt/927aXg2
GGwRqeKRp9XDjBbFzXZYzlAN3Sr0jzvS7in5tEUF5t3Bez4ResmU0uxiqpnNKxmTDA/CDerUzRX9
td/cv03ozZLVa+x32ZWqjvrgr1IrdGB2de1ge6GSFdpdu2tPY+u8fZCyLczB0UXdPFgfpIi4BxRx
chhjCa3V6qSg8/5e0RuSpVNuXvZhUiYTxS888oI3VjGpIBXyeH/NE6SlxEdvziiHmh+2SHDjTS4K
lj2YsGYwzoZ/p25xgGw7Q6R2zPcOUdRV9SyoIGsCIohf3piiJt3Yq966d6vcMWfsBlce4yd+8uAo
IpPt98Xz33NVe7H5O1c2mqzwpK3ZP2FPgbZ/FrtwjpZSsN1vRopF4MDv+vqzzyHq4JH66qAl5kMt
+Fc1JMA9yP8QUGKQ5jSdcPdKv/Y2tpXwr3QzozCbFKvAKuaKd6h+5TT6+yQmG5j3VdvLzVqsOCP+
3N6EeekXNXjlnFr3AXfJbJ7R2Rzp0pFm3mSE0SjUNbELV0HUsvwQon/AOqzbxgNqcoD9l7iJ5w8y
u+Erm5sPurAvhJAwVlSMBFkB/AaN9dEHqfQNdVWpiRcj3TH/PvQWhfZ0VPfKEZ/wpqO051YvJ48/
Ws/JsYRMpvC/j0UMBwKPF7+R7JZO5k2iNtAoigbvXbCy6f8YDJWHHRDHJFq6dXqtQ1Z7lSbkPc+k
zouPzQatL+2+TgV8v1Ruw4OUevhMzLCIHnvNTkeptQTWx8vWRudnt22HPDTm1lZlW4zkU6zEnwXK
BkKIAs0Qi9ZFtr2dDdojPlp9CefZfEUlD3At9oI/hDoVS05ZhoqE6ZQ92Cwdz+d5ImZLLE+YuWFB
0HzOTlNjh2pTlx216oEXT/lneBNsonU9zY0DbzBGzaP7GvmZBvCNLQobPFGfuj3sxTQAunqAY6+R
5GrtIUR1g7+bVP4dD3fBldyYI/LBqaqs/vkEdG6BvFOLabhQvkgLB3CFV9gas4iRe2Ho0WaoLqNG
XdINVRfpUg6joysXUnBjHvOfumiiKgm2SZr4lpFn8+hjUz+3umaqqWBuuBnaVwvVnHResMR3a7/M
IQCxTFVi6HfzmwZDEJw1LBaI6SMPCd1ss1Stf3IPcIS0IUxIie+GITgZDchUcc7xA4rnoHYZKaU/
yEqjGD2d0mxPIyxAU3WjAaYHKh9CHtqhoIljBWtHo1Tg6C9Nr3IAAWwUAJs7hF/+w8OvK4MjrPGe
mYZw/oGIepiNzigwK4kMM71KV+fVnkL9c1pcasq0/SQH62++uW7wFRjqPe5hDCfvX1cw1qOSc9/c
au2ub811FL1GnebtElEeIa9nC8577zvCs4Zu/YHaD0A3X6jX6FOZLlTq2kVglnCIn15I2U0Ts8bA
dwGShMY8jNehiv14q0y+HV30zvpMYcNs37pFd2WUD97rMcRwpzMapJ62Va1CLA5DTzQwuycrK7CG
gdC8qd7zu8UTTUPxhz+cLqwAQSiCcrHHY9h8UTdlx9LPhchPlkAxrRuzV0je1ROSo1Kac0mH5jnb
BpmB1z9pMiWf/zspcmKH0U7TqKaJrB9Pe+7Y/fq99HsSdSO8JD+FR5LG/mLadvb4NDU+OzBgzWuN
BhOIHWDsEnPVJgphT8wJVXLi/x2XqwYnn3JUcXBgeiw7cEI9/EyvC4QuIIQn9me1au+EKlqLmPWo
qNnZAxI4sV6Uc72jCirUjEX2CeKdeSBukvibm7VS3e6eFyJgUUx79z62oN61CN0crFl5t6Ro06N6
SxvdeR/1chWKFWnxT6G69ryxgH+Hisv3yg+9+MY2GYjWKdWp9tM7iExQWglR7zmyYh+RrxwBNGHa
plp0uxiO41ByoKNa446S+twjjBaPNt/Qp7jUU+kbzIb0CxXkg+vRP5mZrIGRuTO2J+oHiwD326sv
D2gCHQmUHAxVeoQEeQ9fd5ps7KUgiI/gFu74u8t2PbH0UDemhSrh8HErgGDSl4QrVVcRqt4W0nOE
gyrqmFjI/RpqDlsnVvVdSfbOqeKiKbRs9884nOPr1YD1VZzKseethtll0McT//pEcxN1h55jvqKk
9uRyNaqAsSG3+AcxmWuWPjIWCGnjJQ7zaaySQmmfJ8dTdAZI+O4WiJ9WQ60MY+wGONIsFC3SzLLb
Oa5ccWANSk7hCFmlOB+Q8D/hkj/TF+pUjvxOcPmHhbMtGM09w+y1A/FYxujbSCVEmw0Yhhm9ekDd
z5E2bAUa4RJGcFMScp08yb9rNVktOS0ONJDkMsGEPu5Kd0Y19YKzuEVFPwT61QLaHVb0G9abyog+
b2jALi/6KiyPjblgdQel8N83KASsKIqTqFUiWmvO6eLSy2jSz0Lz4vb+oC3AYt5mO3Wnm7OfKMVv
ahSM1LZI2m50M0+uzW7Hngjb8EyuTIlc/cDlKB2+e5S8XxT5KemaiDe4kvuVMO//NmfCwEcVqwOn
fce5/RdwzQBWTNguXovbmDAKyksn3s0nl7rQH/xbfyYM1+RvLmkxxXoejnxviUWV8doCy2Q//449
Yq0OwvOm7meb9l9EFm/9XqZcoVJ9caczdONW/au2qursoedC5J/hvNj7/hN8wEYGvGTDMvnMLKr+
RI8Wo+e2mFcwRDM+D7Ahlmw6bNcJ0dquVkXhOguCMOFWehiXNmb9vdDWTDfgQEzHJmhO6Py3Y1g1
5dCWYMM/yTHj9QFwIt7hGmNZvEGGlf3UwBsGROnbugkc6MCwlazow/jH2q4Cfc4Cc1V7T4qMGpKr
siIPC6yc2WgDLFIrvEyl7J66gcKN+cd4sJu9TPXQWLYXh1nwdvm2u/GjOrzPKqz80tVY8mYiez75
/AoXVeYC168Xh3tHKFoUK48wATvBoJt0J0MpX1qkvJbUbX2eCUC8PcZ34Hlbrkh4Ke+awkCpyjbS
j+SvNVrLVYx0lvA01EvHPPenJRsHD8f5N0hTy0iuDRhcB+Dz0P/JUy0D8azx9qGnNaxlIMDPZ2Sz
H/mb2qYEozBrARLrV2JF9GDB8+PaW7yM/WjdFfNSe9yWcIFwU+NvJyfXo8MOkcwqirePE9o4CjmN
RJmsIOuxAS37z0+bOqvfeboTwF9YTP765G4qEBv/XGaeEQSFX1TMM0s/GVfsTjyoGoQVg0z5NGZ+
T9+xz9JbfW2eLpq9e38s4uV52bOq2jpPGhOM24BuvA+UNwk9YS6dEm7Ga2oWdj3WQGz5C5QVqzch
63vQ5Zb+CXQoXLcsCaMLvghfovNuPGYRjIf9X3g6hpIe8Oe0n4lzj9eB63dQcirdpOzO29W7emrB
ogWsIeBjKjpUIa7GWu2oSNmkxmNlqDBCOt3ObmvZu6imhclWuWW68UoplfvGID4FblABWhvvhKwu
iiEGyRS+JCN+RVNK+9cA71sF3fKm9ixPG2dM/PXumF6DJ0kfO534Vd9zTO/s3zj0M1/rmoIc7fNn
1S1h5Vy1L58ViUKSlrDAtu9TBAg+fNuiLyFNdI9Q7o+h0ZXZaP6xJjkq1k0XTXSiPVr8dS2kLMbd
I9Ni/Jj0wESGmOixVHx/mslaOgoumeuJ4uDCPgDNa/W2dGKg5C5v0RFb60uWAna+oayzVN+Erc5J
4k5uLBd9O0R1+gvmXW6xJ11BR2h4jfxrvn53+TNDdck7/sp+JFC/ZPqRCrYGDTwsCaeFWjWmElP1
+nOlnsaUzSZKs9WAMn0GV/xYEu2o0Cl+zZC5edBkJjCLNsyP9kgI7cule03pab5+odaZ4dxfTH8K
g1QfJUc+j16wAyBmOmu4pHCuyhNK/TP/yTuZykmXE/e7ch/HvA+VGZFL0p4jL7lEz+k1xwi8OfuC
Hpnayk8Xj5EWf8v5ZhN4kFMR0jXKzoUbS4+NRKpYk6Fc90qEMyGdc4aLH7Xoe7ZC2qGx+ziLKcIS
7ceFkMF5zQ/cRdKV3yai2dGJFLPOzUKlmKVP5dF900Sg/VDfckReZpvH/Ge0rdeyhcXiqjprQcqj
BCYk5SwRURUbp0q2jTBZtTgHuclrx5PqEmtfDsmC/z3hMMPVSxHCsk7fqKClVucJvD/x1OpVwGZQ
S+MUey5FtrBXsGmu7pHpXybbeWyJLk/U4LDjZu5PZB3abwR6+qMaWYEa5OoCVkwVx6pWgOEfB9KM
8LGB8dpFBbkMZBWdTlJ6xmpnsZ/r5S4KATN5AGbz2SYpkJcx723G4J34osHlxzlkEcwbTKSrPuMA
2MlpDTZFhjOlGnysssfTYXjbUMdin/EjoIoNKNprjFVGY3jJhN0OR0sjSF43Mgnkqgfq0ISMC5yg
/oSXigwisNR8uEUSzQYvBsA4uP5+mDdJOKNJHCnPtPygfssVJen+K/lticfGmT8INa9mkdYrUBV7
UvTKy3xU9eR2VBnm/D29pqqbNmmN4t8g80kc5kC6vn2rFg2X2T1S6Esl1QeV6S0RuhECFCWdYz1w
86iIzU2u33kU/QK3mqv1WpaXdFd1U4uGicPFXxYr055ijPLcWzZa73HcpVNiAAjmb62mr80MvE76
A9iJQyHNcj7ZQfrxdZBsYWzjlodcSgmWoAVtRHOAyP+TOF33R8XbAXfk0BBSCaNeXoenIH3s83XB
e2YWHTcviJDTT3rvbZTudrclF1nhKEd/ZFyj9Q0ZJw6Wc8EvE9EZVtgRlu2p2ICIYZrQS45zrOLv
zWCDTny4EPxPuHK2GI5munPr0CHA3fJRN2AE2vEzYfU5xqzTgCbFAcTCdtr5a7yZ3pwnQE66+DqG
zrS8C1OfiijcsTV9Yvtpg/nKrWUufGaZiWVz5O3lHgic0laCK51AKJQSnhBLwvlFCD1WwNcRu9hQ
x6zgwql2E6nUYUiUJcP3xachaebO9HvRqXcQpcRYN4cNLcSP7SSKp/iEGgZSh27jvt902BKT+UDf
VrOL1POJYr+EFEWrPdr8CWPfKqu+8IFTGcTiIn7W/Njoc8D5fkjQEVLx779/KXEj7a/H9x6WBDH9
BsOTA+KiCcsWldtLdyolobjJmal8DnzCikdZn1BKbkEcivFg6/r0WRLKpwQ1TUSs5cJRmByzpdkq
jym84egB7n5g1/UuHQVQNyFXhYCYSkQL4wcm6pSE1mHh5PeW8pQ1B9aLzHglJBAFgBvot6eBmtA6
NpRiFriTAiwPaHdmzyPhuux2Z5x0TVV24LesZ26fGGfH7Mp52OGmqsFPtUmgxuV4oFmFfWF9dIzY
3GaJVwnMldZXQyKPnGNJpW3vh91KEwbAyHlAHu7mfODImHrzHYAMRgsXkTtPjZUPUxH+gPoTqQ/L
eUiH4xXS+h46Zn75uABQo7434dzqYo2bdlr+tm/sIQYboYyBATG+uDrclZqYsXhd+QlMhC2WcTrI
WYrw8MWxgtg17xhPriiQKEJUlXA7rKMn9NWOY5bvX9YD82oApWougDx1yqtCiBcBEgF/zJM/W1aI
6s8gEA/XIOrVJGFa1vbrZhW6aF7LaBaWLle1K3m2qgdrpOW5LmVkKilgOWExNGzWYR821lUNpVIu
Gz9PAchwnC8naYUbzXIGD/GvHcLzeJrJorvOGctOxnScNZsABLsHC32rFLtwZzLOw4Oyc3Wqvf+k
6z6Ai7qpPhaYieO1sG2IfMo8G9NQUVs+EknoSSyFFSJiHOOydqnkEjuxpG2kcs04CpwtIKd4dxGg
JIuSiZBujBrfUG+ppTdoo6R+CPUTZqysY/JhoniJ803orMNDDgcLhrCc5LvMGug1CW5TboAOAemy
PbKLNcWjG+dItMU5yNjnzQWSH43TiW83RiydwWO7ofqSODNMr1mHdZ8N4tZwWUL866Q/W8MLZXFJ
h80QBSECRSbvbVmUvYV/Scpe6pGKjtvoIwgEW3u9cTRijfwqbKQefSOVR3JlgFj3uWHm//ko6lHI
91bN3rZJuTKMKpQpKAefyBFSrTH5ftfTu8s9YJVhRfAJ9T+o1s/Q4ItwhZQIeGLY17UQ+0FnWWQ1
sHQyhBuNZkkNLca4027nS/QKzkAiXLZIgI2RNOlMFAWtDMe2lRI+4WB1qw38H/flOHFAJ3hwbELd
FqWP0o+5KjfK9u68swtXhGZp5N9urh2jDCI4EBaGhCDsO6/WyL04IhVRR1IKmq/es0O1bd3uBLuP
bVhYb518J3DgkZAAIaINTcwm9IgHBFL96N2sjzQpkF+apkxpK0jS49+p1s4o1XTj+WXHf+1rE6TK
nC4deJUYoNTLExS7Jz4pWgdh53T3uzhT118UMiH4cSWy7yM0ViiL+Hn+DkTohFrXJogC6kAl13Pp
oJL24URChzeEa7rxNHBOoxiKLCFZsT0Fz6T2VhtXmN0By40rvmq5iL+UGJQiGUdtok5+t2f93L+b
E+uw2aor/O4/2o0MWKYHLXlf8ZfgTcub0Zeli1WZVECV3fYw6V+hJnDnytR0Yxc2q8/ckPvQNmp+
vfEuH5tTNnU90gM8fLbBtYcLCSFK2IPrL5LVe5TLemFSQKO0F+QW2RudcTkbQnYPGfzqi5Yz/7of
ypwvK8QRqrR6xV/8lq01jrqJAWNsWy6ZlX1GsrXAPE9zjy4bqlmoZuk2jjObuGfjqhkm8xLRYkJ1
U/ZneehCsHxertm5FazG/cVenzGud4RP48CBXUoWP98jcA3Xg9LcnIec+ALT/VrGmZQ9Zode6Wz8
hwVncHLyYaAD33PsQzVpdPhs3N3DLYmE3lIBNKu5gTPsuPa1/K/JCX0BP/DhYe4EFTXzH2Xj5pKj
0s86elMNVsUmeGdYBJpW9kq5y+YvRMFg1llvLuCyYp6K2mcU0aZWF7dWxjCWPExsc8H+9klUBO1u
AfEH4tx0oIIjnMdIGQzg1Nr2lb2Ih8fazsq2A6IFk8Mfrb6zYtCfPAafXBLXoY9dbVsWBaKgtPTs
GGf8dWXVjWlSzJB1LAVOPWhhZzWAW78rDU9xgO7FTQUvWWrZ4zVIvfJ9OA8m7YWRBlFmhi6vhhSX
3c6pExnzChpCBQzLSNDqQePlsKjHBgBMpEkVg7aHf5qZkj32GORA1qEKYlThNUznoBqinxwh5+aZ
YaJgF8ghjQB5qVsZCECUssiESQaZdIMqFlVPThAtdMa396BJSFM4fYriqnFTZhPA5qhcUsqW0Mi/
w58m0sxQanxkNj/rXyUaRqF3d2UeYfX57H+JGGbW5nDyDyr+o6qsqzSGfwykUdJLpAlXc4Y5as33
iW1rfcDzY1C5wM1vPAlv0ViAb6KINgwjXb43j/Af/7hN/P7SpwNsO1ue8c4vbYqfCDdHx4/gDx/D
pPLkMTRBMxn9keVsOIgPiWkt9E2pglyr2dkbq55h7V8M03rCYjU1iyndM4jQZtZk6YUiaOnBmwtX
j1k/xsap/in9VLBI9h0aI7JAnoFfiwu87wbrPPw/JYCPb6R2KNELdg45Jmep62ZQvAK7mS8Z+Awu
lcoUnsFs2Nb1xW+3fTjMJC/jdYdW+B/ASSfG5nzsioCgVeMD5+hYes3P5tt/nCbdqyFwF0q3Jx0U
Ej+EtkMd3MN2cTFK5rYxj1MxgBSHGQeukDm3sNYmyuN4Z2EK78WAYYlT9Ih48cHHalNOLZSRRmLI
iAbnJm+OA3BDvpzXPjTRRuJ2Pqk2BHi47ManLqifMlvjd67d2sJA4Q8/SVe1QESlvwMfHfkfk8uj
TEhh8zZGeEyBSwMJBxy5EJXV4MliFNaXy7NaQHYpfRIID23b/GFZxjnNNwcK6mRqn6+7J2PHXhtY
p26hqiEFOE6TWVUO6I6EV/EOHm+yv1BdZ37ac5z4vLUSPIfT4RUBO9Ul9xbTvH9imhlktlIVSjb2
5okY4v5EIO0xQcNxFsWx3wTnoNRwISBEcNHLl0LVM2rCZUhbT8GkarYp3GKecZxGN9RRLpwKbQ09
8Ek6PG7MXgFlPHTBFOq7dDPcUwQupdt509cylKiyfcyLefRScM1G+zgjuUFaZ5pEa8iISJRYIlSf
1S+eY1mVNYs3G1GrlcJxjFB3zJ2oaNdSP+TqUn5n/Dv4N8eoypYzUFv4OfYzfU0GnB0A3DJFz/w2
WcAd6+JhcAjA9GPfJhGlVZdVjDoj/KvaBqL/jtklkNNcFOChIg06TkCT6Z2tlCgsfzIIyi7JhMMa
orHJPiCBSvezCKQilKpJrFS3qlSz8l/0LngdR1SJ2WzyDmghZitPSwCOnOP8PxSbflRMS5MEaoO5
1ZFcNdEn3VNKQsYtpEdJ+PbBal9XTL5BrMhYuGHhJna456DNzftwDU4cyNYEtZ8KbURHcyXOysFM
i1t7tZjSthLgO9DIb7ut1h/GmsYvZS+BZEvli+liK2AEADE0jKBZxpvjjG98/L3ceoZNfvDxgBRS
l79sBHHT2njrc4FDxbnCDlbM5UIHg2NEuJNBi3YT0LYCh4DiAbn66AQYQ6Q0vbqZZ97jM3OcHO5w
oh9G7YEPYtfaVo7d80sKsDGnWhX0sj7WPloZHriWKMMaGCNQLJSaIjuebVJHc6iYDgodOCuvjvBN
0N9SVc62Yh6Kwf/+eVUDP1/5uR0X3t6VIBxEhxywu2BubJJcl2E1xLzto57wiMe+vy3uYfI54XLE
wAYt+76xWUBWQFkPoemm8AUa5LCraIoQzi56cLH3/ZBiq9cg83d4tS/V2Q4YVN2iDfAkDy1DPDG1
9NUlXcxdEHDk/5qiN2X6hrmti8IpuJqvaJiMjTTy2YHEglUWVrd09tppW+EbI7HAiGOiLXG9qcsk
m8ujPFCg/NtRQX6eobeVMAlb+B80/eFfPNmCYYMxHpqbRiXTssC6RlezybOlC9p4RBKkr5fuTGzx
ZD0JrRxS4CCpY7RthVgEtr2dwjWx2V1SaYq9ATQ/tGWqtqGD8Z6HbrtbFj6DM6ZRtXGiJ4JinWtJ
+mE90e5NNzoR5EUc/j046nhCPZfvttS0AsDrxCTFE/UvOqI+5Df+8zpVotMg12wkhdqBe4iRzOvb
DpwqKBRWcpi4x7YB7sW6GA0OL584IABfkn6ZlEQCVtG5iFsF3t8zkTrsVXafOaF64uFqm6Lllm0h
xnfgqsat8zxSu9Ko7KAIFCCMe5l0UiJMLScaRImBsydUVB5w6zERpifsSyWyGLGdhYRgzhDPayDg
FjNPaz/EORnKO6MXWpEKXOQ3ax2vcecFymFuXkKqvcISL2wE6DRMpO2OhvtQ+EXwGGdoop+vXe3p
BhbjwLqjekYoBHNiFRjNCd8jvBAKYENvceQ6CJ0oYaKW1eoAvoncri+u0pg0M9Wi36c8WjVJm0Q0
4YoaB5s0AHgHDmWcd7FAWEsT+NIDSzuPwaUMivYgt26qQctw1tQy6hg6giBxdGsR+IlLHIifwsEU
GE8oBM+29+8sGPPiEutt2dz67K65+bH6ClWqT9bGZsJjVQ2/CEQgotBbnVVsf8Cg5FlpKvfi6rjj
yGmjOl3eB7vsqDZYR/OYDB2Qy7jUCr1MXeaoicKqV1bhK2+D+Ahv16cP+nJptYbw7FSpcS5IH1Ks
uKg4aEaKgID3BLotPnIRqNJbTmva/6M+t1qZilueow11XqdqYUv0Da24Yr7D/EbVSrPOKaoGrZ+9
PN6Xga+cmRmRH4dS4l9SE5gk148ZJRz62v1SaX6S4G028XTxDeth5bzth1BC9/7VPLBFXMSP8Ih5
BNckf++yqDeTBVWQaSSANdhaHdCpNNYU6jestuZw9xFrFrBbkUlAGLxbbt7as4uIYlilkH+99pkx
24NgPlD5OLa/QZr+2pjdE46c+/13XuxWMKwJSfvJFC+iS9SNylWiVq96ppLqhRZJJB76dBNyZ+tj
Zi6spH/XGumNLdQI7ufnQuTWSRlC0SzXPT+NXDTQbjgj0uMMa5oOQdI4aJ9qMpXH8tzjzRVpn8YU
aMzJ1R1B141nUXqgeePVkpBFOiTammXdxim2zGjmpsxIPiLYvV3xi8E7EZIZGEXMEjxDkZoteszu
8z+lrh8XBMmbrCuLoCIMH7WD4jBJXeqZ9yxnoLnx58qKoxMBP96f0l1bhfZtDYuZuAUCOMzrjbXZ
txgf4T78ImgM6p4YfK6ZoXIXNFgyzAvBQUnaNClwvxse3weJN0/XeWwkhLq6t20/g0SODxfFzvFL
VCgA05qhI32uO/gDVsKDMippsdBul+t3PfWA8pyrOUTfsTJwNy+APYGR/BE1ual3OF/Dfd8H2GeR
9WDR3lxkYX0wwRoBFV3CDa6LtjHP5w+kWAlUxe+pgUBLXwq5DxBSJWOeizD2+o350ZN/RwoAMoKh
EeleqkVncRIV1d1/VKYV53CLVWWbke/jGf9l9hzu8t/n4+4d9888wSdeBmxgyPQcKkuDQQg6FPG9
3ENxVAou1BaoFHkML+rL34Gux7MTA+mj9QmDMhYjzamruNNcMj/JKYIOskM43QFQHVuiPpxc9QcP
/zHucb5aRGe9hERos54UC6ro0PJBD3KYS8SYcyYG0x2NqFwks9Ho/h0CxGpGs6YOwSYHLat4OKoK
NqrwniK1iDimTIXyIy4roBBbj1su98g1a0FmgEGX34beGiYLTxmiccZ/jEuwPci6xs4yKoY50VOM
I7fz7jWuLYog/0+zcJnc9sFHAu/qM9Xj7Gp+joF0xAWog6upEHSGVofinbki1mpXQZRkR5VSM6Hs
6Lb1w9da02ngecptaVK8XxX0VmL6KLrfSoNj4Su3t5yQ8X5B4CLFL/93k5G011QhGAf7dOqFtENK
mIrpWE6kOykX9NIEgk+DcOMTJNS6LuiacCpQA/HHto5vMFA8NO1+zZg1Hozs053IwgDqhRSbiEzJ
UzeJbRrAdpQFQ6HC5XF+sNW0AcYbW6rfkaADBw5Ur2UXjjHzteLjfNWrUmZJlutSF6ASJ/8Aqnya
5PMLm/IiGByr485Qu1wsS4LUWfa8QISw8U59/tNJP+teTN3W/SIAhKFRDODS2SuxlyqbMOlaZx03
65HvrOJziSKyGMLAvaMHOa0j1CpGWABIQ0znNrSAsTaoqlZcR5pdzrK9GAkmSiNbzQ5v2eMLbBYC
6rc82JrVv9PFh5Fzp6v4S9gsJEXt/NW2r4UcMSoNKHWe5ZVVPrGWTfdp0uXNhiZPG6fK/kBohDzA
KSBsI/9HJM514lFVL6+ZMe+ymVFqhhvCd8xiYnrUsOaJsVGVvKEdz5wOMPstGraa6KIFfs2FAVEO
Aqi+O1P2zZ7eLouzFBw0hEru3L7dSM8lqIlvfSDfz2WK5DXz0bJPb65WjqT4Bzq3BUvPmelDQvTd
iCmkoafw49ZSyiBQeGq3EQb+29kWK1sYV5lkqCgtFF6aAej979aOmYWqj3ptNKcRACYaBxd9PUnu
VhwhxcjnFv8AI2c5Dgy1vQfSeEpxJCvInKIJKricu6mr0JbVhFEWNY6bCvjOzKz84M8Qdv+ICWPA
8Re10bfk2uO/P802B8qt//DtNBvpdP6gEZGAnuT7YpMTbszzmKPr9qkI6D9OpfbPXNXqpzTwM2FG
UaQxkwYV5TysooHrVuNjLaAHr0faprgsWLfQehllFLpaofVXErdZr7jpFd4lwbTZt06MkMCwgzdm
dD7TcTruEik+HwQwDmBxigmk3xqPHsVcvUXDhMhcrpqZSKPb1aNHmZkTC0J8BV/T3KEsiYcFVYQ7
Ge/fM1CbRTV6OSrZ3PPsMMnzGUuBpua9Jh+pPaHeSy7z+0ZoKjJm+FIomroAFx6IVEKg5HsRicN3
lXDzoYgdLSNYct7JAiTFJ2AVsQCojTLbAJEFBGyD9U+DdDvdB+pb3iWIB6nSUcboGHAdkwv0mJtD
1rfdfgRfGw52rPHC8zLeCD36bhz8cOOgCL2KYWdQQ9Zc9Fxp86z/AY8/3lpsiGjkUaK011KtTT0R
Lkv+XgJjE3nxTIFXl/+vyp6/pBO/fi/G9s/suezVKtlLCBqQSVTbc52etAbRPBzFFy9oQ3SdbQE/
pDsup/cNEKyvPMn0V6CRxkU6wCgIvUMwcXKj7hGTmDLAxrL3BA0kyQbbugyaLJI3csrdqsj95S10
ew+fJP9NRLLYHg9T05egT6zInWcyz2Gets6TjKvywg6mwY7r1eDnRc24XxLCj4/UCpyJEeJ5IKpI
mOhTpKEfoDbo6xg30lPJ86h4tiWZz+8dR/eRybo3scYiF1m7e+NncriS+cnT3lrEw8iSDoC7H/eK
zWGVya5XQN+fkyaurvMWSHjRE28T2UTVL5LoV+jAs9CVrHQ/eirpkycMATwtrFJb+zECrusuESZ6
+bvwC9gSshQQK0kbI42CKX1PRS9NErtmvsYaTrK6PRFi1ohVbm2Tp7F69zkMk9r2/XyBvmW033xY
D82qjbLHwt5mLB6EyJX+2pt3Xveq+vQL+lTCmidShi7+zxVU91tpn9eWpFNzoG1C7XQ4mXsbC9eQ
+jEUj+DBdVVE+0IXc1up6e+hgKkBlGp91A87X+Lklpy97qoAZZdz2TCwcK5PKv4yepDFoTNwIj6k
nKrSApts6CYUBS8drfAwD+4EARy8x5R8zFyZsOtXOoAzU2/cYO1LZYf9qeiPuDbuEc/a1ck0a3YG
UZ6nTYXZVlybl9scjZf7fjNurc1QL2FLJQpUGxW8nL/ktDiXw3NyUNYB2qjtWHlYYT++Ma9AL8ui
nEdMl6/Kxvm4pkbaYS2XNiTPInpku06LrSYYK0u6mMkj00wFqM16gr+8BJpUvggp22hafEgyQh26
SZ2O3oXDQze7MkJhMTVyLByV5rHB4U1yCtXO0fn6tNiQfDMJTnomrQwVrSlrY/B/KKhlPhmofSfz
CrvIWLvU037brw8ozdf5R5vZaPVL5/F2A5yiUbUfbgwKZn615bWV0Ux3giaaT1VssERt3T632zrk
ftz06FuY2i7JWEawrRKTDCzbPUc6CUMVSrOiJoR1JIMBxQ5VpiVfCz6+Gkn6JM8PmIFwHRKm8Jc+
HeTII0O9BB5fV96Fsfa/Z9xJVkCmdsc2Bc0pbXd4uOlwrI5ZgGhx3H6KZiNkbPJMxLK3QShRYzv3
z7snAMJQpYCoGenjfz9MAO7XMxwYNh9An5FTNboP735sCxPePI9HRnE3BUSGHJzR9FkueTkARVVG
6sirsAk7OD3dXYwNowfH3bNRQYgszb0euKaJtx7HHjewJ9ftewwxJTDf6iu7PfBo29AafQYCjz7d
52jJiiTjy/FNH/8ZoH6KkHKMOaXtnVTNurLRBXaafHpiD5cP2iekRMtfqPSCmNQ3m9AuCCdEorys
uryWzR9Emk7mLEvQjiUXjdNMCnw/z6XVChtoIrUtipAAPw11Q1/xHqLODLYyYMXqfNT4fJLKP1Tc
40ExeroFeqqnzWyA8DbVTm2Q7+KmlAwZDr/TvUCUGJw1uY09aEzw5MFiL38h92F5+cvpID/aQrcR
7vRoyYO0WdxiZ/W2NnDGJWfxv6HJ8tqbW0KBZb/Oz/Cc7tbjGwkg09S95pws42h8/najY9EzwZ/D
jbqDCUm4BTj9+dE8krKd2bo4usYMmdfQASsSNW5XjLIN6LQ4ycDyyRsNsYS/y7v0Jlm7NuqKK1Dx
HI2e4SAezI7X4rvuvU4smvVUKKumWCG2q2F+PcQ4/e4BS2xH/cMIVIqZp/SHMHuG3oNKNw/do4o0
txiaMNM4vXpFlpSd5x80CgiPs/ucfj3Z6kx/R7Fn4HcTFOU77a2R4t2uRC4a28xjc7i1qXNkV93x
ZVwlVP/Mq0xiDQ/J8dvOujzJ1smS0rWHNVDBDAHeGB2BR08PW5MxFhnuIpUPzEC87GN6brwu+GaD
/gTH9B4iyam2DrXtBy8V8gq9traksSx91p+koyyL7+DiDuDGwiAFXVECXPBoxB64z9P4Dj+P4Xbg
hZsHYAIQ+doZBT5V3x9VH29unSY2YGhlwMHipR+3dHvx3GYjyb6/M/OWm0roR4S8fm+y2Ms0qxKB
UIKFd5Tk8YzRBvB/6sgZd5sgfsBaGOulH1QH+ZqLLHtGj2vlCStRRXU9xaX3ohr0DM7fLfx+UaZ3
3moEbb2VT98mqRWEtInxmx9mAKz1gtn/zAeHKGta0kUp1vCM1TDNy7oXefEPDGoFOTIn31FYunBj
dkcr9DEhxqAiPFn6zf0uUTcNXw9DP7G/TE9pqN3HWklOFnlxo/v0SBU0x/t2uM1o0Phws53F+6rn
lVI40mIHHJkrc9vLxE3ZfYjAvwkcCFnq69CpPKIklJ7Wy+ky6Ji+vBAmRWypR65ZpjvIakVw6Gg2
hfzX2ftNFdA4DUViB8c//igj7FZ/T00rcXY+85BcYyBi1tIUj3daQFW1Yi5S8JZlVL3sB1XOEYCJ
fWQeKf67UYPv+kQFgwZZT/7CfaZqoszOZvF5ctTh5E+ZoqYDHXcTV7uge3A+qnce+fpM/5hqoEuw
LUj4Sa3SApKmAdimllQIG8dnpKW9eD43PU2kvHc/6gYYZI9Mf4/iG849s/KkbjPOSIS8bIAeC8Re
Tzku4mPjfXEH5Yl8QkYXUUoqrFStedW89Y7yThQ1zVxXmIHGNgqUmUgPi2kiOptbGXWdiXnd8n8F
jRkmHwrBpwwcDpJydUZVCF1TRf5d6qH4ReS4VuC9Cb7iru1dbxlGeWy8U6Pm7Hw7QKolnsbqMn0w
lF4LPM31Y//+05nerRZ+QJ2F8X/QXMvY3UISWTNLW52X+oz9nISpIuT33xMUqeTnfdP06wFyOSWR
yEpGGlefi6k0GfyMKkGqqDXzYjW58xaSLickuahe6UNY2lB1v8TAGwaC4m+pbAdmstdMtnxDYHuZ
TPUZExoRfGbxnN6ZgMmko4iRfi1UByW+IbrrttSLo5XvqeDFZcjd+Mi9nPtkS8T9u/LZT9co9g/s
p9gmIk924GhaeVx9xbDDpCuG4sWFSAqGdGUAfgleRhR4rI6DLyExUImtuz+1olBxcA41yZ6LzggB
26ZrufhbaoqDy+vaQgwgU2Mnuk52Wr5Meqc/Fi/T5f++E4JY2mUSujpekb5EYN3j+7oN3mFNHEEU
7T6VWRz3VjkPqzyR0SL1rp5gP8nsd9LMiCBuxmMtADUKImLe1tNh+rOy6Wl/ab6UrhRSlEHQ5Uke
ioomAJGwbO5CQd7cihxmMaJ5GYHzdoRBwjQg2fE7c9sK9svOlnflLQP2rXHtPReGB7Zfn5WoTYqI
KvxVVKnJxScEmDAQrkauTg13NLu5zdr5mef7dzCT6PavqI+MPGlNirGL/VDWuVa4UZAf+ZH+hDSl
gfJHaBrT2VtrdF6s3MZ2qvV+LBzO6Nc+rcz/NyX/PCFPt1pMiv+wZwwEoluYSAyzJyV2NQixQba0
UX7PeE8ed/rUKK5OOafR+9+oD530ISWXXepqhm90OOOB1tjmIWzojun2gEfxsrxuI5QpoRnrFeqg
qBi6VPafTXyxS6z+e/UgVQsvYuRxfsla4dDgcW4LksJdXbbqhHRu4l127Y4mAmDQVMKiEtMD/K+I
GOyqfV4TbYg4UZfvQ9+6gKqsiMYCqqvtS88QV3pxCXFyaXddyGOD2EVfd104RFDsmLVQFjM/PMof
+p/JSMgxJcwOHX4y6gRIZQBKXY4sw9pMXJ4xEXSMm8mKd/ovyXYZm2V/JIpdDGQwD4Gnc8+AWDv1
NpZKwj12BsM2+JKVlv3X56RyAWrMCf21bYfjHe4llqLyjCNT9VXhYZe2DbWcV+8MpTByG0GqgO/q
IytYyjo7gFr7QMmfcIkTWBUJ9ussRGu2xy7tjGFS6F6/T1i5+NlgBiewxMhioCv+LjfOEQ6Z3nPr
paiht2sRC00igz7EMh3BVCzUMlJMyJ36l3XbqfoVK/27E8Bbe7yB9bgpyHO2mpkdeoe8ioY9R5OQ
wxNFbEEvS8RINXOygE4/3j2gL6bG5Xo14QOO5psM2WIeSYlYbG6qXijA+W072iiUxsG51u0ENhyE
UpuLsFsTV97uIBHrarQnr6UFSsIdN3LJkcJq0OLTTLOOGlbviY5GD36C9pA5Nc9Uhs4YTMIdeIjY
yALj8u3sRvqerfE0ggJqZXCEbh4TB5/DauAqU/kKYdAJygS1v5ToAjXquY2VfqWdJgcK1eNJTnvK
/hCB56ir+wMVpfXOMnhyg3eSn17TQHH11OIrI3LVv3eWXewQmppFVv7KtLd2aJLbhh4pdLvhSWzs
CZUbDXYwjvOccdmkn+4LJGEX+nnlPqGuzd8R4Jd5PQ0F9oMH47GQQGFHEOBkHl/zoliGPp50dKP+
ve76H8uoHG3G/d3mLrZNOV8lP9xV5nQ6vIM0y9bAucSOUCFD1nN3OwwZusw7mzQ35S3EosnNHP+x
GcGdUjyx2n0eXcLGd5gijc2/5gZj/M+MHHuePsEs4TXiaeYx/QKSB5xdbMDWDXP0scTBFBfpk4Xx
EHWRrV+AuXDBPpVsJOHwPqOtTqOFiwqV76K9Cx+1Dn9VhPBmWdFfmszYR73/GZ9iNC9otl5mYpBk
dXvHRYIPcO2snmgWWzHF1G98Q/Qbg8bKoZn7n5Z1AW+ndmjl3bjyHDBYhnLsGEOEZGXRgc8+539g
YdBB++2fkogTaB2E7UGLO77pZgjzW1ngjCnQV0pcznHdLVThP+xUL5QfjwzUxE/yvGsJVNefJ1Zp
1TcvQx1no8DB/h3/8R68jHI4xgeKpwHW4Sor84T/vKpEYpjwLmPY72R9J4YMFMHFJ15ILMg2fybe
kHzLPHIK4j+ZulnEZdqNGjP/XWH9kgqfuPPQTcgnCcHMXSMvLhk+F1Q+A18mKBx55H+0RKacKQFs
yKIeBloLRR423IhEQbV1MjFR8CbV8LifY2oMbYfJBujKxMy+4iF5IZ7yCFhmF4/Mb8VKchl3TfmI
lcxfQXfSU6fh++U106ST3xyZnqfR7X4Wy6xJuFbe0vqmlNxerx9nAqAjIOGkXjFux4azz5FKjyzt
IqU2RGvqpsfL6beklaQiAqRGAbHPq7oUSrzr60QcZSH8qFY/iuQYzrThj4odbGppEqGhcp/ueFFG
kL39RJTwimnigSlfEKzuMkgtWW70jk6FlZ6gEjuQhueuYyjKxrWkZBSJDdQYDl1jJVXNr/p5v8Z4
Hxzu8+yzywhqqbds7sB8gaCEjSwgLtBAJ6q2jUU0MOjZEBorOqC12UVU99GKNurw8y8RxEdrHDHL
X7CPLgxGDdh2JkMGHYhgNCfUaFc+rdQjBacfdjPWzEOeb11x2CB8FPOToxJ2xqmc0P3VySveWXVb
pk4XJQ6dwO6kRIQeQwduFBmx78XoUAfY+LsdftrD9fI+HnAwGNqpi5hFtK9FuPlXGG/S2qUduZUa
BJM+aHuiuRCSDhKuUDcs5nbcvw1eDDtwNpkdFgMkMuZKkqZx+cyhBn38+GcLcADRmtqanNXugzET
e5Orl5wO6EXME7lauRLMAu+ZO9Nu9UOQhTdA9868XWd2ofEhNDfXi/XL/dCSJuwyJi/8ZxabBcA0
ocvoYCDE1qMND8I76hLv+NaJ87oMYPxAKM173hhDOq6ehjibm3s/Ujvya7ycPUI+VCIOfwoQ6ODE
zcj4qEaX4kIwPt6LZTbKcGabwmDtZM227a3SyHmZyxC4Urc/XeFEs7I6iYxXQgYn06EQqa1HIx8Q
vvcyM9OS2mec4P/IQzXINNxb3QShkNSq6CPWm9jbuNrLzlOJCeW2QLuoIJx7OQ15Qz23tf8ETtw5
Bpf+9ENkYu0nHrlZ1i4GMBDV0ZjZ9tNweV97WXl6tpQrykgC687ExnGoMIb/XYHaDLAKtMD1xKY8
0hhjm4ANtAXPz5zNi+kbO0xS0b/OaQ5F73aQzPdTCVT8JpYBPXqpyaPIo8yXCcjE5Mxbb/DepWXa
qGTqhx06QdBwVruzdRI+vLtKeujwdlkpeOM0AKHyMoh8LqL4q7w0ljMQaVQ8+jJE763mnjxckmT8
HrS2/WpLgsuoHNjPeFuKNDKrehUuunGph/GeXAvhA2RvPoOFlgeXWHSKMnq4BgUiWIfvuUEjM+Z7
qnpM7eCArOPwCjcwLnyEMGFYZBeX4fGXRjQAuei9N2nKjmnN0xrLDNmJq6pFDiQxez7/OA7DEq63
ojv5Fx/4ZsyrehzvRudb4FHTEcrwm7yhgpS7/Mntd/iGfB+jhLMVIj17Dte9kUz69eL6OqDLEO1B
UDDK9U0yUEagac+3RkWp88nQjHhscemj/m7lODb9EQ0tLRz5bLo8qNgcc2HNH2SKImqhNdIA/QnJ
Qbg5GMdHb5J9gEk+kh4aVllRZYjWemV8w/G2MrvEyShKFPS4vqnuia7yAMd+2McffIXQpzwzOUIg
+TT8T8/siMfL9FyoJTDQrfEMe3ioS96NHgRKrYiVRTTryb9VUTb9zsPUJEhj2KlpboBIOISCCymk
lmAkqV2KCV5QWlQn4UGDPzwkrhAAni+WmdVf968i0qXjZ53pWnIQS0LY45dNtFgEG/dTME6154cs
04Zs0pP/TX7INQqRM6qDgDFb9tSnNU6GInWou+mSkbeKEyQkj7VFoh/w8Qe4S2w3ppYTXaf/wPtw
4/J++mzmOyov6J38CGnOChAVATfDtqVM2b+NFII8WcKAMOlGmKuY/iIkiJoGNCYcgS5OtdCn1Idz
lw+dx5exJRhQ8nt3FVeTp8Ep276UtrSd5YF/18H+dq0OqCTqDnntkpMb7YfHYcN9K4Qh9rgAhaqp
JpRiVUJS2VzSLk6f4mopEufDrnCP92ie9TCCrjOpR0G9dkZgKNeDvfBrWPemF8jWSDxWzRbTl3J1
7uB7q1CfDwdrp27LpG1jT6XZFfpRM0zYhkbmrexmwF0Tv5HBY6fBHpirzqfXAe991G3oqf3+mKjX
Lh+ADN2b419No6pvpr9pBI8NMnPeoL4YHkq6Uw6DWxDCq9EggWl1NGQQsrL+8vroMB+DwGHsxdn9
3TSd9qkv3Z5EYAfQzE4V694QA6A6lQGU5w9HPFzgigUK+3JtlvlOkPfyrnCHRz8L4fNrHK/gPW+l
HEVOgg8UBycg+18IpIxWHBxR6yyadb8yNDzGhv/xEqe9zP7NODeILJBfLmysFKL99zJEiVCcMIBo
vZdhY7RW4509dchgU3xkPGiVbNZOdmswT6xNOVlGEW4ke/zNgyiVGuWBR3xZm645Ko8soxTK0qQR
P2aVeAoXHLY8rnbaQ3dad3HRIVAudab4uGB4psquXio7Mn0HViuyN0dmtm/J0axikmqfd3bD84IJ
bPFjiohobRMdOjkldYKPb08IGBbds/SaZx2CeeVN6Yv+XMovsEZAa93uqIj5ybKZ44IfR2mFLFSQ
MgjQ0ieTNCO7pao6lxmrryzTQijSlpdgjM3CAnEfTJhcvvRVGet2LIv5GzXepzuASgWG94glDvM5
D3VJDbe2WIKXjzgkt11DiX2gekqXRvV1W8NCifH+Rh2VYFizANrBMfVAN47aqF2VSPmgTp/oqbOn
wu1nBsmiM6xGBTmsha8uddqhQVps+GqzWcnI0kiWQQx5Puz1l844IligxhCcuO0dmmUX6RhD93A3
H68vUxbBxpMDizsr3XCRzLQa3knneR/9UwiHQR35TrpsLLcx0mvIsVh2UPFFQqGHua1khIGq0bUq
M/wfE62GS7vU4907jl0qj7hkQOm4rwRZRz1tNMGlletv4NRu8m9TGkAOXHi8WLNCaMxvo8ZFCEjC
IcLt5U6iT9P8tiwL8wTzgLh6vr1Za38Uyf+xIjctz4qZIYj63DqloyiCpNRaSGKJmskJyB8lYEqu
HISuppIAa5LwwPpK6HI/M9BkeyI5L3WEt9eUbWl6SLm5N1g0ccC/gXR2KGTZ1dWm/vX/h7SC6NHS
ND1ebiCcrkPY1FJPyGYSf6/xuVOL9hh/Yk8HTcZG1xSvpIR19VPlO0tmajNOoF5vsrIkwGANoFlC
IyxlgAdVHT4JenxnFDG1fT9STRh1Cu0xL14zLVNDi10NWALa3xAZPm6IAIbx0oeFdzTP/sZc0Kpd
r5iiF/Jt/PKZVUsUXfBpsIuBcz2NXznZtIClPydPKJJxA09JX5TDJuilrW+zGnfsH7fSwhnVkfhB
ZU53pYw70wFBhLJv1eJmNaiYzhEoVJd8p8tr8Qod01rHF2f+jyCwm06VbIOE2h1riJakepWGQ9rn
OBziy5WU9pYGo/X3mNu0x3BZOL3cEPaU5Wo48lEurdV0EaKWRbHJ+YeVFpUcqBN3PYX9L/Nl0c73
oeB3o4lmcrQyvlLSy/WF10zR1ti+RPQ/xL3QSdZc1zcNXEd0tahwpw7rP8hKGwmSqbZ1dvYJBD6Z
QbEb3wEn8hZnt0uyEcqM7OFANJqHpg79Ac1f3YPHm1V7dLA2kSLyPWuqE1t1p4u84tUu8LW1Jgp7
65Lew+ECmLCHHreRNohd2Ize6E06p2x9zStkRKrXM9Wn6yGjgC8A8KTTF/VCwyNS0pSjy5/xB8D9
pKVENJhwymhhW3kVapjhapTBYQMz3aKfbEGeyBd7oU+lCR0WZibdO3LRdrNHiUtHwoLXEeimGvBM
L7H74Sj5Hv+kKNpN44JgR2KCm1ZA9qC+raIqJSvOokVS24JEYrnXIR2MMiVTzmdEsu68Kd6evHrs
2lH6fAk9RfI+/w7KSVQqReOPXXt5mtUoYyTZXmNRY7hjNCkZm8NhECjizz1dUxSFInJcCiOkW9T2
poU29Mu4KhOSJEIVypiqnnZf1CdpUEUMfTBZTw1eMVCeyxvhlve+c2R896lKZjNdplVvmLjbAJx9
00ChfLakupqyV9QMXnAr3bvclTD5fKzVp1EeGagefOUmeygBiGaKYMFT3XW7fR8oui0w7lFpFQ/7
PxGfBkrrzuD0Vfwbvb2O+a7yiXJDW/2qRU4o/Hjz6DCqZ5C64/UOUWAsOleoKylmkg7mBdyKp0kx
LKzuhAP2vDg8jJbpnLIuLv5zFKeL0c/KnDHxOvWI6+++o4khMol2kto2fSdCmRfJ/E6tAdYD9ZA1
69b1QHbPOsXgJp2x/hKTkX/7EZHQ8TeFTW21dgNYwF3rxqdxG5RsNzhRii8ZRye+8pIhq8uNfk56
+RWBZoCapns5ddf2loNSK0kixqGiwRzdxWAGezDEyaI5SyHlgnzmeFHHB18G5cWj09DDVIO2ywni
X9trthZnu/drYnbbo+69V5db/u7GX4Kei7MbhvRR0BrpyY82beVVh4Bh+7cwj9q95DUeWgKtodus
jX3ogbEizkKl1YqLBjrPKtdKaVgzlTxDDZNjNNLePcYSEEvi5hbsCKLmBkcNKJ9Y3bXVKR8K7w/B
8TWK5W5lfR9p0gcU7Rg/4T0bXLQVbIOtmJXDSpEBCmKrNjCADuskQ/iudwEU7qbUmwird9xQOPz4
IHIvUiLUMO3hbs4KeAE0m0n1M/jR+McpDTPMPXKe5vlQ4WmcINgYPFV475FdwppBW4TKygps1erW
hGIJJHiclAlP4mD7bCmBH6Ip/LFr5EfuDqMi0EHF4yjr3kRz6/RDUUKBxwC46XVgAAhl+MOAI718
BkQluNl9mb91zPLg+F44IHTvCbTpvrqcbuZqCqNotEaDSI1RcqHlN8pQeyct4l6PSEUIdsSR4dYR
V6FvqEYhXiz7UMHsXjjBMpu6hh36YaTLEYvMcm65L9BIYy7+FfSbKmeJgVdacDLQvuko7gPbtqTF
wCExHzPDAOvaRlHxX385vi84UVPR4z0WAG+mRmaxMctcqPlXp6qtd7qV4Rsz+TfWwvNM7pTJzjJG
AGgNoSLACLns1Y6Tre15b8Q0BCoePeclJ2ZP368hMxdrV79ioTYMqDZz+p41QrQ+B2dgj9boBf2c
QpxwZzZftx6l0itTjwTegKBNhM2t3Hg6r0zeYmA3WR+je4KanpD9SGl1enYD51witH7/BtQ3nTCg
x4fvwLWFAbYwf64jBXBmvHnsF8p78pVN4pkc/T3aAwSrlftZWywmxP2gcfSBbSUI+C60zJAcodWo
xQ/ptXmJ9f6jsl83NZ3nbbpYZA6lzXb5mP7bG/t1IGuMvWn0tSUvuc96Q5Y7SPXTJD3cW0oPHJB7
v+tJGmZYOUrtEQyF7TZ+r9XgLqY01Px7yL770pLScQMXlijv4W3HpV087jLPOQFEbzqlslWWo+m3
HrnyPQVr9D6CiQB8+KVu45uQntQwMZBNKCdTMlI6Q/g70abElZBd5Uo9qlAeKaLj1i3rHEdTq9Jo
XiySvxAQiRe+TDcihiymZVebIYVs1oShMaMps/MccRqgJn0bBcGxT6XsEyU4DAKKqRzidvIWxKTt
wz1CButnkW1rUaBb7obmfv4TTMF8f7r+saZOr4qMoNHDakgJgQ78Pg9PBxsXic1l5+h1Odm275Ms
HOvxuj/woxLbMZKWmO6eHo+8FCR+vqoDYfNhD0IUe8NjUXCdg9UPQRghn8T6l2M0ow2P77xNR/bo
JZ9KjHvjHlR3nrisVAtkoeKGszVD1HDq4RBm/wN8mx8XkjavAsqhEEVSdLDvzhuLZJh1pqpv3/Do
SWET+jEc3MZuRii2neoZY/nzB5pUHVdd9CIwJFXOVCACJ3Hj+pJEQ82m/Z+C34MBypIgkefFvPgr
ew+dHGaTYvUGg6I5qPXWFtvewR+MJ6EQdH3Y0Z1ncaEcG18sgXvYrCgSAjzO6BXskl16VQ03JEin
lGz6TzG3UZMcYcUlQl1ocCWPAZdIfyNdmFwla3cKliZO8m6Ke9sK/wopZEcZpc+nxYeGgMwZbXQx
Vfw207r0lEU3KuOOf56hSlveaE3knbgcg6hkdpGuIb0qMxHtHeNtF4vF/2SN09IZhHPsGoXIPOHe
Q4wIUnxNyB1MuirgRxuYrAsOB1CmdTPDaX6+daYvwzE6VN8c+v7qwAcs0jsHNRUDavkI1WaNTrbE
//Ejcuj+1jU1Op+JDXrZG/046h+T16tDuFJI98bxnN0RFzj6cAjxUnCOD5k0pv8/RzpQ2MPrn/LK
DWwdtChxi5I9vGVoXUBHNJB5lkDISyoT8Y6OnUQtgVxpOCB6d8+tY7+nUULhqt2nUdYXSHyCGDWI
UnTQigJtISjEc0Bg80JZabnmD6yyjvhZko+mG1Z0ZpU5tcUH6YoaSi96pl/JzxjjACwI6ViiUHDF
1NI2wzRah242P/SmvmFTaOTbQOPncEms20sAybFRo9F0MxGJvQDXyIoFjHTz0GYiKrpbHAZhujtI
3cyxogAI4BdgICxRjdy5K9SqB+eD8hXWrAhk2R0nhHs/c5Btbruw2XFNTJ6vyU65rOIrWftjP8Oh
W8Ey6vh1qD7tDzG3cRM8KA48l0T6c42l6RQoGM6xcMMk81eP/Zv68mYuhlpMht+Fe4ydSiqQLAyi
qBXJHKoXiwP0iKL4Ip2TsBZFdXyawmlOu6WXJBpfRmqpI5QMn1i4zgxrYCgJs+8cqy0NxDYreYf1
zDu8+JkdVCNdW2/8tNPTMCO81ff1WKInBAtVVYcbUmsKC1Z9kQ+Dcn+vwFvHxz/+FZAKB47C7kY5
OrZnk8tetrITvVu1EYUbS6ZQBzFDC/VQWkFoTpEjJdEICS2iwlLloy2xvMWnbZMk8EouuOleUvqZ
IgJa0jUkX/tV501Gu/Sw4UrZzYQbF4HbhCfoqMlYbFpKQ2QL6wHynd++V+G6F2Zrek+qmtPt+WtE
r/PcTwuI2e8AtYUOL9Oh2RHfa4KhfG7eB2p1h53jiLBolGo7uHMi7ibPiZSKkEcRBjsTXaog+1FN
s1ZLal2FZV1GOyB1uxbELXOPYFeQc5Iy3ErBeKxIZlAqfes9QQcuZ/I7jBuriDvkBnNNN0zfv0yW
P8CD7CO1C4sKCac+y3se+l6a5NetnZU7keDGzueXL8ULmBSKVi2Cdrs1r/r4jpDCWEVu82n1oNLu
hrVzYwB3zyeMqd/yb+5107hGUAiHgq62igMqCVlUnFv6vpFDOQF/t3aLq/qKIgWJ6nvFFYup/c9y
BYTvKLsoLupDY+9cu9A4sRj2w2WwfQ4cuArNq9qIDztwS+g/H1LYG+O77sA89yPU9Maj/SBBs71Z
klYe2TzRIVbI37P4MUh1r1hUzeXJaOb+2fD2Pwtt29w34KmY9DOQU3wYkZHlCbpNsK3D4x5cGeV2
rQ2FJOPGirGBctSqd/W6DRkRWw/7VQHkMIMI4DPuzGepqBVn1hA1YEWanD9/p7KJBgHAa86DI8pO
2GdmSLRhAPYdhaLOSdgZMWZiMp/fWi4S0ABI+UjDahUrJoPFxV57ATRa1EmuwfROv6wT9rc1jbmr
NAzWo0iU0lptsdUmq4umS+gHUwEKCiYYkeKCqP6TPhiTxKWL2AFX4wlQ6IrOWRkydSR4knBO78p8
JleSKDx3RKOo+rUkgY5/1yuxJ/+Ra4FpqvHS5GwNrE6liGmGbYbtLMlC+S23WCN1H49cOnTdykH0
4BVNiO5rCPa7loFSQ7QO4r7PVq6xSwlpv2pcZB1X6RTwXytnlTXuF+efTm8E9H0AEGx7L1/qc72J
ka57tecNjFkjjEk/Uq2YLjYPlG2SA6zxBqD0X1suYWfA9PCMh5u9wxJZuFZPPVM1Zh0RkQEhYu4m
0V2oHY8OI2Nk5HAQtk0CYDAo7okXb8U/Vc5Fq4JhGAWlF/aqjlm5Rp8jYdKSJ1CBLI1NNw6qzebw
f9OwzMK/2eC8ArkS04Xq9GXwkyZPT7DSHhlgMwdw344csOmRnxTYxBp8TOGTTn6KW9pvfOnfT2vL
4wo8Up2WT4fL8MyOUWMhKl8X7v3sUTrra43oRzgMyGEe1GdUlkj/yJVa7IT5PfBsU1UFpxonmXYR
Agxh1wKkNkuzx4Z2Fmwk819cHNRUEQU3QSr20tl49qIeckWtmJN9yZAbfuKBUSqKa7m6kOKJy6yw
NaFYBJv0KWFhs8PPx328BoOQgXROZmNT+5u9UBWadix5NQPyf8oXC1Ipi0/st4wWg3vEtnZ0cW3t
JLi+q2rTIROUH0sUuMjXO3ZULdeiyk01pC8q6PQSzaE/LWBp4qVNCjpUGqeC2e83D5ZtP9rV16JK
Plk3nDUZu4yK06/2Yge/HylFajFTIvk6FTUiu7y+7KqbBsTdNV/twMeRg4fGdmH3du9CqJ9oZBiL
3B0ibpch3V97B77lauS/vINtqEPEtF7Div/oTLMb+W9LSMiQqhkgi9imCkVjrRmcD7gIpj3TgxJM
1PmIn/FDhtWcw22aZuyKqILlGUYP+iL87kyIK6vJWlZWfW7PoiJpgUH+Ez5fLiVWieengCtglHi0
EYTGMMsh/t1/pycVHR39Wlncs16YgelqCmoSts5yIJEOSQzB5e1iuva38X9FGMyFaM8YA2ksuL12
fVWn+M+FA662iW1fwHh3SfYwhFH62PrYgPofM5w0kTaCBxYktFK4hft47+PhIQkIB1XBHS4zipc6
s6vFF4FGhgwjJ81gJmqsCaIWkmgu5pro9p4XWuxBatYKWEBMFpy52R//WQipFoRzB04PbCdBseUU
f1fJ+NOvbquBnjhf7BXamknceddzcgN30xvUdl/My2HZp5KY6AVVq5wJSUeZMw99KX6BtCT5ukYT
/3HNs2d3wiHl0Lxopr7WuE+wm0gdIbiAkr9qLOz5wsKJCuMs2PfHMaz2Z5qDVta0019ojc+MSR4F
IPPRC9WZR69oO+nPrxsSGqHeGv5wpZd74bErv8z8sUGyb66MKvQ8V1Dot4lWw1x80tmxrrz2DbyU
6R0F/JTcbBld8s68qCzGBTvTtqfdG5VWjrYDDL47+RqQNEjmojzxsYRWkWWf3SiOYxQXZ6lG3Roz
Qbl+bKN3dLRya+0YspQAimU+plP0b1EYIWo/KdeNk9oA+yCq/J5grR21HNNMTMFke8pVMkJ3m0TA
IQhHUWuqQYESEJoFj1pjizQYvRpsSlPQ7Y7EBlql4k/AqOW35oUjoJ3UhvCzVlB5OcZkFEJnevGw
XsXtxBcA4Y6bOuViyFFCkoqWsde62YzAet47W8YcrCGhiw4jJfcACF4/un4Qd1Qr7UnTUvimDMfn
GMyQHwfPTi177Rb/6Gdnc9R27FekfwZpy0dmwj7m3ET1Vxzb9LaFjX8pBUY2KKLJrLVz75hWKFxo
aAjnX4yiVbYSxdkeynwqaP2YK1mMY2iu7IuY8EHlUqhDwDBESoy9TAFkyomk3lPXdMaTef0G7xNd
E6xYHXcGrdaH16AihfZiNKne65wkxOaghL5sPKnouOL3TsYi4VY/zeFBVENsuK1Aeb8q6CR1quvN
wZduXeD3zsMREdfHlacl9kyauy8jf3N7GGveU6lbJsH3u1z+c4Hc5vLbnooBDDfWzafpw7P/0ilJ
esUG3rta3OJrW5h34olpri92pBZqDOBgq4fBycsUqUIP1ErNbBMyQJoskj9K/1lRi2o5A9Z0SRxB
mTxq3f8ZQto4Mn/fZlorxAsyOflXdso7uOvgOm2QEmLDlSGvk7r7HttsCjtt1osZtHrwcdKKHDyn
8vs7MtwmF+gFH2YJXUINQ5wsMhT6PKo5e4oDf5ui5LP4cJSUPpPlXfw0tvGoFIFJKBntlj6kSLiZ
E+dHLEnnxkg+DSwdAlVrwVr/CM/zaoZbCWOY/Ibc8f+K1XTpDt50j1OvsKRFrsqLhFIf/1ug4xU/
IwjhHJ+qyusdyqjp3s3fd0/PNLZEi6QwNtNXxZ8Iedsnh7ddf/zgnOfLn1OFLi7RxR3PyHsX9LHC
kyFkp2vwTTHYaGyzvUx9kMfm3NHLJGcYzlzqje+yDhtJEuQV+/BLRrc4g+fC26Q7/rEr7Yce1oQj
UFQLRZ9WvqXfXSraZnfaNM11sT1sNLO5QstbVuynf+DEoO/pSOTzzSJVB4vu95GBR0rdSNKRHR70
mg/Cl1+w8+Px2ae3HzjM87oX9Pu4/A5vfvM6wu1eAelyw3tRObfJtX/6e5Tn8NCz2EOjiPkB+49N
+ElVQ5Yuc2SWUEEtDwKPa7u78bnU4JTd4IoO1B99TeHQiiWfN0Ugr6PD/ITnluv4O5DJJsj44fKo
clvIsnVpd78o9uI+hqz7YtbUOpcJjtFX1wWNA68fB5bUXNy7rPnLOlLGLo9LfMLs88+BA3XHEqQ2
O4etEo8yTO6+HmPMeWeYowoOk6OXzfP69gqCIJoThb/RBHIkuF2F9Bc0Nren1IQE8U667yhx7k/h
+SX1rwhPPUspUUbdn0NMZyF48Hzfx7ZDrwBnMX0OC2WPJUfwVBDLVjWgUMiohkaNepF81ikIcw7H
BvvAVCcfbRnSR6iSqWEoW6uvvNWyHVaIy9E6fukc/RNRdHgOxaxowzptk10UFLPLaYE3Qwsj857k
8S+NaSmEMcoU9TsCPR5aO3ygnI+QMNB1IJIn6AypfLcc0lH9lqPuWNvOesT3J31Vt50wStrKvlk9
jCIPDxo+etfvzbuY/aUPawdSDDdtqAMxe62n/PAuV3J/cL8csJpQEo9U2zyy6US1N5vn/8N5W7d/
KfoH8kTYfEZm4I7LGFg0IPzYnFCOG40uw7UJzQoffP1D1+VXHdPD3IxV+HqRDZTygjR8xNBbaF/Y
WxZ2yrD1CCbchZ8cV66mNGkggl5fgqmH0lVOt1SU4q+gTMb08O4vuJ+tz1q6H6ouJUUUO9zD5824
fU+E2CYnlssfL/XlaPhoK/7w8qAUgwryQYhaTNM2cMGdkW/MoHXQqXZDWbm0wkCuJq8u/izi2L98
btbKzmCB4RZ5aOmHr1h57lfAV1iSpCJ5kPfYUWjH0KjRp/SblRbjT9SRsn+4kb/QGs3oDJQC0TM9
DR4zeljjeSG3N3UO1sfbX9Q5UGL2IiGb2YEUX+abitE62N6kXGBYPKpOylKgRmJNoY5U2LBgBtji
GifpLg7IhFZRt7smtp0MrYc3oqJbsbCCEr1d4PB6SnRib686DroChNu0F8ZST4ZauwabxmVSLvBq
+Exf74GIiIAjnK7CK+1L13tuypppO98c/KEF7QgAbnF4xcFxtE8fIGiVGv/ukwuILlAw95LTxV8R
AqB8c91znHjBL8IY43X5YnfWwIViu8V8pHYvzxrUYdWwGwU6fgxkvfpUG+tpJNQkbYjBNzEVkMdO
e2uBC4ixNH/128YKuQnJYyCuT6W7eFGCC1+rdkSYcGv8K928w5MDa3wchY2BqnQILxKIKZ0j4dHM
hfZ0vlFoBuufdISb0RpMX0qlpH0RQwp+7xc1jkmpS0Nqah+ItkUs2qgKnL89yVzRwgOka0mk4kqZ
gUnoQkwzNf9Kl6HWfyryijXxHRLxm5wDMGY3n+OVFDXGreVEXbQKEje5U7MvdhW/6+YOAMvwsofG
ZmzEn+Syh98J9fhbKfhJWaDxQI1zbHFlpci5RMC0EN3iNmA/stPt34CNCaRzDPTxB5jF5mbHZ30p
3T4o1if5FEDxbMir1YVVNXUgKm/8mV2QayuU2vA6c3CpylDVkVz5XQ8I7YA5ELfs2zKvLFaCAbQL
Ootu7cFm1fywtXj0TXx8SuaYQ2Ql8fh/mUBD/N+1xO7pBfut+7Cqz4GWXzUwb63QqKqj5W0u7isx
e4xbszw8cCXyjOVa1MeutVUSLPe3M20VGIq8tODIDpm+2ijLys1A33M/mIP2NOKMzkrlKIlsvJQ+
Ci/M4B9cM35Ic+bKk6p0Pj+MQeVuGwFO/3KQIVFJ6VHFHFB1r0uQu7HBNLRThU4wgPvVt8B6UQgT
vQSrMXLXWwmhakGuA580VAAPVw08O4v223LZ1ZTxzHcdxUvAHVOhfj9YBaOoBSZSWwUczoiko7tH
Ob9n+UPK+W/OKGROgvUk+LbeFuhbT8kD2eKT0B8Wmp0neseqadtO472Wf81NmCc401uLg1/H/fJs
oHflpJGslwwRjvI24RSCu2bW2TkzrUzjIT9ytIyZU5i9HsxdWUGk76364Dem5RMtUmLwyQGtHPE7
J4ix7LYDiOxYiwsnnSSV0aAeTScD3J9xLgoHszBJFli0KW12VALtAUxcDF72euAHiV5ZJb+GWLa1
f4EYQUo8j9IG4O2t0uNOqJgV9ptTMzTB+yiixFFdfM6IVcqCuF81dA1B6XUzTrDbbxDTMiqgdTvM
lPu2ezDFqjfLFyD6s1UnmIptD/nI0taXQ0FHMeDGXIKEMm/Li7nlNSO1pNi8wmRK35zIt81NuDo/
edvex2NciAxCEbvPRptS4s2mCM93/BJwKxaeMilSUZK87qnPjT1zrrzfQvAUqKDIhvChDjR3ibW1
XTYwTIAfMe0xqbcxPGxVkYYzD8j2oWV3uaPWxKwl4LiepaDewwhhSKSr2lXPX9zdO0pGE3poXWzV
TobAmPtwa6D5aNZINvKqqPv0MHKWJw6gBj60DmxYh4glBnn2ZxKp0T7/B8G6KAQ9QjVw+g2CS+Dl
M7cSVrbN72I2yDK1OtikMaCxDxW7N/oFmfekogQi0RJzuK4qFuYPdV3JU6n5Bt2bpqRDjrDpcUC4
lP1+1B31uYepBKWnZ4ae1a1A8GBBvSBkTLfAmAd39uVPCc81GPjviMhxhoY9L+4vXICHqIQptWxj
4/28YhqLATRaf2mlxS+zeMGafRHomh6E2Ic2vTV/So7NCyu02Vv4tKfJMslWP0q10NLaIIrldfgm
HYInbDuumT5nM6eWMKjqXwygpvs5KMoXqN8hlqx7BGPFpJJ3Szss2C3yOxwOcKqV1vzTzxVKeBtj
vXEWTo1tlQ/RP9cr/3mJabs+8Ao+7I3eVMf5/T7kRjxTeX8tr0hLKyEZg4A9irSCa3cdTeuTj9LK
YU/i6m7OJq+sMUJC+7lUPVE1DtS+J/2eekrd1V/Jtb6qTiAHxrBNES9RFT1YDzVysC2vecw7APOv
LqG7KU80qyr62hMKjbloIESP+ardOZCvYgbtGCMor913lEpG8YOKidoZRbTxB/+pIFXi+8y8bJRo
cKorRbB4JHF/cfPdvGMXAj2KrTKR5KpktfrG74u+IzUSxbM6DyIzvQ0ceGGpxyZo3sBUZFfrV0bY
FPCi6JGH9MzXNn2As18LrYFH1EDKUQVe6IBW78mY8UCpeYNPpp3ezUBDGdNybuZnHiT3nvq/aeXB
MiF+wJJQBwQ1PwEHoEk/KbA5peCBCO6oMvIDq0WRnBI3MWo+6oMtdqR0aBc4lG9fwZWr95UBItLV
cOBpA0yFEgaJkgJPZm93TwUXSoX7RwcB7tFPR2V36EtktIMcUfSFSBnLA3puEH7qkAcWYs/sLdrM
nKwnGYFvJYiUmLBl6Yx0asiJNomwb6qj2BVSy13j3mt9laNd+4lC+XE65tMd4nJPbFekETvSN8lT
obWdnZrXn2fIJ562AvX8yxn3hNfdcHdm3Zx5B5kJbzAk888CV2IOMTuhKJh62/xo5SW+3bbWNkGk
Y0sncUhJ4jUqxww8PjZ5djfknNGl2IY+IgYMlHGBgGj0t8zVuap7IWdm0rQLk7zYixWBz2u0iQ9V
KuiVE1zDN3cmv+X3wX8n5aDyRokxJvyheavjk/5qUzwOosusRH/Yb0Mttf38nIkhXR00REjB1b0M
LsmVZKGxf7DxXnSVp88PCA15e34zMEgxuijRi2Jeo/h9osRSQwiCfru7wwuoJ72wCViEsHQ1riIx
9XVpO7KTipMSSdDBRVF7ZHHDDyQEfqNOmVcZluSgu4K8RBUZ66Bz4bHD8S3NsTaJCJUxnOfZhTOr
yOVgbZfxv7yQnSWcdoJOF8vBb5thGue1k/ivQqWlDl/Yc7jfCJsWfY7hTgLvGiTGpupka9l021P3
BHr9rOxbHKqmdTsr36DL1b/S2fuL85TMUbi/0Od9UPGLzEagn/MlRRPeQ4Tstd1UcsVdYi9OadM7
83kfWV7yWOJMQmrfJlWTINfnJM2eyf7ad60T6aXEEasy/qM4gGfTson4tNDRfNGCQ4l4C2Jxysvl
JiVwM/CF4qG/ZnKER8/aSDie2lazPvkp/KIeRDCgrcQBFIa4j7LhTr0sSHOYrd83Z+aqoEuZbjCI
yb1kePB2HyFQ49ZNuRObJa9jOVLYprv1Moq4AyM0VGLFulKWi7oTToRCv5I4jZ/wxWzlQM9wayOp
6X32H983P5STU0WFJymnZJ//BdkEMOtwHvoGoZVQrVZfin/S7tmTeFimixUjzZeWif3k4aaavbpf
DH/3fMhZwOeqOS+PXxW6SEXYW+aXNtsXjdqpEZtzwokE0hYu3CpEoQvNCd3ypQAoaej0VapuJuwN
PKNPMfGrijC1A+JZWkmVeTAL31eJnz6JuniueXsiQEhYg/qmm41+MEkiX+GaIB4S/bAq6CGwofrP
GPbWlxAJK0hpk5ygqYdqCnD2XD42kICpnnABULZfRDbS1SUuSfKop7sn4knwnJUaQJ+Ll15fllFX
ZqKkq/g1j0RRw4AD4v4ou3xWhLqcY8UAX+nHe3S19dInHVrPITrfYh3X7hKOA7Fv0dSAg88wfQ8Y
hIbYJ09dQn6XW+DaFp4CRzGoUmEXMaj07jQh7x0PAwQ9zfS4pPOscYjqAS5I5XKu+9avsziEwU3A
/VMLzIbD49jbHASuGBi+oN3QoXGk4VApb2MoV7UZjuLTKKbHJ1RNmpHxKxN66uxWhqKNK54HVIK5
CVtK73Ci5rSnoIXhODwd5bKMYSz7IPwIFmSWWbHA0V3GkVR3mn4A9Ch5L2s/mV1fOpIyaVFxkXOC
tDXVZYEAQTgVahvA5lUYbZRuj45KPQgu9Kcw6Sdg93GDbYO/qqIbu1lXA/4UtEM3Gne8ZjCu5iY/
i5lQ+DHbLkgc81sIEqXg0+vir5B3HFaqDDWHJP2Q6Xsvi037mNZI6iHCZgfXN2nYeMO0dOBWaNB/
f35E7k/1yqWfkY3bm70X7Tto4k0XfKQj+WlwcDokbDjUHhS7iM3WKX7nGCie8QZBTGyEcMhIb47S
A+FSOBDZj0TY6KGx1MAO2XDseU0aJszNc55aiN/YrhndjX0yGI8poGgq/vB9V0jxlkZEJA84FZFO
pKEjUqExAwoYsdwupY/YRLldwWzqnZSwZ5NEPIEfZb0o8s4xCw108Ct+ca8/oLzQnA9/mx07uQ4F
BTp5SpsTozxRKvW1bW77iIQ7+NXPgNh5XY0kX5Qo4q0b78Z95aQ2yPRaUC2k9hcE6oya4bnp86iY
1yRYwqKnKCRbSLdFiJblEa3U/DuSL8ZncHIzd0DMxkLORrlArxlNdalajCeQUDZ4h+xU3mVYORkj
u6iDdVWjHWs2T4GA1Crs6X0phdov0UpLTHIrBEMQ06/W8gNraNQtGXgFhTZeUOV+u46xTKEdM8oJ
hNEjC0SG2/Z/2Nze/1Rf5lMA0Dvkef9ZSXdvx9ByArXY1YSkgsVRA8lpywMfyr45+MDmwYH/42zM
FRCYr30W6J1k/jw+x3xrGU/95yCTdVh7+rETfgK4oFpN63k04S86HkutPqgk/JTQR1pvjsB8fSie
+tEV5YppEXqjfHcJW1JCTTHFghP7HNV6l15b6bgMmay/bQ6Hw81gvNL7vcnAMQx7zAo7tKadljxk
pCtTau7MAnb4GcVqSJzpo5zsK7oMU3xXenvVcUYyccRBOKgSpPb+XmbV8dlOAZJm4afhzfUkdMOZ
5dpVg9RNcqojiN5X1DHzZSeQJGoo++RpkmsWqNt/N8bqWsq1ClFQlpgr1IYkFDYR0bxVaAgdl9D8
qep2sbn9/F9nnIk62AjnUiR4GPjBCh6oI792pOn3gDlCStVSE8rvyxNzSWK5pSWH8hbIEgIDjn4N
MA+JcN7IWIZwx7WQoBY6Z9FczXrBVQ0f0YpdKnJvfeDUCW+shQT1W07scy1Nb7limfhSF/CplCmr
R0QHyDX5/s522x+qozLuR24q0tzbOXGUVAepFePUbXqBC5xzg2p6hX/VEmLMMh4LN0W9mUYONWoQ
nfqp+VtywMpMOhGorPqhf0zhv++OUH1vbUDK05Dq3mk0fGxGW/QeVLlGhc44QOtOZdlR0XB8v+gH
SxDPOaJmTomJaSAlMRqHRBpFNbRiOWLmmGLesGH9oaKcBpn0g/+rPITeCmwcmUak0tfcTBbLne1O
ATT1qn3EozjMQEokoSCW1kZ5pq/vIwYZsFFF+EifQeCIzigPIzAENFIaG23rvVCxrJG+qZ4rsOMH
m35nWsSd+INUTPybjIk1H54y9Hl4Vz+Id+wIhMdrkXq6kpkDW2rFq/IOPm86FoLxfJ8AP0cASSi3
/a1BRd1eJCraf0/Yde7ZD+LkRqv5Iy0kEpy4u7wHg/5JpMZ3ieNjChBl7r9x2j5H5ZnyIWVmKvrk
TrJYbRTQf8axg28TeCtVkhWDwyCh0j+pD3epr95/boEcUr6cwOU3s/iovH6FEmKe/SdTidC0kfeH
q44awcgYm/nn721yD8aJObuP9K+Kq+ISY+54qm4un8ucwOV1jky67WrnVmeoxxRGsoZGQE0uBKhc
VFmXlLnIuEpEkNDm1b30cONAA9EZDXJSqrLDwGs3wWAaUUJIbgFtu7K50CCZcbfdNom3Eieb5XSM
oEM9uHHLeNVXKx7bJA0TgYuB/fmwwaF396M4vfgUSJzJOBhTIHlqtgoIidariPUVYxIuNbkiccc1
ynHypw9gtAzfqLDNGyujgoMiudboc6C3OBDOGcLVMDLub1v+rCJJm8I9HOkgVkmNTjwCbUiSUP+V
pEQuvitZ7VdA4ZWOvjI441YS+1bEg/Zgcxre/UW5TJAuGwiVn14JVbZzrHBmHotCR3g/g8+6cop1
nzhXE6ScoG/0cJgiUtr0OPRzT87A9yVLuMo281WXjdMFWs7Ma/0fqUSvnjkGSt2I733YDM7CaQti
0+ygDmDNfsT9C3QmGxYByk/HsSd6/ofIAmcTpdS9LQfORk/3H9NsUnkyo4SGTSoH6GQRyAa/uHTI
1/GvPUKXvpOGkjsnx8gDq5g3zFG55d8X+YhKCFsyMBvjJz4k02s8F0aiL35dXoIEcDKDId7jlp21
pfJ934tgup9fUAdCiV+icyj0wMam1G7iH4ca8Y+1peSYhggBRSTHMBPBVEoi0ngHnsIgk+D90Evr
Dd2bpo9Lq0wQZp42jr47jLHDEgWAvmEneY6RvyEzVE+V9etjK91zBU6r0zLTNP71zAxUsn00Aw0B
ycObrbIG/biytxnQ47f7R2nYEKXhcu9iEuhnP31GCJQAC0RFDSBj+j4d018bbHAEFmJT5JAqshk7
GfzeIVwrJFFgcE18ozWaxaFgg+/RiRktySUw/nrATVCU4ngBw8Xjv+BkQtf/WkBc0mVwXs3dosMV
r8h+Hu8Qj2pFXt8wEFccPNXLAC9HISb5z/d9UDztbdOu/xqZqvbJiwZbbJZdFC3GWEKF9MGQWSQf
8xquu/RzXXXjedh+oN38ypY1ZIEQHrF7ugy02eWW5At42Pb7hAYv5BDnzvFTqxAQNx1wsN39iI+4
QCfkndxQt2AmsMtw13xfbPAUuIbSSGTcsi18WhRemYvIbbks8H6lHWmKfjoxpy2PW3FRxYXGMHvt
CErns1szVNucC9glAr9yE9rk5zmlEw/dApsRQ8XCXHdlJIZiCpxQNbwfFCGDm0+Xz9r7sHcikFYb
FmLbO09AA5IQMfgEOv6O61owfEcr0MlcZdCWJ3/mDdrAZuOzZW+jxxaQzXckOBhCPgh/97bE4Az5
hr47jLbOD/XRqMjBGURcve7/QWf8k/kd9BRNIWn1RmtvgyHf+KVd2FRDu3VGRwWnatrvnyKW2NO8
iTrbo7N0SMikHeLVOvhX7tZGTc++fsSEoASXQb4KA5C4aI3jIqEAK5qf9Qf0KYc2qJvhPCOqP/Ws
wBs2AQP4RKvee9dIPriUkebUtBg6M0I3k0e/miNJAk0LrvYI9/nuVpLAvyCsEmWY9YGa/bp9bfeC
WqEWkI4GdZenrAAQ19bfzCz0FYpo0RiNnl7WXniFYyOc2QmRoxpazoXXq9omg+ukTfet7wtgBmec
n6rsObQr6tXWmn/lijiQDzN8fqaNBBHnjMMQMY6gkdmQyHd6u5/m4m+YOS2TtuWosA+YSVbwKGCd
aGSr2rRa8P0bqUXBhvsSddmjzLmsoth7kj7L4Et9mDZj1Ick1S6/CyNvwMvukGyiNPDvjeb3o4mT
eCjh646IqN+rYzzAG9zu8e46GBjivXW8aYF9rjfkaFthfo5piL8BMfKmzRjltsVxWePDYIYZFA+9
FV8akS4F2+gInSIp+Z06VkoCZpJ2RrV+MgbwsgNAxihE52YAp0HgoCJUWcMySGZtDqcjYJ9ti3uK
pHE/3WtUw94mg52y6j1fUyohYC0lrTin3fiBABXqo6kGrWfkvtkQ6m0QHTf/4vPjS0N57A+uTrh5
CQ5WBrWQLiAYtwjWa2HP8VT8dq82gcFLPLVZ0LiD/tViVpwkEY9EuuFpssQSub4tUpejsNLRLeqL
XluzVoPtmLwqvmd2ouCQNdF1ejbtKk1KWbIXq+TPW6RQ9No9R9SDOxiJ40oboSOiM42uvL9gFjIS
3jzor2kbAV2sQuZPslKlLoM/B0vT/0zJN9QpgptuLa6T1bIUOQoROOVNChLUPCPE1k8TYNss20X2
f26C4sWT8Q8VSZ4ERO/WHNaVGF44bnBM2/AuNCP8yaEQJInQu5sGegxvl303zxRLiRqE8A6F92jA
LR7uDF3piBa39keS4tUmpKsqMYWSttymOHZ1VzwdKymDmLYLOidGfQAFSgizqSywmeUIQAqpv5FD
1Y1u4sE3avaQPGqu9OstH9fyDG/E8sVIOLUW1kRJu45OqMdLbOjIxbXVmtoU6LykJPGlmJYz4OEO
UAUHBiEbIGtZY+1KVma5JAbg9IgzNapzvwGfYCnktx/qwoeeKjbTDOi6f5MqBR/CQASfo+6jlkpR
XWUaxmBD5kk/o9EhKbw1LYpKV/kaluZPm854aAVSe6nR9+ugZeUT/jH9XgIaui7POGbENm1IR1g8
bGncNgUVZSvL5vnilagcZqifDUok4VjZ5LoAq0yP0rerFD2jE4a+/G+hAlBDyc0T08sAx9FVnsLS
UQvLz78kXUayUllEDmLdJnw63W/oM2vDfcpK//cZhqfP41zQM98m7BtPw7UWn8ej/dLjukegHZAk
nodd3BhL/3ia0c/xorVSDa92V81+k173K83Ky4b1DBSHfNkpqNxSCGZk0WkfZB8RCkiKLQtFEG4X
UXc+Dw4vfM2XyrCPzDhW93KYQx28b8Tc6URWPAmbRjaaeMzjgePuALkKbmRC3F9LPyfuItBFxbnT
8TsPvM5QsDsEDhP/pZ+jfTryauC9JOdHQNLXQ8SCNhGH+5NBc6dvhOWqIqaPrX05R34rkOcL3gg4
S61k93UmIT+lTu0Vnf5Pbqkr2hlXl+vuuJrKxXDoDFl6UwHrF8PkGmv2VwHiOK1cegqBOB/lVTNf
mZNjK8V+Ruy2J/rijo/wZI+R044Bp876M+Pb4eBhiJsEYyQPMu+k2wJ1NV5ha/16tmmpeF9CNtEo
rD23VRubE6ByIWfbWg+b+XrC1GRs3iwjnXOFTVi1a4TK+CXH0xBBEzAmvg5E1+OuuHik1g0OkDCB
3lfw/LxUaO0qT0LiXVXG7nLxBzv0GMDztVRrPVZ5BsNPunW2ALgm0e9QH5+Srme6m+bId6VaQR4/
DMOXNlocnSfso8AeexfhQeFN27S9AjmIdD9iDDqWGCF4Zw1+pqdD2ULDDD/h1Id08LRe6ZkA3jJ3
5Lzyk8n0DG/eTJp2w5hpbTUl/1sNWECdlF2FB8GYydirzyWB/3ZhOXTrX7OxVq87BK4F/KwLbME+
cArDsB8738qUpgwClk1Su80z9qMkl0M14AnpkgBfr+8Y/QSTsJiumMNlgxFP05mjIbrCxxqX8RJB
0Oyln+Vtl4sT9CRM8gmXk4WkHy3Nw+mFzbqurja/+LdAx3acDA/dnnFv5Ov5So0RNEcL4AbwoxEs
BHxoyp7H+szkKwOvf0xs3htUEBcaillBcAPrwB+qRsphujDWYixX/MvspQoxXO3IwdezpMO9bMKt
yOGFy3+qAOZNPNAN3E6oExmhEbeHg0tSlHPBxtdZZIxsXy9AxOLjsNsauhkqPXWWRE6esCvEK6jj
NGjwAZ9D2R99mlJ4YnxOZqWPFw4ZfLOZ1ZJeKiDk6lfRWZVrKO/EELaH5uAvOPWPeZHEMM8PG4aP
CguxVMAK3S3crM9kAMN59J9BuOSYG7tI2X5M5uEh+zjS0DRR0du5P/1jJMj88XszRijrJ1tHqk2N
rw72TTD4PqURtN+5JhQaawnuTrLIDtJknCt9B+li4RW+0pO54n52w+/95YQx5q1apsEwCFAZIn41
FVqX2tFuCQuDlROGFduY2H2YnTUhhEI6YylEXf0kY78EPwT+sAGniWgdhsjQjROmByErZZQnA8xl
Pb5iYJNTpyXY+NQhDXoVbn8qf0BTWd8L+XVPwIJaQTkCcmcu7l8zfzc/aDaGHEN4dL+9+G9egG6m
IALITL7MiaclTeEdmbfHuH2uZ0gzJCkZUA4xz2eEEHHASvHQQsOyLticQcoFOb5pGbwz4GHiyB0Y
g2lcOWb+wI5ElOrVrrsS2s2VB/xgnWVWMkgm7tfIsEVwvvHuaHpQLaEaHLQD+GUTvTt/+di982Hb
0LIsTfuWhQZM/tDX7ZOpvlI7+rJK/zgAgXhlCPDh+jfCmF4tASrccdc7YimWeyr7AhDNsTs2FARW
2ZuOaLRkR50b9nj1/3ONFQP2gvCKs5S1Z9NKOhxoBdK/vFyBJPoZvSsiiwU8Vlq2vSUxqt8kD6U8
5Xh9SlGJ95BIkE9FiyAIGZYBp4nbhdDP355n8dZ/E7sxxP56pKWvUtiEwnvXTK4y4zpLmM0367Fo
C6DT8lFmJwSg09hOxCEpmPGPvDGLn8z1OTI1CPhJEX/1oz2XhLF3Chr3ACxkHvA21bpYggzHtwf0
7v55PldqrSkiCKDq4xVLA+eJ92mmJknbmq8VSp1SvkUDjykUtVhsmHtbmPhvL8TG0AvEfh1bia/v
GHGivEevSCEdbWQzGlYDzUYeygetwKtcYpoIIl3HqbGeGDARWe4s6wKrdScTezn4Z/3CCySmV36S
9dMcQaA3XdIfsU75FU9Ac4Y4j/Nrd4FDTH++0cbre3lKKd05lzbSPZfDOizonYu1Bvf+J5yiETHy
MSMV86AzFTPMuO7TXiof5B50Oa71cwWPmUwabyzW0GQDAAm8GoZbzYLrl4Ot5ExPpIi0HDt51AH/
6xLFuYswDCR0+gRSXCg2ka4HC9/1vR7LOdEWrqGwvScVdbv6QBXslHYHsx2/4s6GUGFKYrdmYYJI
1P6VFW3JIAXtu3JH13Tnlit5ASDc2LxqO9+LHda55Sq5OSJGwHb+UwpIuZqqn7IkakHUqo1fbSSA
x8AygYQyDSutmfX7e0/x6iddWaHuJCERY6iLZXqCbdG3vNnDOgcAZ5lzY/v1GB8j/QHxm2JygID4
k/7eXuIN0zgw0Fi2+3AkycN7wBtbtOzlDxWQxwCrJ6lQkSsekchEnjIbBX783dGySgUmi7JVjvX+
CdH193aSOznAVgUxyJPZVtja1TutglqQMXOY0Jy4s3gXjperxfvsWAT2sc0pmEOTsJNnqfla+q9J
8nrMdoppzEVupeXkk3E6rK2aASGrTiKudkZoFK+2H7HinZrMh4is3CvpburFbDIIB5lkCH54hQMR
cV2Hn6gh8Grllm4I26TRxkF8QLSQgcgp886zGv8bK6ycA/ug9mlEfd19EdMGIKh6x+eP09Dl3Frt
4bGOpKmUXPxS4TGaa7q1R3O8avoOsrHsdFJoNGPxglM+6WlLENlwTCrq//RqXTYyTQ20ZDpwbmcm
8WWmIEZjELdvLm0XeCsD8sXLm5DD3Kw7xTlIsmjfOZr9h65o0dNzkAW5CI5OffQUNvaITTG55sFq
XCr8toqwGIyndZ9SK4x1+196byusztHtB7SsfgrmoyADcyRzLAVqcFyqtgCWE49sl1e+UjwAKliM
+6CeH+lrAuBPSUDsJ+RG/oLMACMLAMBcdqYjEVR4BnkF8idkKHN2/lMjP7Ju8UBbFOMX25iA1z1B
P6Zpv722lJSfmnMUcc7FUugeUhAn7GVAEo+EMyyIxBCctifwaqf2euZf6RGCNJUXyt4ZAbl3Wa+L
ABIf3vdSSpIsIr5gpFz/MSichcuOlSj8FVLrezaU5He+65fmK7HZVmdPSr4XnwM4nj+Wyg8gS36c
UE0pnH9wRFnCZkhaXNpdrGMiRZNJCo3b0lDJbZp2HJ2EkJKYGjN2V4m33DrQ/PrQObDVTmRsieH5
2fKqgQ1vP0GvW8yRGIsQUxmSG+oBaNNOCozQfel/XaKIDCnToSAQsRNS6gdUn3sa6qLwNp7FHWia
QwC8kw3iAn+JMtVAu7MOU2zPwLmBXIQc6fbxEOv3QgYtnLSPgA3B+2pJ5uIsmym+N62AlwkT2XdP
WIOp87Mm2HfH+vQgtNgGwAaM9Q1ts3c5Zbhe7uPVcI1CwLReq5RtdAx8pMuuVInQ3P3Rw7VbDIWD
8rLCOCaZmp4s2Wzr3YW30DtGw6b76WjtaLm25tDg4HfKftTSavJezAOxEvgEhaeCWnsxM1M/07Jt
WS1t/Oyk67FTcacP7MWWav8vtD7+W/mgnQWPX4X5Bm8Q3lTloCDaYERgunvLcV9A+FH47uEuyeb4
Wn8Kow9ft6E6WqcpARUXVkdQ+3g2h2VwiYX/Y5mInTq0/XxjSWhIs8fMN3M/kX3g7E5LigOsLWXF
JjT4qMSC3bfnwUfyI8ERX0Cy/PtTC0S83DalbmxUbG8xQJOki0tPz6rdnNZ/heqAHsWD+K/nA4mC
RLWfNyEVhHB89aL64v89ZkNkHjG3QKmjLWL2buM5nkFeCPd5XcmW0FICsnn4cUSn8094oVB2c8dj
aqXgKsJhwSVcZOo5YFN4Sm8luczL5pzKsWtnAGGAYcznKYc9cBIJcIBw498yzE6atzjwE3m7SJp5
0iZvczbsPQa5XjFTvDcSJfHxcv9OyjfgI/8PdEfZM4s1/VISIOOexkJgK08XdAVkrLS17HBLDNPi
h8vg4OzvXY0T/oEZuBW7MbHVq7uvenRbiNnyJmmzzZUD7W6h+YEx9hJ/QFFaU6XRPJ9N43WjXk1e
W0sh+0a31yWxJvPkBxm4w7pm0Uiv9ls85QbdlrwOmP6K8wg33ARpnMmsbPNCODCI55xct04Td03Z
6qAeoJkY20XZCJ6vJ9/aiaHXdXvl8Ibs8Bh4dBkmb34knHhwHVi4pmUuJHZ3qgHx+QXAFjuWcngI
rAS3/VZC/6taoV/l2ioMN9So8OgXzkFKLoNO0zUkCAkPAs/fVNSZeWpz8FqM8cOXF4xRTYJnh1D4
Q2bsUJf0druThr6xTsv/a+3ByuUStr8ICkw2gjMeN3ouOx8wjUP2RINsxCOsw++qAH8DajeQe0zm
zEGr+sQJy2PPhqVz8mlc/3qyN7wvGAb6r+mB7zNbDaYOxQ4GaKwP+1taJXQthzSU/WBI5UFB2YtG
7S7VXgSzvbHPvXYNeeLFMP6nWPHvGsXDaqH8JtQY65Q12g4WmWGC3wNeyUxnH3aq2+TfYVv8vBtI
hQN16pdRtNrh3OqcSEdsukjbo7ZqMKTS90AS8TryM/60D+Bz5dCuOqW3kPKQ/zhSdaoAx4BD7fXd
ux55Az696i8Cfwlrs3QY9w/l0HoSCpy6Dq7xV5CvG+Yl2ZD2IrNCZV3ea2k/6oMiki0m1smMN/2j
J3tFU73WPjc3scXdAN9XJ6uRn0n120LHYEP+8dTB3y5x5yn5fIsUTqny44xVcAk3bdfLIQrgtUUo
KW0y8Omv+rmGScWHLN2ACnoItVm6vKhc1DbIjBgC7xk+mcRWeau7hxAkbfelxWtUuXXiLupXRqOH
L+Uha1H1fAW/wyhTiaBZhs9lt9tPt6yCGXgcdbtuoJ4zEwS1bfSB0Mk2TUPxmL6e+PN/g8WYoTLa
YOHMPb5CcCjLe8ThcT9h+G8tpdsLDGECrJbEYnx0xFCy8675IFvKirmH4fOoN8nUXxGloBSJSfzI
JxpkmGa45AVqMyBvK1tb7K6xLghsLJRtfbRy47UCqvTB5kzsj5HGj7bxS7VmGvY9Xb1XndDrqFNi
WGUrHH3Q/oPo3OZ8q7FrFFVaTFY9wRGkdYl8jkI5qo0oyLgNTKbnLyCFQq0f6PJqtT6NPTCbso87
U3j/I1O6gCbdWH7GN6/e5sMnvVUxjsCQuUBvPeKZAL0Os33Io8nqiXEg0b84YCyXYaOyh7Wk41eh
6I+hBSGYlgPyjEKRUbm3GK1PaCTb39DQxwIOo9riG81YUITkzWdpmf+UO4ERh+rqio27DLOmSvDY
oolZhhj3pajg+xRjAKLhA5o2dGe6CUfjwNBfq3qaygEc++kvSo0qQlws3eE/OKsZBhbBwdf9LKSD
ah2eq22J/D+HC/P+I03KH93CJPBucT03I6a1ab4JgFYJcNI+P9EkLko8u7/O9Not/ylTeodYw9iT
M4a5wRRR8vX7CZy3VSaS4z13LLrghNH+q1q2MTbcU6n4LNFoctwF8GwR0LxaAoH9vyBfnjr9QqpQ
5cp3lNsnSAvpTVJrhxWH7+C69vG8O35c5fzvNvoAjS4lTUfCl4VGdnig34IyQR3ZEkoCyN/o/HoF
QOmArr91aMzcE0AcxwD75hNZe+pg4ZzUr+k+gnnB6GtuPAWThamVO6FGrqOpI65+BYtf4eZg0hr0
QoyuZU8xyUzLroc/A+z4IG5bkBTaySe0rQd6YldXu2F6VkhJZgXSzjy/1zGLzx8gKxEnH9pZfcOw
joFXo86xJ6poE4LC3A1cC1NyI8ru4phGQdHPLSsVKAzoTBqxnOIVud3L43QazunSlGefKeUvvDGI
mrE6K3Uwz4IHhomzDVxg9DnHyXRXbmqf20EQP220Mj8Ojbl+Y5XCDOFdTYRox+3a6Y6msspnTWIl
RlPN9jTB512nG/9O4olGaoPAcAU7JHXhObNV58oyJBdNSEQI5yT1LJ1DvjO4z3P8Xe4w3BwEzrXp
zZ1nsVL++yi6g56tKzbXt0yzsnr2isnK6Da1FuuHhxSOkrGi9dvk2qKzY8VH5LVQ92JgZLG3rSs7
E8C8rm/lCIdS2LBWsa+NPuZf+dUHIJBBC56lFf4UrEP58YyVJ2kKgXY0K2KQwcVb+P2dK1La/sBI
je+Ww/AQR+DEBrw6qMdMFlzjOdIjiXmkRvcYyQmUWmdcxYoVFXaSJp5on3HUP4VckwQZgjZxB3Fv
2yRFD+xf5PcNxP0LVjv7v93eP54jTXxo6Lma+dfw7ZRRtzSK+sYw0jZAzmPEZU0UVELqbeBpBFdW
QxWz6k6C/8/xkeDsE4siS+aUEOHNRWNlKNzCrzfQSW/r0cdhauryWUcZLwsAqZHPJGWkrkuTf631
nbvkZUBSUi7GQH4vpvG+aAO6ZCwB9KHOGCjz8XhIUuTRmFBUpsC8ggfxYxu15VVPQTAraSg8KRlD
h3jkP42Ipv/4JL9DIVOtT4/eOh8GJ6dyaAKOUatP4SIdUJRBMWdZ8gfvKzCycRTuTVdNwDJe9DAP
+MxI6NPVFpNo6nRzzdPrkrWsroM6nzbmr19+iFqWY+MhOxYmp1uG3v91bLfYg8nHF5azOrWP40f9
skHVipI8au+72W7TOUdBolIEuaMCtXcFwl69dONmpKuUJUfLHCrAlzPf3OPnYm04R4wSvnREajjt
jYr2fcPP6/HZVgyv7tz6oafL65jfmjH6Pr6/39MQhiAz9FbWqemWYY7jkLtsgh2NKJLnrtNX56Cp
1j+xIKryv5s2udD8UaGs6YqSv6dUoFGhhI3aOjfPS2BMR3BfZRbxU9oZ/yPpqzgYwRhsmXftM1qo
J1jGaZmEEYFrd5wgAhE2iugOeCpfnYCNPtVZGyNqkPym3KRl1nMIotqlHkcnDbTE5l3U5Ruf93ZB
F6YIAgEZLse+CSBc8Rf4xJel0zeVGMQoGSrKJweLQm0Y9h4XT81zJnzyFF/rEPj4mS0tN/pw6VXS
1pdbFyKiAMhS2JidiXO51eMdEeJlULSPTvwkJUzzf3ngv4c/m6facMq/5jDwODRaqJwJ4cAOabww
F+p97KfWM/uAMlFJJvb1m13LJMkCAk1vMF3x/NwWWc2iZIzoaiscXdR7+1TepMXjvOK1GwWyYvXO
PmdgLO5XhJF9Ce+sF5xjboYy5G1hGVWfmpumJFtd55nuOvpIe5HJvxIDvoQyyrK7aVPLvGNm/ifx
tNsRSFvurzPQ0qf/rF7f/7ox7hy/cgjgqhvdJHtsNqkTP+z0DJMY7rg3f4/glE3g10RZmuIa6+tS
B+uWQUFXgABWbCk47n+axbC83Xb7qJRHWqkFsnNaLXsS3sixVI0S8NeXXk+WYByLOZbvg0hRsyF6
BDWdYYWWZcW+M8CJGadsVaX5K3eNyOoKVD6Fx/Cc2+WvN7kWFTLQjzprOqerzTvqPq9UNCw94YpU
5k6o7LRttreONt5wXso9gcaVi2u+rAdnJSjz59H1ZWHV8rceS/TGlzmarIpE3IR6KePbz4eS+t4p
QmxlwJaqEULKvIVuyeyDVo8oMKcbIb3KLTWQkvpsbwGiN+TjA2KOG8DNWL0dg6dLYgzEguWssKWQ
sffxqi9jPXC3ZuG12IQbWLspNE6qhHuStoBq6bBP4/ubDH/y3xr7afgxEVUkRKpVSAh0PA4sJi9W
bvUd7ZkdU/ueWW6a1wolbNSAaadFI6ey+TwOGqpBx8AiQXJZryLhMV/iad3cQttKfxDzJliOQuiq
fuVgkVDiA+E/SHLEMiEH7q1SQR70PfsLA3kW7ZfA/i1DAwr9+FpzLbCrry1ZpilNgQgmt6ZdV66t
roIXtNZ2m677d8546y66+aWvNy3Acn+WdK9B7/G51Eew9Atwws8UzcTmdLOApCVEKW9DhlkWeMPO
4ZL+sS/znniHZ5+Fv8Q2nFsRXoX0nH7DbMbtW4c/nuQKk6ZD97q0EEUokMx158GvtfpU6F1UXUiX
E08C6u5nrt21fq/2r6NHlundGd5DMDBSrWg52dh/uKQVuCSC+H3T7oZuqEHRgX9O0Wpo9HvvUMo1
+KvPhtjJ8ubmE5v5BZqhQHaiHHocXH4qJPms0GcH5pgPmlqk0+vAXC5K3vET9K7SqWSCOkOfAUJH
0zKSV1yXzZxUAQhqo1OM48M8bIhYCLW+AQAAY+1UANFXwhhiZQRwwjvVhm9SlUWBSBo+3wJfvSN6
+M4FosMGDnTWmakMR9iqjKay1thC05KphwwsdczEqc/r2lPRGZV6I6W1ukplEh3t/uAADwFmhatl
GjHyxURiSLqnFpQe3+neO8/IChGxS+Ta8HMsyV9rjmycxPHRj6arxoxq7Ly/S8iw3lcsJzrCT9fz
g6O9pUOCuJLRNpGsYcxNKE7Mo7nAhK38L73jIe+qkbbOTdBMrABfMNBBwgFCEjJ8V+8YywqbvK1z
jbqaL4qaVXnxQUTYjwlJMz8EI6nBEjx+dDyFRo0cAUp3Lawik3HOoZr6hwDFEVixkJoqo54VAIMG
fsLzDEOzC3M+yY2NpseUaEQ7gVIwORUWUQHSWJ/R7m5t6owDymEpPIWy9XMhP2igCZBVB9tnnR9B
y86rijSdk0j9s52UaFgDfeaQfMYkNTkYyJo39dZeuGNOltoznrQTmTbyXgbjo2DMvOAFZJS9Ev95
qPviMtgQrriPR014hLZzWDe0dv1fq6l1R8/n4wwvKdZ4JgVMVES9mSxrD34KjoJKHfERpPKisQi/
+meWaYkrDQhlKvQ9a3v/2/MmIxaTVj1UdZzxfZsGuTwFjVLzqS9qgoKycOgOuJgmoTgUPzJanJI8
V3AGa8KkpZnL/48g51Btv2F3sYnbfQ4Fle1Xszwe4/XkXws1+KoRAIqAns0U6zAMoAU3WRCnFxY9
fWqdUbE/lGJ7MnzXOkPIWpeTCy8FcWscdsK4gSR1eLruW4roa3mOMC+9vKXqDm99IPXIwPwdJtPW
+DYXoHVzcXzov1MGXA9NAI2lyvpUCL8CoQWj+O7wMBr3MFOsPtmfHWj7FybXNL3QgUgyfVE4cNR1
PkY/5Xhse70+3Thzttu01eO+Pc6fwyUkhYp09ueUO8ttD9Q1zh70csvfXaKulP1d3zXod0BHQcyj
wQwRLcq8cwV+Mh512bnbV70AR3P37p3qGqStpqy6Ugaz/4QN4ax7ePRT9ox+dAUOcV69/a+rXsN2
AtVfvAmUz8TAxXHwM4PLPEDTWnOu/EIiiawe1EuIi1JFmxGZnHm9WKfeOEE+659oonTrTQM78UNS
QqOfYRKDd8rzqOMqT5t1XcCTOFTBXBwR8uF1Pg+HprizzU7C5to+QlSsumW56WEjVI3LzNgr9nmT
rdZwZYAm5ABogOx3UhnYzIExiuXM/uZZTowXipNh0/q32GSAaGhtSFo3uC36XXL+EF4i2ibrEMCh
mSMgwESLOBlMqsaqgvPbIAcQrhE/3hsLl1nQgOxkgQQ2VJqx8bukQiEVc770oy4jJYs+CBZ8QSBf
VSfza2o3OYrBo9UMJNxgUz9lS9Y+v1WyMjgKU3BZifxm6if5Mo0aWbLCaKXqw+kPaLIIRBiK9vwq
TZbaqU28rPeRFMo1vuo2iRwnGCRMmXspMHcgzgSW2spguEerx3JMCWXR8zC5dnae4eNdFxsVLLsp
GHcow9gjnVfVMcuIVgOiPItCOx2jHXYZhna9G3EbnPHydUgaKR7Ve5AOgYCh8D8PVa6tDaRUp/T5
VnvZtgnWLUPhZ/wsaoenSwws2skuVvK0GZ3pRWpjPxU1tnaB0uMqoLyxWrt0D2jjryF7g7O0I5kI
8UYwA+sj4QbS3MNIJLIgPfKUVyhntlhlTgzHH0IifDFSWukTGk8rUaVHio2m4J748ugvUh+bQCiE
IXl9LCnF/KtCdf/D019lKWl4/oNin5OeYjLqdvI/VLXVqdcgNnAG+aovZNOyx61f2FoMxDT8rKCR
rUs0t2obK3F9d8CXOVurPy/cPUyDO9TB/R+dU3PvI1f7Yw0LOlpXrzq4Eku9tbryDAi/uvaVE2Cs
vsAFxtBIexRs6uCqlu1+LZN7t7Ny3/Yzfil/rcbAMoOpsid0jzBVV5s7+RPOe66xo4BtZ3Fy+lXe
rXbaM3iTVyEgDLMB+YpEqWvkRVlsndy0GJp+d/5Ee2/o/Ad4mGo6m+D2IDQU6Pj8T6SFtABmuqSh
Tg4VR5ejd6EYzC+0wiRuIqIviN/d05LhWt/rZ6/++3XYnKzR3x1tZUmaVRqVi4a56fwst7JTnY6/
4X/V6GgRAhaj0SSNmtHklPKXXH1QJH9CJD5fD0yac4FQyK0eBZLa24dglVATX19MIaE1l8scuDAB
FzndTct8EV6Eqv0SsIQqq1FhiS6vErUKsWiZKkZxgtbWNfe1xOeEWhUTYEu7H5YEHsrfTyUaCeeJ
GpONpeu21z5cLkZO++WcEgpF5QthSCVjYUH8HgVgM06GhHnKnuJmJhzVJJ73v/rh3C374zDcjP0Z
1tN9QsGhAGKNsEuM98oDoN1Y82kpoH5nmfRE0FnlOq9UlHWaFLS0dLx1AzAQNfKVoGnM+e9V+h9g
EKfF6PXmTbW83aYtNbd4tvtIudtAWS25soHWTj4wIDXF0zvo+dep0sF693wIDLbRvK0Xx/kuhVfQ
aDcggnMwDrDQAPyVIn5TccbdHQmn31j2YOph85Y2I7xhmDm1y102XbNf1UlRraUNJ6QjSxKKmcjJ
Hs4HueK3lylqyQhua/UkXGEZhqZrKj5I/GAm17AZqIvJcTiazVurtaczo/7BZGbq7szghI+J4uL2
fqdt6YyDBI08GJ+016buQWmTwdt4zMgJB7ilDS9NnFirH0IROfB2DTIlSsR6wvfjdSk6OtqReMFM
NeI6T/N/wLM9JrH9kpMCAjooZqgB73XCUYHY+97b5XClh29ySL4RfUXM/Gg6D5BviXMg+UDHBzUe
aPYRTUgRe0gaPg+wJNjkSPZbil+lIdMkTOLHBSOI3A0LHJ29UJUThg7DpJiLCqGmpGszNo043am2
lu/06lQoSfqFWYWrJkod/cLkk6lfqTo9oQrWdBxYXtIEFRcqddx92MbXrEniPZyA26i46CHDk1Ie
3wCZys+F4a0nw8TmWwcQyy9BYI7sEXfnVh9t0tSrznouiFY6abMQI+h4Hv+HdS4du6c1CukzCqX5
xnp+6XayFGEU/ZZC8or89CklaKwds9HLBhDWeBjoVxait27U2WW7LPMLL1cj8txfuCHK2h5m4757
3DTGVKezLVZvV/bzRwT43a7fh40COx5MhSMrUd9K2UcDetz/IpSJiUE+yXBLMLNVpycvhYU98y+1
hiWRpjCk7+IIkLSIXPAmy5IGZXodtYXNYElMQCvGiOnHj1iBuk80XHW6FVSaiv8waly1M8vSet2x
/3lTwyE8pSapuy/NkQ2zH8fFm4oD0dAcE6gzUK9A0WIGzfQLJMNWQLiPpgCJuYJYR/PuHG+voBIM
FH7y6w/igK1t0niHeqgmMDurwHcA3kYLWP4+YtHkb7BFg+S7ZTzIxv0s5qDsZpL7BPKU88pvsYKZ
PWpWBoPmJ0HRnEg9fpu8Kddcgr9KupL2H6zr5+E06UGA8AGL0ANy9WTrTAlV90uvJtdtJLjcFUIX
l8SEL6DZSoAiUcJPzFEIxmvd4CV1sHviqS9Rdq09bSTLPAdWcv56JfXnqjvwuVZHkeqSzxi4Ad6u
Xk0W0tqmN4xJFEqxsyWVQCQUbrxXlFJXfID18AFbaA6772F9C30Tc3A0UD++uLao84rfcAnzZjTh
2xNslnfAHn94c+AETogncbie/xhQVk/oPrzvGPEMmKJ06Z6flldUDbH6wwLeyHhp7K29TPOsQqZ9
Kv7FFVJ3ld9Eo7CDewy3Ma0o38KDjbjfUXrwOf2Odb4EUSlDdlO+W3SPONIum9z+uyBLuIllC8uO
BNtXS/+qB6/A8eZHKTW1QYfn2K5dG6Qw8agQJhADGMgSbwa6r16MqJmiveNjQLbxkarwmlXRHWad
9h65lFHZDsHU2J/OAmBoOgsaarca+lQd+XmKhqgVDXV2Kk7IXLLBZIqeHhv0/Xk9hNaW7MjaELsP
8uOBYAI2/k+j/fYe+X4eMNMsTJlwxz+ZgXyq0rpyCaj9tzzzWWR4JHa6gn/i4XVe9wGONSLGlJut
KUAED24SL4EHkczSJ07QC0eRvsazqLFfYIicbswacG5AKKGUi5aVFQn8BJNbGujXdEaFTh29HS99
X+qAL1dTP5gOHCBw9rn6RyYM4xh3wOCdJ+YHKoJquJY5mfIk1SWsqYcoRjdRBZfdDoBxoWkldyxV
RPkgixlVlrllzXK3Q/rpQitUgDR35h1hVxhZ8xoJllasL6HKFa7WjqQ0ZX16P4hAmALAjWmODfO6
Isz+Vst6IP3VGtOxvHAb7IPxMq5VHiOqfYO2p3o33lMrKSLc2t7Lr7wiBgrulMjj65LTbjBL3zBE
D3kIGbzX7n8Ve3An4AJwAczMdfwS9bWNe8HCY6fNw+tZUAAWWVouP7SaoGkB6KDihDtg6zVM6UZa
MJhmhyGcbc+1aJgTo8wuNBwJ/rvUeTGDsKkTGqOFZVszMkc/2elA8QL5DFbxnEDkfhUDdFK3EwG9
k8EexcU8WT+lxhOxIwI8W6vuAf/0Yr5op4BwlB7/NHtCCxdKvP/YP8VMQHc0Hsj0k3mWvyo9lKmq
RY/rwZ1NaJXE4rgUbbuVHeBmigIIqd9wDfdF4BHIaxoB7CJ2HHk+1XvZdQ+emRztxnKDTpKTpFZZ
ujHxiXXBQ1V/xJBRcYLKN693Hyk2asFmBtmChDxdeo4Gi3l3Tjn2AeTMhz7j17dfMqslNySA7php
bZtrq0koFMfh8UamzekBRdVbll4F7KK85E9hFq1ozk3S6voqBIIhNQT8jiOmz3t4q9A2n0+pblSM
l78NuUtCEdaLbrx37wSwZQCpIDNHm5dCF4Mh/HtxKXnNnsM7bScd/U2x0W5hhaxzaxsVaW8Jynjz
jmHIRRpmA18PCTyCZ56t0p4Ug5mUfoGWnjpufqjAjk3Yn6GFH3GCgWapl9P6mzvLmB0bYvPSdje+
r7R9Rnc7Gw3Vi7Fb+1hq9B1kalM1pWzPIz3Aib8cNgoiRaXmCChy3QEEEuDx5ED+sRHdURnhkUhH
DXomTuxcvJrtunZrTXRXFXO8n8dKPa+mm7GT7y7Zh/UUFRxHAL5hJRsInfFxfeCrOpb37Z+5322w
W/KCPVAEObZzEb+uBZG/UUoMyPQA/GyRRUuuS2U+SNahYxAPpG7HKis+YDeDWMefb+06b2YJxjuw
6tExGZ3oxvaAfJP/qryoBY8yupFg4I4L1ZV7k4INe7vtzqVck6OF1Ou8sDzGpwMiS9FmW9dKRhU8
0ZHvJ9IYjjr4quUvW7pj9wUMlP7zDKbr/Wd8p1bKNbipGHwQJIez7/29SdTL2ZPncjNjcLF9SUzq
zwCnOdAliEOakjWY/6MjQW7JyQF6Wu1lQTPjXGJeaCVhfvWlxUcV2B+LOfKE7pkh9RmKgrxdsLry
+z36pBivkOGIarGccupy1gsnbCEuMljmf8GxD8+kpR6OCbSTppjDXs9yfOfYvkncGYabNHZ8175x
G1YthXC4KUWo5Zh3fZK4p7kHbt/M0IA/cGKNv5jLlHVX4INUG07myXq01ay5CFnIr83m+YRSmY/U
nueQAzSSTUZhxOKfRFwqL+7LI1zjFF4ftJ8TLecdg612LLUWKnwy44Nh9rDDxv/WB3t0+giue6YK
n6C1PYbftG7m6yo7pTCV3CrzlhwqmwxRtbtye8Bp1FzaX5Bci/BUzcedatzdqf3ubnoaUKZKsC8J
/qusuZWWhp90vp89XzuHIpdiDmyOK8xVHlNbofFBLS2TAfN7bcywYgg5+3F3tcleSlIhQD7mjh0B
7rW69gqk0GpaKTJ/z2tj3b1DBkwYt2nKZ87ubDKOkrSbOL0mpZF/qfx6Hezzap54oLFvH1TwFYwv
bTvdshS87y62cAZ1xwDtRjng6Y39cEuVmhZ7dAFZrrDLDdinwIZavNZ2Z8qgXLtXCaQg2OgKZjFu
xpIK5liW2zXxvAU8+gz1LvfDofdVz0msrr1/L72Xh1C8kOMwuayfDXEqKurwS4TdN+oY8xtCIYYY
g2eAucpCS73rIxxrtblNeflWAnFPbN6I7bH+6R0tc5Xlk7YomBT80WHICWjRf1WbNvFVzMs1BAqT
bKhSkefU7cPKuJEakF/dRUFjbaIgEGXQXWWI7cC6p8fu99UiEoFJWBqwUJza07xYHBrr3oTd4eUH
uWNkhN7sUxyxBs63RnDeV+64r4CA/kK9Qas/roDmpbWwuoQg/QcD7XP8WWM4TKVr0bpNyqpoovsI
f/n93dKOHtfiwBz5s0RlistrdrxCheeTUUQHV/7KCvjS63IbEWjJRqIqxciYP5tl4le09rL64h6J
zmrotcYjfDx+nB73wGLMfd/Aoqr3c3aD0GFQ0rvD9D1jJxpP90FkdDfVpb+8Hqx5wQ4HbkSX7VWy
CEblMCbtRsLJLFxqRWBo1e1UOsKEj5zl2vTkJZqnXw7FDVtDXvX/5uXarfdqm9nf2JORkhhkdJoh
Kq9TmTFja5cxV5tJNj8klmospamZShA4huY0KJ56Tg9SFcbce0d6936vUENBagFtOp+hKMQvaDk7
oKWGltBewQKQoriu+EANPbcby1kw0x7WkhyW+BR23JW7uxoEo5cirKggt4mEe343whorlFEoAioj
I2wNUudHacbF8qnOGTj8hboOP6vm99rpDhW58bJqF11gIoXRcEVUpIW6MgGI6NwkSUZPNWjAUoYg
i0Ve5z1j+qxSeH6/uq6LRYfS4MNWC96SXgLLCGeKFcQpgWcrb5XWB/Jb5xLpNpkRYIbOZHnHeBrp
eipgmeWMxyoMfckZjv4OPD5S8boAgsxVwsMwEe92iHl3VFEj6Ok04TCpHIKMb48QNLSBAE+kH67O
8xT3Rjf3EJoyfIbtmCH1a8MA89SgifYndCDVoZtSo7ja8Z6N6WBszA6fkipZ59ZSedg/x+TRaDae
jMFe3LQJQy3sAcNHpou7WOHEnZIFsazdQZRp+4ez5mbKhQf8SvWnFVSdBYx/vj2H/OQy+XdDHp6e
XFb6wWBPlHA8XyI2wXpw8mmdIxvHwJPZ2r02qjwqk/xeObLUuMDVE93GNmhUf2q0cz8sW41/3AER
hQZO1YeBKPsZ4i/OL9eXJ56IXQbpCRByd7YtXN63UvN5s6v6yvxoI/MrXs00ZrGKwG1e+DSNoKpy
S0yFYsq0Tlw7segj+htZR9RWojcvMythnWxuVfJV8DIsl0bwkC9XIVNRlE3wlIFCjPBV9BhBd4Uc
7D1NfkugbYUZPNgbDm9WObF1XZG6iYPUjuL8nOfCs128IcJo9wvxVgCX/MThX/K3hQCHj+kvi3WA
C4ZFF5N8mPDAJsheSONbQr8Fu3XuYQvRiSJcAyEqTTrpFho4QjZ6BWUeS6BN5RsKM9yN+Gc+pWE/
zouk3mOCotGR7kR1VkddI9kNZGBSy5zx3YTQx0XCPGJN/rJbpTmFgvdshIb869llnqoMxer3rW3Z
XokAGhW9ERO/YZciGYarPKe/4rFwtrzPRfjALyh3JC6eVoVE/WuQNXre/f4GiivGTZ+Nl7H+6hlS
zIvz5SDPKNiSHcRri35MkWhfafGugllKvIga7yLTEbEXly0vdrwhKSo7jDCXE+XnKlLUK+zPhnQd
gyGKfx7a8CYeIQYVL2/+0xSd35H4xWDS6Qj3A/aIeHBxluDB5hV0p19u1zMSVJ451Q9/srhhRo0D
6GPkR9zUB1vHWX5WDdt3vwtUgdT461aBxe8DE6mrCSzxZeGtW8MYzecyhHsAIgQ2SmKX85hgC8Bh
PUMIZ/Lqey/PfO37/cToCxFQb1uKsvPFbdOIkTOZdfAGiQ2Xp4vkN0iCP8vaZr+llm3FUQRvM1PX
Bj7UhhRUdrD/BuatAS/aIQ0/8XU+h4MGI0mlhZssNIgl90G7oH7WZhpjzB5qv4ncTfTd4r/rfUAD
P7eMSK2NmKnsjCT5w1llrtGc7YG3GMLURJwKY6GrWR6NcJMLRUXIXf3u0FSvo6mS48H0nIg5ocSX
VYV6zjTblDonaUonKwTFKHy/tAs/tOB3c8BG185BQbZhHiQMW4d8lB2WkMbbtyl6jJDSZz4lK4Qp
d7NLaC/J8IMe8Y5Nz8V3Noy7BxDKB8+eco84JtKck0XcUxH2kZmq3t9waRAyXiVJHHJOYkqDtI3g
LYjUsMAswY+gDNa8s/nRwURD2VwXxRjjNcC38v4V6QSVVyLs57X71bi1HIGmzqNJWkdm/Vxgv3hO
2gcp6tZFzX/MzUAR3ObckgpZzAiesGsLXeOabdQUCLvwSX/ZICoiG9YXIdQpyxXueF7Xx23eiVf0
jMhiiALErh1fTuFKRYQPxMT+lFbk2sbbjA7YyOX65VCGjIgz4FcEr4YvNLg0SgPalqo/9RgXudQF
gBXls2WpB5zIl5AaT3N8ZzgT96T7R5fh08jSgkYTb2v/nLcy5l35hTtS5Wgup/WHWeQNc6CKYkmy
kg15ERliRaVMB8VhYMVYUbYCdX73bAuzz0gUko8O1ultyy/MiBrvDyPqyOONvbpdto/dIndK6wzO
4VFeiYIQC9bZVXe/gN01+yF8Aj+ulMZ9Zr0o6sIcGypeXhjfmTLq8/qNnnVElNoih8IoyBP338Jx
KTUQqeIP/QfXr7jkXsVAk4NgQ5Jq4xt5p+cHVV55FhQUfQPZe8FUTYWSlSKtt+pu/7l+cb0khYez
x6N1hjsYI2zEOqOd95xwtxut03MNBPQ/57vzWYE632ygf8CAGEIX2ivoYQNurdJJ3Mr0Q6BpoEKj
bPsNiS2k5wd4JWL8J/WwP6sKqWsVzxx+Mx56uDM+iFZyD6Us3T7Ez9DR7vIdkYRFsd6S+ZGO7tAw
9afmD64u/QEcfm2PmsffvKJnDOeJwvvq0KUz0bfwgni8SL3wGbNUZtUyUjIl9Vy740SFgww3mAoR
eFPIoJi1DNoBCJo0OjtCgeXVOdwtBOrM2rXH9rygisr9ToUlvkrcIILmZuXfFYWZg2ACweV+oVn6
tH5+Mps8j0dAvJHqxV4vyaFevvTWkfI37dHQ1QXVs1TcmcQ57BS7swcHISniCR6IfyullMEfJC7l
CoOEKkU9CE1BjaPtH/2tpR9jw/LRkcDJVnjfsYznr1snlHvmz+kx6JA4EmnPUSNFwQwraIosmwrh
HGVzuJZ0Mmm4SPxV4Lbj/ahvALSowPYPGLJdX2mw0+fHbx/QjjoBJ3yZM5MvZYneK2KcRdN/5yGd
ucNCyzV3bJ527NKdIu4SnpKkwi/VhDuGahoxgYXKISyC8LvBWkyvRr1nLLA0gYjZf7HRxfi54XBH
vfDs/p4TVJvSUxb18rIS9SAR/O3u8o9ap114GpCEah1Td5AbVPyx0LeCJani67etEH7XsnZ66T0c
3DGSYzKJn2rtsaLrUrBczP5epACSw8iRaYw7Tj1Olk9nfJ+Vxun1QRPy0bsGL6K0PFLEAm6mBO0+
QYTikPYvkDmMBuKyAFQzQ8C6dYnH8FgVLHYGuGnyOCoyzg5TE4c0i+Yilx4pI3k+/oC8aPOhwQ8H
+1NiC6KPr/x7WxN7z1WRvJJllPbnA9WkpEf/z+rT4eVQfrW2GLc/2mzpdeiF6+avyxVbcH2cpedD
nAyknHqOj6a1urBgUCO4/Uf4Xut61nA15CHO4l0f7aulI4zKn/22D8z2ajM5c23GP2A9WJYrHVlJ
8+2XLA0xiwckfwzN93MJO5wTX1CqzvUVyotiyzPWgrD267M9OVmfAu0CJ1WgLxULAIUwykvMTEAg
wZYTzbf1ryNKwXXeGDrWnTBTSMzO8ofzvIKm0B4+a9Lv5+Y5FYyRlNjdQG2K5qHi7dDPEjXx1Hnh
3qrqUfz3wAnFGlDQfWPdhiXaniG8MNIQGq80ZJ09q3Xi7rp4xdASdoO800zFihzdHqX2kEag4fTl
N0WGrPJy6ppalHwaHxjko/P25bjUHG6p0plxcDhJxnA4dB8FrSG7Adgvby9pjkDJq2sMtGY/LveR
2y6ViqKDyzCtBmf0kPlhSd7CN/jkAg0nRJEtJuRruzzCOni5qSsvicvjGMhq3BKubGmgqwn0YMdg
LD1N0t//q2ycMv6XIgoH7RD4fp9cNLCdqztyQBzRV3jGM8rJJF4DHLwrK9ewC5zPm3S6NQay7Mn2
Dxz6iUt03CjAZ04iI/QWSvQQkplcdOYM+OnIEDhTyiU/AOTWPM6D7Oz6amMF1wSRmDcyXEuVWCJG
z1VM9T+Li376G4IEgOdmMBRxW1kzofYbloq1JSIjcKhzxetLqaZLVUPj1yOGVkLbhwrZ0Q7a7k15
qwA0AbArWSm4TuijelDD+osQXi9ee1z9DHu567KGRjbjYdw7ZKAKDYhB8+ivzTnSAe5odZCmt219
KNfjFdsLyjByxagKTEajhqZ9RisY7je1Ljy61HvfnLOaUZ8BXgFK8GO7h0haH4RHPwkSl/awDZPO
K3728LehChfHE9Jpb3H/3swCGrcqAtxc4nZ4wWE06HYKduEwzavKIf1Ib3sO5ZApvTzrgA8i1Giv
w8WTP0lQecEdYfK6y3gydKB56ISZTDdd2EPoqsZsud+ihQ+TieTiTo4wHCz9W6I2jDwKahiqO5Fz
8GK7WPuWPRkYL8YZEorKX+0kJuHU09+uqKMF78ONkWVtLMx+T8hYyh2dea0S6SdgT3mHSKGwSm58
PBKOJZEmvh4WoeEdsbbeXauDFiFhi8/2G0vDH8dtP/zEEiEvBTWgLs52MpZzwzy1OTi7Ebkv95Xw
TzQiYGjFTw4I/IEqAXWPOyrT5WrU2q9dhIBuvV7Bn573E1pbPgAJO5J6pSYPOSjqBxfIZxE7dgkN
IdrVlis6P3svsRYmDnIZvTXwinA/3WHbDvfo8/KzLlylr7bcfqSxKCg/yr3anUalafOh+mKD4VXs
VosIqBbUYBWdSreE/Kk1UVihDf7PMiOpw26XX3X2RBwssVVlki+7laNHh/yFgW2bglMaaJcc8qZ+
MqgYz+7Ew73WeLeaMH5vJxyejyv1NuBMxvIDnN9TD4cW4ER9RWURLtnPT7qfRdqHhOhUUv/faoqi
fOp2JI105h4vTkyQezb1rZYO372bOpAdztCi+MdzkQVzpsaGqxQ2oJLC7NDhQoeeEqlSKnRslEvC
5R8a8qxrq0ScxoCkFVvbCI4QdE382A+7h3/YLO2KipQSeycM1Qwzd5+8uPQ6TX0+vPZwYOc+Uk9l
Ofka2zumOTIkg4lqJqYk8IGAhnIefeINLYrezgQaQRqTpGov2n05gmYh+NmIMqXbxL1bdTHbWpee
Xx9JaMacz1QA3mTovYW63vEt6Zt5uINi+M+lmxc4DaJJHBhqhcAMnb9Y4nbUQqYBrw0RnZvWaiV0
4pKab6TBqnPOLdQsfY5GesRtxplA0Ikk1dlMYhRUupt9V1EK4/Zij3gzy9H7KXFiJQk2KUeqQfjv
SyPysisqcFH57EauTbRWKzG9ANbOc6ppdkIGzp8KFN7OARHAmXLnRIkuVs+FUu8q6hDSbOtbpKD5
nG2uKonwouW3I8QytyRDJXj+Kh0BJJobBLvgdIb45A169yzY9bf1RWWpJrPOAJFd+wPNJ4X/eQ6j
pWwU6Nv/4AVkpPRAUQeu4I96oJgPDdsTagzbFk/OOT+EcppeRmGlEyWaNMsyKyzuLkBD0fYkd9r1
oD4XaQh/LZbERYOMHsHiUVOcgCN0vMwSu5fjPS2MrJ6GDmJRclc7xnl0i1/R3P5SXIUnSr9o9zqK
bRwUnWFPY1E3b4reiTa4EiviuZMrOa9X0i4OvNQB9LbDdVJZg8VaWuY5giFRyr297ZDXoGBVWlPx
zotWJv46ycjtLUtQ0CTJ9KjiI/ecnGCOXc/zStpB7Q8U1sSeAI4DMvlIUUzmfdWY8KIq7M+n8/Do
S3EqdVd199ECP+qZUGpKMzcsRNFxTaX+xjuwRNFx4XnPyFVFs1S6wEOGhtdJx7VHmVEDbt7JSgUa
qhvPf9LPXlb+PQAX0/zA0vvvHzviuYLhz1VhtzQRwk4MD4Pm9ttkqAUzF7d4uSnG/saM2yyOHRB0
23PVAvfF/1qeh0kZbfyVUrRe5b+6fYCCpwrJrL4idj63DS46bqNpTIeP8exoNoqwyClwFoiS3TOP
zmsNDbzfwHfSb8+k9DRMtyKBWWI/JtqWvcPjzWWUdS8aARZ1Bj+mDcHRffLtJ8rgxfIqlyT6D0oU
fLApvrqOJumTLtO98qvppZMqXW5LNeM4fS21rXVF+eFGs/q1wupBscHL12XyzDkt3zLZRjRQPfCP
6dv3frfNMJ7+V491xdAT2MCXQEC4u7/3v/efuhAUhp0wQjZjRc1KWck33uaF4qK/kZln/iGxKv3B
FyQ7CQT+JS5oR7QaB10YjczQGMRPtWb873n09jgV4yypQ8w09nokujruRwIsI0zp2mgEd6DhBX1V
W6BhqoVgAfIWOokwMhCvHElZElMi/h3ddorzwDAx7q6hpO54qmz9wBJRQnMm57i25U98W8nrl7RO
ozsxW1woRMHyw8jOzN2VEQkp6sGj4TAGbCavpONyuCSawABI+8vyEy68W+9sb41+aSstZpG5BtGR
M+zEM0v1dRyHh/JIgJ+ktJAtyVz2rhfsrAjA+fhj0VNE/KMKoV/9c5DeSvofUln+eujEx2+QMWco
iv3lzRcPabAbEatArnMPthziNjeawV5henGXKa1LXfeCvNwIqvsSiWesHu7LZrdgeezdtA07OLF3
kLQICh2ncIOrLwtr45RjcXd73e8md4a90P9itWwjR1e047NVq57M8qwNQhKbLA73GUZj8xQwImOm
F/UZAx9l3hh+jLt3ta9szNEWLrTMeyUii2tMWryu8qsru8M3LZ+slG17LaFEEELce1rWig4fgle0
ZJL/5MaRbW+kRIgB+jeF9lPeaBHzDUc3p3ejeLn65tlq60ONBN84e7mc0FyX4e89Ts3QRBKEjDBj
aD2YVy3VlxyjsMseCE28uTILpUpzXNZATtFdFDbJLTh5x+czKyDi2YBdxd0lki4MaxJhh4AV7pyz
OouWB5AYRsLi0AjOyoNCYpYS6jC9zgNH8iHP09RUXWo+padn89P0BujYRaiIKoLJFT8w55lRGdUQ
j0n2EqxO1Qa6cY3I3NzlkohSO+NNCxN3XcfBKieGRbqDNvJin7KXWe0c/IzkqmQ7QOa8I7EfZFlH
sv6KBowoz0HoVXJROTCu2DXmaqg8XX7tijgLP9DG2/lY1sCueTSsxy8FxDzJ2PFGKFjFTQBldNS6
+JG6BY9RsqjWTS1ane2aTYn9z1pPPzR+YCuMe5n/rHbT+wcOaDMubwJjtklb8uIn4gU7If73kSzi
WiuQyUsgMVynZvZc6RZtrtTP08Gjn5YXSf7m7IKfE5AQ+oka980CXov9tagronaDl59pTN5ARIAb
PmNnCqvCOjE/jALxm3JUsVqvx8N1BTmSlxmL95XNL15CWzyTDQMHdZWvr/vxeOY0Du9MSwPbf4Ov
PsLKE1RcE2cYqGsRuJrLeNEPIRyuGOwBVeAZKfo1p6O8jAGn8y93FxRU1vBgfHEdRRVQabDOkneY
GsFCbBgVzXubFZC9diM6YteNPg8Q590aEVozAmR/dO+6Mpu69SAK/le0iPVgKIDuV84Isx0RiCmb
LxFoPAZw1D+bj2SrHd8F5Cv309Jhq+O+uz3GzftptCjJF0u60fr8hnV/6C5u9Wd3lKpTTHDO4JG1
1EK3oiwWJhBqeyBjtWplYWIK9muAHw3gb/ICgbc1MveDDgVz7151qAktLpofyfD3Ug1TpG/nZnge
zbyOp+R6is08uHyoyIiUO3SRVibuF+blhDn4EW/lYsB2HmbnXQTtX+2Vm91fuaUdCEikU1ap+pU7
D8cLaudsTWZeYjRf8NpSGBzqdMsR4MnHNFwnK8igGYDvtagpQnOgrVSfRBQpaf0X+oXmpotQMiK9
TrTzjguslCK/8jhEQWsZP7srLWEx32TOKvQfJAoxMUZzyx/loKgf2cmIGhaL+HQEWi1Z7hsz+TVm
J4Kq76Va2rZTyCo4XZhRRPjv3a0FXXQxirQ4I7xMlRtdjfvuUc8R6z8/vhqte1GZrVJrE1LJs5Q6
2GsN/Tzie09mpMwUrgPNWNY3smW/orOqRfIh9LuNeN4vFS8TFMXlKA+OlSyQnN26yq52+rieSfy+
8tpA6BnlRu5Ke8HaVZNirUNaL7HIk7j+CmZ0YbNH5/Tl6esK/W6O79C/vyOdBfPsB+HYxhyfNZF4
SWeU5AVkX831z7wm0p0BLFjDm5WnnYa+60TzSAdfcit5AmIKWg0CF8uyqQXKzEDaVPfJ4cQfA6ZP
E5yzSqK3kDjXmKuI06RYuE4BgueDWUsQ33T2U1KSgRtm+qGQHt1/W+dUwcY43wOhnAMuJ3MJqk6i
jT/k5wLxl8mWpNqz1J9WRHdYwTq48pF4JEYQPvOyr2//QBDgdk6jiOtAs84oz7Oi5A/AZvlV1Hvu
hZRiG4h/vbhYUKu2mtHQjeRFeHGZocavMLJJKjjZLs5dsXFTywiUkw1Bt/7zK9ll4i+ZNxZVH7E8
p8q5tTXfqx0SPAhCwHY0+fCD1R2duqpOU27pbb/ACTyy1GBbnzY4vgCq3C2sUTiCXPiB9DwBaR8p
lVtvaTkzjkAhhu2lonEcFjtdfgAuggWcGmhB1ewh+suaE7rnOpJoOKtrROdH4ORaqfxCCPx5MWfh
ttjnhnJcntux+DerKxaapsXQ9FY5PlVipH+dJ+Wr/l7NZDDsn7A6ZiqjSr+KfbZYoSO3ar8UPm0r
ea5Ehcb9ChAdx+OhmyOveSHwrrsFSc5kDq90nRLJIuMpCKqotNwpxqKheiA9b62arFFfGhJMsFKy
9XsmePImu5Rk4lOQFP7iiJcFxBBqIJ+updpCGFzld4/+K8x/yLf63WO1k6wA/nmDH15YDPoBnEv8
O7rJE16EE8rDlNHasyoNqYtGorhQYGZ9qarfXNdSFzbQrAeAAwHPMblWwAGFHuxOofbZ1rldT8dn
axeZo6uzkQ64VE5SSNsuhn7FnmPDIZ2BJ6QHFvRpJtnwzQI1/OEn/sW4VcljfKyX1bZcdH4Ex9YG
NCiG4gqMsRKA+PAvK+LAJ9tEnnjgfVWcH71gKQOMJTSjdKxldQjIBEhUXL8D8oM/PgOEa6PzxQKg
e8MT6hKeVWjObdidnGVynWB7QoQRCx9QH8zHTFkjZE2TG30gxXX34MK2jXh3/AgDhT9b3nn0RnA7
M/beQ/VkTw8dlSyTXpjaTBCIKVkOKxW4O0Py35JYeaxhZD4CHCGeUff2yCGJFQ8nDMgKduIbFOdv
SWLZPlwxaTDg+9MjYPimdeqOfWBNhIbn1agEA1vHKVX1C/MGYKkZLml2+iGoI5rxsQPPanvw9dJP
d9v0JI/xqcmCaegBqGoMploCBXiLvpc/nQY+58c7DXSgYklWoVfujLw6GkwugXKupXPoizcXRrlR
z64lEOF0XXsx7I2LAklfGBZqI+Bhr9r0e+9foHtWeyYdH/KzLQ76cBHRiW7FZYDcsyvLr7OrE3qO
WIBpaeciY2eWivWOesVBLSsTYB64b+OHyylLJWTCM2O0p2oJKwybMFRIf6RgoJdTfrviWQU0AxP4
HJcuYD06L2dmbKrSbaVMrtjYZ2Di9se982c++MsPap2TL23zu4JZC9eSgR7JjXt+2DmmOiL23PsE
LnhI//z3UkhTEneJngnNXD0KDy2eR6zrwiaPC5uayYQMVS7rLIkIcjxlM5Lz8ZiULMqEH4ZW/M5N
BqlGZ8jddx2S/spApL5UjVBJUAP/h4r7/kO2pdZV4z5u9gc8UqPRYBRa5cJG9n4F4yy+kyHKaTRd
i2KhDLVNLi2UMKhgarvfVzz+tVpwLDjgmYk+tspLcAZNxXUVUxXjVyMzkM2VIJwye4NJnwmjmecQ
nR0JWJWeOe4Ssqr33XwcOqkDKvnkiztl3nMqzFrOoxE9WA5KbeYbv0Le+W3sWOkuBB10w2aO88oF
pL6HfjRYEhck9ho3G8JX6L5osF0Dp+iRJhU7eN7LV5KXnIrWjj9kN7IEMIqS6xcKVSwNLQJqyg9u
VnD0ysDkdnOBNQM0nOtf0W7/YL3DovsXUKdnCfS76IMZSRWtr0E1C7/hzW8Ap/hJXNLS+8t5yv9T
QnSPqtArvIt+EMV2x4WVGw0l/PsTcdvFO52F5t723u8qKE5lZ9HFn4kGzXzf23byZIt7CVif0A04
GT6++59Hrsz1EbKie5+W4UtzQIE5XNEyUzouOlnoNWcV44B5qVx4OcaClDmQI6aLoOzSO/8xZ6eZ
fr3XG1M1Ku/e+a8S8uDllfkpWiaiOAErv7gOsOqHEJZ5fzD20SminC5Y+vZKNvEr9k7J9KVyDb5/
OcSE15tbC/+Q+Xn9Hu9+oFJnUmRxOsShiAUbAqMai3VhflmqAchSARVQlkM6F3pdrSJvos+TdFA7
gSjhmzHrDBftOSBp3BpA4aOb9pwpIPX3SjtiBZZ6olUbcldPNUK7e7ABL9MMoYzrUTrFdj22azXx
87xXRcI9283/vAOCPdXXuta/tp6CZXkKui3akrOHgl2JVxgmh9hMQC4V2o4OKQo1hNymaYdDaRld
F5948a+SHTzeLYITWXtPZlQET5eFhLNnaE/uur07N3e68Sc6+8unrSN55C7aCU+7oqPCmlCarpFc
gSIlztHu7BGC1/qReaAz3HyJwoj7sVgE1x5kYmaJL2qP/b9ylJISo7x+PMDzrSK6iHJ61JryJkGd
39PszyF30P4rRKNnt2tumEgDpuVMiK7TgaQjVSVFiK1iLvCkY4eAXD2dkXXokXlxcJPjpmCBnf1J
oy5KM7G+jjHtxBaiNEV6SjXOBNtsqGBsJuwQJ7CCAV3pA9cLgSTuNJu+wPwreBM2KxKZrxiSa61D
GyKLUXdkCJ2zbf8qIFApbPYTef8g2Au/a2lskBXERCkeXk8sQyaSVREW5Vc8qmzU7H/7X1ZlTkgD
DClHknvoAblSe6RQP6yFzK/sNjnj8w5fzfRhffTMLR9aXgQLbf9e5v3QYr0bQn66zYr72NhLMOG1
/XH8PlL2u3mUGOyEOv5Je9mS9tgvFXtPbLfvZ0KmNCAwPNU3cZ2l66V3VOb7PD/QOeN0m2zZx0C5
0tc5vG+4mJBKakoiCa3zHOthE4qckHGmVjTLhlyQ8DaHpKwzkOAXOfwnC2vUxdL/zecccQZZH5TD
Q1NtpxDFBNtLi5FXBGgvv1qqS7+8VZyQAuEMj9T3b411OUk/MNcNXIWafwFAcynssv2hK6iCSoxW
ulJq4gZZGzuPy+NadKcB1xDOPkexYYQFKNNugAQDTftYn5//W2qo1AjjYIfY2HVsnQFRjc8NuyeZ
um8lJ7FFT7VsTQKxEufCHa7vQY7mmmGkwcby+gsrKIOaAVUNxLqUhjmA6+8oU8ScdezPc89jT1ol
Qs30hi8wL+6t8Drwf+4dquKzQaQvZFvWkCOlAszcemo6fjmasD5lrpkpaUAEltxnJtYG57v0XMYz
xiEWVmADTNj3+pkncCS7P2HklVvpwdUXBbR1D3XB0eXnSTJbVBI9Xc+JHkWRIisACNgkHwdgiJVd
DqNxqkjovgE4EnwV7YlTHH8l1BQTcLpZx2WxluO69EYWIlRekB128pPPsqKo9wF1YOxwDNDOmdkZ
GP3oT9LD3+iCZgBK8nuxA7pOd2qq9HbjoL2QlP/p1j83ATKcfbn9Fa6mQmMgxZe+yTvqiOjCF7QL
24gY9CD1wrhTPTY739icKq+QdJQvm2Ec9xYDzZ3YgqvmyJp8QIbm3cdoTNQ91JCHsfOpQ9KC+X4h
V5EEs0uUq7clGnb6xU6O+VFyNPnJlr/jfjVkSVjtH2aLZjsokfN/M3aNE63cSwGH6PLYhtAXgNOs
/DlL9Xp/AXmFHyeXeZf6Dp2VNzf+FGrrtDDqNp5W5ua4G6Buty4c7JdzWRk6u30rSAjL9K2KEqtm
ZcPxlDqVf22fa45qcuADRI3AcnnQsGX04lW56XLgmEY/14zDgdyBwp59F865jBASVl7AWV47Zmun
mXN0SOnkGWAChgof8peC3ULr/NV4vg1v5SiVqfdp4raB7A4YXw/RVZgrsgaIW87b7wm5Yq4RIJzq
fhJ9L7vDNU6QAcuDtfOglya4TbsShqHxIjN8qgVZBXBU07anNUYzUy1DXNCRzDzoGV6cD88woocs
7TmkSIGnREA3WU0FxgJfevWix4o7P60VS1mBS+UZnvc+b3EhJS9u6+E/fyQwsLHgkNE8jgB7ch05
5HR/ImK2QNbFAwQD00P922bpEvYl7iUxBSm4CFvLaSjq13+JxPw4ifF7N2AVXpoznGRHFiX/S/Ca
ZniD0V21FGwoVPwvE2/42Qn4KO3AoLjm9NcIyTmlDTVesVcj9UItwHWPhcAghT+/o7opMxLCQghP
wX2vBR72PX026dY7TEICIe2waU7YBwJreQl65Z2Z4NmCn1/B5+GrQQ+OXmsG2RSMlORfP/9Ja0CU
U76p23+w8i7ZWFZNszRMraHyAZGR/5B4fCDXbup+Hw8JAa6izWtkpdwdms92z5krZGN7z/vG/H56
NrznONgD8rkni2GbEhrR+oC18ZhWJpJFuVzlkcTPWb24EtuLOQFUjTEdtJBJ4Ou67Lh7gPAQnWXe
87N/3zFrySBYcySjOKeyhKsPCWqtLCm9JIKs7JmQ+eTP7Mvabc2LnQND9VhdP79DElZILqtHZLay
ADX8t9Pl6GL76a8PfFcL0BsZ6GqsC1zPShoWgXBrYFi0Nt7mQMKRIp68DdE3yolgwCZZyr6hK39m
w7Fl7c+eqwkowOE2f+LbAsmhyCh98Zom8jL7g77oGZ06Ivw9RI7Ncjapo5cWhbPXKEOccT2fBBM4
GV1RptybVSyRjWI1yq1mejTiCyrQCyH3U8BE1BivWbvwgkuR0XhYUuDaJzIEV8jwsYkWOWc6B3mo
atCxRYTwHIRj2IljHxiMfq3Wjjzj9d+kUqUplHEz3mOOt022PWUdotrX5QGudqeyk+vgArRpUDix
sFJFoZwbXc1YoAG7L/UjLTQCdLVgWKzTXPjPv39ezgbyZL6gmgrIKFj04StYqyVJVm13G0cRPuxJ
5EuYUvjUJIi9fZtpAGgsfeVobM+L/TcNMARua2th5PwsdSp5SRuoZUpQ7SEKjw3/Qno47CaiqO64
5sqFfNVP3yXeuvtWO4cjZKJg/1wQ696xVhAZjm/SKxdWfTZWAB6Tueo1Q3YaEByxPOIswwmsITPJ
i1xn3PvuHXQCLKFhPaBTco99pcAXzXW2eH9TrVjm8pJj1cCXs63tz+i6Y0VGh4ea4p8eG++3iu2F
pHEyQC8q9rblCrBxYINeUYrWFcQlyY4D1cfbH9/JAQMqqFZNP3dnJNgIP2ui5RcuSrHGonzKgGO1
qkgYQsqhOoToqx2YnT9bfuyg5/AudX1UMoPJyzQ3/eI5VDj0xGpBDJl5rI/W+l6XW9b1vW47+A2g
uBJszqs+Xsst7AYByakBuFkfiXEhz9nKm9KvuK2k/CrrxQfgFAN5Wz9fBiXaMyJfZrkzojqOjHWa
JvQnChnaYsyTmRcVHaKvicwO5aTCZW7a8yTRy9ece4zeCakkA850z0RDHdhQ3dhuK60xFmk8R2V4
3yaFsO7kh0fticZ+0AFdF6zZT0Q9soKiyxxvtojxJs9w4J0wpFqDRlrlJKM43P69jPKE4VowkPiY
0CZ/GORkNgdTYAhTOn6cm75zOD2fnpF1TuZWNrV01h5khI4oWgvik5SGfFsYa53m61FzXA1Dtt8H
bOApna6zBxzXxzsc623u5k1m/bO5YMioOrJVm/QZR5q9ocaGCWH3DI3OiMBzzWEZv33yL/psczdX
mu4py288pqBTYXtJCVz2gAMVwAWGutY32a8Vk/UdgESUAEUdF5bh7uZ6JyX0EVSKxZvEf/3Z1slc
t8wRB+ooYclRUvroFlgxdHUMDOV9068pyhI7R5XaJUTXqkKesPGz3EyTY5VdUKoWzfK7Y8jwzxKD
H3j7BPXuY0iVKw6kTqdrqWqyzL15pKcn/yQBj6RavEn18ZoVsCiMV1v5vDdBYd04kfLHbMdkXPo8
sysXXVyGo/00cKlEuunqjJreKrpTD3iCxQ+jQiD6An/YV8p461ZcyzkW8AOqueBsfLbwBUu1tcJR
4f1Q84V6AN7rqW9p08PhWpE93N6RRfw07iB7B/8+Hysep9pCf4juoeDG2VIjXkwnSF9mokn+ZXjH
IhJQBgflVpchh0N9aopvY3sDS9EM2x6gbTLl63Zb54Spq+iC2AeABTd2rPiMF1cyWrIxl3bD9gc6
UyGRip9tAyV3KCeaNelMZvy9OYqRSYzqJ7yYrk6hy/kqMA97iruEFazy/jHrJvjoXrRpLYPzYjwo
+ekh47dwBkj/hjeb5CH3I3D7qVnUBRHSDK3eYVEbUHZsGGDhR5IL7nOEzIhFM84lyCtUDUKHaZzA
7ycw+qqTfkmEqpxbQ4eNWt9qKGZKTj6/V3Bvi+59E9J92LaDnJuvtYWrX6hDKtd3fD0B0lgXE7+m
B6kKdL0K29MMeKeBqvrCg+kJP0gN21HTCw22dQGzxogOEAyvl7SZ2NrMnOhp+1k469N5B4f+XD1A
ok7W1/B64s2NM9/L1HPrPDllKMolNfXWdZp1hW8Zu0hdL85zF9fVi9tzMsjeI7kzg7x4Y8ef/JIP
1G0BSLAOuSmTMWgB+FnhZBwTL+xIYk/LrT/UCroT5Ew6NEZ6BVXMJH7x8kqQz5kX5a0xEpaDq/Fn
65EJ+YFE7ES90WsAAWVMeiMdeoKWANW4CnxEFQsUQWfAdS1tN1aTsUNwK25dQEO8r6UeSKpp29JP
TVCvS8AXQe4n3hN5QuBSKCYTwPXO1i29JQCCB7ozuyMnlXSDxtH2YFBcrFHBsXnY6xJskPSgmIaj
HUXkHNvBQQeKGTbMxpio8+mt8q6E+vI6IpQzDICimhcQ4u5I65QjzxkYZap7i/eF0DN5ramlUUWc
3mkvoWyA+0b9vh5uAOszc+QZaIX8gpeh67b9/d10ycWkiSR+DV2WeFyPe9ySmqXpY8NGsS2HamMH
/EMUByebAJPr7vu4xHGNPeUZCbaFhmk6NN60PmcfHbmalX6TaNpb5yvuiUbaobZLL0xCWU1gSveL
ytqAjAE+wv/kN0pTMXhEqlKZtKxd6xs2PmwcncxZN71W9VjWaNVNh1XuaFymEYu9puF5BhkIWP/z
IEJA0ed1k3O5zgQK+ZOks/Q2RWbGGoT+5F6rJxVeYZK/R4iJwUGUVVa1sx/oi5TML771vKZRdBgI
Lb6WKgVZAoYHQ2FpNa1C14adjRwnci0JdnB3BKV0yql0Nw+zaJuB0nyuhKHKrRb9a//LS7TKgfPZ
BsnWJDOwd8sMqTE8f8NsnazT7RQ8ov/uIjVKqqp751FNFuyb559/ht5o5QHhbNuxlIt4BdILlvW7
r/5JcFhCp2exR+oTqJcm+GGVycfKJansOeVSM6DQv9MOXu7swNcPeR9TvmcN2YvdEyuDNucjDAtm
ee+UPvmGAObG9jBOcmkP+q9Eppm1E3ag75lUuJ81Ep1R0rZuwaQvFZCjlrtkAtz/LPmF/GJHETEt
qltw0PELwn8x5zkgOcU4dDTMB1xqq6Dcrkz/kZAA/2i2wsJwlTbXGiGUTXFwrPay1VjaRWLEX5ti
U9Fub+k1ZqONbA/i9yl2b8RevEVvlW67j0K1+Bebixjm835VMMib0Fm9NL9b77BCeHnVW8wC5Ojg
G6mM+cdUWYfzJLnV5ndMf5wIqmLD027USbMAPyvFk5PKZAY5hw22Mx50U9IqKY2BK2Am5vyh+M1u
g8elAui5RQwBlwdYDccwob4I9O6IJwbTeaDbNn1zln1Z5gF6wI3u9mYTpLsvE64sYdSiTgkFR1Ja
OoehRBDtIOkrpzXjP4Pui3eI8G1CMeFzEP+GEdc/uSvEk05HQ+gPphjnqpNcJlkXPoN6UaO2unqT
6O35mnPPWgXVaQRkXRV50MNrXcJyDvdDIL8OCdfEoLw9NGLsc5IO1Gf0BhPTV3m+D4J87BOtdTpN
hbtsKOS/Hm1EbIeor3tns8W+nuxSq+6BBoMeAa2DKoWpTYG7xm9EkjQJv5AXywIyXZRaQi5goYtx
SAxoXrZ0UlC2Z/+qs43OFKw3MGAolJhGOugK9WGby+0tMMA0mkf5HR1Ea/qut8Lo33F9TnY6AwD5
w2zRNnIWwRlvZEsuwEy6bDY6zPtTdB4SPlH8QDjp4mX1RnZOEmL9jp06ppv+T/kLB0sLCCdtPzev
tEs8szlC0DHbdlvmQ0d7tg1sgKimeDLroIrqXP+FKcvRy3C6/9Go/cLV/NP8+G6TnETBfRkrDsiK
hKhecztKQruRUpEbletBaJ25ZYbuo+0KRZ1RfP01/elkus92vIXr/k0XjxMlz6fbfoRkfBqYkd2z
FWnxn6q4J9JJv9dZCD+NaMfpqts9reAEnw8HYCPw/Gu2z/ubhyRIoH+NsEqfDxBVQgJ16twJu0e9
gbjxANomIKPhxAc0GN03jHjfsaxihDNxuw9bdGtLBMz2Vl51ezBqeQalIWDVNzgbPvqwrgkx1xDV
8uMBkHvhUZ7GOqDQO+jc8uat3MXPiwO62uEEznDY74b1gn98pn4kxuXco0tmIGnrLj8EM8xiNRbb
Nh4ZM23OyEMzIgqoNhB9Ndc0xxHaSt/V7htHIfuwcxjzSbwlLWfom3Eo4ZK6KLi3PipqssaIEAHz
O6AkHIn53d6LpoOblg0MS/hRuEbAK6xiDUEKhC0NOYLJ+CrO0f+W1rOw+JH9yxNAQfC4HJCWcU2X
LHbSYEmLAibi1P7VHBMQMIsAJVZTv4/NjZf5FNoHgU2nI6PyRpJguqU0CA0wvVDaucAWO/BsYqLF
wpdbn1HSTKWjavDQZlglp2tIj8HQN78vxSWaTR2ywvqfms9ERQ2/+P/mvy8nijhG7u3Xe5AWrK9G
D/Py7UZ147vlbrFpQ9Vrosku6B1PDyLY8Q/sRTOG65xKuxmm3IRyyVZHkRPY20ATVqr45yHzrtQ+
548Yacn8brJ3sSxRImyby76e4T9Krd4HmM4UdYIRC+w8VFgSs4d4FBpJiAra1c/PBSHbzU7zY6jP
FEabWtr3IQoQCqqn+pKr5Tnxdko9YJH17+SDpbXlOk6oWS6CCvkuicnMR0Qyigg4HjNnpScOyhO3
yhgN6ICT18yz5OoNgnyJozoigSRKH82aeyoNf/q2kYDtRIp5bRmZH/URJa9j5PMmY0wxQeAN0BE2
7MksJk21XirrLTNxJ/a+CJg5i0YCUw2xHTS+/jCma3g332pXLOTctmAS3U99MjVfjvGM7BBEmzCV
di18KaZRhfu5er+/0JlgYgNCsL+Z+bPrR+Wh/ajKNfN2mI9Nb+shKRaP9ycrG5Q9oN9OlOSE1c9y
CxOzqqUWv1EodkS/a0iQR5R6tsH/gx2xv30H5ftGgmtDswXxEzS7EEWmQmsKANUCMbrmspkUgGdQ
lypSWnvyjHkjBvR3btFQQMBPPBHeVnyoCUTWl6IZDoWUCGK5CRMZA0Tbb5x+CUMnE7ZqP/XyFyL1
GzsSkVL19Wdr2KR0Q2bOIeHjRZNWMyauq9CNzG1E1LkyrKjSwurKgk/v7GJGiaMA7UNxYMNNFnb6
ezV7F3L/FAJ27qMeuisgaoL+QncE5Y4gH7W+oEJfDVCJCV7YRJXaCIJ4sRIavpHuAdbcG0ZBKhy/
wjFL7kxMqKYBT4JG3hd/Wuj7zVVgL/xb4yajFDzKc8W07NsdKx19e/id02YTEnUIeoYw8Xgpu3nZ
d+A31xSBCcMFOJmb4BbFfcneqwm84Ob61LxjWAtwGaWTt/GUt7fMEUJhduJNnH8HTQFtYfNdZ1fk
xGlG4EqA7RZImFkch6E1UePZgo8fct6o2LmndmOsFEe3ZNzp3TRjurC6pkKPz3m4CUNXe+guUV30
KVyaidU//m6i3PU5AZZz1uUK5xqq9cGIc91ioV+SuDZ69y6CaeGDEqXQkoeWpHnihQ5BoA5WDMo9
zkvownwvcUOnDo5ss6wnzLTsB2ixRfJWG6pU71XIVEaaaN6vFkpqsWARmsosx7e5msg0fw3FRYSm
EiLfE3F791rVbiXSouAnYXbwQJX0fq6a6tsHKgKUIiD4gNyftl3UAG9rnpHyMEXVS+JgJXQJ1v+x
GZRLUOyafcZK5LRg/LaiR+NiZn3ZV6CD5st9RPWe4LNH2w/YP/jj52KTEwD8rOMgrJN1EfwG3GJU
bmCt9eXebXySTGnhK67hdn8PgiiQ+Z1vYachHzEFtpuYNkGxOBGN1xkESbWYp6FIHjUOa9A5X9cL
0Id2kdVpUV6+dq513OT4MbQude8LgBE9kIxM0ckVQ1szDoTRMQQ72HD0PJN/hhDwakc1TB9zxIW+
NBvlxUywKe6L9k3qNHOXW754n6ejzqRDla2GqLQUDqHD/INZW11WYyQm4dexK5nXeH91n6loEflQ
nFnJG2EaWeevcAKoxO7SU1k/Np4KgNmCinA3bH1UHfhcjAeHniLnkpOlGJodHKdq2LhfjobOTh+q
rlQCAOKR0BkX5zaWyuQM/7J9JG7srJos0bbo6tA+yE8ITyFH3iPqZbiC0COsDykypJp+6WvVz42S
SNeMx1PN+yp5cAtghm5s3LWe1wQVDX03sKnV/wcYNU8j5uZZG4g4nSRYDOzsSv6o8y1FodOQEdpS
E0zzcIY3VQS2rUFxoc9LfQkuLj54taGbpqTKbswqEp8cK+Vmki73Ls9/eP5eTLVzt9GhzK488B53
rSk9rKPOc4/iH2dG8wmMP6QemHucSO7ayJela363ZIkJ3NdH8z4i5tQVw9R5XjO4AGi23LBoWPZi
2p9bR4h5SWFo6EGUGI+pH713rYXZptoOMnY5xaHVid6YPRdr2EbzlTHLty3T3F35bM6PyOeH8AQD
zcQvs68zTmvzbvkTWLLX9fKUw6cQiEXI/UxfsiBLEb0LYEUN/k92+nQdn5V8fo1r3wyJN8q6SOuX
d0J3wf18QNo1L4SxlYDwXPpaXK4ok57OhLeMT5C+WIojP3bvgyHaqx4QYb5cwLlZnNHPkrmXlKJQ
TpvIrr+BxunPRSaMlQvvGmNzYEu22LbbguzjsHx7vmR4eh5WeaDP0kgBq2stpvvZ1bzLir1Vja/Z
BQ5l7hKN92f06ADlF38WmBHCAtEC9x4reilpYkOEBWKIurv4Z2Xh09C5EQ9vu9Srm3J0YOSNA+bo
uQQMfeMhvuWhRrU+Jxahh4oce4mhWkf2pHiRTrDUXyqZsa/EwKIR8n9WG4KicK1dH89p+Cv0CtZQ
TqeK6Rd63ZPF9J2aSx3pqR7mwv4dBUMvAuhZIfyCqWz0EnnxliIOalV4GRftIKUfhAwfpKQ/Nn1n
d4T16MDKYHvGypBRnoieMfBnmrxkMLVOgulNKBcQA43VykxhzL2ErWIcurIvMuANoJtdEZthelZh
RP3x5XaAqANp108ZE1Q3eZnnMBcOpsp1+IlO9Vf25lf7GCUUADsZWSITzxBpMsm3a/Ur2bE7kkuo
5E1myppqA1g5PK0u2Dzetd0XQMNDFaFzP+7AfqfMWQHLZpBooH477WkLoRRTnAKyOOJYYbptu2/I
DObyvfkx9RGK2TlF2N+W/hBf13CpipOo5dpTrR/B8alsJfxJeUXLVprL0kqKqo3I1RjXEXKALfyR
arSZcHcCmNMB9mAH/TAWs2HdeaV2pIfLo96gcMPjK5KNihYKZQnMGfU6PMx1hORVBw8xiPOz3M31
fjH+sEbJYOJ/KXdTObqYMGW5HWlyGc1CnYE8e6R0KthBvsIr1EoAXmBQ5vHskXEDanXXbyl6y/G+
ZZ57hAwDWbD2OCWgITdrxD9y7/fQsANEehB84/eiDSSwA71hevzIfwCwWWu9syrgrCzMLs4nJUKp
QeOfUT/dIQ+odgSOtsskck/kBj8MLLWMUKci2J2FXn9gcyxs7MYyRyJJSr/3GXrK9zj8GlnTsoF0
RqYhTw5S8yIKjS6wxSnnBf7pnlWi85RX/Ob6RQNllMgG0bHJ7G2qfXt4JnP59Bfy6RwGPYCOqzh2
KDSW1XUXafIZMCzertvp2rFFGIxM5vs+MK5FJeVxMUsiwTxPGVTaEFgEnEBZCG7y6fyZfWU2UAaT
3/A/sxV0+cMqpAOK3bV4XyulZs1s+RlvDFRELZD1UdjQElnEVzwtOWVYnBSqchjQY5NfHaulQVwT
H7q3CMU/LihHR7CflYaSRv8FYnNRhAcQ1ZGAiuHzA+TXxVW05wnxJtbSzFTOPKhLibvDOC9XZ+02
720nSY06GGRDVktcguHIySiYdHdRNUiPie7Ifr5Mt+huLp6PzwLgN/gRlyVQquejosir810rPoI5
qZbxUQUVbrGCSmkG76M3mt2IxCmn3w67h7AmyET7jl5s/Uv9A6sYyNq8RzTYZBjkBmLDhnVUj5OJ
zwsIDGA+7TcEp4d8pOpITSFylnUXy82A5/YRsHYemNb9G6bbBzX4Wupc+FUAugNQA8ArQDZ8/x4Y
SCjuKuE2tV5+NX08+meOt+bJ10SM97kI3zkDOcKWF3lsjvuhXleNYh38p6z+vqfsvAKTaXFeTN9J
LPFMGHWouuaKV7EVpjd2l+mSE3y56ErgtltGwnLtS4ZzKeHcBcW3/tMOItcE9pRYDBemT+88GgJA
7Kvho22hVBvLK1JicjGgxOZacF8tokKAPzf29QBwn/Ev/fmPDkvHV+PvPXjodXZbSDl/BUxh9JmC
blAVC2PyIoV45u/ljc87M5C5krnesMyUF3c8zksZhwbrApvGoMqGlAib04QZS+9WL9JvbbPBnrqn
ZJlUSuD9r7/zELxrG9meSzGkuyL9GHUJL9KbyGQvxhx4cAymLFm0QSu9erI0dTg7MjzqkECEIOf1
QO5QcrOzK7vsbiPAvyCQQSWQ8a52Z9ousHIn9RoM33cR4k4ig0DfJWBOEJAI8v+c6E4QbXUSdzHY
dnFcterpK4QFVL1oLyJNzpXSvpoiO8DUKI4hICIvGfY2VIA69ZkZXyRKB3dZx/8sr6FlZ65YxxGL
3hV8cYDplRIp+1SQ2q9xF1pYV10uP5D+RS0UydfYlZNGlPDx5+jxrAFy+hnF5kJ5vq3pTQvcjsJI
VjBDZtp1Ik1A9BAxcBO3FpbvkeEoerOCBLzhBMFXCDRXl8c/AwfN/HpnSyw2QUeSIKUFXPsczU3O
sZu6FQc7bDVCf+d+dQZ1qEK0vQch/pDlI7VO51L+fxOZ4pX3GusP/B9MGNuIqoDNEI5Hqkpb/26m
8iD3Q5MXnlWmlwBerB1AO6fo57ou+RKrDwbhHzbMsFAjNqhtGYLHQ8v25M9ebIxlqVqRdqYyP/c+
fJ297qrSJikRf1BCgQBJx5rVmMR+IpOfp0lXXRNGYFm/gJLt9sV7EL1kiDbL4J5jdH0tmae1Pc6y
MWR9Nb+y8yzM3PpNOdFy7lU8Sbz/YC1Fci8hd0UiPg6v1FLD734M9ePJBDekPcBK2c7D+HtK7JXy
ddQMPaHbACuk6qFrrxUnNbX2Fn6+Zk1fwDgOGpPdcMr6G0LlcyqRbKV9cEkgu6VGp6Y0nC2kAS63
M7x9dP20oGKmdur74TjzNIMpxT04DvV9oYmD2XbqEr/PUTFnNlLUb9mh8AMO16lUQ1yHQP3p1AX5
R96GpRkGLiRnAUU8O/K456YYRxzhBdnKw3Nqz0XKVj1HoyiFWEHTWq7Z7Y0ccJJijGj2hWFl1Kmb
huXTmy7VqeeOAwJsUhXhAClnXz/WnVK5s8VUP+8rC7ijB+VDLGW6GCbwQsu6pcJuzQ8FkTzbQLhB
nMgwOWxHy1pfYvfLtdRWnOf3+V7Pbl24UY4IQawKZhK1ycWsgcr5SHTPvLfL+u4L0yQMVgo20Khm
+vOcjv7J++i+kM2kbnKN7ZBXgKnIKLZYmy4dVJmp/gmVViERdqADvdPsnAzVMx+U20Jytq+/4Y4L
DSWXI6QdXcnfnO+UZLbJhcSxUsAVXQxgPWgBbytbp3ahCTr5i/JFYFwB7xpfoU0IT5FVOoxJqKtK
jmR+x64gF/alJyHgYryEDXDCojo4pM4FO0mDIFV946wgO0O+m3EngTv+5KcgRBx5rQFiQGWdwLpI
Ca3BNyh891CahMH1QY98Vq9PmD0pWnUdckkGtpssnot6uIBq9dx/XbDt3xEeTCYY0DupnHGZXbKr
/EdaM7a0cEqwSN4VVPF6blJMj7Gw6LrMjEWtp5gVyTV3WQmSk4bNyKiTTh41Act9cnsiu0PMLgiP
JaVa/ssKXhFk5DxOEcenxEwhrldTDzZiXe0tb/TlycGQHE/+Z8VKZwwFmFFwcqc86VeYGXAS8wEm
6QxJYfvxOuYgcDtak54+AxTaLSyo+rPiReD3aTH7igDG+pX+8ZBEu2L/BSRfHcEwhOGmHwCgdc/Q
BVsvdBZbesC034t3/1BAV4UmuBHu67PRHf4qSl7rHZ+RQ1CDMSV/Sr/W/MgzzVUiBFkAm6AHW2Nd
4Fpl60EMbOPZAbDXb5jlj+WWmQhzio2IXtz1fdVyxtldk23k0UU5wLhN7de2wX+0zruJgItUvnOt
lsKqPb1n1oWVPG7fVZs2ZKojBnrQhUMvr5SOHpRifMSMr9aRX42SghhpBO+4e9C/40S4a98BehOQ
NzVGnVFV4zv3T20uNaDmc1xYWo8Tj0FYVANb7mhzq9MwxUnmRRJTUCA7oZkUfTiK5fNKgw6Pkizh
wrfCbSLC0NFWjxksJNAZ8qRR+pprThGqVtel1b5/dI6JOCPskiSbdJCvy3MFhVydDLvjWoRLd9C/
AGdZcN0nu5/ME70ZgfFUv8O3RwD7/uu5iAo+j3FEAxydrha35EDdNe94xoTbDdA3YF6s/iP/77+U
7olbNOdtROsCpMkZ7vlwlIu30rDvhi2ySDnF+RkpF1Fr4vcX4iiCeoXqRUWzncPWogOOiwRleefz
R3OkcPXwsnsC2PyPcfrh1Y8eLDOsf3tCKSdDLrV+81Hvd0YjfLlxCI0FK9TlHUrQn9SA/FADXgaS
ih+MPh+mxx+nmQol1RZtorpW7cg62QRmPcbOil0amvOuOZE+3/CTs/NvTwHMCca+l7vywdy74haj
DO2Q4/nm4zLptmos7tYv3nEuoeFgb/tLBXyXOojoWAMqE/vFkwMlz/6vvAiBWIa9WcIFgLS0vu5R
70O2qIhMoQU2t12NaFvsqaHYt5HsZUtJIHS+ALnmdD6dlsyhyouJLVQXKg4qWHsLcDKp6QkXgtnn
5D0k+dc8bVrpYXEVfcjeOndmqWauDWpE/Bc7mu6c5tvlW0bg5Dky+mKEGaE+6DqdTbgJ3CvrUNvy
r4Crqk3qzGndDkfe4qQY9GiDT2G7uDZQbtohuxPhOVsEbrIKd4msDVOVGJlwvQpDr61u51S+SgV0
JLndfmuoouapD+HYINXxn2jjCou+rzzHXjseV22/d9wEUOPXFbEgwaXOv8nsdpGdxGoIGJ7+fzW4
Xm0ioT7COzmTXyzKte6xI9nz4BPwrunRs5sOPtNyJU+qUgL+JFE5Q4NT0ZCul7dqYEVUk7KbQoOQ
yfqkci7rmFnuSHYmeTT4Rmg1DR6GQxyNzsqWz7Pq46tRYWjUY6M8yMIdiGXFq/Mv8d89cpt7sq2c
kMZDG4j7vYz0z+NFqbmm4McDScaCb+ingpdcChZQepvNTp4bix3i/NxRm806z49MuIsCz+88fdKU
m17oZKggDanA1C+CI+5XEkLViOKl+r4YXgSVWG0wjvDrRHlpwyDuHEGTa0I78dFWLLuOQPHhRITI
ENsLRtvaW+Wr+9ey9gj98OwzyZ+BIbWjzMX+JoPF7eXwEnCrKbRXMzENKB5QZ5azmxehqpWQVno9
liriRK4zpVycK8f6ODMANZT40hyy/Q74ql8dWnynqOHpQISCox0jYWEqLFbO5hZS338Ef6sDnwA9
oJ+gaPOt6aK7KLH0boX7sPodu+3ZA2MIh1I9TPpdegAPfPTG+6PQvtp3GoYtuh/X6VdeqZwb7N/x
iWoUFgMJg7oZTCJh88d6t5hJRB9xK5ajemgEhJdv8InXjEYzXmiEMdypUjClHv3RfL2vIqhVg1as
a5hb5w4WlDNVB8TDtqGqK9xiPKLbd4FhUQKabioxgrqbxVgAuRfwv8JRZr4JAqWNnU2PTqLM8D2C
1ib878dl08IP8km0xLz/33fGthbx0LwJ7pxQZ4U0TAzLDRWlUj+P7pHnzwSrp6rKdgipE7UtbNaw
RtYSIi43FCsiUUFxt3vmh36WwQpkDjk7f++uvxdMY88mKujY5Upy0cEN1hT6XbqeL+MJSyyZ6hqX
kIQ2vhvMf3cEwIIrWY3MC8zIBRU/Z1MnkBE6bCl2C0WID3nkpnTpCgJlM1dpSsT3Z7KPxM4B4iNV
h3n6TGn3VKiXWrxZvcHFtlkNCgU737dWo3tvQ5qyHGnN+VJHanTOJsj456dtKGvM1ASZf9bEpWJk
odwGPh6We4RqU2INF3zxq1B+Dzz8eaQBYCeGgnPzDCtaXf14T79gRd78g8S+l/f+sP56lVL8grSq
LgXsJvLncfxye2bdRuG6Vf47QgnXeFVRXv3JoV2opGASavziP/VxET+xwCqdLfT3zoTCA4B/VcW1
tYX0a1jBGJB7A/v89OpK0dptmeEqQS0sQqprOgK75zw10QnpCQCBqbfMO6fNGxRAqQV+GoQ96esj
2BCwdqnhMD6OQ1gsN8/A2qT77sDZ7AN0TZRgP9+FSVyGBDbZ/b3DIJxPs4lOgJPUfm2WYoE+k9H2
BpUcYTlO8V9NESMpDGQ3s6OaZK4P0cikt8d0S+pHBow37QNBnKF82ei2bhnz8q4YCfCPXoJoObKF
mXp53NXfZm/lk1mmZtS0iCb92FQuSM27F4bRb45MVRwLtsjrEpzNa1fF2nUyhFu9rHjyGXxOvv3R
vKO9ZlnlZp/SmoR+Fq0zTjuEBHtM/sLyYJmJxiG9tdgwb1PGfq0Qr9/gVArKLwzOPljZk/Nq6uK8
PoJDiFHM5dJy91jgq0bk07EmBOBqOSuFnvH8U/6TbY1wo95I9kmS/p/4t8IkycTEHicjkDV/YasN
OoJ6CV6rZcWGx1Carp2twPZ+sd5nYPoJoIittEeqD4ABopuOTeZr6vPACS+IEwYLh9Sr1bPp2Rge
kQ40ARQl5GqoiRA4v4Dw5bpMPtEznk6RRfVc6+6+C5I1JzTFqZLWQL+StZTX3I/GzE8H0i6TMGxY
Wq6gKhBnXOh9ZsFE3pRWRq8luQ+KXZeOEkb53VCnHp6r6p+lY/wKcweMaQGyR6bULx1/ca+u/o1p
BGE7CT5TKzOc7ougZHBlPq4ougdrdd5se2QD3OZt/DcVAIga45JEcz3i0JT6gRlMhjLUy0s0NxYN
qRWSvxlyZSF6gk+lnk6rL/2Ofni9BuYHLPn+FOOttEMyxgY7Fyb6yS5odEOC3iqP10sdV1P1iPWJ
C4YQON9ahLD6oNII+4+cR3HgKBG9Jp2CTgr3IHqa3ZdZ1BkaSVY3PyQ5TYeMkZfxMhUYKQLgSmYo
ItBsxEd+PVTyDTtAuwuiUq2m7JORc8EjecgqkJsLcs4dXwguN73aWWFZfYBHHFyMGFf9I7Ykxsln
R02cGRuFapgyOIQnY9YcqnpKOGTX/YS/D3GEjUqb3h2P8sOQwoVFfmHRyfQMbaHqnRZMQv5sWfPH
OrljBiMQLeLyJhQ6/kHwrnZ8gqEo2XXolkm28JKioTybAMLsS3h6BSnjNB1rdU0PJZQ40fSBB2Ft
56VfrUA4WmGxy3kR4QOoa6+Q34cP/R2KFmK5um+2O7/wCKT4v4aO5TMESF0R1O3cgx+tzZ15+tiN
qbuIxXI61w+VCBFWLuVoUSDOULYzjZc+VAuGZZncwB3JPrqXXL1vlXAdYq3Dici0knHwt/s0glxr
XE4kgFliXVVDp75/TRJfI0c+nvNtPOwshyURkfPgV6vbVJxxVUX9fKmSuXrY4mNZVL+puLolC1Gf
4OD4Ob3hU2IjdkArvqzbMo7IDnWy0EQXPvb2OZWzLzu0yYNUrzBZo8RbQ03KxygpDtYUZpZIWXq0
kl4ypWi2h9Yl+Mp+1NyE1oD9vKLCgBvy7aM1Zp5CUlwME/bKAFZlqdjy90K36R20e4ei5EgAvlDJ
UcQaeAid0B+//Mw/5Gnvfj8JOL5Yf4aEkb2ZyJ1MWi1SnKHnWWyGZiti3AoCW+377h8HxYw0fOUC
u+QEy59sWbArknEFEY/274YzgfYi1z4hbNd/RKQpo9ELLYhgpsSu5lZYLPCeN223Qs71SkEz4uGd
y+8ab8cLSgZ0vFuXU4ighfsWgJUqleRxfZkGDrUuBlwgSsQKAwr5RedHa0DjDyl3uzzgn4uyDX/n
Mnq2lMIvjPoFr2EVGih0F/j4yAcfBxo8WHlFHxMiI2yPxpnt7e0NR10bhRwgHuor6uWuQItJWzpr
+q5DkEs+6FUmR3A/BA+dCm7PClMC5ex07lWXyqVqYom5C+X0MpICpyzv9I8b6tY8oUALiEwRl2e1
6D2dfdIB+15qLNKe3kn6+6OL0wyXsrrQvr4MYqBSDOHut0kqHoJ0SbE8yAc2BMZSJw/sQ8HMGMlE
YKJaNGjPLTU0+UH4tCfj1jwD1mDOzgKvo2UP36pGi6o+dVvK0PLzohaQST6yAwlQFNLevDXhRTsf
LLSy0M5g2NMv1Be+w4Zzs21U7fiXWsg1/Bdr4u3qFwivoQYonlqaL6g6bC+i6fvL8eQEeXHDKpKn
a8qbSLW555ycKnB7yZLxJfMZfcCuAyMgzA7u7Tscpq9AypP1wCMjItYZofX+JI/mSQMI3x+Ha5m6
jm9QcBZq/cm+Ibbk5KPHcuBSRyy7VLuwN9YJKoXsEjrAHWxsupQwHuCvwBqiBIaxZ05JTTkNdvfw
0tbOp94qgQSEenzbiDwLrg7guSdJH0eGS31yAtxS4yGq4GnQMKmpJp6Xobt/t5e/IaEtR6pLUMOb
2Q5ufGtRtX1OYMUKla3dFlIfAOeDrYf1b/186JoRr9pTJlt0YUTghCggy0v5b+GrtJQgk3Ql0gq8
3UEEkNVzn6ZwH8Zedy1DGEWW3PPobwWPmvoigoYFJIrHTp51dqFBj3ZMppA2J15ySDiV9P6T/NDr
e5bvUJbe76ZlKPiRmfbhqxQ1rNZjkGXXFz10iqKLprcRpDJWr9NwkBcx5liigdMm7DP8z2UVFisH
WZizX5tlYPEVcALK/BaNjPgFjD7+201+jw/LPcJK4+5IUeuEV61j9pzCNOvo1c4aXNPbIbLmZsYe
L1GNlEcfZbxdsioFVhO4Qf+IHDoiJ9JKcaTiDJHtREDZpSkqS37pDgf5e4Kd1unTMCpR8WNil5nT
ffBme0XKlBXGajyx/aIh9WAzhEFceNrY2R3uX99iLyy2jUzPYFbLug3wutsTHzA/aTlshdaUUV3C
AGd7ej+Ysq6/4XK6BhUHpMviHU780BPBkv5f/K8q5W1CrSt+qXp2y8tmQnObc8oAUGR3wdmhBESO
1LcdygkpGnjesx/5LOGbO9x5hrjt/WLyFbdlaMayxIpD727e8OErOZN0kkcuTG9Jc54MUe7r2aG0
7Eq1Aq7viDnKYj7GeUSqqPWdu/b0VRcHAvbMnY195ofxXZGOMrXtx5cc6dxCKq3f/kTj9KHYqdzC
UiqyhWaCG8Anf1rbdkGUGx4rKb7urs0QsusaBjQt3n0mcIfE6qAdPsRaaj6CK183PCFBeZNlSah3
VPKl8kSQ0UXMriC4fFK+psnk1r/7nxz8AqPd0me83CfNDhjq/XbbYduD2d/cZeX+DxCjyE1H5yqs
kdxZC/YY4hhPGho8UwYCfGLtVIEgS6FVNE24XoJmM9XYYz9aF999E03dGlRZNDSqYx8bp0Bt6SVx
jMPEBLwR2sQ0mVioMiUDOF7Wy5Ofod5K4XSGtJlpy9xJgVJKhZ+oOz9ygFB85NjfWyaKgCl0l3Tk
9xNjidEMxJBctJZPTqNKsw2L7IVRjBQIWbSVyhUVeDOcgRqcpEWTtyq4kU2u1ZA4phy4Itd+ZqtJ
nCE+zYzAeYM7rVRVYz3wCsIQzUbcLPkLMlnupVD02FsvPA9keK1A/W3Av/VD7286pMYdQZrTyFff
3/8JZBLjAOWnkH8cLyC4RoNxyjNxw9W3u6qrx9woJsZvB3VayClBxJwZYJsFl0Sj8LKsKUtc7vm/
B76YR8kd26gRFcHmqPylgYLqgBmbxm4nLU3b3m4l9ADp7aDgIEaI0E7o+qlCiyyGR5sSM0cDDPbI
BTCEhzRzsNjxuQIQls8Xv5NRbmobJITx64THQLhKszKOcb2Zs/xAcOJtuMs00mcICfg/TAeAS/5l
BOIY8YB9ARx3ls8jn8G5Sg1+flJTUs3Z6381RGRAk0xH8FgJWR2+6MC0OXbdDOzzG6ghXyyb0yZx
znlxutYVP4jXb9F0S5EOGRqE8gtfZFURRDLIev6oAEfMthObx99X0colRHPgoZF5paZRYTbTOoEP
3caJowBtm/qVQ2kpUxjTqXWO9t1n6e8AKUhVXMKX03QUqpI0aHWGLETghif7Hw4BREPY3QouHzCS
FBkslVANXQckacEMTT6KhOcmkclkJ5xyzcu2lGp46bfKmRPrPO43RJNvTU2M4vogCEpT5z30tj3T
M6KmHVCl907zQ76qn8GdHqYBCx+U4p3YEXVC0w0ivg7rtT6ghhzDq4vh9j1DZ+fIu/cTaBq3NMKt
brdgqAxYvcAR7hiQ3Ak8wDVeAyzjo4IpBPO/ngkXtU4CGixA7pn90K+Fgy0bOLZhE3/vKb6deywP
FBl/zyvOrMmbotV7ku8KfFFE4BI5fxVyp0mANrjsVQFsKIHAaLNpY7X3sZfn2RegBlT3IFVFh2Wl
T1KvibbFlB8nytckPmQJtw9feQXMTasKvN7HjGCfDaEobNML6ioRmGMdmwya8npPKvbByFS8ND+e
Gpqk/9dTMksqTs10hT3SPoUGwnq2JtssofydpTJnuxRR07P+gru5J6oUDiPDowSAk5Kulh6kF/aJ
xwJTQ96MZrAeOrs+jhvqLsX6SEQZ4ERXY/o3Xbmm45XnMvLwIAdxwTQebfX6iNEZSoVUj+c/P81+
T2YfR5WC8sh2VcSIpcebS/6PFfkBNeEhCxwzLakNZFuDOC+xl4k/kiIrEi1e21N94e4H0HIZWvgr
Z+3+mji1pk30nx7sSz8RjIPvEAbWHzKVID0SXlC9MJoLMPMJQAOKjkYGxugVuO9QaOf+U/rOwxxg
fG4uxfntA39o/RFXLZG5Iki+4t0sheV1/CQHKxJUVbm+tk56U5ZOJXQdUuMlsSqtCOg5agdZ5HFA
5sRNloLU940xwWWmtSbafkeNHjE7Bh+tSiXaIgaWFoxBEGiIulrVRT0uNupVVSfQxXOT2y+hrnKt
2r1wDfnYwtt2nfSzYJLUD4goVq9rVeXly9wP3eijIXdZEkNZaNn414npqx91SHQ5DUcYYVLGV/t3
AnTY/KIXMLCrsJvE4Zp+fVUdYOv68oUnQI+JQY8dRl5JPopLyatIWhtgv1SN1LDQlBJiaQCjb/m8
1OnFCRm63AqS/zg3/Kf+ufcGD0roYRfKw1rfjtuhb7luwGcIOoRFY4wrA9tsAFb6PCb2nyY/lIYp
Nqb72yZ+v55zGMR1kbjKWFDOC0+dc0GP1j0prgA41jyAcDGLnl7qx/6TRPY3uOuQdvl0BX5ikNcW
uAQ7ZJIzLHly4777Yb2VvUTQsq5LY2C+5PITAE4eXfBtJ5joRRZ3QO2ZCQVk/gHPT7xfVenFPFMg
FG5swdevqxNncNkj6zdOkjn3uuXahYGGKeOhBolg7nH5wAPDGnBkQLnWIvAZm07wOSs27JqNWYOJ
iTOQTrMcgs1AqtFdPwLVuIktn8rcrMiCJ8SnkeULwrVOPcDEggkqVCUkH/CNkdG4AFqPsjjGzcC3
iYQvfWi2/xZEym3w48wDPBWiRoDw5wt7OemRUpdyIwTSbrS89m66LPgKTVeQEZF04xBBo/ZB3+5l
6D5Ha1WuLoETn618QRefLZ/wQrTIIigyNvP31qcE+aqHEDpOqAzor8MLUkqdQ6yq8b603cykywf3
DNUcT6RgmU/DCEJiHjF4/hTBlKTNun5tNdS/NdZgcQ641qp/ejeqw6GXf1cV6QWZLfZuxoFQIHBX
KeSE0smDwPbaulLUo2ZIQsriHLlzaPzrOCZVfo/Vhondjr1pTFWozIxnK279k7nyuR9W10RZ47Jw
Ydhr+2o+q52cvxUfQhEePiWAHGeJ2XpltGV21U6cQKkvDfk2R0HUvFn18T9wDgDqJtMijWbotnFc
AwCWiBqmzdHaocHReXT1UJS4RBVMJ8T2zV+PNnuORZOP5E3LyB9BBcjTyCV3N/lYFHGzJ+hNNtgM
koSZkuW8CV8ETiiRpWkqIlzKIJM/MwYG9yh6gLFbGJyySDixlgcuiVc2zmtTFEQy1sdOIb8ynER3
Vv8oR+2h4yxZusVIVG9cwKxx+T77TJjwqPsg3Nr9IiheWxzMfDjXcpedkKQZBeK9Mc3huLBuroYb
e88BCs0gY0kn90AurN9Qt9maQpkk8NHbEjTejhM6L+sINMxzX2DYe4Uh1XNMLDVWfgTM00D6HS78
g9tqKamW/kA/IVKKEKqKlmbeoGlY0o6kD6K2prbr2P/T6kOQ36SoHy5JwDOz0XRMpE3776SLpIrR
ZWMKYwB2WdnOa5wKZmXYNCzIF/9UILeGlVCgow7lMJZq5c5IbWRO5knWspDXNzSj1ZUsqrnfjfKs
4Ll2/tURiMwvDqWbG/F7vqSkLEEPdccdYc+kaAS8gc+9xY9Ni3OiRdQI3rjv/UiF5Y3mefWxnsa+
VRknAIVyGRo22lhoYChhBqbT6pNky4SWmFwkBXzWHy6WrAoXzF8wNHe7P0HXwUQ0AMRdlSAvq4lI
7tGKOtVNjGQfP8MsSrCXaUksKYliuugMJXtOj/ZXnGaEAtVO4e3moPIeBAawCnXC1ojteL+iwy03
FSG25UtLRgzcEs4cUJi+HJ6lZzUgHgs9TwdSFHRRF+iSx5QFYZ5qWaIZWt76c1u8uCe48+6yZKFP
XLX7UJPN8Am+eTxhS34kOGuY8gNeBglx0EJjJ///h5yUVJfYcLjyuL0DxegHXY9dpiZhj3Wd+eam
vct9VLCC1tnEuvA0jRNNUh0nmYMKAVcvYafdK9zzP7ypyeS35Qz25AZiy2Cb5fl46ORXdsrpVwn9
SzM6euM5MFXN9TeoulfhVX2ICl05H1E3iXCnzoTbFp9KXtJLa9o4RqUpbKX197nL/srxYP84xaBJ
vLjW+/1J7E2vfLYIYFBhkZhPutNfXy8RKERFWIsfXznakYUyhCwtJqTf8yHMkz4kgaceRukBh3Ay
niEacD/KB7il2LCahOhHIEFivX5P4CFtBckrH/H4bqG/v4PDHkFOLNYdUIGB39z5dxVM8te1dJ5M
0OIZ2/wGM7u+4/92zfp8+4De8Yv2xmGbjTwzEJI9zZrv7UDngx9eWu8n89/mEdT7pJ5EUuXdn5ry
1POAo4jX/0BZfGfosM4fcVpWLZRPWGV+aTnnG1vuBThCUgKFrympkUUJd6Zblym+RMWnSmH4/lgQ
pO4Ev8KjWNDUOPBExTvIK4CpKdb3o2ZsmNUCCLFU5V05vE9aPu2gSUluxz2qjDVSfpDDpkm9exfY
RwQXtNIb/wEsqxAyTYjOlj+c5udzsJX3buLzT3jNK8Soa/eXcNCaWTPs2tEmoM2f4mtZoBatnum3
EDVwUBChS1WFGtcStsI+cHw+7iki5VmsqhqBJCu2IGo0Tw1VHDxmg/whZUBmXP7fZjJR98IrgbeN
ADCZccp2Y+RL15kF1rYrXfKeXj7htGzZDzfHxZx89TUmunN5O646+WNWIcgCHOy+qFJWx5If5nqM
OqW3S+803akA3zVKvB8n2fjLoIpt8fo3DB+IatMDBsQ+pufuhEy1Rom0627zYcRcjx3XxB8YtK7m
9IxkcYYPrsMWUfbjGlujO1N/GB/CwnLfJD70dDHGfDYv5Y4tpEcgjLXIirQuPTCYRxA0yBH6C8qE
dG8OrgpXIscDbbf4gVKf7iKO1TAfXjtK+mguj4uJGrySrxziaa7Ccl+Usp9bQpWsj0/IU2MFmW0l
F8X6+jz2WJUgaxitnOEwgAF8UBx2ZLvtJousgFx8OlDA7G7Bc+wNjcIU3r+0WgsAx3gEzGBUoulm
oYPA2ud2Z3Q1NSVs54dmJYk4CIjysDU8ONVOJmIQZaCI8k+8ii3nitGhoyVKCrin9l2m49oM4URI
tz0tiAyczkMY6nTLG7dbgqr9lNjDB0PfC4JgoCLOleT5gRXeSyNt4X66Zw9ZLbAaE4wtsJQ/njcg
aCKVEncthdrBa4nKwdNY7idowkr5kRpeEpXq7nQWG01dYYG5gwpktbjr988LXDq+qgL63Upqv0LD
5jZlQcKVbvHztbaP/0IfP6kCtTUaJgpCgYTdLzyjSdyrF1S6eLQDo7RqIhV6AOYIxAVfxfaLgVer
VwGvxaGOoRQmWC4qDyTB8gklG36o3g8Jb4f7sAyW0DyvH/c3dM8Eo5Tz3/PWhATm8ovCPE27JzeL
urpcZqYrS5aiCBHATCdLHyTc/+rSU6QphY9leGU7e6/Irbx9xJJq/l0yJxB8V8RKK/ZFLMJu/n+j
wWuLgd/el0UJMdtSCH+/7cGFYijKkAokui0NC+Sy8klvB8s87zijqkWP8xYlYJ3xv727mM1xZd7r
KZlnj+gONBEb9Tdjt652jDb8Z0XaTVtSlVRZONG4d2PYdU0FBo1ZgKooJNARBqE2fsTVO0+syBZA
KXSQrQows5ahAwFRr07QASlkMU188JjW1FooOBEgrG1f8HJQnpqtEDvGYjVuksdFy5TQehfLhqH2
QKMLYsMYxYCpyDhHLfFqiTZbZuZHCGdBQap8BdF7sq7IphR0qbwTpy6EwlvmQiuP8l3TpAznDHos
fpMQMk9R8IBFixaS4BFc865c4w3tpip66QUgOw4gedUfa+nXCPchB9gkxjFefPtM7kmurqzKnXOD
wE9F/rVHw0m/59708J8QoJrq9uurWCgbSjbse7afb0YYhKg3Fhn36Yuu83mlR4dEbtHRMPlNRB6K
Nawyx/wL279Q87f7QVVupWm5vi+T0PnCKWmaTpY6XtCzbBEfKDg9HbjP3HazdzbnBaNHxQOhzFJW
v3iAijetU9jZDM5Qt/uO7v/sL1oSUO7WiI9C781LNXLUsJH+QSlRTfA7jddOKYPvOZCSZA0N8ZV4
BSHyEOJ5VSPDauy1PQJWfm1rkwgWzBfVDpWpclS3woWyrbInRR4RTIkiG0fLLsFipkI3/xAroR1k
sZ1K2iUOCXjmQBnVlA7XqU3GOh+K8THjf4DqwbLNH+vqFfaFbcJY1vJwH1UFXg9OYLgFYN+ClRaj
71G5jk5TR4QYjtGtpwg7R8doI8fwoWWy4xheFCXouSAgv4D1im/0LewnfZwmKs1wDAQ0LciNdup9
IrXIEB1VkGMSjNjfQnzCLXL6i+oVNq7GeuaNCv/mY6ce7RND/RtA25mNCfzqqoHyY9piV5DkHNkn
OkZRcKvtkEkSvHrxDgeNefN0mP3seEO77amSOT3voXdZDiwouxw8K7RFfils2oP2yYuxh8mrPUyY
lquLs29pU1ZPQX1G8oh0MvpYeYV6kIweQOPVXMC9gHa8I3wNx8nQ6uO66CGhjYbAduA/104KNqoS
kjQA3xv+ehAs4hoU8ic/uJOoJK4kTj0TKSqvXClJsIW7nBPlT/OeVrqLx8H04AwBrsHup/+bF2EJ
ihPr94G1B7K2hEHRN0c32E+etl4nnuRpYTAWAasAwxNrj3RT0xCn7Ze1FXYC6RK/1pAoJq2q0LUg
AeMctWMbAmo2u1We8EDkMqtGODtXHDqydznOWopLGy4YqvrrNt73S5HcU7f4U+IeEXEb3nJioPTV
fJ43GECXdxscGLDuPmcTO+3A81RQKvjRknIIGOXtYx7o6r/HzXV1hzYWemrXNYoMRdVb4BxQqNg2
itwzOn9sd/wGtV4Fml/YNa5grl7ld7Y9rlo9Xn7sOherfo8IVMpv5uT8eHzjO9V9R70FATT/KX55
IUVk+u6es40rWFeoKGWSKJHNX5ttRQDSWDrfGicz9rPCojRZA99kKoDCRnoIgdVMHHD4Cqv3o9vg
1HKEyHvik2QTsItsc2SYG1to6xLvkIVVoWpBAwNGlgeS3MA420rl5C+OlbqIVV5AgxzHfXPBcOkQ
BCaXxHElyxFsEabPZUDoLMKCS/auM8HQjNj8nLKAPKTufWE1A6hYyHj22qF4DDhiycV6XtS1d/+a
Atlg0HHgcg819tR/orrGbYqEqtwbmcBgDm5VvPsWaoYsmQKrZB/nuWLfKuWiLI/JFpJMNS4vlEsF
rRF8JzW+luHmFDmayBtb88HWP38JRmpQcw+h5eHZ1uz8xLDgfYfOYyTxb6wfkBEJzlqwQBANehLv
ex50dcdOh6LIuLSz0VylHI3dsrvl9GjXo2nYbLJEampIbCcUrJogkm03qB2jnqs4SnxcNv3LYhvG
wr53kWTsUB68lLKTMxt5FnH8aZLfDtgBb3m25tXe+D2Znun5h6y7hP2jQe+EFZMuWAFQwGvvlzRI
L4v1tUzjOsFwd1lhejcpJyeBT7C1R61SMOhUG3ZFmDnQE9sNW2r0cUO4tcCxj8fCaoVnOIQN8Nd4
1jHih0VqpqIuoDKNwDjsJfIBw1s/m2KZb50j1BR6pnYJDZztnnNckBHpv3DrqHrRK9XR0IgWP6nP
tyjJbaKAvz6xrf9yAQCKR7Wx321hvjhBpK9UK5WMNmSuy1WrwsUaQWg3B+swYsgdzE5IBel7RfTn
u/etYGEKSgHk0ZzQS+vnDm8dELcTPh068fF/k5GpFWU5rE4LZvN0qOJG92yt0Tgt7zM9B+ofmIHa
26ZY0rcIJ2yIXhtWWqz40TlFms9Na5PMPVHiLu1t0R0EELDYhM0XIVx/g+TRj2Xum3DUyHjmH/Z0
nYiM2TYZvSs8rq8wHDSlqPiVIRvJTW1iLlVnlQIaJuc9X0XlxNJFF55SlumptB8KZOha//ekeMVS
gu+yIRhsEvD6GmTt8YFvzwmGwS9Wlzl6aTudfe71Zl7q4ZREGddy84GqX5QGdaGblmZ4ijxpxBv9
vWELN2Ir3UebPNFs3J+c7LvrWFTTV2YZ3ygSctYzVGM8oso9Fu3Oa/bi9Sjq2pq0Jk8mctIMWBMI
lKDi8qsfrsTmaijhlXT5IXPI107+qHF8OuWMl+4UPC8OdYbo/VVGUWXq/RfOLoyQQFPSiCmkd/G7
gWZkw9hJmYAIYfSCdlZ1horInnhn4MiXZqbm4KoeDgeT5T9Z1Et8e933FeCn9i8pFimZ/3XtDQEQ
Bp/uixD5rc+9rgQelJdizAYJ/idRJc3IbIah0LD/ZGeYqdeAxZbUCOIFjdJ4bnHTvasOJWFJ7IKH
D4TaEET2vI1YkZgvutX2D4K9SoIWUzvAxHN9UkFQUOPnXz6L2K8JqmxudUf3421Tmu2mXsDRhinU
lefRv/T8BVp6AGVKXoOvup8BiFAL60YTq7ZyzIoIO22LSDivT/hmbHm/Tab7RY6IHSHN3TB2P00I
Qxz210UhbQ9nMhCr+1o/4dCD+zOil7sRpnrB07f6/DsN4C3+4mI1cVodejWO4QMauGsKzfz8c6TG
xN88MM9Ik1dWmPA3vpwNKzfJQNh/ACTwlZEuv0v9X+EmP38aMtP9cSNczhYCtMJ2UhcMbuQS/5m5
gpzjnkpRtcb8oBCPwbbHiy2aItdF4Kw8YB2UIPK+UvUg/FMgP6R3IcWrRueby9+6JBQcEa2MFDSA
8VFCipqGWYLIWA7HfVYeRMSZHpr6jsC3tdgJhBLvyv8OCTpPTWSSIAF7AySWXExwsO4fOlPNDfrB
w5DLQfuow8aeMBE6Fs6XaHvKqCDHNbTTZo41hcbJQFbrMQo+OOyAONdvG8AdTZcb8TcoAc3VstTD
tIZlrs46L+bsaYopVpeG+beWYAx10C9aFkN/eidkwhysbUBkRwWvR4JqAeOQkxpAqZcAUQx/F2Rw
4KJPZHJaMu8VpH/eQyp8OGtbWx0C76got5Q8DaJI861Eq2M+WRwo4nY5dX9Dbl1+WFztMoaksMmh
WEKIELU1ruiwsQ0jJ8uOt9Y2gVTxXBf0VtdqRIxDsEIZTiWBS7OvlZDt3Qd4WyBoycDg5KANebWG
MNDRgzOrywMgfwDPbK0MZBVM5SqW6+bgoaJB+ZNi8IHcRiuq9LLuEy1Ya24BiDd5mOWgLKrmeC7H
WWeBH0QyQX3lKQpHnORUVrbs14SQ3GZJqfDFVN1E0vUtqqDsEAYGOzU9tVgezOmuZQewMPwYoubu
IcDDGbv/rZOXlXYg0fidiPNpUKlGYvbYVvpZH4/1ryzeG0SRZcME7GB5ZSN1SV/gPYTTQLJ/0U+b
kdmp4yJ4DaXXD53WBm6j0IJoAfxM8BOm0RVF2+u1pyigEx1h1gCQi+lI+znGwDuQz+sEzee9WFam
DtDgz8aUd0OT+vngqEgGTTrHba3Dy5VnW8uYsz2hNdSXlnj02pzjQ7+kD0m/K7qwicx/5SN6mOSC
CCPLIIXNkW+bvCeJ7qfwY//d4P905LlteTKwBCn9sW96X9L7/0Rk43YSGKmSfwH4/sx8igCxqPUF
2jx3XUL1fVMZaojXQz0G3igSvyHote2tWRoZU4NsyRGCPBhHuWnUt03XOZMCQ8fqWNHRPa2Qv4en
Z+ip3fLUejgT9C51eEWcJ6nNuJ0j21qkuMawb4XcKu+fzewZ/h1Q7BuddM55lwkYNRNlj6glIjTj
L5zKCj8MYQQx50qe7hUy1gliw6ur7BazOsd/aw+DtQRLsmzqmTSrMupxX9MZz2PKkL0T/TgtO6s+
d/7rWMGT8kL5iIN97zCcM1G+BNSJyUOwbWNFq81wfg0QqxoWJy+dfp3aKZ7h6+jgZhqUSHCPPuTy
f4It5+pQyFKUg6RLVrFlhz01bc7rbnFIKF2hqBA6X3Mu9Ysq6jFNvkdP46QLDVM3ZgKTCJ7H/pEA
3SoCr3lzBP+IUbg9if25eZF+EovYYrs60+Sgx+6NUMbLXn96+77TEjNkHnUmItd0twP+jIaau/7Y
UjyJgzOkSTKwhztGJHTiRXb921Zh27u8fDL+Ffyr26LlDPvjbqdJ4Gy/1c4LZbbTXfgUQI1jiYRW
M919SkGNm5XZv7CHzOtX9SJbL457Fhq6ZrQMTXP+skWaO6VNlxOJ7mw8djIqN1zsdcjSLzo2SM8s
GMekv9cYXseTHTkYleiUnndBaMBZR0V263H2l3zRnFQqGnRsNSNGpf/93LjRYVfCXrm8bVlr/2T3
HfqySMQJFhSHrZ0C2/J12bas/fBfpCHxhLXLD/sUUW+SMRr/BUsycmn3ynosBq3CFBSRZFvTVeUn
sLQDQFr4diUqzacLqsfwlcLTUGULyRtvxs8bq1mt6+1xmZ1paKei0qpfAkswimmFgRj0NzCA1eTn
Yl5v1EP1Et0/JJIaaT9SW5W9o6EIg62EMSsGN+wmriDJnjFVuq36WOy4sMGXrdBbgm+EeuTf7aLl
VCiIkKGRoPtU55kn2pLsStVSYuc30iKYLXq1NUHw9JepAMVdn9hlsW4ehgn+ZHYJQPZ+X2jo1W1Z
Iwy4RPD36VsGgzAQngBuV2IdzTRfjg+fPFQFgvc6dpxbig8fG2k3LJOhSjmFhi88qpH+4y0jj+Td
rs/I2OGvNzjxQDnUAv7wfVqvW7haNyqeay05Yi+l0tl8yHs3JACBJPdATbVNk7UaI2b2yFixsueR
MZLE9I76j2DbOz7TrMxz0WH+KaxCK6srDSH+/f0WkjHxgiMQS1Wh8mOZQdnaUveXJiRVJalKmY8x
jJKDY70cSaDfKxptrYQY3pa7/VGbfAz0s6IXlhJV1nyPqtob+mrC8+IoTKwqH7f12q4S6frwFYXm
ARdsjiElcU/sCe3t/Qm0T0Q/Yp9J+2wd7KkctOzbGnI/SLEhi6GobW4vRdHTsddbXdk/HgZpQKDL
BU5sUcovv5n4yzLjO5RcrVUvoTlYSDhNVXEJdbqr3zCuQgqhOsT+HhJgsyLCceEbEEzy8y14crYf
kUf1anXg8ooQ/jp84sCUr9K7Hgi0AE6CmK2xcFCdFC0cjr9dtcJXJs2l3XLnN9Hc34gXhKbY0vYc
XIRPYdpXxEjJ0PPC5XUw0WfEO+HvDjJodIQTWnn9kOedqQ7c4P0j9vLceLEPT7jrPZjSutcCyiUG
fDaXpnVcnMBjkz2Mm1XpVOWzYZZcftwNdZ5TJumVwM/NIIpcHeq6tXdTI+++FDGv6Epe9s4j+sju
+izRbjeqJX+p4zyeErKuPsZWfOgTSWBG/Lq3BuPnlkieT3g0M3+5WGEzjrF9otcW2+uagSVjJYEw
ta7XgmWAQuYexTzj/gWzt/1vPBe4C0Qx1weZ19MsnyttZgI52L7G9XitTTf+1M3uULCGL/ysNczB
L5O2MCcmWu1MzbU6KZhM8+SEq3+m8OjalNzUkdBNqBSw6KLJh1bRHlfamk1A/5Abb1AyM1t+PSQj
i4W2rIRpP/KAmnPcypLFxji4KotMP1ENEnEIbZMXZ5NN5bA2aK7WDrcEf4WHZPzC4pM/FMQnmZ5F
lZoGRJukoZ1vKQGBtZEbPsmEnK0UPel6vmXUkDQF4w57d2eKblz4QG28i9NVdeJl/OcqsVK0aNC3
w6S+Jwr0pfYRcxfr0URFNV43vw9Da20Dy8fOCkphygNw5jMX1lL92KBRHge3es0YwJTKQ+Sl61Az
Q9YaJKBG6BxQOqBAiRUsmAT3jkPdFcMFywzfTGPgARX1zpRjyb46e1NIRIMzuLFf1fobvEiFRnqx
f//LoTWxctYULbO674cfs/guWFFVuShs1heLz895T+uuIpp3n3mYAdLwjyOrjlSnkFvw/g/bZtp7
WpTi+hA72n8Isx7qQjvNBQoFje3sOoV6/yxIP4C4jzORwRLDIf/hp6z32EfDy8YHKNiu6EyNJ/X3
kRb5WRufwX9EvCKoAVzMc+8MZke8YqLfaZtbDFqjxXpcz9y+CBxRhLSr9q+sasFW9C3sjG2UH/j3
8BlhRwK0KsuQ21kF2iTJugvkKxXrRpDzbxUu0pQB81F0vJWcy0SiqJBrISc1+LxNfND6GmoJg6qj
vZX5eOBHhOgl7PqrgaFN5IDzFcndkpyBoiyTgjZc2QWuSGDITCNufAUJXiGNzSxe+eGoyX6JoNy8
ML6vHAiCOvNsNhbieROxMvXO/Ua9G702btnAQrI8Ls26BpQdhJ3Ez9be4DiwHSMoYe6keH74cIq+
eK6wqj1cj77CSTU/cEuBOnCgeGLpWErkqTy7kIUOx2YZzq8kFkpqVX2fjQnJ1K7SE/OVoxm+dghf
JPoVAZE9dIuIbWv4mOZ0RoYXBYZIOLV49cqKU4Q2Hwb/4i0o9aMjvqJOm6mW5/I0HZPy2+YvOgAu
c2OWo4RgWKqln9lw656LOMmaRLbGuyCdpo9qMufY9Rms8EkjWc9TNbAT3vxwfqAIwEUsvouqCwhj
dpyAcErWTlJ+zD3s6mYg4ux/+Ub9FRHBBrf9sTqRGqdvNllY2bPqUkVTH+/DQfpjdTJYIQWHw1nq
2WvRyxIBxOA+hk20utEIPlqOliYhV0kVLEtgmtoqRCvJxPLsN2NJkb3KfKHZZaSQK3xq76HKdk1v
HtH4xF+2Mg51Y7yjodI/RayBiu78htfXtVlJto/9XkM1W65+AAmYtiO/hZkERpp7TBl9lCQP20tx
7uP+oq/i0KhXG7h1+11UBjvdMD95cEWMWJGl4GIoHDcyCgUlbX5I73FzPfe+fHjV90OMQlIStsQx
RQXlGBbBYG0URopXpSUtMkmX4Hlqa5sM15//T4dBUToT1jiribIyE/8anxJ4otVrt7kahCFk8dnp
yhCDpmFV6NwGE3zbUq/tN4q17Q1k/hCfXv4taLKO4omPTbTvI/um+IyDqprLNwb34cvJrQltaRff
ha2sgsaBv81T6n8b2WjG2H9+KtA9QYXU1YSjpYYlqXR5Bil/pTCgoGLNiHlUi1omf6maXbi0yME+
E7Mo7vrIPAYHSp8m2JdnhyHUUIsQguN0Gwlmd/nvjWzhP8Ujar3a0Yur2mnfdcTqMkao+2yNhRYK
zBJuT0uUkJM+jfIn+iUF0BuLh9+2mF5hwRlx0ETJWJqdcHpsLZVHAcGtWxlIhozU0wW0TjIBx201
kCI8iv7nIpycykOk5kEcenrVsv6yoQG+LyvSPE8mcf87KJdGV/NwXkndW9ZZXfG1MOCfAV2RTjaJ
OM2io23zxeJp6lG/AmdqyJ+Id1VpTL9/2eUSkJSYA/sVNcfV2HyLP/jV0UfwkFpjUwcGgzotAG8b
6j14x7/uC4UH3RYsaHauX5NHRa6jsxJV1q0W8bWUlGewhrnOoDzhF3XYgXLPy3Rvz9fOIcxvA4g9
KFSSrncGXxT0QxWdeTXj/ConTi/diqUzJlz84XwHGDoXE9o1w53JLnZe9WSGbsDtrlGm6zDzTyDA
lQw34ZhAK49y29aj9v9/7HhFr11lSFwHyh3kzvhwBdhSM4PUZad2ASvq2BMpxGA9Qtl7ftYUk/Xd
vUVGizV8jZ03kLSydQJ3l/AuX4PZ/3Yw0LMH4NrVMhiVfGAKrJpmJaCOnHDRz9kYsJWeuvWoxPQs
qjCXiqOMioNiN8gAODRyywzQNRZjeLdGIH9eJHsWBzlmmRihmTnGd3ZebGVWXxRwbrsM6QYwgaMU
P5Aiv3N7dvIZVqBMdbc7vNpO6O9tFWZWybwRbK3bgIXTyKirUrL+xyaSD6mg/MW6KLhKROv2l4ah
JW4EqMgeL+OuGaJIJ2Ko0yg4j8aRnJun+lGVTeVoLx0sV/UbbZqyYsZPUjVQrYoB6OWlQYTpNM2U
0Y0JNn6pLBnKVl7sufPVhCAYS8GTx1iFFOyY5OkG6uZuJRH68wLPU7He1JX/le3CU/JHkxU5ZSXX
nVMfmp+7+Fj1Y53c7aTCnHiu58Y3Xq1zE9tvEVyNCOVDZ0dTGsXTJfxBMayjxdBDP1Fwwk9nEQRI
CV0kf2Cl3mmOZr0BHWUdTzq1zHeZruM8llsDMW7Vbs0suu+13y9haPwvbzOO0l2g+bU+vAt8MDpq
lcEnXA1bds+1LF3yLfkgOOm5j4vGTFHckhPcwfdIFqPJiyL8Kt+rkj/f29iOiyw1f7luHiU/N4eJ
ZGs0P9l0FUzcfLtzdzPyGcJm4ORSj6/2i1+fUDQuQTMd9pJ9aAiAvQ5GM1xC2kN1CN4FpFqyZ5jj
0154NRGuxytutAhu2AKV32OlqCvzC2JILtQK9wSg+IT/r27U8kPdYtHaKHLNoeK7J7Iditn9KFTB
Ie1s7a//w6TgUb1HwZu9owexmcFl9/D1ui8Mlv2uAogU0P+h1oMoQn+spGM7n0/SgjHRhwdN+3ja
T+W9vBowtJ4R4zzR3bSaQqRjswxwO8xhgnK0opEAFdnqFeDKNykN5u6RAdENcj1Ruoh9LexVDLhD
F7r3QEa5WyD32/C0xfFoWhh0c2zw+jORocWFqeu/DZsFIuF1xK7P00OEC6rMC5/t3mosGeC//yWE
nCwinacTzrcLojEWhuGpHQMC32uo1eIeOMHY1oetD0oUVTuyuXiyi4taLuN72AGgzfNJJMe5qahR
Iw+0rE0YTvs3SfKXg6ulamEmfFX3SMqRHUWmGmyTa21NSYqX2m2X6mBcCG5WGXgFZIs5zuQZU9g/
VtfWZHVlyQ+J0HcT32j0CV6IacCdG/jdfk1pTva/10KJ4E1IC71nrjKj1cjFsrgE03Bd1WrPy5yI
kd+Ug/kznLniv4ysbqefqZabBz75QPoGoCZMhORHGamnlns/IoWc+PgwhkRbXYj8sszjiSIvlPDE
+t4U5IE5RdCnZjOIYBi4lNuM+duXWfHQOMDO3dAkVr9v32R60zGK1UsGdajFEj6uQI5nHtHQJixJ
/4gZ94CHfgRKsZCletRx5IGJowZZDcCgEBvdt0g0RPxPAB/FZTrridomu79jv5fvBibXdPbZOn4u
kM0XN4Iiqt5x9XLxGttvkyieDiVzNUbe87yf89Ka+zDjjMpIjiOcHmz7y+iWhhS0xUkEGv9mZNpu
HY0xN571+cziEcIIT5AUtKd/zZaY2A8pUoKW69a0FfTja+0AzaqHRViAiyayyxYcXHEglKbPKwiF
RLhS8gkMf0sdXNSw/TXRo5uFKJrYKe2ic0Pdz/pv+ZJgstyCh1BLtKPMeOc4KCZoIhk0v4Lrh0+a
wh6f/5UfK+gMFh2hrVZmuRQYCo8SrV9WxY8NKyQ99R7dSoXDQ/odC+dEkLcmvYhxst5HQ1FkjmRp
ci6p1k1fLiCVWKmbjNt/uM7lo9LTxwfTHmZcyVoa6damT8JdiBM/xq71S4M8U7KjzkoGDCrMRTLk
mzJ2DJMG/CRPLA3kiOdxWjVSo/C4/VXBIodH4HSMGgMp3aKthvWI8DfkP+uc1UW2kT4WXboX5XED
n6FVaQ7SDtP76WfbwTxP22aAAOMsl4qjaeUeqF8psFH8opP1vMuCEYkjAGv5DzwBGDwIpSpm1bUF
Y2Ip+IfPJRNm7suBIFbY6WN1MqJFS0nE865+r/915W91XAEnfn0Qhem6Rcue/6cfxCXzg0g/jVa3
Vx1Cwgug29Ypiq45oV9i42cZJC/UTtMWe5XmgmSRSKyD9Z8tg23Kd4f9OgRUvXmRND9ZUw/qDdsu
KgIDmWniYDgJpoXyu9UxMa2LMRCwFVV/W5LrDDlRdmVtmp1xHF/xp1oHp45X0D/tAjOHJ9IbAKvU
Fh6B1UsrUONI8ynUTY4utvSjuW8SwgjLxnI6HfzxuOe/fdsbOQe06w9s70Gf3NX6Fu+rL5/gt+hr
PXimGrF00C8HYToBB2QuHSwQtsim88FSZBu0cvx5ar1j+pRkD+x+LWCtVQmDTqGd7QVe2nE5d6hV
WArF//lmAKWD9vsuUFJVBosfmk7oYsf7O3rynKwvf70lguDDaZSUR5BULkMl/FcVq4vIx+Vzq3qz
iaOUQoTvjFsiwutVQbIWdyvPXl4HO7NplcvS9l83Z3bXKLStcHilLcnBP3qQkwgD9bSHUJPhlNmw
mJcrksp185+rKr9Hzw0IWM/O7HWl74KlmWO4kpnyPl74QM10U5Ph2y+qFI+8XDohIqoLpI6u3RMs
YGI5EGWD7svgP/mk4pXFcE7bXtUKF8yuruQUPp4BVJ29jVyvQdK9ORrSWhH1wiyBgbhgcQ0iIA85
1yfZIMS2y9WC9hlXia+jYZRIr6ENgBUlDvX7ltlqvio0n8MVPnZs3tgfO2uaxOgEbPDJ2e/B5tQ0
+pTtdMYKq2uviDllIjPYyOJODgTCPEsezU3UXFjnJMwpcbxfdPhW7UxbWFocfC2fwHAzRwZ0IcTH
fXKiYyA1Xp0utIZGLBdwcdn+CaDC65zdezhlcV0Y5zJom4l8nXLj6KEYDEcmXJq7+8h0RilGw9uN
9FvOtJQtkRaQtpkFua17EWJsQGbojoJhgi8Vxn17JN1Bd1ojGu/Hb8t+suhWwRHO94/TtSaUsVEG
9XkuWhMsHmfGrXWAfwV3qfii15PqA+sl81iJJjvti76pqwCxjMLzfNFN2lV8yc2MYfSSG5/YGc/z
l0L+tSb4kUFxB1dNQowf0/I3/lnjU80vNDl4Tcj6NSN4+0r3ebc/Oggep0zU7eQKw6nopNKA4qBj
uvD1V2fPOU/BA3SKOXuZ/KyqCOtl/K6kdQdwuoruD924mpV2HgLRT6E0KQ0r9S4OH5+2tcJeUldQ
OZCNfRq9k7M1X+2zH2fjnMMNb2pUPP4erXA/c3wMCjZGk3I3fWa/adpzCiZgLSLwlFlgmCu87qup
OBeeCcegbrrplpZC10FtdkP7VQL8et7yAPU3UdmBDBZq1J4v0xOVLt43IDe30ss0f0tBgga0VCOK
ezVNj42d4i5zL9i1DIRt6XaDd49z4Hg5G7UnfWCu5Ksv/lEmHv+fk1/ky4TWjtRRUyWHvSeTe4OE
l+TGzVoxMf47bHrXJdCQkXyNoh7FhKjc2RcpbGr8eYOHmWNVuAuiO/shkUvLTfNUgR1XDt7rE5qn
MCr1h2x2tJx2U9xrrSubYRIoLifOiJ6R8qFFCYU7CnDjfJ14vxAZ0YrjAUvc8kgct5KqxHEd+anL
ats7vWwRNbHlALE+eEF9bFni3IRkiD845YmrM33VWK7L/Z4WO4++vYQ6GrvwZr/XXZeVzA5RHlVi
KYXqsxCRyF5samzF4MM1Kov6CFHniZKDHeOPRMNZclkt9eDXyIOOfLH7W9yvPtjK2BqhnSEYhV5M
j30LeFQY1fKJi3NkMoQWOyHUNrb81l17HOjSzvZ/vP3aq6u8x9eRvtOAmfNHxFp45uHAkkMvfX+3
KRtIexZmzZ4+s38rLjQu2b7ok0TMyiKS2AHQX2a740SVTo7GexI8g4gztKCrL5zmz8qHwW2DL7Il
Wxa4Af+8LW1bFzPodr2RCzRje0DstmOWdsDv4e/mMOGgDH81IqRpFapVNkce0BRbOTgTMTjErPUs
DxBgiFoYQ9US6iaJVcOtYvkwYjpXrJtp89A3Dp0DTxhZZI5NZ/uH9Bx6gPl+zsOCTsXx0BFEC+Cc
/5ld0g750LWaWAulTsmcUGVEA0ZTALkwOXbiil9sw1jVUYnL2V89Ihjd3YsAlvnbEA0kzG4Fmhug
gt0ubWcC6VkjvaiiQlr+ik/UYKejKzKUt+GV9jyFR7HJPBO+3GnBwtHc9mW3EymIfixXYfGtCxpG
ZlKWnJGOiASNW4uND1s1NwgiR66HTMD8FDCqsV+CokiIOxVl61rLrPdPHO/7A1HVRb8XUgxIkW9y
/V5KCA9lxodVSquvQvhr3+YWtEtOAy11lRPAG/pHy2py8JihKYgyBoBXWySxuHAghAqJLaUwsqTv
7lNNdwAe+cNcJJyRhxv/gPOzWRmvx1afZFzQdudoC4qX2Y/+tt928QkaqXD4Wcj+cs9XESI6zjFH
Nq1hMRWounqzMIf7i1DRK3rW0rEHqq2aPAl5yABcAwD/ZGrX6kIFhc/BQBcleEnDgxxKB4IUh9Bq
Ez//x2jtWSt29qAr9jw75adtILEOGA+1qcqvGLLAwN7WEe+Cy3lC9q5JV+uqrDT54q3X6hDGKKoM
cXqOLWOaMWQR4v6pAFJ0qu7lIongGfe2HpoPOkXVEhEX9nz6w7/bjWsnL/aycfdpYO1hU+ywYpES
OSDZvWqTCFd4GOmIyiV5bwbO53poVh9IP+gIZGsVxxVgmjedZdLxcouJxd85G0C/4pEY1HSu7usB
NATWtNRIg1lOuueiP1MTOccde/UXXABJjhQTxCt4KOMcGirZRowrGAKPlH/gw+6C1ppX0IBhmvN3
tCVa8HP0QfIMnsCBU+g3dCd/ZEZvBSMaLSTNR3pJXBC6fmwRwjiQCH64i5Y4T4DN28P+UZdJq4Px
Ao0U4TBFzdq9cPBrRDDWirGqC25wAgPbsmmZ1baQ5dtJuh3FHqmo3flGOWjcPW3TJ4RKBhubKHox
0r7BOmue+wOtxjbrUr40gpiPH6m3EGpd0SWie5Uz/oKu/ZFJzNTJnnbB2C8Nb8cjub/a50xeB3bN
Jo8HPUsvlWSPTW+4ZgftU2fclUFg3CnCvcIHc3XXXd0eeLB46CAKehS9cTyK+hOobTdRIjJSgUEP
ykLGXlRr05lecitraXRooDFO5f6Iw1RXfdAL1Hny3enmNVp4KwIDM0bXHTPL8WRC3XpGsz2goZYN
jGR7QHbeh89nCNr6OogxX0DaXFSuvMl/lTLy7fP4ODBnkWCESkBxULt1ncAeUq5WowdS9E3Dg15i
pCfS+p3uU24UHZrvjL3Z+tt5C0Rb5OsHHP2EoatPAR85m1ZPcRAWFooDPbstP5ZHXctS7kJ5We61
BVuVO++I9Z1agHc+rT8ULllpv0YvusHy3FsU09s4GYt/1P8xHQ3odkhiqqMeA/ZSiegJEKQ6Dufd
iKS7/+Cx1im4kmS31gSpxRiH4gK9pkSqTm7IdWUxllByaSxaUvcJyv9V9q6X7g4xjyMTkoznftrj
47nagu2DlE3Q/u+bsvhNffwg45jXswF/XFLirt+yo29JjE4npT5gpnD5DTqG/pnc/YQ34rYzz4Gq
pIQrbJlul7Th+ta1yyGCqOln9pk0k/ywZ/IH9C4MuwHrgdWD7G8sDO3WyiT+fyBxpd/oQB2Dwuby
c/caLKuny1Sfr7j2+yXGyyoP2XjQCjSyJ63EaCywq4QrD+Y6xTseCVaWd42WTdyJHBISkUszDin8
gm5dx0lTBs91nu0MOosYlPrV464rgkdi9pHRR7nNnLXtDuQS4vDTWkMickRrYDK1POOC6dmwj6ec
ir6HnvwaQcYO326NxEXpme0AKVclvjHJFJpB9uBd27wAD3R3okwXc2Nl8WRBn5vTEWEKQpSLXEtV
GFk3Si3ez07S+RBmTtBNhWMsf4vNbCWLwEq+xbhnODYkj+Vn8nPGAe/mxaIYerTcOBzVSr0U1rle
L3RZBQsIt19JYqe4d78a6LEzVS4C7wHc/UNIGISh02Z6EG/OUPHnN9C8dJnqY5z4+AYdTI9YkKxH
CZ1qRoheexm7RoXc/QPPCnbLh58OZbjUKQ5k7a0qc9xPBIJ2uD4xEhuhR1zFDl/X+4liEjcwXOXc
NaMwr+TrRKQBdPzz5zPzf3ddBYi7T6ZfNXTU8tKwK/YclJSD/ORgcK43nYKrM+YQWs2Xxmsrd6aO
eeAiB2RC4cW9nJMLOaUMR8xJVx+6q7PlSO++EPwojLT0HV9zd5ZY70eUG/lpXBPop3US7LCjRWaZ
LTF4oN/S10dBKr+FIs/sR1HcDCpAATZ8kMIc3WeTvvNoH1VTRNNWse7OE091t5ANeTxIf6QdusDJ
Q2RpehnWnwhhXqgiKjY5eIjB4p+/+LkZLRFmjdpk7FbiU+6/yW1wSzBo8BB37GFq6poKfiH5380q
TzBC6tEeUgO7xbF2Ps6RVOz/UNubneYRFU/109NLGTOSEo/9fH2SbTINBKyiYXTthj2qc2rgtEqe
RwTL7jxuCILlGHdLqDusmeeCWcDnqEm3K7wDTwIWlnwn4SxUKScnlk+pRGWbFsGb7xFEhO5xTFi3
L0x+s6JnKxPc4ElxXPzJa8/p743sNNfsIvHS+gcVV26vzzNnbNfrzLO+HkMSFu4MO5KpUwZM9HHB
TSLf6xY6/J/MiNcmz0aYa9Yor6bNpN41ypXeDR4g6hwjXFC3TUkCIP074LSNeca9Vja0ibTDMSLl
GTy0tDbilOA4xnsPC+2t+jlh2CUqtL6O23xzfYWlVqg2WkRNDC4r9zbmF/+GTBy7BMHC6scoqz36
Wi1o5hb1j7zILhnRUbA+qs/AzznsjoUEaPcWGvCx7n7S4WniLYaCjS6uS4iOomxLAzQ0NMXMsi5W
2F8CBEQJQ+ytEjPuMUhjXU8KIw34CRSnokagNaSs9fz918yk0e5m/h9Lyl3CkNL/ALMJHBpdqyy+
ggUuS2HZZDK/CEXIInItx/WGThjGlNvoTW0Mz+MYldhZBYEMmUvhNq0NPb1dmQVbzdGdzv6H9gt1
dZeFEHrJVn9KZlba+Bz7fplVZykuJ/UDIGiW306ZwPj8cGoL80faFx7yLz7ZahPfayiqFfB/eezB
nPNKF+Tn0LnUMOFrkihZfpLs8FdaoTdIrEFA5kTcFv2UWgH106uAPsIlyD9B+USONdzxIfly1AbS
M9X9Olw23jwHFZecgag8ynVliYbiPqpdLREadqIeef2Iy1Tqv42MiJOgw6gCVsGoriLamYkFJ+Ry
PX7Wy1vEEWKJ72WFUBZAl6SMYsSmz8ZyhDWjxGhIAInIU8DjiZM3Iu32CD7/jrn5NRU9puHWrv8k
fpbteiD6a0tgg7HcPHazJDxhg7XqWhcrG+c6ko2Tv/QlEU5CCEkiVAqbwyHJY+SDXy08a284WLeE
gcxOK2q01+4JCkwDtz97MjeoXkCYAUah+sngeAw2e751ysdZSKbT40XeOpcMfbIUHhnQ7pFJcbQ6
ZCZ3t4Q94fM3S5rK+DXge7XQwEP5c9lsnCi/Rlm5wg+ty/XdeMJzK1Q2GiLGDWgl42X9NcxlQNNi
fxEAFM+mUD/eX86FMY8R+L+Olyb3rjpEHJE07Lw657PpopSQmyAVrX2SZTcMk4EBJ0DFtCq6z8To
y2PR4wnLn/gTXFI/DvoF/ETbYnWdiqNSg/QP3Exrf0hQQXQHx7Uor893ea9PEOrrNskivVgW1Av4
X+VHxIHCPy12CenPJOi7tGbQEBKbDzI9LfPupCN0+9H1N4v1uBGGyIVGHO5bttzv7W8cJg91ZY76
OoVMSDQM0ybEGzCQUjxn252/LiSgmbzjtHSBu3ItIJf4UKTmMAE72y+TXj9RqPghWRs3jBXkZ4td
58c9/Jc19OSRphBFN/SqA4xyob/OzKsqBhmbfejt3ExgTipl9+aVDc+YFgD3Uzqfg85GacU+YL+m
ET8PfFl+/DMf3dGD+TkYKMRasQPefDgZyuHmb/WIvjJFWrVXBksCvutONkKTXqgz6dqttXcv+exf
5Z/aoOZ0doUoQ8zcFF5F8Hih1f1iVOfDmnn1SjTTazPqqdSspdvK7DE1UoZ+/yuvinczqEkCabxu
Mf82smUcFsnb2f51lLW4cELtYIPE3y5NPAPjJq901EL1xjK7GE4mUNB4kHpbCxphTS+ebbO8U/mi
4XdQY8aTBXguAnzQMOD8H6gK57ODyOLiQk+uY08mBYBongGrgOFt6R8tWi4+H8NPOB98gKEgVbma
voqgTBm3EOSSiWuYVph/6eheazMPiGfNpVolcQ4ElRTXO6PII8rYOqNKcngT4IGI9CHpsfw55L6D
6EqVXb/sZqIy5mBw5jiB7TsnoO5NiBnOagsBDwXFT6c7NT5+JstzebWm7j0hLfnlLBTzxdoxPkAr
eupZc45AcKK4nzoWKK3matm1vxqrnHODcX6dgN8AiNPcsdliukO+x9ISlzPfN8i+bQMTbGG2RkrA
pp49DbJTFc5HgkWu9tbZyvu1exwXhLNd51zDGio7ArZ2Aan72Q3UsFS7lugETu+iNw3nPALWTNT+
3mq0IJ/3p2+OQ3TTiioF4ODQHjLb7cVA2350vlFzwoATb1RVOGhoJVwi0Pceo+mX824tLUbs2V22
OTUH5Q7LIqBU+uyMeHDgJN6l/0l8YFmV5xpV0OqdRI00FDo8bGiH2LOS7xmqQrNmX4Tqa1Z+WRyz
xnLZTLW4vaDqV06ZAPipKq9PeXyq3agiO8DiMTdLW8eHyj5tZ2SxAztOSljP5VDAfMHbli8QPwO4
lsIA+C/HK4E/gdJnhE/5lFP1Pk2j8Yc5sX02BCvljvl7WBHqFIIOPDuCEVqfNPv9IX4WkhEo3Zla
4sWWGTudGetheWtsg6Pf58t8s5YNtS5ywUvNDTUDNmfKwbz80IU0AdM8y9LIW6vF+z5Y2b47o/S2
2DllZqXFycklMms3qTvJyccf8GECT9famjcqnnOZphP/zIvfyX392qbBC+6tYB70ci5tBF15AxwO
r05rbpS0G2umz/zE3SP4LaO6eTnI6qZFgOl5HUHlR0gjLUAf3PdO6dPyl28Jn70M+U6lC5VjWdFc
jd8cgfvB25RuDHGlHFRlVhjO24ZMa9JJ3OXrBoU1Ep7sbJDKrA2Syv5zImrMH4f5a40hxko4w9yY
GqqNM33DsZBklhbZb2IathjneqP/TE48pacuy4I+fi/FQQ5h+3+1u5W4L7WNSML/vBYMtU80QiRW
LIp4yz3X8lFtBlbLnw1LOntK0qSifbGOVausL+MOBlTYKYkg2uDQ2j61PlPOOTTLbJzmR+mn7oYf
PuSkEeurXl+6KLTF4NAVhJyc9rsU/uMvOGqnmTIuDpq663VTipQDvKgNMVH7uG44KO8Dm8hf+O03
xKeoiJfgPpEp8Bz1EpICz41r89RMIjg35pL9clOaID5Q02P4/P/PF1Ryfh7QrDq769oy97zQh7Pi
xfJLRnFimHj1ewcpf1MFDuOtIqCZ98obfzo8QQkyvsmhwIt2o+fHWkmwFMrsh4oG2wdzJLO9Bu6H
9/pCN/PNMJ4XRHmE70uscu7ySI7mxmjWJ0BK9eLG7eiieyZNmGEqjUyCsbtOA/r8vkppwSkJoEb+
XMjdI+pYIvHe3ZzVTespKASyClmbzsZlR647yHgtgSebQ848LiMiMXMC+pY8P/7mwz5gxpaTVH98
8H5nmxyTAScFYBReONg8eyrVwBlTFdF3mJYw1teXDS6aEceYlwqdQTnbcLwLaNUD3O4/1OUMbqhR
tWUJzz6naeApHbKAOTb9dH6co96377cGOWVTCsDzFKtdhYuZRQ8sLFVAkCGFPCfNRU2g1NdUlqwb
bhCFzWhd5/5Rf8IAt5hIwuYqmrUXMEx3b2oDjUo1kYYUJxpvpK8+uqyVIOdkPkCcQA/vIL9UIzYI
s10RbF0i36rpuT/T3GtGEHW6zTfJjnRkCS5YcduVIXzOc8bYCRb2d9JC4HhimVp1of492Up5J27X
IYzClHo6G2xUHuTqkPDKaFsqSMQMJqCcFQxEcpRbY6gwFug9rIWvvptEYAF6KeeYd5MWYMj1hd9U
PaucXYq8cdFlDga486b6tRl6g7Sa7jqxuZvuvNMSMvSD/UqCLylAS/mRxPgwVUgH1quRK2KxOVDM
oSxPo4tHJwLT6ROQaATOngWX6g1X/VcEgE5i2ySczR/Gy0eH/l+C4MyKbX6ELSkzOTfjPRmOef7b
e8y4Y6QbOa1MKjIn6Ia73hid5DpjegwcV+atu4ztmhq0DZ6jP3VUB6ne0eZIY6dJdMl0s19pqNuf
nOmZlY/3gL6yjmxUCM+FVLClYhyD+0jAYnl7ysqjpWXu96aES/5UdXWWfhsTMcyK9fklfXidNh+U
IvyWtRyev6EDoAPlBaQhM2C0BJccu2QhVVngxe7T2QRyj1FNoKWu2dnxeFEdysNbrOFGgX9pxXnZ
JHYWXAZhuA1NfLf3V0npHRfpoUcryI6+vQtn1EYkozkWGs4ABqmLCKtDhc3SHnc+w+9izW2R//ts
/oimol+I5CH0+FlrllA940hbArLYMBeCSnhJRsvQtPLGBGsfYYOoZWS3hfGzvOWCKS+Pg0R27YhM
jP8BDmwKKxm6rEZYRGAiev95qTGZQFKVQi91vrRVR9LR4Q/xNTSwOymOfwiOf29tL1yJUuthcZ50
0/8J7ldGMKj8MUI3BWOn8SJv1kd7NmoZEfVwCmGm0dH2aJdjxalXj6UqBXoNkRDCHEGFSzOgVYF4
2liG/+cmD7QvPjPk6soTnAd8Gkmote0FfUpKn5KH0avRHbP6SxugQ3Gn103NFqx1mwRt8lnEDthK
RSpCGORk1on8miKWw3IxpCQ5LC0ncDbd6tyLGl2LL0GRXgWPMyqDVOQgbZlpbPyM2tSj11CbsfwE
iVtgm092LMzTAovuqkBV4HPa1YVdxUzatmfORHU3Yhu1t1Q8xQQ/MyJHnittL0a7nXJKD4Tm8NUP
yiENg4IWYRtvfrnEQs0liNovkVXyg+qK5z+SSWNEyFfiXa4P3zF7ospTL4k2tImg1COhfkfJApx1
Myzn6sfbXbUsxXyK/igIFIRYXADw+OaaNurP+NSdGLGo2aJ8wuFylQlpivA+Y950e1jgWRq/OLHk
va3NhbKMztRe9yyI4t9GbDX0/IQVPA5klCL/QuiEzA9rPKmfQwLZdyeYpWXI2IIHf/J5xUUVMahF
TlBiui2UPqI7Gs74KpYK8micrp9VYIj/4F6Xl8S8xzdyhcGcSKeJZqmCJolze5sTFAOcrmzTpSJP
yL0U3tncj6jUVd0+vUAbL+iEZkmiYl8pn1R510+wfQ2LL5HgTEUyv8rTUcmSjWd6snN/NQYPGWH+
0ygk9kAOXscKE4GwJfMWlEO8cjPvTl0t/cJdN4/aMvr+18VTP6SJ4ZOpkaD/YduxbbjAB8Wwthz9
YOnuFlVQZj0Q0CpsB1Gv/JHXCKOFypUo07fMQ5kkD7gdRSq6QCDUA3pekjMFNWojPFu6K7k7ezAB
+q7y0L+Y64Mvwg0bs+LiLcRxFuo69LBNVc42Sl/p+2iIj/frqFIcmBECVfKLqqOqsrfzghsb607F
RvIMBr0F2D++9CfftvStuBju87BYGwmfG0S+I4fvtSXxb/Lv6kirq0UiMEqzyVEBNEUxNGylBc/B
MJ8AFXK/uSBE9/Ym32Md/ZwxlrProp1Y5/Rm0fWYJVq3bjo4O5OsaNopVWf2hkqD2ZGnQg03bllF
wJhWKrhSRKhJVXr0CRsTrUYGkUV2XcO6BBIQPfQG1X2jJqb+7dD6yBU6CUzwr4J2gL+FNZan8WKC
oZeeUBs2EQrjLqFR6LzxR8i+9IeAwzAJNc9a47rqWkAxQeesFx/h8s2rS8yz8nA3VrB4VnIMys4t
l/0qqSnZnkWSPz5361NIrVs9BskbMY32nq7h+SfjGZsRX99Uxi109m8e70R941VF9K+OzZQByGVM
1LPeczxMXbAyOk1YQYISgWPlhmsWdlFCsQBf4nr9N0VMpsS/nXCUW2hiKKjy4L5lH14cu/0+8QWN
34WK9CvCn8Or0pJ2iJjBaIJr8A0fWhRWf4NMeuAAVPiXNIUwUngPGNuXBN1jUpOzIiW12PeoiTOY
ygN3s7vcPZ1DKx/+ejByfNp8XG9+Xa/dH66ICsjgIheRIruUiQyCZfZBiRk8Ow7VeoecYYXMKrXT
WA2f+gYr9GbffsDzYqKlJRBE9RW5Gt1ZAtVwU4gBOwxar18k5wLnvqSxhrf3cDr1yzkZe6QTaqD1
Qya+IXQecVZHkwmO5M1UDIYUXedg98zmdVRzy8D4+b80f55KL88Z/FZrL4b4SQJlirDVYb2hKE8c
2LtLL7KBPOGj8/RELMIEfumb2zavak5uYRlfGfpK2i/5RYOp29zl3q1od0TiEtI1Bj5hH0tfJJSc
MR8Q+/rvsAhkuSDEXGVBF0K98OvL3UU+YerySCrXsaD57PPE8AF//b8s5ke/n+0uVHPaQqB8Nf0N
cP3aK5GPA6/j7RaFdfGYTf2RvS6rcUgb6TS3KAZPGq+H/Mh6fpd337KJrw+KR+gdzqzWWVYti9Y5
iStymREZu2/RHkc8lvoYRVE/c948Nc8RT4XRlXFTFsgT7C6SjGIA+hwGT3ZUjYsvuc5Kh0sH1R3C
iBnkml6g3d6rF3XSndH7AMTaxedclD2tnrSZlp5Ix3161Z+hIyhFXSvQMU4Z58tI4eRR3DQPhp/W
Gr0tGi/3/2pJTFuGU7McWlyhEyiVNnypfeKcAZdIr7/xcl8IopTOyL15QNAnE3E3s+MzKS3arwHs
Htv+5CSdmIEQ7apS0rUOs/UJ3bJxjbNqRX54IRvHkg5D7hamLEPdOHqvP1jqzYLnggZm1ZLIprcy
84S38RovY612KmBDEthZU+nfBEab2QywNorzYrg69mEqNsXb55CZP7piXyxVb+slh7V3/fJqAoFO
zPaVeWrKLEOVLSLDXLoFdbS3Gzz6Xyy82L8R3b/QffLQMjmHqH0SjVm6llvIcaGu/UgZYx+7PoOA
dxK3kScfUW2PMJU4r/QRBnq3xeEwISTytamHC+PygxbL2eB+oheLA740jemwf5zYiQXOdhyyrb9w
7u14co9x3bbOrkaMe0VCsF99Bik9W+Y8DifpB5Pih1VlWPxuJwekQnwdhMiGwrNmRBJNCbziOlxw
90uaWtQSEAv6Ipe8jBSEpv+Xw0VXzH9k2i0rPhfHyboMPOL56avPMkMfDWKVbQ9L7zzyXhLj82eW
3x6EoJQ6SF+KBQ2kzCvnVxhTULuhHYENZW1UYTF0gKhqSEyWKOCaOQJHM7qw9LW1vhGTRSHt3XZx
4/zWHgIqw2q9vHpcAhNIZXOTf7sHQTpcRXEn7aQKz6XnGS1+8D3N5nsOZymaied50XRnlEmPU71/
7P9JUTGw1tDNba9gydhXUWTwvezT8UZjGXkIwvjSjm9p6JYkjpqCmXq5z9/ar//zuRRqLK3ieiG+
Xv/kJncWO50HturtwcTnGKjgdRup7aRHMebTEOifobnlCTy+PD48q84NfsYfQx4yjFWIhWxtzi9F
4TLSW0vOJUC19bMAqawXry8snwdZyIsYjhQJNDAY+sakIhkUMd5kBIldRdxOFwuzV1x5RBpAIYlD
tkVkdPJ3hjedPOUt40D0gJL/2AlZ0xqzX6ol1JgFPxIPyLHMP+/5pU2ues+lu8ZS8xb9XLnlwgvk
nEH2PzYiVSu2wETfaMZNzsfpgUS0BL6ttHO7ZOtT8CSSipTai8rajcd3yn7VMc+q/ArmCmhfxkTM
40H7pwQ7iuJOTeKS5BdKsyyvDMutvMu/N/L9NtzBWR5I3mL1+B3F0GOjMm4SBrs5FGI+KHJkrbh/
+gyiwoVkNxEI6OHFQuUt74mhSYo+7VCq/+CJ7QWpMCwOv0PjPfM4F+tBt9+2JyCVlkNj6iVIJQ+b
unq9IqPOv3SN9go0v4vPOwikl35V2JI8kCJBC6yfj9/yUXloaC91cx2a/mtU56Qw7T8r9KzAwu17
zBoO6Y30XiVVQd3VhQyppy/ko987sxu3HUaAbRDEH3hQAtt21Cp0RnIAcHyxUWKme4+/IvqkmxyL
xyLt3aeN+iF3wV2RU7j2Pr1HygEL2SFhRVmEs8kSY1BXPLgDCaEyIQ5LSt0zZ/jRS+VTPQ5onkFf
fpy3v0X0ybyjbefTdRktM0hldeUephLmx1ksX8yG8aMDuzgUY+YYfQFC3UlolPoCLRyPy0EeRD2E
iuE05zb6Um2uXATPHlZgu1yKYhiqctZcJ/YM0MGntKUWfWa6mrGGV1ygBYrPCGbibS03osJC6Z57
8IjGJszgt5XGy7IE9svFqeZiNWf4TaXi4ovO3z7pHG7Qse+G1uN1sxCB38FnZLM6dogxHWKmGhUa
Bps0OACsUD5sBZGllxX6vUAyWC7fy3Hdl+ofGJgyu6sPP+GlASaI+HESjOgDgFgu1d7umMGJ4s20
FGC/yseHCJVc67OJC1chSLLgbrkVfVJ+ENze7QsefbBP32Sc5JC1E8Fji7e0579EYtuXWz+AzrTJ
nNF9tuSA+aTU/pjQYiSckJ1eOyi5JZcS6tDvQZ+muTf9EogghWlLom4YVYbp/jTKHYG5M1K1qh+6
YrvaF2dxPhXublpqQ30T8oMqjFBfnneFxo8H8TsyGAVA9NZ96e9qWC3gONlVdoKNBGoBLyp9t4In
JfHjtN6B0/3MZkR9+mtUiM3Wive9AmakI8+MNCn+kNSPdiECi4mYpAShMQNBMWmpx0cTFuTaLsvg
44+4qfc1l6lz1Lp0tWR5kTph9c8teB5JYgCNfHPRvdiNrRqEx0tI6swWqpfgagJNcluGU8Har2Gl
azT1jL+xGvhqYq83z9FwWqkm3JrTqRZNxaV1tFz3m7Jtfnvu8sTSyPh9/vOx2ri8f98ou5vOdJyd
D2X5cFNDzGHWCe7B4V2QxOIpRee83vblUdWypZYfQnsQC19lVPv26eCcn3ks42kHXOCxGdigJiwy
pYlx9QMbBa3Rqbb+8H9eMovFIOAkg5Rt1u+PspGlpUJTfGJDuRbriOeTbR+VH+gjFyk+WLkYPhIM
WSL9YUcOSPW90apqUtZV8ahN+CpwP2gNsFfv/apmPDnc8CHYbGZISZt2QyyqUnO27+/ykQmmmfZV
v4VoqX/WKmA4PU7m1R52Tv5jgtylxbp39VSeq5m0a82K71aOnSBTfeUKHQ4HlWe6iHNuxeYo2k1e
G5W+IHQvVd4anm7H56LDZ+ojKtfCjW3RyDHIrSxcaKmeutogTn/GY8WIMGctSiUOnxt+KzXb6JXY
QkpS2rbOlZbG72Nf5LcDqJsKag+Org3uoJhq/7mTte6qFjOmw8Y9wokDw/+5Vo8+SQkegrAW0rxK
ImOYkNJ0oiCjsbUyyfSo6HXJDSllersBnmsT4PmejCs5RyI8JGzgmjZcBWe0d/s4rOGrncOCfp8U
6ZDlw/8mYI3A8wqHXH4HZQsK5NwmgVgFyPzLDjXfpPZ7fgIZ8+V54XIYMLu6l/zf8rY4ioSRJwJT
rU0gztuB7EFFDsCFB5ok5Yp7AIoPYx5ZFdDDvKQTrsacIYwmz3+ToVJkC8WzExOrq2jptB6cuGRR
Rzp4pXMVZdz5XT+fjCGGIGAMKjuszQrKsGvcR9+0hmsuv5b9GWP/qudZ3g6KHzAqVslYsbhjlsG0
mHQQf9mma3GL9CJSaTQsFYNJM19jEW49ZfNKSDGEF6+ApbhHY5Yrw3RPkN1lJLuHTfwnb7ZBZAmt
m8ZhZMYt4yRoH8sZtcXROuPH0zcnWBZM1CAwDwYZXy79aFND2/4FaOB0xT/gTwfGSLGALfIVVZza
pkmjYwbDE+T8WSt6KtP+7d3aeF04IdfjtB3DbKZ+eVx2xDxPOmwFi7g5dQxs4vc0yhm3YW97WQdb
cKnloPZZ7aBq5B/z4bqXwOyEkymyHwVIZsFQgYuQcW8P3kG7Lgxna0A1NSS8FCeN6fetOOjAEWqa
s4gh3ktvstmCyTY13KqI8qY6F4DV0CsoHLEG6A5+8VZIq1HQNBh+uUbGrAP/qlVWmNCXy2vHSp9p
MIlAlRjgUV+KbGPL4aHeCoEGvpn0j1UdXqzifGI0SLyw+sbUAHPgE7TlhY7Kimn/0PuQ3il9VAHD
vympbpDrVzmXd0RnAtZxuMCLN0r7cukJ7erGOPFcB3UjL2Vzt61qm4FDWDezQH45vJZyXhkpihvG
57lgcLFzaFmZFjOuX6da+LqLy5ca2tV3GxojwL0ZadI45lRtRLJAEGSqFKT+ZlewvZoD+kSSCmF4
lpBnJ6h+dz5GQqvsiDOVMp7bTOGo80e9xS4BMpNp+yxcQd7wgUJELk+w4qAZJmnJQkqyMcWpNdg3
9DA9yho660of4FvtXvKwd+hK3X8y75++m7MIsV/5NIbmzrzUvCKyjo3uoWt74A/C0umKjjBcIt1j
ZA7ACKosg24zWLDP97xSwFqIhb/tbtJ6zk/cGXTn0T1A0al4Fp+dBSEXLfQVXOpxsC6zYaOUSDmq
DnHYXqI9ebK5W69exhoAOhzOn80bwJNOGFT4602+8VGv52gtB+wP9zRZd5cHLQSNNm5KmMVjj3vo
Gg1SXR8CVCZR3gaenJPWz2Yx+OQlzZkXnx2sMddI2q9LRUHhma72fCEXIM/YB0Q+6sN/BRFpLZu8
RNAVQDyC1R65+jIsa/iIxcdAK4BtrF/iDgNeI7jyFYT9nzf3Sm+YfdJgLFKO4i56+pFPb8SUdgZY
a1VoriulF0orsQTzUNEPLdAe7m5yJfZJRoKeSQJZP2CMH9dzU9meIIODFs4IsxCMv7Q4po2jIezz
NBY3TQnD328H09xWBIepYRHGnTBB9jvp1Yd2P9f/EWoNW+46MAA0ZUB8n8G9pAUOxX+n3OOUlmbR
+WtPG6Y2yx6LA8QkofolwYd34YQLqcK5ImQdXjlxTGrFf6cet7ss2VD86a2hY737lBmahM2E/kQ8
uJ3KClxmMUAarHILL+RRj7NgFhTSHkLhQwWCTEv1H6JodiB4r8rRpGZakOFdlybuJisbogWeg1Nz
rBcCrkbWBgikfsUK7cPWIxSHpvx+7R3CRR1sn5YMWRKq6mKS14gO4nqcIL/kwxOLWBoPtT87rSO/
Ao2+CrAalpebBThrTUvCqRe8Ex0ne76Fo7jNpKGuzV4IfZQXKWPWCPHQxqOjrThOKB0wCVv4fqL1
V7U7bCuJ632fcDIvyZKPwCdX7nem1rfH40fuVahtcO/r+E/6K6dBFOQtzwRATmMpeGC3bN8Pn2kD
aCRtTzZ9dhTkWrr+6yzWipOVI9clwti0+hzo5JPy9kewnljrrYkeSoAJ3gJ9HXJZS4zBWfQZ3LLK
ndUQVF4FkMw6fjtoYn6jiR67W6GK6FClcyoLCPvTzmf5oLlUZCHP4OhXvPHiUiVN9sYI5BpjewmL
fG3r73pt9NVJeq5yWRlqhZJqFO/MWHyZPclQzzchTsqBGxTesHOMFF8Kg/73YhSktvIFIr3EpMnx
A/EuLj12HOdqFPxj/2l9xbrbz8a/1wo34bUpIdrQkCAVJoEiuJyAXMovsJbYYbMbU1h+eOs0u2xi
MHbQl4wzP95FbQB4Rao4p70KOKn06tzuT+JRE5xXjXjLvJQXs6SisRr63wVFPU9lGZPc2mQ/bHnJ
ptNvSBJptoLrB7Hbr63oIjyqZRJP4u28ghGHuueFnrRWwNE7PFpoV2ZYfc5DQY2d0k0ts392pb6l
gc9LFOpPxkvYSzJWL+X1Zi0g5ApJYQSrufSTQ61RGYd2xTTtWoD3rTI56YdiyNnDaA6jow3b57Wo
+fN1Rw5kOMJ8dWGopHBwg1MAcHKTciptEnhfH0a/g2Lt9CTiLYhVKA6iucqBqXqjCPfbapmzkEb8
6ZebZO4NwAarIytOIICHwl+pCRsXBxXVzk7yDSQdE+H3ZLlmHv8w610IiTANPelJt2J8khByGS6/
Ssk1BVdEXI+/WkavtA0daIMKnzMDeXeQNhCKNWmsYvie+j/C8QlEhlfkEz2JwPwwRYRp43om3Sx5
mO+uTGX6gJORkOPeDwnwrj+UfF4I1RqJxiABQlrYGZJ0UfgHIpPg/CJ2Z8nb5m7V5m9mwPjFWwvC
hoHVafMYgayv4PW9uvHdtTXmPRsdgBdNau0zy5S/GFayluUNj0vpu8PEDFWtsbdmT19bkWpHumuN
WhNsdfCw+6QkAOmfrAb79p95TEGVpW4yyGHI2XfP2cm1t9e3vNVnMrUGs9PfzPASQlk2h07GehkM
EFUxVCLF635vghQwdiSzQbxGMBrbAqD6ydTbiHhCOhd9AawCeGsq8mvxLLnlzDrtCf18aXlcb3lv
tx4KH5aROzKSZ+EBWfDsWN3eZ05K48ac6ZEoMwlxad3CbBwxLdqkbkE6Pf9veaCwjRNmHzX1CZia
x837xpcOSsv8Wlq/991qaUFO2xKulXxXvaQ1kc5ernPvFdwXuqRoq5Hjtco14n0hwC8jzpm09pYe
nf1ypwoyydaCZCixjuq80uLticePCqhnsk5fDNu6IQnMAhmMGbWlWXWiYtW+3yCXANXbG9Rc5Hy8
eBbypd9gFDaH8126VKu30C2fdWJEcdI6b1BBcwImLO+n5wQnMA4diTMISjF3q7/S2rLxctiTcCp+
lu+2booE6GofK75oHO2n1HX+L8/6fCfI1O2FWYqOcnWOSQhvcLIoYSh5T1Qn1PuAKVJyi1nMyXhf
w3PO0eR98YAA024eR12c8ibN3e/DUSoX/CcI75R9uM26JHnD+l4zSIx4L9bFc++TqlnpHgc6Mh+g
M2fDizOeHB7ji5D7p+yB5zy9lMHj1UUC+Z0fs9/n2rfNOBPc9k+HHPQed1O77Nd03UmbYLNPMHJQ
lPia9C/5/Xbth6ZFrdPFwNkQC8/WffucCXwrIyCOXXsZmMM0xznFkkjHTrQLIGKhqHtEAf7oCpdK
B3cCU5/MMtC9rUZH4DoxLH1vf14cgRHaPZteC/QfZK8uGgHxEkWPUn6N0iv9T124F2Il8lWVf1do
I0AVxpapUIyZ8luGvnuSNezhUISt5baf/VRsQts6XlYKyRR3qgtQ44rcvTRQ4/jgq1xuTe72XuDX
20iZzFBeGXo2gCk/pKHlMq1rQb0kThOjV6aFX1mBMJu9W2DC3KV+ghX/DtCllavV/d1YEK/+d3lq
kotImPHYWVHTDwbjKgzpCJEjTwrWAaCBXADm9Lw+oOvr0w97mqzsDUfdfsUK48ohLHVL6QEdzxHe
F+mZ5fZGP2hsQwrQtp6eK0+NfJELuvJV6tkQnFu5JiV+TYOgpIovVuUX2A1SZyhV/XffUgzUUswF
FHIi5Nt07r1KNOtgBq8duDMbiijL4T4ysoRmUZHW9Qi+XRg07G8XqANnd7YfxZWtMcpBzlahAZY2
x+7cw7qYrXhvn02z67QEzIxi9Gk0QA4hN8+Sp2kJsHlO37MPCWlnzj7OUxMBk8MdlXrOTfenQJc5
e9dj2gqNzqvQuG0VYi3KcV4tS7T6sPnQfZP+6A788ndwbIWGddxVV3mL8TCS1NIRatLMFYo4k7I6
0mW3bRTxkxmc9+7CC2cAcmcHlyKfRf0HXGl+po/byHYm2bQFYHNVjXXkDJDBNd4fDy7Q7fJmqbBX
zabbD4SC1PL+ZrIswvzlohutfIQQt9IFBQFXsUFi92M62PsXnmtOJfGV4cnHSE62p0tPFWIFgL/G
NNCnigUL7BJQPNPQorRdXnCoLzLiKi73cGhKK+TQRMIy9pP9+IUNv6UeIE2merlGSg3nKdE3vcZ0
v9A8u4Pl5uXVhDhDTIRi2G81XwkGl14v2Da5r/scYy+6bPb7Qv9u+Olx7HN6T73U9egXyP9nIK8F
UHTS44BNwLZ3N3r5TM7LbTcoGPtN/hJKzKFQxJ/Z0wiCJjoCTG/tnXfqUF2wcupkdjT0E1M7Zq7u
RXvMkGJNSgyRCuZMegObo6GJcb0bj4qczBYNtcI6sQAPKKnCjd6RcnqzvnigOwTm/ZiBo89uUADE
QVLXO/yy4XBMpvM03i0eDde9lPdqBV1cHsFn0FSsNfbeakJLzP/UeyT6NCaEUazh0J5SVrWNrP4e
fDybUSPoPP4NbrDydkjIHA7ZkYBBwVRLr+kiGUqHEqsm3UKuvPR82rJz8AMxhbmPLj5aQbuY1yzv
KZlI9f4l/uqlQDP61QY5ESnJ/ZcWWAdKhzgwWDRqUmnMIrzZZr/c3wU5MHEL7aQbIMip8XCnkX7K
XhsWcNtf+Wgb1l6T/C93nKOT629ylKEc/xW2ULbCUUJcs3Xz4kgX3TYKDkwShSeo0hlqUDO94Lvl
id6+Pz9wVJkAXwMXaYbCoQR/6u/heJmfq0xD87cwfN0k3y4Ut5fA36BHmELsOf9pqa80uGQixgkC
AnjIBspP8eELEOussqFuqgHVCvh3DQ3pgsFk5/YSFJqxsGc44kjxncdUhP+FQR34SVwgHEISBRHl
rc6PFYd5Hwii1sNxyxMA04mtP3MR8LmTs2W24tuxypneYvE2JB5FyUWVrn90fJxdEV0isv27OZHY
DfA8+dQajyspjXh5pU7jOe6ldYEN+UE7kYgFNTyzhqfkGDy4dVO8w/ytfggvImHf34+bC+RvyVgF
WHZWk5jDg9+qN01nLyS6RpF/cJcKFD6IvQ9GZuAs3FLX/x7VJHHmNz61p1s4Ga+xmo1h0g6C8Y+J
NrRRC3uj8OR8obEy1Gb5wCmR1EqV49vaZ6ujuv/hLeX/JtimJRYx8rqst/nORoPujAGEOT9JAq8T
hM11o8kTk4+ZHvDW4dnbSQWITLVbeAMO6A5YV31ZwnkwIPsOrnjXaKS7RscXa+yh8sadltH6lDru
42+/x6U6j0Q0vCYbvbH4Or9+qVWzobNxt7nM3cL9FM+3gv5agFtuP2o+BO2Yq43o37aCnpyZG63L
yxI93yFDXucWY5b7kaZ2vLi44s6pn1XqqgxwgYni1eBwnHWymmgGYWC30wg08I+11hKU6cSZFoc6
bDhxBYE8T8NDpTAyEsoa7f+PKXFTWpzY//XTfXCrtxzjR8YT60ueTlVJFDYFhD+rArLzZZAvTZ0y
PG8nskOXiwWVgow0EQOy9Olka/SBdBAyE5G589TdM630BteX36krH7i0IDdOr7qfM8nWNDpRUtP5
TQRh2QxCXWp/NaslqNrRZMEOpbYiCWHng960Asq+KWnoQAZjqB5m8en/USDjjbjH1YLgUPNSOy/x
E8Y78GZhpE6l6UhtdjKqEJYGY/VHWLyaAG+DDzapgF0Pg6EdfPkUOq81ZmQ8D2ZHUxZaKJDiDivJ
WYi+FMhW3EvDFkSfJj+7kEAvmjI8Yvj7gVHEgX5Cw5mvuSaf+XANe5TBUszLn0Uw0FQLLZyyk4m3
fhvgVckPXQCcyOaDgDgVgQfGJA6oQggxedpKUpU68zwAIhAYrhIxSvh/m/1c0gLsm17OoKpQtUwY
nE1EtRvG+MpL65IfezHGRVltwwz/jeqmDA5hq4KpQTfLKl2R0Dta/4L918pdMEUbppZMloYN1xBF
9XCj8Xn9XCbPHKMMBMydq7NgUzMcUcYe7ss8A9JPKTkkxm9m5+ug9NDe9ZWZ+O96omTx8CvNr/sY
5xhTou/ytT5W/NrhIE9Glz/QKH34LWICH3QC9p+S9IpJiys/pmbJ3nYO61Z+9+5Sj74nhEqPzVb0
pVulxUzvNZ1wF4TvWuEdbB3B4lobji8fiLJKtO8605aARuYMJ89JnBt32m5p42nSl1dcg/UIcxxA
lOCdFzauwxXpRC9YQSlCUwYZcvG+erYYIHNH+z+J+Va2rmrZQ+jGurz0G026oRmj3GwN4uh1sG1N
Dz/hR2mXs8I74JZVjGRif8+R52QpELeOUeREIacJQB/bGpIrAO+qMG7uJqenaT9+BWJH+6q0+WSO
BUggX6rHH2DCF+nEiIw8elzmhCIG9VIg/2XsgDdv3JSc2cqCllI510uz7vt31sY7ut5VhUQMUalN
Q/xhW4pA5eRLG+gR2tJ5KoS+dfu3JQ7EVCLebkhmiSsIqn1BRT6Vx+JAP1XRcCDmtRgCYjPvXmla
yKC9tyehU3Imx/YwE/kMgKvxbyEen60hGBGK88+ZdjH0CmoYksk4aOf0ScFaSrDONVOY8MratmYm
AsipVIZpFbwIeNQqUl9vKzAK7TFmHSAoPjpIZ/7+6BwyTpDM9OTPtfDDrrl0NawAgD3UIFpFCaWf
qmiIjg287X94aKZC0hQeaVwbLVtZ8TTxDWT+gO8AI8P6ufeHpaHfha6iOtSmtUxmIXm+lCT6WiXa
948lTRli4sxU6zeN7oF2XepipqDUfgxU7OSixeTRHMp3Sr9q9QMHDd7/puQkC+yc7NdP+O5SP9EL
VJmH1QVwq8U+DCMICvxOHoYZwIpt3+YvoxJFqSLpvlu495/WoMkwBJ6S3aN9JQ7hNXlmo0QGtdME
XMkuBo4OP1UN+47VGqpAGWHZzlwLxaTPE1Svdj790grKSYKV+8lz5PNqDhZa6lELfCG1gXOJ5say
FUeYm88as9GH1fhznHmMyCzCv5hAcxIwhEuvSrlV1cfhqB6ZwYvES5h0vZcal566Mp6xyhs9JyOB
sLyK3CEJMRDzvHDB1UxB93kfvjUwfmhApiFyDmefWxzBKQa/U4kkh0w3oQ5JxsN+okyzRflCCwPs
E/IHD6xGyF1eYRvHp/3ztthctT5QrvvitbMfEU4jSXv0/AjGPLL9gv658VThab+tj5Qb3ExQi18G
bTWcVsFmdCgLNfN41gI0tp2e89oGsX7acFgoDlHMqg+/ipMpW3cnQ8wjKXWo/+QpTcY8wq4oKOT0
KpmQad7hrDd+e+3100DcVxyRemCtLzhoSrYr2BPqe+7WjRnAL1XJSXqHIrrHISpGJIUBcqRZ62Sx
cu2vknN+qg889SP2KIqnq48c3dn8nVJiS8RI9dck4w4zAZ2CDP6pFq5tjDc1pUVPASUmBEa4jbrO
vMEjBv3lj3BYgIfMR9O02O4ISAcKE9ZwYwyQfSQndEqEBGLU8ENCWyMWSE+dq5wX4Md8tLI3394x
rd49j+lErTx849cbGFKIk1OyIYRigNqOvYEPKV1f/t3FBNUspMBTyYju224jnwI1d1dpeWLKVNN7
ZWQxmXoVKWPDGKASN5Q6C5x9Hmd8u569YXC7aKSbi1BVoP58+wShtaqmR/AJFECRuvg/LsujGslC
0/tnhe6AfCdlHeBnQtFtW6w9TzYJEdznMu3vjW9OipEDHSdGsxC6hss5OojrKU+JZBXr0w3rKXL8
xwGpcNX0hy3waldp31H81NZ5naJo4y27ojQQSBmE73l8VSNU/y6S2v0SB/bM2Dvq2hQtzc1QN8m1
TLvM1OZc+UP8Gw8HK3vrDCAL0m1zpFIYtncb/oEvll/S1HbLKaNno8t1SyiY+I9Via8hREsEzkxk
YVxSM5mzwGAIgWjqReV1ajNqywag23a6kmQPHwoOkqx/QOZtSyYhd2NHWRi5z+9A4qbKh/SlBeHz
mjHYHgGo0pCy2Sn75vHsr1M7wtNG2t0tI7x0f04SZFMkkguAoiEJJiumxmyhhPtRUOov3EUJR1+Y
XRm4jp6vy4PYbBeAk3y5uXYTDHh7UyQ6cRtdN84eMcjMPix6DPA5HcHoUVUu0yElv0gq3fYLBORT
wr6s7uOe8Rm1ybI7pQ9SeUIwSutq9zDdaOVguOzeWX2qNyC7V/N3KMKarF6wN78dMJLd7+mTdAFu
XOR9SOgeNq/eTX2+/7iVUE3iX63HrFoZnHZ/1lVM6Mob5oNY1cb1S1h6ibhPkmqGq9CTP+Bu4UJM
YPlDOrySxNNJIzzHz751oDbxGOVaIKsuub8Kjkry/rDcJhKgjT70+I/Ylsk7nmw5UyGaVdFkuHnq
YjnSEJJnlhWnfRbPpb8phUlDo92jQs4zY4ESgWyxXbsK1PHUh/JTjq9zHGyAXmlBQYYbFmKFlFuR
EXNyl06jVmP0ZupD2UM56YbB+A149mWrFAzIAXhIY67wytCdJlYkO3jXtccUQvsIVZh58Tixu/uU
P3uWruOaamvnx3VUDz/uFWeWS3kBUn2F+kaRTqIJbK3y3MPuyteoA1J/gKMKoBo+6iLsu9WQSAEL
yOKGRFkYPJsyZipj1YBJTJfBwC8tUjR3POuvX0jaj3skB/jwKoIrDsNfVJ8eek+isMxU9LgKv2UE
MkCxuKSOioH6pnoc1mlHIpaRlc+E7+jKMQIzq0R5Bsms4uv8QwJ0AAAZ3T9Inc92QmBQKP55BeTY
Phl0ZGCNq1br9LolM1oilLrjtXcrSKuzP/WuOK7j7UfI/+fEoK0lYNmT/SH4CvHoMRMChJJ9bk2y
DZnI4cjQzt4DGkP43kS/sLMmT8mvW3zIafSplRtEQNJPRd/TdheVfy8dT1ucKzItcB4CmlNrxl/D
MwKRVUGf+GoSl7UeekyuX2+vDQFbvf25LBVvXdwGholDreKkWDvd41O3sXyRWH7zti7piTUP5AC6
8vHSgZunHIAo4tJmK4ehss4pmpoERf1LiCQE1rz8V7F4iZxoS20Ev+WwcSpC7hq7vQHuWb+/PyIc
SxKd0i/Ne3eVDTq/RSrb85sht40QwYRJItalOJHPrN3NLa0Sc8DqH8YqjsD75MHRW2SNkq56uhQi
E+qK5anhuOPvaVdu5SlAdhgMI1dj8l33NIhQq82m9O/DU1WwcL2a1mtNcNW8NBE2JecRLa92OQdm
/Y9KAmJD+9iiPQSroQhwV3WesJrOMLRsvnmum4LdVd8CzscPJ8eB4GoRByMjbpYNI3VjJ3bgQ815
Jl2CvuUtU55L8uyTKx4hA+72ybfLAGmew+TBi3jv02RFAeEE+9dY77Uh07TDMEIpRoc/4GFa+Ve1
rYIVwCh2xDPl13eQcO57OZEPaKmv/5U84j1ipLvKG562THCvlSJo91BH3p7a3aL93kzYZudgsFoF
oDJAeoveGBW2sPaqE4Fs2wJ51ud6Ck9UPdrc2XtnqnOTtgY2fgZVxqGWwGe8n+lMUiQCP4qQP67l
bZfA5bCafMBNc/1gvG+8toM2caiT3b3nLcUz3DFXRf31EV73UJPjBOBJEs0GoHCvZqssIBcAjk8s
2/UIYRY+ZAogwBESsSOysyeMZyv4iisoweCYuzWg4G5QpkLZ9XcaqH6v5if1ghh5pX6d0vw+NOfV
ahHXAEGSBjTcAglaCVM2AzlVB37btrTm15YFgjcNt1OPnvB+b0KyF5v5huW2DSJFUeKKENojWT6d
Zj7IXvaBmEa8MhsZnJ7MGPk5YGcpNl9ky6kuBFNPv4ElTlpeU/Kjt/PtWOHvK9Xk84rXyULsJTn9
CaY2YewMpnuvM0mM6NiUMWU7xJn03IpEzzkgnLhez4QD67uPQXHyYCyUIGKnzGDjBpRkBBuRmerf
OIlcknVvO5CSkXScwLlo/e1soha1w1B7A4KTPGSBPtTF7XP7AnZM1b0q/zdVWfElU7TjVhRpBh9P
Yy62YlS8bkC+UG7SfPCpcuwHZp4VMtcA6rhhK2nfepSI4w2E7nbu5AK44cLTgdyecf9GtHuo4YaA
9LJC8dBUUg9AGvZvWZzWGpzs9CAa0AC4tyQsRmLy8QPENQa1afCgK2iihcWxTpQ/HubZdBE3mwir
VA26T4FlKRwywKzv5aW5yvk1HyLuA+k6JjizKgrfqleGuJh2arGyQW4flH9zs1zqc2rP4xhg4N86
DviFead5lG+d251VeFV02RV9dTI1wyXlZSjBB9xEcg1AbW75yCfhekBa1oDTCup2Cko78Rkd26eR
cSqwQlw/G08vmPmVlZyMyOioIbikTAhgqknOtdIe6yH9ch5jMThNeRsBnyqBXIz6YejGNKYzsKMX
1bsMv7RazAA5PWhIEM6hVgUDQBqYEJ5auNsiKCGu3URLfJv1PDHk7G3KHTL4/xwiscnf6TW5D+7u
X47RcbVLOy7b4kkEJUbuszfXNlrLnf7j5HmqYMah/N7ruUNaZBq7GJeD0/9hkz3ZD764rctbWSo8
trmY8NsV8xUaztkB+5/oRd+ZV98XqMhPPhbjrsapvJLCA5CdXLv9HVZB6i4lXfAVmzttEzSKqycJ
K+sIwqk/Hy/9ODfsyrQxaxS12QQjjo2/PsE9L3y5fcRZEwcvAw7gnzNjr+yeqmeqOlLqJoFIvDOK
TtGXP8xqcaWX5M4gDz29wZ7BizpWTxHSJx0qLv6h8tpr+Ujd0OFvFGU+Ts2aL1740QTAkOMq49P6
aCwBYByxXi/Pls+WY+4RQDu6Y4yjXtYxFCpD8YsNcj+gJvXMh6zBhyRKH9+r7tXsEZpp1I+J2UvG
JwDKX6rbRvkg7eZuDT1wSslOGdVlOu6k/RgiCLQ1XiXit79uF3PpWxyaNdUBGLD94OHP5+5hr6nZ
yA/vz/7CV0GBzmCpDZN0tYxbJ0fa9egKtljTiU54qzdQKzESMNdady5WR+vwYpXKEFSSGSv0gCv8
PLq7hBTE+yx/Dj/qXyjpO5whDdej9xKf7Kmc9iLjT8bYOB616ZbY2/tF9uQejNkIyqL5DgJe9wHS
fWn3uexEUT2dvXncY1fwxHWD6ZuJRBxHDeKQ8qVCVkaUf14t8QTddiZ+lx+Ns1BwdCpHV6+grq/i
UoL/OiX8kmOFxSu9APD+nQRHjfRcZevMIWCzMlv/3VOs4bVkBTkgyj4xIJqAckhUQ9Ng4y/2XDAR
LEJbSIXv7UD/yS3996o9igD4mo4ejvDcovJn94s9EYq9V7tZMvPf3BGw3rMj4Q72uHGxvJ7QUkKK
fKoQmgI9be04ZxOQbBrP/LAwXdkubn7ahfsUCSToLRgJXQE3nmeInYzFcNVMrXMpIsJqucN+aHJx
8S2vNCLgak6RzVkqdmxd6l+MIKXnC4ZGrZ/JmCs+20ki+P7x1IP5/+263IggQYOB5ijXKjsVgXlQ
eDHMT4G0CfcQH9UqQ+TLNsXDSZNI6+vlm/iV+ruLx+5ljYI3ct/D/pPdKtpPX17CG7HAiZagTbay
YKWWXbrw+u0/i2jSl71gTon5DBy+qDACOppeGyl5X0uBUDUMh6PtYwTdhqJLSGnFXLgVfomHWyn6
20pNn5/kE9sn+ktG2DGl8TMv8vgJ8VUXlseBF5tiEqVTVREWMYnG4gpHM+rgyu3+BFkvAbugAdj0
TjmRu4TN17ZD+egELEZPA81KFk7pZgFx1PrtN4zjGod574z7e+3yhrLEYukQRiDa+hSc8++hkhJK
tm4NpR0rqQwDFU2gzrmxToE7jqO2Amm1rkC6V8UiCs3d2uPo3Bb2IlNqugB2ppff4pellBKVGOq0
LfYvRXrg7rAlZ1naMkl4U26bsopDpkQgjP9JI9DwkfrjU3LzeZ/M46bRek2eysIt92yZp/j3MUGn
uf99dwHhAlkA3bLYefExYTl/YTB/4l8G/KqnBUGeXA159Q0rywAFQbENDJCgq+02eUNTVEuLrMIf
aLKdot4R7eL9ifxX+BLU7xFT8YyZD8FT+ifiEXRvzMj+awWnvvUdnuQukugC4sM0W8gnHn+gGfHL
R8Lzy1VlS55sljStLX3Of6CyGANWj90ldv0Np7Sx90lrf5HlhhnDXYRvjgaV4jmJNBUfkirgqr67
v2UdctAFVEb7maxrIwrIJGW0CHb4Uw268ZAPA1ma/T3jfRcOsRcPQpr6aTBCn+04Co95Db/uNXyY
Awrzm/9ppr82eR0XSTU3XlrINKd5GYZgh7+QF5Wr0SCfwk8gBjIo86Z6ND2Q+gUwtGKBMv5zPDb+
nwOF2/uiJe271udJWtnSD4y8lKA+OQ37ogdffcKiM/okux0wWTBJPsGzisbnxhdz4FbQp0MSnh10
QK5ic8hjMSdsr68r0rvA3kU860ms6dy2RohC6UKTSaCRAA9QsY58x3aR4+jF7eb3uq5hLgBRHAqS
lAqPXw/BgUIQjRv4K7b1Xkvwg1gKUt8ojZ3BAKgpbxr/tYJCTujjtBIlwamvVgWooKj0Flg9VfjC
aigK6AAzIV3e9/tRVHga4QGl7cBWv3bUcDlzTSjggX6p1BX6src/UsGK/YtBLCcLmrUVu0jSUarw
ckHgcgdUAnKdOpSUlvmiQehOjIocQT+D/xBffa7Nq2dtIowl4nVEQ0DyCtU2rnGalAqTjixeV8az
g5pNRYT7Ac73nvqs8yP3qouJa1JM1AyVY6i3icGYk4KT1T//nFvvyHX2PrmA5aemUTuZ/5HzwER2
/8I4sue8XlvqadsnkpweP6c9Ds7rphJi3u6aFTkMFiygIzmMuqMvaAJubsRRFc3zSUV53rRCaljv
yIHt05BCWQPva8wNlzIeiFujFQt5NyPGviivyhMWh7HhBGmcY/rZoei5AtHRzkxHeJ8aUZP20oCs
XanK276w+7A4Kuxx3tUq/LrDxuEo7Cbqp8qaPHmKszrGhNtkk+BRV/B40PZuhaBedpGj/02Qznwr
0vTSbEuaMVtMNrDm1kRZPseEQwr73+Ugju102oDyA1XnmVBBGhMYIP4uvL//uKIfJxK+/HUFi2OO
O2F2OVM2u3tiLeVMoNY9R5QwzvbkifTYBreDYJnRDLeActl3SBytip+VhXGW13VG4SD9lF+SPKkG
BIvH8zH2acjOoqj4iMXsqs1HrDU+ojHuJGXR80L7nSaUB6anKVGOFrDlKTUayIdJxirAsDj54NLC
q0cqORMVyO9aVQrshtruirnWT0RCOAVSI263xh8V6Sj80bBelfilQfPHyczEt7JT0ty4FnOFxZPc
Br+8dML4CTdr9JxfNf4RR4cuVkGVrX08xka57Ia2JDLldL6MwRyVCK0h9el8ECQ72OKIGtaL1nPp
FayDa7+nVNIGkpzfvJBIWpw/fy4jzeviq5+e7/FoQagzc33a9pY306I2NRweN18BOhn+6n67ur11
0qoQVpuf5aKjf5Nu9GPj6cIthneNa6/ZKBKdfMnUrCgLrZMMWXTrmiZgjgKxFd/ixjpOWFUndtfS
plGHnKVmdzlun2ROqgnmrhrmqtSieE6GWmuREf58GZo4lWjCpzKjqr5GqlKOdZJanJka8YZ+nH/g
twM589JhmJ/7TpF0N7y1mzhKyW532Oz0pWe4nYIcC0OYOmzdYvu04VXssPlJE30yh8cTyIh2dPtG
jjF+9NDEu78GuW/vxsrxBuR0x+qlgyqjBLWCh0lNz1Wqstpllyn7fCmgaUCbiw1mPtXFvGEkJDO6
sOHJ2hHIwGup4IWAZr3PV8Yw6neEjEOzEadGc9xAJPOrzTeSUNqNQ6PCheCx+rPRqv64wDqt9me4
OelDEjJNlpuswTUY2zlAx1vS846xaL1DzdAN3znTI7XTZdkYYbRc6uQFDtmUYXIJVQ26fks58HqH
E+dbhyQHHyOYh4EXsDok5ZAWIYEfsxGOSX20xU0+eO2xSXOPRbnVP67F1pJMMEzt3gR9C47FuCKR
9W4YgHDNRCvS/wsXy4mu4smDYq0NBoYZEY6OXrjLnLU15As51jpmyFrTMzU6C2UTmL2JCJjI93ft
ImXLe0WQ/jjyj1soih33FGksvO3uAPM7CWuwUyJP4bl0yyP7EW74i8NGvn83nu66Wi6Du5/oW4LG
aPjpHfHu8LvizVhLwYFbQ4mbL7MR+1POodNN3Ghz4Xn0K9QDtJgMyaTh5mR6PlGApGojc+hdklxt
y47yv+13AXw21wp9lXLu/e1B8ZDds37t+asIjlYByoZ0KsvFQgpP32otfQhOZVZODqcmG+VONmpx
eXCEmRkZFxghYwLZxsGu0SRA4uDvcetWVm5OidAbAytAsPbN+rqzUBBlp59M2RKxO2S5Y+X8kfbG
YNFAKnX/ZN7qtvtfeGlPZvBZoJDMmEwexnM7sE3jvU1wrl54s/4KK2CKlVDzeWW4Bozytr+TDg9m
QbOIg0pvJINU+3xmjmfmuNh1pMylRPdwi5QUL0bvofWsl3i82F8Y9bkyvgQXCe2aI3ZkM89Hu+pH
Mxrjt+3CPhET42Y56QK/qcisX11UNWehgsm7uR08n+qnH1CGINYarlIlOWVsZGt/pPq00WkixGm8
kP5pHCHG6XYzc/WbMTb9pUdPVcTTmWEBvLsm//JF8AahCCi6mfDsXqQnums08VIxjwQcYEtcy721
i+cue65vt+FadgoQCqxYWomUAFy/0viaoGQ+7O4bX2aEMKg3v9/yfCRKKX1uRk2LL+dxQof7oucX
12bMHx1rUj5TcUIOWfgy/EZs6DneW9PfonqSu7kHIxUOAR2V0JsvoK4z2NbTV7M/53hJH0HNp+h2
/xDBNM4SphN/IQr7omW18BgkB8HjZvBVa5F+0jfzB3G9oQocxhWxNzAeJ8dxBnHmf5Nwqd/u4mN7
vxs90oC+O5eGKgTV1o+WjAzaBdrbdouHfRTumfFPFj+Hzo3YqJQFMHJE3+Rq+vBcw4oDAvO/sb0s
3QunyLMUJDtuJbHHqTFegNUQ8fztJEDAVR8REU06s3nhu5Td+naQIfp+8ECaOovj1PRiH/403Q3N
xupgwbaED69aQYNX8fXgBdPUL895O2TWbdLWuMh35CeSEv6rsRhXls0yNc5wFj/Kjv1Y7HxcMumb
jG0HSYF/RJgvyJjFXsl1evF6HQW2C31yCdBW4eNvb0YkiHgKcTamtjRaF1pGO0TB/ZV/0TZ1E69s
Y/v+pCXU0ZfQDy1rpvTFaVH+guYqT7Ws7+b+qyWNG8ut8BW7jk3rYB+lUxFB/NpzK1uVQJpdIJqZ
b5H5hboNozdcKQb7UZitpVatEB65asTs7S2oQ0c/G4sNdVsxudGOdOaJbZQDqExyRuehxNnbpgsC
unFdEjOqM+Kr7ffuzw0M3r2ZkV7Kf2q2VqebVXneiRk9yWbaRTWBn9r+KoWPerOzShW0eshlvgWe
gmSILQZ2e9nzmRILv34/Cswe9sgKH84XP6b3hizcxzK2edBXcxTc7SN26tPcyeVoVTX9hzOcxKzZ
M5ZtX80TaZTdCrtFB+ltOqPqdSn4wpoRIVDwXXA/wqLMu28LBTBe2VsP24fXwRn/rP32Sjtq5QZS
sKnjon0c+KHoNSQFbyFGfladxeBO1ZG93hna04ndGYuQFei63m/E9iMt3jAxxQX7wTfc9llQF76X
g8vhTtHayL4xmHGrRYmfFzuJeU2lVixImDa5O6MiKvlNmrF+d3GbKi+OU/BWh1QqjotIqZJ5pe/z
SxfdRcAB0Lhyq1Rwsp1cxva7S42uXDHtBlOmtIwP/l1ESvVV+6JEY1ABsBVw30y+k+SdYQjuFwkM
0h/grEVLj45etW1M34f+tD5RjsIDgScW0XBul1rOljwNcZSLnDKou9MPx4rgc/Iouz4ozmY/0tWI
R4qjrWauTbv30MtDbFktbIef/K8nQU4QKG0lLIsnlRmcGVdEN6dUS+4svtw+f+XzOJuLwDm5+2p2
iEoUbouiTUUn722OyHv0i0YamETT/14TOk+rDgdXRAPNDY8sqJX1vBShCszBiOJ8NBrn9j8piLug
yUyEoVEEqTma0/P8EsxgwmiQg7dMtH8j4rcQ3RRB69atSvX5pZXFMK4BP1Mdjpis6hrmM6q5fFJy
VQviwyA79icLpkSY2zpiBdIx8kuwzcMhXTczd1tNhRlwVO1kVuD+UjqR1R4Fn0ESHPw2AL8XcHCu
F4DSbQREnJH/gYbV1IScVaKWssDhC0nA+as2aC0R5m/EBnnEdrMJb8bD/6rYpJGz/USFQNc4RB5O
uMUIRR4P1xeZASIBIX9/aSsn4J50jsO8HyJuScbX/HWR9lzmLEa/Fx1zdypYkuR7MaM6fr3sCDqm
3TyD0x+RaMJvaD9hLBIC1tSb9ovVyOA0tIsVm9SQ62QB+inFCYOinvNNk7BiMEyfazB2A24YOjCA
kN5lZR00lYq3HCHeikJq7n7JduOzHFbDVxSKcZTU4kq1IeYEVXJVaXI0p80nHow69t8v1c34IVP4
1YXIFKVnTYmNh+Ftj87AzHMTwgScs4EHdJ2Z/DcdBznHy918UsaVpsnMOzSt6gitF3IiIMDTrNcW
tEz3hrFavyYgdKfStAh/Y2aTnOhnPAfIKsN/XFMa1C3dL2SStGDGCposp9Q5m1KzzDuW1B5fRgHm
ZbpwprY4DRR0kkIQnz6gZ+s19Z8xsiKsMs+fOM2S5jWj/jOhZQqXa6x8wL+eJYln38L68jjxDJQb
tRW17vdVhvTq3Sq52NnAahmEFlG17scXTmySHXFJQfHgxUlXpslmKel5p2ke8vH76hQfCEs02U/B
yaxAskuuGdOvTTwBvrhMtrlOE1HNWfdq39VI9UsgOpfFoE0zOGRw9TgguOGrq/sO1BehvGhhVnu1
MzPyJbaSb8Dgh1JIclKcL7PGuEL+6JK1dSRK/c9GxCyUiArfBw4QrV6vxcVAfkH0S0cUrF17q12p
Y5jEq7fZmgtI7gt1Hqt14ee7hvZgDvTrHQUKaPKgs6QlSFCe+wzwkroqCuEXOvLXCk9cebRJs53C
cBgYm0z38KdkpjyMTMmht+N4Bn7nBmUO+54KuqntxxC1zXMTIMAVCZkphdSUSQmSQRnDNhDNGiIc
x0ctYYPSnSXyGuJ6r3qDpi0cOtUkhka8v+iQ1ASfPAwPTyKV3/HsEmNZdTKeEav0JgeGPNCHvIK7
TgDxuiDifnXdA4B/1HuuPF6GscwBk3ecVYM/Qv5Udj75cKd3u6c0FNF1DXjcbhNix1pA4l2ff1Cc
YrP6Dal52vOD1Tk6eqT07XhhYUGGM8sh9pALzDsTXGzT/5mwNeMZjVDDSR0Y9fSdrwCcya8vWeNw
S7OZfuUJ9DLDP8HiCWvduRPbrPNwDlQYUTNTV5cg04KB1A/VoBwR0NjLHdWuBZzqQlflmxjsLW5E
1Ri3iGFViytDTjWHj5/WiYt426dTT3Qj4HdHAFezb5hAMFEVAXyn4nOPEKJBDVxRCBkntiwldiS1
yGDqQdJdXYIs+93RGGoKBL5qKiY6ppXwz4q3Gonhmyoy32KtJnpiN2W9fOywht5MNpqh2atgRHTc
IjOg2SJoWhGbb2gun9kTIggZ6GzXanQCpUiOWc1tJcaXrl09TO8GeT1W9xmiRakRuSAAnXKFebdH
ZfsCcmVlr+FjrmlcRCSH/SuGdrPXsoYjpmDnPXu3r7at6GQkVkRcMfwyE1SDrIFBfzKBDp7stYvV
CJNKR7AKuqVF+lSPl03a9MU+kwEroToH7AxR3nInhsi38vZ+I9sE6gln8hhtE8SshDVD3YSX1xYt
ZQXeFRJk6niLa9ZVoe0aEjAqhqRads0n+69yjZtLwwmsdyRem+so/e+gaAUMw+e7sNUY23Gomd+S
vIGLRLdS97o63/2v05HyPHeOvk8ZbmYpZyPh0zYdtBbvWsnzhusg8aa7giXPCE35WgGe/pq6Fbvi
ESSxkSlyzit8K3Pz8SAFVvs7SIao3r6/SrqLYJjR1GFX5GwBM/06AJhgO4IrC4MyXQIz/W3+zemt
vfA2y4ievScpwq496PfPgM1FiN6wXudHNZ65dtJzJh+N4zsGVyCgS21T6bU1dN5WKpRSPB1/zhxu
CJIPWicUJAHwQuHcnmvtcG1fW3egVJVX1kOi4IRBK712rC9aqyMHXRp7FhsA2sM3qJ3BzFPm+lu7
wEmXWWoDxepjUV/iJCTc+dmCf1DKuJQ+yghVsKowpMZg0RfmGriEpEpO6zAHLdm1oXkKYJiRpgJo
WGFYmCr5ZCcr6KaWFaEj3A8F4ygUvhki7oWMjm4xmwRgeX/4nqmcr7i8zJ8jy3e7t4NQFbzpU6br
HwKZPYc8IHwrJzdN6aXJGflYqjJuH566xGBYh81+X7mZF1Ep06EOiQ7uFDf0RP+zOTp8X/IvgPM3
c/mRzoy2yGst+EzdHSwICbj1Zqx9AFAghhs7mgp18Pvs3bjV5GTgsLqjQoqjvPrgFMW7SYjsqFui
Tu3PZxvWGNaJn+AyEPN+K15rBcNSgGvr+BOWzp1mIhEM4URN4U9AWbkIP/nKkGfYN5f3LcA5tAHL
fVqwgwpYsFAinwt5HoZwxl6DFZa61aEOeY5cLj65ievcRfZ1qJdS3u9K3gvTL6oFovIiMSmasAyE
tSaHJXE+5Bz0Ue0voaiR1Q9Azih5R0AZ4QcNy2dCZjX4IP6jhtSIgsRopCJDpWZtaaIXxnEPXJi4
8BnQGAmms+ohCrez5q1taeb1tm0pepXSaACdchdZMjroeI4sq3TBSZwMICFkuOFe2z11SGOAKt9/
NTVt0wixbOEPcHgDdBo0MK+C801S6eab+IgsaMfrmU7dhnkxhveNrsTo/4M9Q1y+sn65tBoTtzRW
O4+3n6F54TmdFR6rpGXYMHyBckUNLPQVfNXZwruB/632i0AW3+C9egIGT+hkUbt0yqfhYcbNVHwr
pQCXpxmbquMkng/R/SobBF+ZQ2LiHfp4AZfSmsWGvpBf5YBfMCknxit167dlsqxml82ykz5+/iwX
Ch9WjeYIlhU0AauucnWVuFjeooPqmYxWHM3MTKQLDyRXPBcv8bB6iKgSl6mqkKzBM/S47hvPR+hA
DRejkcRfNMNXWJO0LvmgHFR/TFcwxGYBQfMTiYY6FddHkv5NTEVxzqkNEqqiJ/2mYnjqeb6hhCD/
o8Bg9iUFDvC1+I1MwG1itzWvfeXLXek0aLyc/vTyeYjy7Yymv43s7bxSf1PpsP3bonXhExkjoukA
6czvz9tJsfQs0oSivsTL8y8rwr02fvK2I5WYH+S9Q1KYr6Gce+EBiIXaFp991oIy+u+lE9X2b9ab
+AjGgM6FbWisMopO1AZfkAuFN0mooyziSkKG4sjW/eSxooR3/j/IHyqauBMsHLJgI3S4pjzQJQvZ
t4rn6OOhdYNB3q83xMEswl2bjj+rJ9Lf15dCFa2uIKT3jV6EsDzwBmniNHTxKEhZSe/UPke6Lt/c
sNmtSTvoDiVOZbtCfyxdOvWsdPCr2TCKUqJAN2iASbXyy2w0G5jb6ivafsIbloGgTlNSBR+8yZ8P
Ss6QPDQJcy+W7loYwuIjWxZBjnhZBK0D4vpw8Sqswhh2P9CH0weh/OIZvmOSYenz99qpQ927EWnm
18+tSfzbKm5k2kB0x3jKJ9sqRW+QQX1qdwUmJUaYEhiw4NC9hA6MT7DBsnKQ2h4RSjkft3av0OMi
KFVMuPYYn5VdVQODpugPi0w1g0Rp/2uskjht+aAWKTWU2d1qh7GGJq5yzEONt08myn2UxHW9iuRQ
e3yKv6arGZqIb5VgrFwTj7noPPIrwnGbQu7QeZNcYTsOzLTNYhGHXvt4SGl8p8Nbxkrz5WEMFIOI
nDm7XwPWqiGreqZhWclSZWcUKy3XFQDHBDifP2YBC8xfAvmou6h5rrlWgMWkRHgk/3C3RT52dryA
IP6mpbdDfBEqLRLUYA/R1s4yVvNcYedCexxaPrHRB16u+043Lhx6iW82BOQTeuQs3h5D4xLjrByy
eijBuYnYESNT8cvl6rso76xTXB3eiVkoOhA9Zv3PCmM86ZYRX/gw7c5hrxaus7fabNwIJBRmrBlY
Y4FkYn1zoeoDCEn/0IMv6SRzV6zMoupOQGLHjKNczDC/z+tQ+fWqYr7ChHY3C0mHiORNcy1SdA6c
P5CPfEbuoIr+JI1QiUgxtz7W0g+f+S9j/LXMfElH/AG1fYCqCkEYIFsMwsNcF/kfMjiYJ0eW5Icz
qVm2GlktCGlBj2GVLwkFibb/zetsvs4AWYMUFSAaMVOMO3Ji4FRExI7A/chu+0Si98XtQHKF2KbA
Zhv1LT/aJXfjlMqUi+hE8TG5tLm0RURIg977t0+MTJj3zCRA/+aePgjxjdXci9CMSBsFL/A6lnno
FsyFaWw19UAQ6a1jdbsF0ysPOMHrN1cIl6+bxkZkDt3NUu6bvVdYatp1Cx1li701OP9zQnOxqLSU
t5zkd314gsYJ2XOemP8+HOIQhmLi2itScbrsgYzQIfPLiP/y/LiITQ87MGX7FxfgbqN0X3DK11CU
wtmn75CQe0yTzMB1mEwFsN5of+WLFvufIlez89HbGZ0mOyI/trgjCmcbXep3N5hhyvsIYvam27Bn
55f549zrrxzWMNUobVhTMJoFCQjclQBEKhX+PbkfWCXdB9MhJGHCiP76KII64+IxJACWp2zbGDex
jj7NrgoxQXOAvDbzhl/UJKU+Xlc8VgkAmwCbrLBi1/fFR6htmFQ2FgkWEz+CNKd9URtFmZxarafv
ZoUFxfAOv4kJanucCgBPjodT862tohAsw5E6G6z/WegboSVh0ebQy2CfDweWU9LJCQ0QQlu/SZGd
rVUGlzAia5vigJnUFivRLCmRuIOqlq6SAnXxp1WL0xU1+goFyIJG1Ci6HWUn1k+ROh4nWyGJIY4i
P7yvXNg8gBsWadB1LVKOOBFSg6gzVGHEcLU5MFoSWTZKVKbSJLBigzfQAcwEd4bwpTranSDNt38e
gap8VakC89Qw2dclSFt4VpA58f392a8lG6aT/9VHAnjlfZx15fpzy8BAjYmsaVp2K2GQy7Q5bdA8
Ipk+6AjRz96D9Y4g56LvejylSUUCADAHfP5zeCHvzM0nD6zhgyjWEmK5zgI8/Lp+T8Sh3dU7sIt/
uaHPMLdYhWflSDhtlfuOgiBCnIjoVbCMm9sDB2LfAwq+W6l3wp0Q72TTUN60YraYexX+v63Sx3bx
haI1x2x2fkRqfVFyDYrjHQ/1JTRlV84P6sdDXZdGFHzeAdRpU/kx1mFLrOwaJIo0vq6cTtQUoJ4d
fGMT0BmwkpFP2BqPcI4iPECtAZ52Km7839fvOBx/DqZkc5Fjj4tR42BYdi1cH+kapCELL9/btk6L
1k3i1An7M4cCJPncGy18iQxHfaQBYIPLCY5BcGL7xJ/XB1ncBdWUPV3u1skmRsijExVghbrmD2Oe
oKB8wajySFCJQGdXW3dTQQb3KUIrQKqfndGL68hBd15QL/AjqlAaA+Y00Cczy/jJnwv0jC7CiMdF
kPxE0qKrIeoo5kTM4OPi8j2lOUY8zj4h8lMAUedYG49WSa4cnOzVXcVtDY1xT7JGNFwYF2cnpSMn
3PxrYpuTfPn6mYRvjjMcLcEstgP4UIfr1JXCNk/oDjlgyUJOL82cUAd9pSu/BDtr6hYt4BFEa1ZL
XbZTK1zcE0hCBOI7xr9nfjYZ8VQwuaIlk5PNDzKMDxNhvZaWyPIVXA5aP4HagKKn29jvVvoRcomJ
zlv+q9yEUrV3fdHf+se8TmA9vTxr03ipA13b1S4+agW83MPplQXc+JaCqgOsDBzyFF3k0XYcFhlO
XYzh7kY5Ie7K5Vvdu8MTV5vjJ7AX9ETUGiu6aNovj2+Msf3oeXkKyiDMt8uF9oyin5E8j8Y4ZAzN
/fuZfT0XyD/0Pg9ZGlQQ7R2jkG+3fCznl5kcZNnGj61OA5CUZJfb/r449TafdGCt++OBfAh9fQ8l
A93lZhSWzqOru+d7dK4ii4rjSsoMB27HwtDOOHFxTHNQs2Kdsnqw3/TT/bZV9PkTq8QMISMYOoKF
FeAf5Xg/8w9sPYf4JqJw98F4QEtuCcXgLh30GEakNhgTllooNyBnpwxKRAOjP67pVRQVjuiQekZU
76zTB536m8tDXwuIquYVPxrBcTVK9RAym5/jFk6yYBL6Wdw0BN9wAHGMWZJ+MYIrgdefgJLtz7Nm
hTonUyWJcUamlhFZ6WrTXqAhIQbTIc6QZP4o2/ovOUL+t95srPYsv5OHxXchh58C1c2+dsxoyATj
fnnXsKX/eOcz9HIQjW0xF4dZrDcoLrDTMxbhh1UeRTS/B7Xg9AwMF2IaTJgGGjoQoyLOAyx21+x9
1Bfnc6udhexrA4aLUm2lc/qW2T9whDpeHVTKkX3vgwZEWiKrgMvIvUmQFn3zwLvsXgEUMxAyOgkx
VeH3mMlgumIUuk9OHN00ZkmGzSi4jyIK1KX6PDq3N2J0lhOqTs5UAyD8IW95ICV0mDotyicW7Vbg
C5BFW05KMPSTEXR+qchYQAODwIOp6tmW6nlhYmUQaDsUs962P4KAgjKursp+XHu4jra9fGPmM2Zd
b56ZGiEfTRK32/LuniWfARSPlK1C0T8dc46XIK3Gvn3eCipDGmuJdySOuRkdF9WawMlHNnpToesq
c3QumVG2fV7xxh0DQWXw8h4prrafk0AOfvKjxfZioyy4/mb1uW+MtViQ6NZGmh7uIvgO4lN3X3uA
9VL+TJJG3HFzbRKKzA+7ailTE2ypzMXS69rypAh3Y9Z5IL1Dvtrizuj7A1l9mTKrGW7GWVdHb+E4
+pj46q9Ue5TXcUW7ILG6MuHiWI866Krmi/9p9EhQufY/g7+B5c093XV30CYhSnOtiqmCOePvlNKR
iEldQsfGKI0hrhZwaXht2816EivfD+f7Wv9eBuPQ4X77MBebi4M6mtLfgF1u+kUqb+yabOjSo65G
EGWR53XT4dzryHq2VWD1BqaHDjnRP4+cmpsU73Z/gw2OoyzJNK11LmJ8TyJjfR8DuFCD8f9sxw/2
MESc5Fjqk3qZrr8QLkML2BucFR4h0T7zC+jCl0236paW7Fkd6GT2HqR4wh8lv32COoBItjUo7A+j
wg1vxAGI41o7GV50ZPGxo36zOe3AVq/sCaq45UyANY6/cPtSteAZEBB8oXrxz4pGoWrXCV35Mexq
u3EoyQWoa51A145/n9dyhwG/kVyvWcamh+nQJN6T4eco/6OlTJam/jpwtWNtVx9aQyWIwXMDnqqY
mLwZdQlEaETwalSCpCeZMQ7NBrYwGoviHD7q5QEtjqM+BEXkGHWGDlM8+n4XLPWBKNM1ZvlduUtx
SzbUsKTvB4sXaTcEDbHtotpB30Q/3mzb+hwg6XjPJ1GSQIuYWFTdL3Jc4GrIXhXfm5DWyrCB85tP
V6fAfEuBTUY7SNpyK6RkRJvasu/JcSELvVbR8V2yR3fLmkjuVGcooYTfho0K2DLolsahuPVnJGRK
19acLPLaWw/VqJ9XBRXGstSPmW4hgNdx5+dWRSBGc6IU0qCNaDSZM9Ink/QmOrScOzQCAZesZ918
VMNHFb3zfsI82dK+SgbX/fcqwmMG/gf7SrO/ktzUgdKZrmLiy46nbrr1s5DAcEl6IvIVILb2vsGu
7TFLRWnIfDaTaO47WnkqxUdqxgxJqxCdyg1R1SQxI70/3iQxctGiHmLdgd7X3PFMcFIkS87EIKon
en37ReeeWq2L/UORS6s+aqVk3QQyJ2LszO1pu6fJcw0+1Z3b5vyqPUvjYNhhhLDB/dIBNGPmf1kt
NmnB/llX11aspYa2mLW/xYzAy4WlY+VZwmwojc4WGXSYEdWXaBdM49F2AySAVItW+aDei7jIQ2sx
gHVZgcUnNiziC2pVaZFu929lGxWgsrRSefVNPgAi/SXNF+QCCWoIXzhplMNufDwTi8k/Bk/G1lA+
znbTzCVI59cuVug8a+EteQ5x8iw3DU/Fif8DjEGuThKD8WXA2l7VZYl832eSRnypbAy24rEqL4y9
oIei3uSafIB+XgsGHitp5xUHKTceGS0CD5fncALgevB8JkxTsAVzzxpKSbw/pb6EFsNsMsUlE2Ad
00KtSqojdk22GHbr1mcQ++HO+x7d5SdcfE2veOCHAE4QuAYzinmSyzNDz/6qypoSxg4CXLG5pX4f
Vl9dlbyYl2cJTgvtnO0DVi7tkFLlH0tf0a+JEk2cg/Kw6wQBroAKjjP32MWW6gHM/Jdve8021im3
ZF7wudoNwRS0AxBVIRiaAj1uk0L2nZ+aWpMC6hAqgyI8iojMSfqwdFizbdcvTzM9ZJZrlB0stwgx
YNldwIqy7PsxXSh9pdYGXA6ctRkTGKiW9Y0KQf5VbJ3/pcskkBKyL02xCJt/PRB14bdW3VbREodM
wB127ljUr5q8LgZxwbO7+5vhloQDdPnWXLB9CnDcRDJHBKhR7sb+E1NxUJ4nP9yhhCtSHkwOXoBC
qYjlSKxcS5NXD/14Z0xobLDqtiW7Wq7Bgufz9koSudA5CBaCgpX6YaSxzSiGl6KCFV6TxEcYMOn2
YYN1akKiwODxNrdyyOR2Td29iRdorAw+IgA7QxlJN9o2gmmykMsNwB8Iy5bPXUE0j1jWboMoG0Tg
11AwkWPRK8XOg+X9p21PhX3T2WzqaFAX+EOQ/zZochoxV8dEvKD73cfCCB36eGhgsQxZgHojnGcp
JbghfPJLXRK4Hp8qyZRvN28QH2CpEJadl3Ft16zr0vnOa8VP3CIKDWd4zibarjSqUuQc3i0dr050
Mv0rTRvdlYSwj1dLy5JEN8FFEgtkbnFx8p83JX3BOLUSqrSX5V8lDsDlVJDIImgwk2WYk1VN4jy2
3fSN451zUBZfMGBvvfk1Ilxkn3jODOT7EVVyNsLGDokXj+1emm8WyiwAysalL6+Y4lb3fSSfS/LA
WiHWzZdIUrgRRFTC0Tr5sZoJwEBkOZn+rZYY47i7zp28FpK6VKFCF8H8ZPeyJ6YMv3+WPIY6q6re
7+Jx1AEMmWZ2+aBxPd0uE/82L2PzLSXGJ2ixPst5Cc4UoXwbJKaYMXN8UxjOLlJjm0Cu0Lg8LHU9
xB/wPV1rz9imuvgsw5onsAqSy9En54Px/Bd3c2ipVy/iL3OMPeW8bWLGcHq1Ymrgh6+qlIt1N9kH
hCxbH9VHdc9ywWgs8EBwboSwy6dUwYeKRL9y60q4S+UqzxT8nEB6B91MR7mPWnFYvgSQ6n5Pf7zQ
uffPHeI4F5/WESjujD+rZaBLT/nfrx0ftS3Gy3h/kaeeuX2Z8McUjyNey7RY5qwBVMFwOXuaSQ5O
zhSHCE1uAA2Uo67/tD6bPtxQVswmxupeI+hr0Q1ZHNOQa9R216yGxRuBeOx4z5RrMIRWwbxWIQjU
lWNmLS6aUCd/tXD2gqYURwdWF7aN/5mPqWPNbZ7JU56tBeTdXhY10IIbDt7kIicj1Mf86TcYqu0G
Sc4Z828fTVuWiPmPBwq0qtopktPc8QFk7Y1v/M4gbTNJ3ffPUoT6hm4qLPsxoJ0Vweo/O0bxzwTE
QlOy9pnaaszpxPfethwqUH38EWpGk2n8KbeOZ+UcuDn0i/qbTOkehTfz0DmDxd2tFh6iYoLngXF5
X5+VPhC0eTvSTvsn/5ApTSRT86h9z72uyQ8iduw63Xl/ahJMaL+Ucve8+N13HA2Qe2LbgiIRmNcx
wo12Z3KGJ+ch8X1PIuW9xbv95HqMRZzSIx8TJHhT0aOppd5e2vzigDvdpu0SVWI/nOmaCepaFIbX
pI1vRDa6qdcmzsdBPNMjc4EveX3SP/UwBDpeA17QictUzK0MD5bbPT5F0jVRjYAk3B9Vr10E/c7r
y1lRU+8DNRL22+s276ps3vCXLwfnLYMSOUQ2Z9fgPvGOOTJrST+qxQSv6TotqYM7tE7jVuiBQqWq
YbaUsPeb+jwFNoDO6DDperD0YRpWiEoUSks1T+kU4koyHtqifRVBKY92Ij5aKA6UsFC/mhitisTb
dWeXPTeYb7y8g0t9GvW2kE+RWG0wg3WChgMBtej2mTq4v+5T9H/By2K4gkBcjaBCrQ3LD4IjZc0F
hM/gG78DMxlvYvRLTuN4kxh3I5xAdeklN1iUsV6LrIQAZAvvdQMeMRB65hve7W+GltkPHkJCM1AF
/rsgAfifct26S8zxb0DcC9tiqzLbL4bJPT/exQY3LchTVU+UHNtQiR9hinf87FArQD2D0B+GzZCO
gh2Yl4F/up6vY+FbhzSwdiqUTlNTdXA9ekw/KWbEVHIYdK1phkUEIDDKVKe4mrVLEmfMCgOTBs2H
w62d5rBwiztv8jfA3GvC6HbMnfhvS7bXB2apgET9oo7sXCJmGLCFySloFCzansPFSfEs9O8rsoP/
Tgyz/7fG+m8QAAJvbzcIUoxBHs3KGn72LcZyd/zMGKUYUYUc1f/2vDFsVjKc0zPXhRdedZNI6s76
jv5GgMU9gFvF1KEvg4Bs/ihDX1TFiXDOvzTiHN3WnonH+I6upkeJO/YvuF5bfjqUm1nvxchFqg5u
pLHdPKnj0vxVa51zE2xd/54/qOUO5OhjtQnvknj1xt24iolZIRNYJgl+dlEzsy7bZaOfmRGCPeTv
112iLV4DQdpYB2Y9TuosLGuaL1JwNt472CmFSg/h4cRlwkJZXC2Yce14bPPjE7TtweO9d9tRxuz0
HWSRd/tpE+oCK6WUgqwN8UhfoML3UdMYDGhABmktS7jbt8ZX+PGupiv4w/Swnl8U5qq8iwZXz0CZ
B8+MLpgUsPAeBY5TQd/o+a7bt8hpeVcQarMrnJNALJYdxsQoo8jyrW1Z4kI83OIGaRZRAAgik3ga
0nMMnnVAA+caOijn3rJepx1gmW70VqEZc7R+AnWhmAFpDJkO6gAy0nuvM4dy3w+yWOIlYfibND0X
JH0wq55OqawvYWAayGukYTzwUL4PgZ4buvMww/TX9H5eBQnIFBpjpVRSvgHG6JZ10geLtiSpRcx+
JnrYoxoTJOSGfLUZbxZN0m02RmzqnQ9RY0X26MQ09haCz4paY1e4wiU2Qrb3pdzy1h9PURoFiIwK
K0v+EoXZHeqlCfgRt+0A7ldXFPw26uohz2kAGDaWUgITZhHqOZuMDgfjAmREfDiKXEA8T/BjYwSK
WUedfogkT56n7jURMSVu6/R+OTOELp+Wq86fnpZ5MsF8MTx8a5InCKXtoJ8tgAj6OMahjshb93lQ
KJJ1Oh+BqCDxSTHQZsaOE1IWdLQpamqV5UMoQIS49OHRiDVG1guNUwVkApv/biPsaaxzIxVAQEvE
jE2IRongQGiHam77b6Wwo2miMA7RdD4OFcoEWWpqEXzXblA3tHEBdO5FxQPUrjn6Yj4DKebiYSI2
VyQD/nwHFCf2948Eyjw0WR+RZpujOrIBvReND/EYu21MxpNXrjeopEHwr+XoyGiWfHKpYEIQxMKJ
mzO3L4TXejs0ChN9zxc7llf+/QeXQjXgLNJ7H3ThGSZYOvBqxZ3tR0aQvBshrnonTnW5UCuQpk9r
0As/qU/MKbJ75zLxd1ib8pTzU36LXTcJDmbqYCBKfe+U2L8w9JGUS4KszL7yAJy4i3649i56PNGS
/c+vQS4X3VJhvQX7DPY1Urs5ywg5679nir3Juhsi8dkK9kDBlRsii08xkzSTE0sbMn1ci96R3URA
lGbA5wGhiBoxV9x/ywZr+jtSOzLxOZZ7sxH9kXiQ+Vy/bnFYXU/LgCWWeBQlZKqAKoIwgpxNg80G
VtmhbIp8QRZwxkLwWDsNhbpqSNGmZ4h5Qf5Hlc9+rzWk4FLacIUtaYrYvso4mDEb0F829AScvuv/
UItmlWqJRXvjakjUIaxFJUu52Z9homgyrABpTRBW9ClyUC2XzzXuOLOaXo6t2b+ybnnOWXtHjqqn
myadpMfVA2nibsOPAeJfWI0Ek3mwqakhGzkgTCunsT6PBMWj9AumOYVoAGwjYsiK01qYOQx/Pd+D
7dwjpJZsOR6rXskvx8aWWrU7ZUYNH1siJXKbCQM8xN0bM9X8Es1jTdMOQM1ako3UgSqF14Sovp3v
M9hd8R9IVSS9Q9S72Urpg7QYhH+opxhOBgwCp4c1QETAjxGWWqotDbIogHIk39COkJ0/6ECVpnDo
r+TO63oEAPk31KZ1i0YzstzAZmEXo1sOG5f+uj/zP11y79nBdJZPCLB7Z2hLEdb07+WBiKqN8M3/
6bJDIcQM4OhOA+HIetUBhTTVA4xUud9pv0xQfNrr6Ge7ltgI1paOfO5l7BFON6m+KPlWtsjqpbdN
KTialWAbfq1a+bKMu+MVYYVu/nM37oc78oqKskL8ujWz3gL0k8iNEclQn3WRDHkZDLq62Nghuzj0
FY7imsi5NTWpeKK4G6pfC1HhbRZsV+NrWqbMsrtDP0MXoUmRUVRR99kcmN9lhA+n42qwCFIdOwE6
P2zY1kmYdUmh7TBN+658vNIqmKN+EdkfigIEP71IAYZMPtrdWk5H5j5NuG9gpJqgloffIoBmO9k8
kMrYnoXMpMEUWO2XmFMej3+r3sijowiEKXuw2T0rToJQ+7ybM7hwbWa3VvyhYNFESTrvq2zgvTS6
fzV/Cp4rRKFdHnZF1bQf0Z9BClcDmzg33DYxhmJjcEkoBAkGnGhK/OT+kKvuBWkTYNxFZd9PAHM+
ExXePnKQcLdwUdyKsNYfWOGvyn8Fkzu5v1FBvRgHLsAk923e/LT1SOD2xLyDBnVklxxiOXj5vQre
zXP4mjoFtNKlPSXjFQgd8NCbR/ssnNCSnIQl8X/W4oCdlTXKkPsX0Ek0Hkwy+kpGydkfo3JauZha
XA8Ma3GvPcAG6d8uJoz+gjfduwlxA14BSi4ESo0AIXjPRk0+c8DiyosRFQJsnxl99p8RMyEHWpGU
HWHhhwNiGrSqg5zJ8hW+ZMN2R69a0wMAoWwgpcrDg/eANxyH2vIgd9j4I7xiJrxjtaxWD6Czh5r2
JktWbJvS+HVcnRlun8GpxjxzNtZLjt1/c6b7KJWoq7whpt35JrAkeMQkZydMqXVh0jsTAb/zvi0O
oQIWcxqPrQ00/dIuUFWKrCgENA3QXXbljPicEulV8rTjjyR6nfiArwEqgUFhJnlknqUuaacgTJN0
7tUsZ1x5xBJkw9SoZHS82DXmiCyJ5LYjimsfTNznaLoa07nPYvIpr1RJxrCzK8Mr5b1zjxWQi7KV
tRfuaysuk7+821I3ZJ+QLCi3NZ5h4G6xI9ybYIHFrbar39H9MGUy8dSeMIG6btyeT3b2bgp2aMpi
42rBnISW5/gIoFf78zkiJrv5T5lfvjJaHH4EKg7eAEUcZh7QYzquoULNudsyjySCKEMZ8aIgs7+2
ZS+tgWWe2FR+KK8it72WRGWBK3eMFTrwEJsl9k5a8EVa6nuwc3TSgb+IiP7DXjTvzM0hXSaiFReN
WcyvMNJbKdVnBA6zloN1cVSMZaFQKFc5BvqL5v5wbzegfYaoJ1+H6f1axavVVadfRV2tMP9pisZp
M2IXjUJuQWNt1wE7vtxlhZ18UhpCemMkdMj/gmrhGb/zEniCSKFQBtDJUroqyQ4vOVKojIaY36IR
QloxtQTIodIqyJ0RIEFXmhWIujCc009xGeeCyFO7KJH12BFDi01vAkiTUz9hIYStwc9INmfP/Q8A
//JT/uoeMZ8Gxx4aGRnfWmbQgPDKmXpMckK6kwj1qAOsz4oF9Sao3pqTW+ucDVYvVK8YJyjR3AVM
XUA81h3njRQ6XOsrCovTj8RKy+8dG5ly5ofcktJ5a2qNphGl3J2ZMHKEKqw95H35b0hNk77oXT9h
q7HuHj8kDK9kH+y5JBmm5d8F9i1qGLwwg2jQPLL6L+SP7n8SBZb1FpLDc4DoUoUDP3ER/qhhNyjI
Ru4/fMG9hVL03Z6h+aXyxFMJBQZzNDcgKMu2xpix0J3AloAmnyQLosdCT+r4zY5AUL8g3eu5Fxsj
C2YYXTkcZH68HiNJ1PLNdwDBe251G2lcCxCfB6tu4Fisx429Ata1vwPhJgcl3mrlhrJdmpCD7R3X
fwFL/Q1dmwDo/NY//p9S7rSehl1ITGHl8pWbrw6GaMzik2ZdiZ0ZXLrH1vuo3CwOw2PBDHHyEEFR
VSF4ac2hOF8m9kH+iKfOrA5sD8jSG4Cp/1hRIakNHjnUmDVjI+qNWcvO7Sjqnx68NdamgI2PmRME
lvZbJogpEigXnj6mF1geMBiK6XHg9sSk/5d9Mdaw1cgVB9wJJz9z4sXdvzT9R7JSYEeBZJO7H/zs
S4iwO84ydAU/2/Np2QtIrS326IkhchMXcCiY9qOtHK+m6Qr/TxvmXJcrLgUhHIFhUSGIFbov+2U8
iJwzJtUuDKl7lwtXjpdtH07woPN4lkg5UyiEa6r9BkL1mkc4aplDaX1TcrUK52YmAaMNSf1Vhi1U
/bHG1+q4lI+r6EvOOdWVdKoYaAm0MgLklqoqdsbrLcMZKzopfPWoX6k1Vmio67+meR8foFwyeoW1
K7ekW04+RlMKCn9s8kFsfoclLG94/rNfDbpQYVAjaZNLFdFFIoMfiJfeFpNwZxmCBth909wBQDEm
un3Pebam2BX94osGndB3Me4GhAdL1cZUC9oMy84TlBalXN0upq5GLAfprwXF8UGQTNQV9G4UAEfc
9BvNq2vjoJbZtZprMiIZi3Xgn/wcJ+wZp3G4Jv+wA0y1CFbX7JQwxAsb3gPSxIYCWilWhFlc/r5T
vapMYZeQogX2MxSGPw1m6voFzcGTyqS8hjtpvhZa+qHCr/qxnfx3d6QZwAaenivzQ2ACjDMmGgqy
7lfoIgAhlF4VE8Yn999THKm0VIbMNOQkr5KaD8ZdIh0sHvNshwTj59JoPqA047iLnw26+9Y3SDLM
RUPp4hRDnCPB+75Z7Wyq3s04PemjqR9CZgM4j31UpkksvalnhQ4iRXj6M2ISC5HRESyMIcMF+xT7
wVKoFFSGcN7qA71ySkAmxr+VVAK3MFB1fIjXe1nQwQM7kC/spvrgvS5yGcm7bn7PUn4n3FTBNvmx
Y53dbi4vBDApZExJVzqB94upFOGLrm0xwSmVbzYwwguuWlCdGEqx+Rjor2LvlmTnDbQMNw38t7c2
n3NSK/dmCHWQ/PnkIiews5g9r5KSqaxWc831KUWmmlX0+RJFbNk5numerr3gcSywP7EqZDGgrasm
KMSaQKIbkVDOU1en9hWgwK6PEZeFMUILuNIUlXfwUgt9efbjtSqIS9qUBlpMxoQTGUX31Gj3OvrR
WHnaFDue2WtrrHni/ImnW6xVBud0jf9l0XyydOqjA1Gpc/SlCF+bhCD+FVZXNqtV2dRn060OQOti
wJ+U0ewvEfb2bU5hSYoeblGO28Mxq9X/PkCOx5LGQcp65F5A8K/UwNJBhLEOHOHDzd6D98RXJHYm
UHQwi+fAct+bb4pbMbnLlpM7yTqNAmQ7ph1cmX8IV0GTfRKkm2VtAd77cXFoVACEzDeH2JgSBz4i
1sx9WGef5DZ4825j4CgaTTgYeLa2hd6H7tcVRAhJ7MpurdlqIgQUOh9tmNAhBzYPqTc4ZvT+slhk
P1+0gktTJOE0jN3XuDUQ6BZUf6Myg3Lqe9D25qK/AjXc0azZXp9721/W8G/yFMpOdkAp3dh4gdvv
C/pxZN50PZjkgGIUDCvzUZYA2Mjn+8fuefxv2BbRbTg8Uxo6GzDhNpSbsEaDAXfaX+G+qYrpi3lb
qEnYCDCb+5aLMKChkM3oj4/c8Lkn6LWZ8sjV6qiDasNcX/GdkNFWo1BZPvFTsrSqCiuDgNu50Mas
0e+ySPhjxk2WPIQKh1vHFFhAny2yHeNTxQuF3Lc7vb9INcyVy+4Cgo/7vd4AsKmSYlG8OkOgpanK
gzZPu5yTpTr/AF2veldnkDAW41SOhp8DRzeEeeLDqmxDC8rSpzdykbWSkGMYQW3cJTj6W+wy4zAe
Ygu9FmWTZc4dfRs/2TFxrihf8k/9dJ5pMgTs0DS6d4aAnmLjcfyhKFnLWyayQAH5mydwBOteFGnq
eDT1gGJ/CilwqrJCpRhIj42rlJ5DB2298rqdrLv0ZaI2b6H2Wb6AklFuH3dBpYtsSFp/YpJKYJPV
6GDZpqLF33cqr3WdgnQPluIkcMctyzpN3K9FDdA87zyqTz48bqr0nXnYhmuGvaExcU5gzIiCT9E7
jSDk9fOAM7S216t2z449sMwt2XFXzzbHQEHsreHHKVD7fTp87YgPjEdKda2Dwr3hHzf98Lx37Wns
ebXc4BUEdCQjE4/z1ftk/TpXdC+KkHtIiUulBuTSG8DVoxGLu4q05s1ZfQajtStvxGy6CAq8lggm
S/AB64uEjX6fAX3XP/WNYSNuq0TOcNXtJwjy5ze98ys6OPJX5BCb7M2mPRCmLcvpM/u9BnALZNCA
RpOGyhclOADmyuYOo6wuQqCkhddL6ZE3piP5AKD3ffgalN0CA99Hw+kbvGxgVXsdeSCKgfvgbn9I
iBgWgEIAaYmtHjrXENCrhhfK3QBF2ck/dOls5zad5o3hJZC676Epf5B9aMxs3uKyoNf8MDMLnUTR
W3G96z0gRd323Vab3rQJlafdU3vF3twVwpZbY25Ox1GoXubjSH6HlLh4EHyFIXfktSpuDPrXHufJ
u6ioYqIKsd+npQLzpiQBc8TKhcJOMXNObaCLc4C6HfmCAm5R3eeDSuILmWtUd+5nRJEgNfAnU1cZ
BXmXBh4gh+mBbMM6C3G2vUAzfxm7MQDODatkpe9H+c3EOJSVCjuRyPc5RFCAhnVvpOTyFrBSwFcA
jikCppORApt2G8qNCcPJdkAwOEizurLCljFbNIAC8PRZGQSHTjEwUyjlG1LQ673p6A4rEyvSbT9l
CNs0vXGq5ZfKqv62wK1rONviklcO8GxZK5Z2bQLj0EtZkYURvxYtakahCNmci6CgOx7gnkN+EwmN
xMQILoZzC7DeO83PO+1rtFvN19tE8pR+s8E83HtMG+u17RFA8GwTShOLainyWKxxQ+91geZ2CyuM
zqvp0ytBDuLOtA/jhRM3ISb/oww+NLkYhhU6afgM7ikNx/NpYI3stAHWy7BH4ATGKXXkJkx0zGtL
iShjRQ7q+RhbjqIRM5GQ7Go/KAK7uMrkLmyDj4xitEq/6Qf+PZKSD+ezcwzBrtdaHyiYTszBmvQm
xyIeL3MUPd1d5/+gG/gCLVUnIV0opS8svj1WYOgI3LlFcAymstCKH2thluKZoDJV3EQ7sUrWskKs
bBFt2mcfBx7wU10BAb+SmKiB3RMX13jIIBgacvFpAOYypTwGN6hIVjjjBZoJ+ghecVEo7V+8imNP
+gpBwYJyajWoaMu6HoeZP8ht6k+YJ6+fvZWDXoOy52lArAvDhoVg0VwpEXiwRb7QwicFX9kfud3j
m3FlmRSqYBUyYUea8euqN6U5xKvgHbr7JlpXmIacAF7vymFDzDlNVF+yFFS50Grood+Z69p9TMlf
2/dbVRP7/Q0KC3Fjf5JsJLb/UYMNTREp94Y78LcbeVUwd79/c7ljkmiBkFG1zvfi/270ut9D9jzb
bHHupqRU+bSJJi8BMOVV4bk5DH2TFhXZ8GigdmkR1pafq+a7pVu6FmIq2vZxXfWmhPzk27WIie49
/IwNxjamFNO6Pm/pW34/etucRssh6tNX8GUVpN6pABAiiK62IbkURoogx20VADnVA0Op7Q9FCM2p
w4AiPBwAPGbdO16r57FGuxDg3P7lWkqc107G21oSHxTl9bB+cN/JjPhcjGv2sf7IikPDT25nhi4u
ttrwbUNys7edBIdS0vSug7Ruiv3XaEma21TuDfrEkBju4tpym75wU+UfCiFN4DcvgswoW99/Muq5
nA3NqCQ315GxPWECB4dduK7ZnAUIbKEDBxJvkCaJBEl+Gbic4rmEs4hvaXf6Ujm3nHHt3YuSE97s
+6iaG2c6gvRCeervUta1O15ERKJJWp6HiY1hZJH/6/Jk+MJCX+/BTfSn8IS2PckszE0ie5+ftnc9
CDUdXsfE2bz+eFT/zv98U5w+xtk6v1+t+/M1GvjtAnoqBOPIaKYQTaZ7+vbXnMGmarlKgAO/t9FE
ru6oJecPM9QI9f5iNl7ApCIVMn2FQVE5vSxpdrXzkiutCfNLgEcVog0finDLLCnoClKYO8XCj5wH
gxmfXOdt7RxnbyRmN29/bdFSvL1bRSnvjkVXLsB+evwyfRM7MulS8qWZQ9KF4So7btuG3kdPcvCx
ufalVY6YMZjfqzK0ip9ZvjyrqkOgCjzjjOI1xUfMRIDL9kESvju11vy+wcD84mEcE1pq/6m4Av4V
sTfvGEHiYj218+eYyg0DVS3BDLjRx91RYocmKYNtg8xnVp7pgLf60xg70w16Bty1xRVLUYzTcpXA
DqA9UqDLWhstWbn5m/bGBvcPs3XH/V3akxDMsZC0TJ+OCe+DyCxC4ZT40bfq65pPpkhOpBRM35Mo
QGgG6ZGoVNMR9tW+WjjhDZYugAMePXMRJ2v9NSkIS7p1z8hDmC6MAuXu/UD1o8nnRu1rmDpmuyhs
buE0tPzmgUTZlamDOoNXtVCXmEKnyjHpR1ZcvOz3M+Gr1jIn/jrfH7zxeAKWlg4NSXArh8F8MApx
UiD8ruOTx9HFMbFMdWoVbqJRmn1loOjQaHTKYH20u5Ymp7U2rPF9vUs7+22d6kJqdYbqD69ms+XV
PJvV4C43GD1FtUSPfNl7006s6yNB2uM+JI1lBSz3nLIPWcmmnSY2mMOzGAyBk+KCe/mtKh/u445b
cSpN2xzVbDhNEJtrYvN90Xzv+kUL1Gnecf/e/BWFliULdMgRK+vB3g1lvplYmNUqYNeUf9YZ7Jom
vOYl1gHnHpafQ0tYn8b+AThn0LWxiv6fj/7pwe9C9V175zPP/1DS3QYW49k/fvR6aE5DJSmPI50D
jtJIqfxJD6e5XbX69g4SUJcgFOIlr5S2SxCKA+vBvBKafu+w8/qX4eD4yF6ty/5XjL/pkO6EVA7V
uuoeuwXTJksa5RKkiyGGVrF3KT6HppoGyLeipcah0unoAEAUDkGcM//AV8OoSnQi5O6KdVbKWaq5
c2dYbpOACMKp1BVPjjaXiHYicETQq/CtNKBF2OREUYZVl5cwJNlDCFZ+GIoBN4+62TSB2pWyYQNG
9ObejmZ6mNsRpqO0f0xHMtemuKKdAnKbBItNiemY4inFxUoFBbpobiQhcCP6djsaGzezTgC6qOIy
9CiNluXJuU5xayg3wUzXfVCfQswXXJeRTxq4twqNRvVUrL2tFquD+FTNc8qcoZbuYCxrQg2G/W1H
pfCgG00ljTY2CFFcoIb2dcWUgQ5jQZkDpKYLKUXbCwqTyadLMRjk33bws9fA9hNKsDQQaaPdyofn
+VL4hRQQEn25G6n2OkIdjgsAo1W29jvew8MSEP30KnStnh1dMF0gFL7JGZeQfkxGfOnY+jgv7c8K
J18lFFRVNma2Fh8bjCvrdI7L0a2/iOFT5LI1QXl6lKmnPCHa0A01EiVnR/NFT3RaGgC3zQs+5DXg
Xk6Tfv1M+mpHwHGw5SeoLrtGon0i9tu5GyvgpaUxrlxO6aCWhlQRTBBhfqTwe4Gqe4vyQeDSFNxV
Rp0JeX1yVRtnCRHnnwKg6yG1TwiZggdcaDYu12LjSBUnzRlStG9KiYNHh6Rfg6FYh73W5xot/n26
4o0fzc5TgtXLAn9qhp2S/v7iMWcui0CRLIbZhX8/JhpUTV2nNpf0Hghjmauafef9wfxx7O7iuIAm
yiKFCq4zQ72Zsoa2wzlT7MM3nwZN5ai92lmsuan7gqxtWywn/pKz5BZEpKRYf+h2wshoEDlG8Iw2
Uyzcm2LqztvEYI3TX/McE6zh9AzuWb9cttqeWfIJUnuPu0n9q72JxUEGHp49Ge2Y04hDFk4rFOOQ
ZvmAHsUs4rx/P0qLglVzYjlb5rCIj42nohuOgHCrb7eMsESoWs/FkvklzFoz2tUVSCDvMz8XS7Nx
iRZQe0YqpzVS7R42DUBUIzy6f0bC6mnppArbC7GAD7xOZGKlPB/kN3Kr9up+vC1jTFwj0KSeTpID
xwU7eVXyJADXxWDnXvNX2A4IdHYEtZCW8jp5wWm0FsnQSA5aK2emw6crQvp5L4eNAx2AIuCaxNx2
f1BLcSN2skGXYOgLivn5VS34F+WFwgJC0fCUKzF+d6LfznZ0VHK5VsQqggJw/xgk/7s10GFu9/b7
XKEWfvX7tCJFx+RewJWOKFjekluGyhj/wzwF8GoCpVDzwWbQ29NwCgfqpE6jOqbDxcqulc6q9cgw
zUdSYiF1NSsAtas+EffW7/sRtcfEeXFd2rXx7wl2W8s1AAra2HecDhXy+0R2jtoHn57cn0QndQMR
+ylUZKDvvbRpx4ChoRxCwcESXIHpbgSQnNdgrMhPCezD7G4LxVFDiyAzVdZg4reCFbqiMIFDmF7l
T3kXndOIRyH0i+UlmvpAMgBXa5kMrXigyecbKpEo3ki8z3M2w97dn2Zt5mWWl2E143d5t8MZEvjA
gX42R72HbxR0ceE6oOrR1GBb2KCwaaCGb05Xda4GcjOxOG06iZ8Ny1DodZo9aI6aruWNo7ug5vgQ
fzHF/0UJuy/TH/VoTxOgFWV9l8vT0hF5rvpT03680EyEEZIaKY1iC4rH90b2y3BCjg2ZCYaD+tD1
0eDvGj98HVfnSCyUwS90NeBXMdLc0ea0dNrL5i1t8KTPDgfMKV3tV3hNeW2PBWjpEvAoH23+s1xV
4EcqIzgvYG30xy3mE1BczafbuSTH6ZJX8+9i/wC8ehlusJZxM5NAb3KhPPSo7xWD18wLd8yPlgbQ
/2+ePYusH9NosdccKtzJI6znK+E0uLgwtevALjuw67rbMuL0skvtJfoHvA88aPiJ39BdT/qbKGLk
p5jp6BLCSv8wIBi/LCR0UXOIXSfy4A/g3UJhVi307qIGm8qgtcQGGO/fFv4zwnkET722kUtW5Cl/
t5VYKfD/+fsXrLecmqjoOwZhKlEe8KklI9GADoMgbwmwfG7Nz7PcpHxrREs90bMLWwkY4mXQJm4H
mI6yx+wrfJ2jmEsQWNcA7TvaJM1eFtQbRe+FSVv8IzrnLepRkVG0AkIokAQCKVQkNweiUJj4y+dR
gEnyS98lmqtPPyTFFvzcWGslagG0a8mtaI2k5I6PEQKqAa0HkeP6SJSHFLinbeYxVeodY/KL4pK/
21HuUbVSYbEFXDK0hbN7qnmka2J0Mu+f/aKm3By3wIjyHiPbQDndVcWGDxGk51ti2fq9WWzTiEOM
gSEn9f/mTk56jULd/ljneo6rENrvZrvpcakKXZAz2PdBElTuOy7Qwrptgw37skjRxV9yTf86SZMi
2NUGLotGML0/qnrp5UQb268cfEFs+ZNwWrXI2lQ3oiY0XnWtBZacjP6NzmJG0XTpKSFd/O2P5PX8
j/hoiSvEkyVBABRCgt3vdO+s1c3Z8z5jisHpSI1jkSnrRaSRV5xHPDOACILY6MDQBhFgZ52j5xlG
SfQiD833RYksotwIy1HlEq23Pqziucehvy8H718voYAp2VMLXtPETx32FJw7jXaMsQPbeqtPfZAs
NE9k9AffVATiKK7kXyTBUw6eSk/6fX+RSUOquxY3gxA8fjrXCtk8UX8G5qf9ZZVlK/jwlD25b09e
CscLl2HZibfu95FwKkrb4wgG8CoWpSiSsWmluvHinDzXm9vZ/wFm8uKjW7QKICJ6wEQRhVzusshi
GNoruqowosNELdrNNF8zk9/n7mMPM8RLa4g55JLOEYSEeC83hW7VBsM1AzB2yysZx5f2Hv197atW
+d1o88/M8AKPMOWVKdFKsTR3QJXh0QTicak3vwTC2oHqzchIRrw0z5O3uokNuXyyr9DMJmuwq9YD
UPweAA41Pur7fAigVdLR6tAvCH7hAF8kN4c2kfQkPm1m5qtro9Y/LTQo5eq60AJqgjySfBH5pFNR
+7PizIkU1GhWcNP8UiuFj64+B+Z8WFz5SVnuumxQuVTS/1O8nfdk3aOQD1oDzT4DrFMVbiji5ug6
ofcBeS59n12wSnQAmY8nc5qo1pMpARPwRL4UDGARRyg1jljvo9MrOvOtFu9nr133wcXbyhphtaKl
nv8fCqqJbnrwymerfsKQEyzIE28180p0E1n0gFmNjZ8xvsiGqhQvGjYW8XaJptoCaoAxwp+lgzJi
hAm7S2CFVHUMxvnYxBqCZVzijgO6jb/P79j+0K6Kh2tZ9R3WAO2LknIqEkMnHblJLYcC0U8huS+3
bnD6s+QoZpeb8sU25H2vlPjOBLt5kJ7YrbhjcokyOHxn6gLqCgrYldwPQvYnnxmW5vXvBdkEj3Vx
WT9dCpezuW8/tgha0HeN2l5Mguo9/ZLp5VgVGh/dSh+nQ76Xc1zCGxID/pT3amuZRE/hsctZ/ZLg
Z4x2VDBFv4Y9c9rKz9bymPdqXvom/FBwrJVXclshkwrqydVLACFsGdSH5A8j9i1I32zWFYWMvy79
3r+uWvGJM9QsJLyDpvqJDfp+bd4/ArNwuDjPAQx8Wmylr5/t1Z51LlLRRcE8zVvrgWY+8bZXQb3v
vMirLvvJGV7PmGSttmGBO8KQzvhAEVlgpDrd6WTdXqE5xXGD7fYPeEWI2pOtN9AKMXplDiGoqTNS
p1obdHG+SaqC6zcCGnifZioRv1kU5cLtymLroYzr18t2hSEngBd/L9CEhBIYV/qO3U3OUMB2V3QL
2YKUiRxGb5P/0tLRTguAFFahdyxehTyTMgzdIDjB9m/5L9TQE47EDymEp8Fy0wgzSZNVeNredRSU
e6Cw1+kLXwAXAYPN4USgLCLqr49UCZ0gsB3mS473A4G6sWsxvhbQ04ClGkLJzyZ8WbZl3ljjTPPE
+KQQd2BNOf7AVNsK8+A5Qxaf5QpIdNS4rhllq13ljBj1zFHFk2gGC9iP2mAEqiwFYMlUXWNhJBiD
2iowx6L3fKGLxyBfl+FDmNPNO6nI0N79sSyTLv1mR+2YyhGZeCRFYmcIJ1NVMN3qPnagrjJXNOqB
eceFgBma6LO5JPmzO1ov5zXyVbfn1fw+W6xwBMIcq4fjA4wGbyJfDGi/ksmBFM8HFKVYybIi7YqL
iBRsX8jF9RzE8zUpN0exjoj0u2mchBhxiFbIvsa5+H4qgK9Q5TEAxr+L6HRKP3emF3kqd53ymEi0
PJT0bYVDpEHS3a5RP2mYQS012rmSStB6GErtHpVuWqtl8clD4LJBoTV30d2FNdsFWt0zLeI9z6u1
XJoufkK4F4gaVpb4Ak1wr/hwTZ1lGNVH2zy1RPHxyfhR7Ccs8TqNFeKTqrhsSXWVN9XOXP8xRu/+
0AxzAwBiUHzVF61mlheBA906ObyoatEbflhnJhWuaQR3mOjl1UTJX8oBKVd3XeSHzsUyXEJOejEE
2Vxylg6MNK+trv+xI/Yay2NHnG+As1mHlZCx5Z/Jot0XY6QyCCQVoIakpCBQkkb8KrrUwSZbgxN/
fOmizWWs5roU8REBv5Jv87WeL8rarwnUOBPC8Td2EGgc789kehKcjE2SnBjq4SmMShP18LNBoB+8
vsy82Gxh9RTWdyM6T6osgRtAnAvAyrY817dSO3Kw39xi9/lAgcUvuCtNvP79Jc9SHF0ktV1+DRCx
bA1Rwk8s1VS12vCTCCw6yOPW8vCfRrxVZnLwVA0r7iUp7jGWOgJFZ7uCwquXcKLjniuCEw9wNY9X
u6MbzAxmpv1tDs1eq4eqkd+gbQzE8uxENB3VMOZ3sR7Ii8nbLEWB9hCw366QovBzVfeATUhN16VK
Lf4BiRg3tE14EuVJ28GR87h6uEe24uT58evhd63dr+igBinQPv8tTSA9v5uJSyvgfuOIRKc6V03J
/gXKxJQFjdaZoLuPqGyrqV4yMHMFVw6nEcUakohv79f8gT45pgnlSx/1x/KbcKJbVQC2WVdrndQx
4IJlcYd2SfYd3o7Z1XyBuLTtGPyDshqaTm0DrsJsprGk0EMySVkgJVb2+IXMI56XSeEfgEfS+mrp
DuvslfOO3Hv+WEYmBFKY6rkiimJFv4f8WbCsjH9EmMd3GjbDbSrJt4LSPvlRETtrVT7U+jt/IC8b
yk8MhFdoZf1vOyJrEp0lApgW7MM4TQvQBKiXHn6D/SdnCZdoC66GqRTaGWOe6gnzIRHJxKsOdCfB
VXpwSpV5SmId65zl3zxgjcMZMgwWMiSHCzP1CiZJN1I5bM4zPpA2mLioekWJaTsZgu1tfip1Le8I
uE+xZy/+SFbGT0SpTWE1+UM12mpdzEXm4YGIQwEOuBA8xuOQi6lBCEklxzgsBn8fdbjQXTAD0rit
lOPS6zLo4UtKOYEEsmRB8+FpVgwk6teAVmMHBLyJpBXZlyjo3m3pE+hcfT3gNBK54FAQhmGkLaDR
sIvAXppTpUpcuwGvtjf5rkSZlcB88tkkKFwabPP1ybk5UP2DshPMs2/OrQVqrXMUDSHE+i0NLJa4
YJaIkkienSis5ItiN3XXmbGQ33OVwotmhbzwPE+12nnzr3K0s/hHCen3cmvnyazZf+pkv5tOHioa
hmYB2Thqn+9MNw8XhMOr/rdCXKd5hqZVdtw8rW+5eFOZYmzvCjIsY4D41ua/I7XoTc2Ibi/Ib3D7
ROB5LLGP81H9OVyVSw52lVvRTt8PP7sQRDk3NGjNSNQyjAL7SWL7unNsfruqAgH2spQu+hs53rGO
ktewh2RjK10ZwuhumWZ2jHHJA/ulx4sK3iP+s4XCJz+OSTJwo2/OhWO/zkxI/g/FJXW4CH4M5aZj
ap9wgHAvoTu0u6+bQk1gXFP7oq88o4rTEESHJp7H9gR97Lm/0whjOScbEFNnbuGHw4uKQzYAvUEJ
KmDmirAreRWmqXVjmX3OogPq6nviFpruSMderp8a7i+l/1qmVR0Vd02ZM74Xlb8d6t07iX0MEXPC
51OB3cT19aUDSqWj2sWF7O0q1Wd3MAuIvI6K+pK0nztNSt9XKN95JC8Nj29v7q9eT2/KOoL25DTj
qlZ9OG8w1+o2mTDauRcOVDqyT9YJnloNvWq2ExcxAxs/R7Uu/fuRcB9XE4j6Z3KQRbYVkp6lj0TJ
DPLqYwmhIEzKk154dr0j8JOGiulInVfyiQef4C/MzxMHYpyABaZIG+Ypzn0Yq9Gb42QrLcna6vXR
5KFy5WYXj5SoeFRJxkg88mLk5NxVoBdnFV7H1XJrUT1FabnkEaOSNv3yg8GzMbj0SQKjVW/knbJb
Rrsfr9JFlNy6NHEyct7SFkN3y+aaKNTF9FPv1ndy5MrXBZTDC1I0sO8iT4gmPGKO5NDAuD+K+kDz
ws2MAXoxh8AMgbPhsLq1oRg+Qme+stLrC2H7ftdY0nbMa3u70EeLnx+MJFu4oEvaV0Lh6TIWNFnu
DRcwxYZ+zdlilbDuDy5/sba4LEOSYevmPhghXvN60bGsUs7Qq83DvCH33iEW37po9Trdiffodn3L
kWgjo1XWL1/qwW2+fbdvWpge4RpBFjamjDLcQRVl586tk15/ehCDHlUe2CH8ryNAGpNZfkRVhHUC
dhHDljSWQrO5KJf1MiKgJlzGtavUwM83jat3a2y1adjX/JS/0HdpDpPY5eW5K27PzOvQ6UQkyKGE
3d6LxW+vSvGOTEJCVPgDTqL/52wSzm+n3EY5q5GYx23vF5SMp43ap6P1sJbmayjKLxaAXCcHjo4d
1Kei3HlMDil7AihWAudGvtJy+7m3RtFwg8xYgpO0t3M/pfcF+ytO7zobPrxKsVd4RXcNCwnX6KN1
NJ62eHf4bfsFXAi8zSOh/0dffj9OHQVDOJAdyp4lnqu8T7ekDCProIa2uComyRnGPT3rynfQxmnB
y2Hh9ILN3Nv+YbtgTeNOoyqUG5yD6sYx0/9WtM062JvpzBVScYg+k1zbM7xIy19eCubkqFgf1rGy
crK8x805KD2hPrg+IN7OoaO+/B8DWiIUccrjkpBNRz9ytEy2omu3xoErHh4aJzz8mjHPYfzU9zg8
dp6azYmm2wBNplTrgIZfEYzD2SGiyWjpWN73Acl2q7GE/2iqdXlZbVUB92aMQeICuvNoD4omH+vr
z/n5gcFWHaQmcAaLIKln++lvra2iowjwV3ypd1hoR2NIdESX7mcNLL70N5M45JP1qndMhir+OqoE
cGSHqgDz4MLm4pJfIguqYM7MEjhOecsx+fUoKMvBA3oMlKw4UcE9CXE8IsSL0+m0RexwrSMhAcIZ
5F/dhoYvxx/VFfbVJ8wMYpVhOzryQv5LThG6HGdoU5OfkvNo1wRqdH4+BDKe4edLaeaRd2iEdJ0t
kWc4I7LCDTrBEqphBQu2QE/6uabsfkMbdWt2muqFEzpehn/6z7XhoYzHjBv9m3Vqmm2siWxc73UD
YIjW3urpo7Y55UanSXdnk58QJClO7UR5H0ZhIhvrzM8mBjOTkiX09O5YWDu5fTxO8FOnmkctTNsm
JYXNFDh7dOxDvxr5iSPuWH5a0mQpATk+krSXo78KDecFP79TndTDBJ7tRLTx9zX/sXW/QOfgIOMl
diXnQhLm/bp/1AE2f0GtXS3qEFAQtVSAH3J0TOq4kXkDC28RdeZSnTMiNzVplJN43TGflz8KvG6Y
umKixKlSGFcpKJns5A0JwohhDzpvoPT0v0VbseN6ZwCh/CR3KuTo+hQyNt+9gw/WbVewbsIp9pMo
GI2BdtnFbJnboQIHuvu8mkSg4P82nMYV6HHdFL93pCL6rArKMaHyejm7DNwPbqgtAHn9Lb/Dudxg
cWc3GAC9qHPBlUn0nch0/zk0WRW/Q9JXmtPnDibn68zTaO+nUS8u0CFYCf3+O8OetFkOaDM3F61g
molsh5fUjeEZcUTfjiY/jUJ8+AySEDHO5Feh7z61cgYM63wWIpl1VaF7w9FdxqiV4SBCIZHi89p1
LqlUCIqO0zGgDypaz5fY1xtysW5dDlin/SG/dVwlXRQ4tB3N1lBYhfKYlfOxa+fARxefALZGhTon
URkn4PNx8uBOQBKdX/uMprSleFpZVSlRmRVg5qJKob6aGkmQk+ynUtB2Y9J4Kmlccn4cOzjjto0l
TzVk8/CJkJ10Y0fhMiYtYqnFR1otyU9sjuKNQtnuvVgzJLKaJWEyfDR9g5bSX/gRXBxfIWBefJHv
fX3W4aRGyGVF06ifrY6BVNe3nbjAAEuCEz8pJoo2XUnnROaom7kFry9rqAsD2ynZhkQebus70Nfu
pnwHzJZZ4phMkPLVDRp68+Mb+h+9z32e8uCSXgBlV70hOs/5AIKFcMlm5P7D8K3WUIUYS9DahxYi
Nnn1Bh3owv3mDnJqCTWh43EtxZ/t76U2eFxsbMyzH4tbBCwVNGCQ+HQRWb1T5OygDjOMthe+/P0w
mFJJSIacoSqWKbkf13GHQkLOYEpfHwpB7/MlM07tJcwuTzM4kmQm+h9XPQGzDFWpkUwyjU+P/69E
FqNA4Erm3/AUg+dUGOm2ZGhguWTpPWVvm4FLV07j+V3OsJff5SW/kmxFOI3219HFSNNvPnyTvjJf
v8dYjbl3AZe2aAlTaH+A6BG/sM69BVzBxDfRGqK0N3Q9sWADIZnoIRBG9MmlLgYGofNETeIbAAE2
J5dOK0pvMQXCsSYKCJh2SW2qPsBjoxK8ql/qWSa64G8RIgemhyA2gg6C4+bpZ38vS778MP77lLYr
8rFv61nmo0mgCAlGJuAoH7J+WUz3Q4xsyCAAw/mlk91ywwtzBqW+Po1KFBI2JMtnuw3tmk3EL2eK
A/K4wXZKcOliqJk0snzh3UHBXAJFtoQEm9+28yIB5GEG4SUlJPHMUixTEFnOaxGu4ra8GCjXdEsv
rwuex32EELv6DqXmtClExkeUtjjKgLZECCOgPx2zT54p1/MAzczyeebTJ6EWHpAqq/QGpEdUQ8ys
HaETZCGKU0S4baL6lZ7GRQptvJOXDj0GbfYYyrxiUxwjZkvSx6rFWtPzedmK+GP44W3NnJRAzGUX
Uv1KH8CbVSwU6PTUunFzT989bXn4sQ6cKhTItrred5LwtRW61YdbQb+d45Hqia++95FzEJ0qrsIJ
NqsEFtts8CEK+tmGRjwhIiz21a07Blv1Ltq/HZ9DJoeVZpMpJsD9gPSBPjfEhRCoa+4dPbox7hOV
9msWOjTKXuRmCv9m6D1rj+AMlp5RfrkYpXxGJXLRVYtJp8WY3RhOhy5cn6+CpI19peX/uMfYhd2H
DzOwkLclNFnrNuq7pvNGqJyzsHRF1ltgGQXbq3afxX02ahWnMFzMJSjeC/r5k62DPcgpstHrRdjy
+QUgnnqLn9RbaQfFDFh0WfAJHfmnV9L0q0soJAvW+IdrQXB0fVsY+7XLoCWNKZlYg3ylfb6Ya2At
JjjkhI+EWmbeY02jMuc/YcBIxJJgJsD3fZXxlkuk/QyT67cgpk444Ywj2Gqlw3KXIT6cwxKIrR23
6fGMnODhehqL/7YxtYjnDMCg8NOfj6CxRo2rugTZf9O1MvurkCaJ8pEdIhuQLccjvU21DkKuvm9a
BWwaMURxdecHmFvo5CibO+2qa55JC817PW0T4vqA8ad5LAlYBaGD2pfgnw3FPyi60Sy1VyJAOWjz
kCIOSvA1YNOB0A++aLdQX63s6p0Q2CzEAwlb/12jgGMvkRR+HN0l5TequG8XqPePeGTtL/dL0miR
RjRosw/hPmcYcFiOgpSzRPAESrR/g9nX8JTd3FS+BYKlGdEOrwX4MIsrkaygFNbZ7MUbU1bF0l4E
oIFPVMPBAf7OcUGmGx5HzDULGSih+ryqreK0x9rmghDGC1Sqf3JlVPEjWU6ROfgCvLz654lYK2GA
1fxowrH1LCywb8b5aZw+3mdBCfsRV5JBX8OZLoNIFoUS/5WiiXaSpc8LJBA97/nkOIGRvtUNU/zm
LZTp7YstjifbXSIpAB3WfU23B2wWkczEJhA7SXUyxTb2qBpYcR3Abho2G99GpabRV0kXY4T8bvda
YQNbGSlT+uGvCCaWu083dJpX+lf2l0H+yW3sDuKnKCSlKjHUb6zraS+oes+zpPCv06xFtQiPWC48
r4vm17GYYUHCxUywD4gtaWilFl4jfmkvdqnsp1sFSWa3gNW4d4OJoRXGxphAgEG4EX9Gt2hiN2ln
yKNHSYNf0hbkzFemz4YMBb//ZO8gC1ahX5GYrPr6/PlaEOJoQH5Xznxr53X5DzujtI3r4ol2/9eo
fLt4qOg3612Tyc60tDjMnzMvcAsT1CouktTVl2Mpx5awbURoTMb/UPz4A+ynKs8OVHNvteUWB5aW
bEFn3OyZ38Q532xHdVAkY6icEz4cHXPNN3lphTwkKZpZOY/qHMJxKHbl5E3hK5obAbSZJ7i6hjHc
cw/N1PmswwqsnbCtLT+Td8ljdsGQCg2Uwobc90ofVXFWx9PfTFGwBKBz5dCE0jL9dUG6fvUjvP4N
WxBfRPq9WhvVwMRWM/uyJkwK9hEl9195iJlcSP/iKHY6ChX4e8ahQdVWSOrR7RKmbu2Rfmf5/i5+
Kr+teA5l2bJwRQ1/xVStFLla4zHxAMXX1EdGM3i1IftToqY0TCkOgkn+9LVW0MmSvAp6ABIEuUEn
Ov9+CJdALtI+ZAamD103anZFKfVnzIOv5IGNSAjMSXcofysS59C++QH4U3x3KGezHx6emMOMG1lf
jeAhghBpfkRboparp4hP8ldlC6ZwxyyMrDEKg0pfRPTNycQ6aKJCsrX/613eA5u2iLTyEiInsJuS
rFK4Dh8cvy8MQRLeURVJV8dNM7zmNKN7fNzCU7Jv0wS8PTrVJ8FHyxZeWJ2/Ja0scnMAgT3wADXw
fRqw/axn7qQtKXWfb7OXXRYFIQOwktMA8v1/HC9F509mtZy5q4ct36KcgYx7uotYVXzuYHEee2f8
JdwNgOKNJg6ec6lxNlntko4HavSQQtdKeeuJpxiyTaxxovq3yfmNiMJ3YZu9TJwnTBxedmTh2MsI
CaBmP01eukkLf6092Gf80sP39LjqJykBn74ZTsumQ8BPo0aF73HjsHFd8hpngaODeesxRGJAcQ0A
ts7xK2tgKFzJuxLI3I/1CNpI5OSPLrf4l6FfntQTIR2CuaaxgJ+jx9c1PaDzwA/T6wggA5FFwSqL
yCLd13JVj6rnlheI5sXLzpK8NRQChGi9Cby1bS5OzBI1h+bujpNHCCVTJqd7vaFSb1RRYrx+v1nL
WTV4acqrZCMnYWHo7GblS5fcyAcNc4+Br+5VNf+qHv/qegsaIkfEbhH6qJCXRVUrSosxe2UxiWHC
UERRH2gQkWkDXasgNBFqy+YuN+jAc90VX6Ho+VOOfwyqwwvQZZas8YbWoovvRU4uCEJ20XpVijfJ
653F6+51SKXwQlX8B8EdnlX7hlr0OOJsVPymYm4XdcIYJgai13/z4rNLYVkV8mmQF/yVUJl1MP7M
FCKq1+obanPusSKl+63Q0ch1euRt8iYo4neNbGoW7pKd7hg13zf+ij0cUK9UGor7K6eKAHQp4mr8
nWBp40zGmIf+FATOT350t7UyNn+r4neXNsIu98l5pjX8CgM8ub0mumQP5+sf5bOHUDDUTTxjKDSt
kf+XPgSBz6YSMCh/8kOiadE3NXbWQ3sMucxAxZ/MAcMvMxtnZY8i806E/jxifN3X8DfuxHqrgdCp
i3nKD0LMGEdrCBgoUodJexz3csGO+rn7I4XCq3+oJTeF9IqK36Lf2wXz+XgfElrXebar0ZY5mm2i
CLIF3WqtuQyBgzBofurdBcUZGjAbJdD+fP4k5xpMTUWdaIE0NOtvYiXebUZdgjOzsz3lQrf6/2UU
tx01n0FH/t8ZmNucQJeGxE7EQJgHhLduFGmQPVuPulf/EUHEHJo7O7fr4RQd1Zt43F2jMpkNSnHz
AhmX0LWS+Tlg2F4c41ieXQc7gRS06HnHLtmrUK9xJ5XkO6RKThsXJQWlCqVdxBKyhL6/yGThwfmV
M8I0iHIYo+rG0/pomza+UCpjBeR6LB/nHfgd77xjwyk2oVQOoiA6taNBz8zxWSLKoWwENMSIWTa1
ywdU6tQ7aEzB3MtWs1mjfUwSPuXGB8iWvcFEJyythk+jSxN5ZxM1Y2ETVScAs5cRXvaBXPMzXMbi
htiopnIbab4k4Z9QROKyZi9KnK3CeR8Hl99DGcolu2pBT8abEnwRVxFmEAVqbFSYxxTqXyK11q/f
d2Vi3ZnZqxWqu2J/CQtKN79RzGxVOULLKBDyVC65AOLd7A2pCpO4jdRdaUbTOYPHByoDLjTUJVBB
4lQhQpczR3RMlN2u7XFRYt6VJVeEKOWsbLqnTCKiAzbvgohTJURPb21UH11lgXniv8NK54oq1Eev
OqNJkQAXwsAYEEyeRmf2F/NHQD/55UbiJ7//JWAXInPMCaEQqs4BNFD1j4KxsX9OYlrduyqMegQ7
+UiRPfhT6O5/UkZnt6k16QFhG2pBL+TNm8F5rb936+HTPtMgvkxX/4qritHj+KygMjLXTvpI3IZ6
IcC4li2yvwYNeXQOfEmStNkTG1ePXEiMMimSD164Z5+ZOcH0YGpKOZEO1w2+/NqTx+ugx5NhNL0a
M7MZBsbk68WcmjnFXsfp4xlA8Nxeql3L7Hp1DXYOXgfiJI9CzDrr8iXXPR17VQI0/KMGC1czI83/
8nkKuB9eXi1w5oPee0w8ZgulW7VuSyWBPiWxUWtHtOABx/JdxKf9QZsPUVZVK7Lh1kqJ8M02A2FO
IraruiBOrGhPBrr0p7NiVKKwLT05112oV55tH0y9jzUZ5mGZ6qXD9EXdXiZKwgmHDXhQnGKS95A9
59alxIaUo4WEbgARlH3EcY8k6zWu8/qcqiqgppS6OU7oPzP8eb+Ak9KvCzJF6SiBFLQttiHIm3R0
y1M89ezLNDTSPyrPZ1Q5oc3bSvZUbWohIgHWdAqT20ZA0g4vbztpCM7y5S8s0cmYJ6tYcSTYnCoL
fz2D2WuvRNdZygUgCI/4lf8KzZc+8j6TkxpxLQ2zmKwwGzGHGpVi/0bIzZwwIwPd7lt+X6dFalkC
zWRl+QKqKZJ3YEZaCD2kD5enNa6b0hCuXJ/qjWvhlWnWaOnEkCugYZiowd9prgPrhirymkTkYu5A
qRQsPT8pEf8DKt9gRuk+jCnb3ETPpVYhOTyNwb4qBPtcCM7PREXik/WlwwafAsM/GTv3to6Y2N0a
y8SRq2WFNEioThkQQakrG0eb0m1yqDiS9XOphXsiHwy1ursVJX8eB3mPYjCcOBiOIY0oUQYXvffD
iUNsXjGhctW5XRRu+XsB04k501PSodHpslYdpA/ueR7syZhmp+ZYGuJAqWxcn+k784NybD3+F9wx
7RCyX80gS+E1aJDMWS7w+Tedw2UUE/kPcUNqOssgyTa08+/0hZJeWg17GHjIWj74sNODSuSKLK8I
vMLy0AAyNyPbWsvKrfxmEyb7Ndq8GcII1/OsyqYsxaX0eWbsr/zkaUsChOaZlOy5cKftfn3QaIcZ
vVBUWGRkTbxd2HkMKE170daZSlbpOxuUzBFJWQE5YThxDuhVOnq5V2HZQmo3DklsKlgVCvOwIaUz
jnGZLtzlQu3guet1ncb1u3jtX5XpLVpTiQcuKvGE3cVFZHG9g1n3jZx0DUF3wT1kYX+gzYdv43V1
oaWFtZj3DtwAAfis0kMu9jWhbnEMzBklWlGlCMGtuYkQzilJary0SfYR65B5/QQr1JYRh9udf+jx
UmKr9a4gYPYKbVZ44ra9cDPl6hC7Q75xeC03prXRGeGSaxNOyRly5KnSfjDcY+GjvLdYjj1wdkzK
isyNgyQVQ8dMuJ9Agnf3XGFvVKREUF7wo75hxs6y+wjRuvbnz2/OpqVRJU7uagfUYJEmbIKb0JEp
Ei5EX3y/YYdoCseouVO1NThEXDpeg/9KSpSOen7rLCxWO5gIqrffl8nrF2u41jGP6UDV8TIXKT+g
2Dqoyw6EXVkNxVSFDxZltJ/aXdL7cb/NktcsVfpTQa6TjQaTVt0hdp/QjIC9p3jS5N2q+E2HL+0M
YbgNcxVvjEAOEZTzD42/wHCMu4k5JfDgGfO0zZqJUr9px4O5V0IrFmTfj9yPKfqFOkKbxB+eCEs1
ln3JMN7NFtzhFcX93gSRp0/aVfV3bE40GZleAQdaBeoJjHctWFObx5z+3jXY3wGPLQoTNgKpIhfw
78vORkpREmpGXDF6WhM6EJbNpH6epXN/lhKz0GoqCVlE0G3GI8L+coZ1aTw9Q3ci5x2nElMP6Lsr
I8dk8tD/DjaM2BBXMVxBZgQLgdS33nNsedbY1FrHSS65jiUuMhlRer5rWehsUjTLbPSCQLEVF8SA
Zvv4Vb8SWqKq4mLypfzs10QwB5iG/VB0IUgAlF6UR8d7KrDAasJoHDkcbPcYDWxwJ0TFrpBJn40j
i0kPCJBt8x0dqdPyRfud37ItPbNLH7Cp16f4E5QQZR6FGskPJ4WahQZMDp2mRk+LKadZAMRRWOB+
04982X03MrYdlveFuHSxIv0hkDkA+BfL6+pI5Mr9D7/oVzzH6q6qa05CDmylM140tqmOWjHQi7W/
4t6KfQ38RUO2S5ND3Cs9i2cLaY6nLOXsByqPoGRbefzQQybOPQiB93G/85KZz+d6Lppk5o/LU/OO
6hYINywuN1wIVUyZTXeB7lww9DRIp4WmtodbB87xoBrFYKl4SCkWiWyLKvbqVXs1uLIwA1XWERSJ
VP72TJ8sXl21HgIuztqS5zU7XAAux1Kz30K0EShCqO1Qbuuxr0E3etJye9YwIgSnYdyLmHctpaVD
egfRp4gi0ccG8OZR5TO2ge+WfMxIuh13BsJG6XCRlpmFa8FhU0Rx0G7JmJgWN5RyHhWI3d9+BuSe
k3sCnbg/oIifMuCV6wMKsZ6uiH2T6eWxkYahtzGJWKqU/g4GgLRPUBigU1PgzUKikWsnRvanepBU
zfAkn4fCdZery+6kNvSuEe1CbkjV91ODhABwfxRsd1zSkqACwKjlAEamdKUt4rNEA+XrHeeQcnKV
0I7wmNcdX4k1AmDqUEvW0a5EbK23iFPGXNIpNnbAT3Oj8HSLBA9OG1uFOuhP08vaf0VStVwus8p4
+Iagt1XC3I0g6LBDCptv98d8A135tDedM8GaOKSSVYjbwW6GxnZ3x3LiEVvuVhxmrVtNhu6jkcJ6
RsTH2VKriPTqSuIF5H4KV2ayoqDshbN7csuoUScYnDOS/WwxjxSdOdXgEtOhpgaYpwYnnHOfXLrp
SD8LgJGhR7M9ITMklEJV8mleF75AWIbVDcs+GoAox5muZ4BFgTuzSTn6QSU0DH9n01CrVMVdGHRI
Zh7HLb4qVA8QF3XrIZGxQarDfgRFQX3romGS38vPt3Fk1XHfbNRi7kR+19EGxL+w6nn4PC0bbWkX
KDtqEdMzzGcL8uAzakuPi83AdCEBE0JFyaqS9IA3EhBoZRGcVoWerTaVSeGKMFEWWC8M+vg4jo3w
J0wifXcMX2QGhk92zOU5p26XS/TTQTei2ChzM/EH8OFDGM+F4wyQtvusmzJDe5RatXNLG37o4iII
dshXome3vzj1+fDo4OJkq0/UaKcuGCMJm1eouyif7Ws6FcWZwGLd4ifYOH+Lh4qqJ0rUStK7Ccq6
RBIF5/7N+FO/s3lxBeFOZijq3OSrLuhUwvitR9oh0uLkAcqINomqTBPTYMRfNhJMbf32MmBX0184
/PSiepzdnpCQGwzOQd4xhAYmMCNk1b/Y/IYmlYdRPVVIrqGGb2FFt1Rxhz1UNGiKAgviOhyqsz5C
noV+4x39J0WYdHTUtoLt3fkEEppM7PMMdBMmVUe5Ld1YvHZyWYjIW9lFMgoxmxwohVdR1xQf5wby
G0lmrrRMwOklhtL1zm8grx+swbINsC8Mb3v4sJiW7vfzZMXd8nqAY897DnRpDRRvKzmd5be5ll5u
e0r9lXvHrJJstzBk0O4MKYU8l4q6YfnQHVmwiWjiq0/Rw3d8FgkUX7Yw/eI78yc5iDBKYMykCTab
Hz+FOVx64aUWsMdygB2pUhpZD++vOVTCWbPvONJMBeYMots5pyt1ee4v7hRdhb352vn+hGlpCvI3
dY4dUQYhQj5zgRB4ohY5trAnjVZJRoym7FcvnNWZzmVmc5dLSJILc9+WD4HebML9PKxUqm+QeeKl
potIrbUnGa2F9ASd6jenxZscKHh6VjDlFz2tJZC4dKFm7FVROZyOTLSasazxffkDyqarMiHBf99c
pVuHW+qJwhJpTu5l9WsTtJkUPxKB4gaPOzpfLRbyavn/asa9gpAm+nkylt1n8sEYMNFyUbcb2uey
8XLUHXnUobrg7FGDidvXzTR/kQp/lshf8End/saZVqbEeCC5ICDNY+6N3B3WPWEdruTFYjv2pDxY
8mJWhrpKBoYoqLFuOr6bLSCeWRyXaQGjTzEQqFS0sd8T0YZ0+om3dVI+L8iF7AxIfJYw+GPsF4K7
tVCzYeVETKMSWAWG43wZVTV0cOj0g16+UchBMxbKCUpdOPLaBVeMmslu9XMOG0F+OFcbAuScj6Ty
tV8Y5gS+L3wPUPBfQRjRnk3Rou7gLNxUCYEGRP9cqEpDQrxQ9c+mcbrINYEPd55xJv7ss84xmr6g
DY1bHe3qCmgCFH7rr3OQZzb7098toNwEoJQYili2hjwG9g5a46lAtyPKLuRMorM/9Tg4TfqaWF0U
LNsuBri5lf8nALaVc+vcuHk2AwBTfaYc39Wn5xncqmPLUZZrNVudzHVVqWSyGZNxqfaPfzgjLMvl
BTbjSlFaFrOdkLKsz6fg/8ShbIvvQquhQ3ibg87MVRaHwsOJW8wJQTm3sgompH1921WQDSL0zcEE
RO1We6+6NTtT1fXXJifGz2NUD/IlFwVEJjGbv/NRxelAZ0aKPdINAA7IKoVyz9zNoLoJ3HY5xyjd
K6aGydbLjHuzVcmsspoIiwSJe12SpHCbecAOAKlUa9K8XexDGD+ZGipdEWq6I4JIftDGd74KoP5f
lAG2AsXHELdy3acBZGqeEIGuSCWlUHMbrR+QL3HpUO3A75TCLtwrd4gN+DbYjZK4oOzr36i2lhgj
p6astrKU+ubUZPFieuolTnIMiSy/rNEYzvbhtbm/UCyCWs+tTePUpj4H1NPPGwUxKRg1xPP6TNiG
NT7SoM32owKDYyG8ACdx0NtKQ2+S01pF1PbPK1Icz3Ud+zCpQIB/lOLsBzXHEGKfCK5ZlkE4tz08
LkKezXz5tWI2mMPuF3oGy78ELsbhjaLupxSF6dKbY26er6SaUyHO1d+iTLF/y9Q4uuZ3FfFQdxQx
sUFtw1JrcZ9K3bd4HL+26ylyiYeyBvOPkXETFzRFHdR+NLVOAEXc1y6P6MEulu0IL6kSl2VTCokp
bhbfr/xFvrzO5Uio9hAxQra/0CShQRZLT+ykIcv0aME8tVBHjCuBA4EGMxh4VD5x3TGtY23081W3
xzfGMPWoGJtKwP900kjpOabyZXBtj8VYeCOJadIK3npvd8gb46wxCNqinZfzA+ObHW7g3JWvxeSz
Qyfe/KO8lq5Bw1sw31clHqcfzdfZstiy4yd8ertT/VTblrHrJaj3gVOVVV+J52fiF4KmDDVKpJp9
jWUKQGXlqQKHrUyp5K2kHmY3c3DLWPFuxsXfDll3sazxPI/STho/0KhBpVOBZ69qt8YiF+/qPgym
E9tql7DLtofs65adplc2rbSFwMYns3DlnXFDvQNhTVz8zg2iQ+VdxCJhz/wRQY8tkee1OxA3PH6q
JztdC/l71nQU+VnOEhNcH52Xi3cRmUYP12gt6YrMeG7NoZ1sKM4k4TajLfTkiedFAe6PE2px1ORf
zNC1n9ROkY6ceBbdZ2Pv6RmsSiWdUQPOQpqnH5e9mmQtG6cYGpy6XJ/wIrb48ISUazWqrpH6oU1c
sD9QpxqoLm4LREet5oO2dJfXb4/UsII87W3+/Q4IRpdpw+FxaAJIrnDkQ8nwXYdvzUb8651UQO73
pkqre/upYupJFg8QqR5EqRAyAVsP8SE7FWEc3Snz75cMAr7T7YBTJAM41ZJ6VtrqhYRpCXvQK6Cs
+1ZDfPccOkjY7ETnJARaEDVSY/AUWuLkmtj4nSdkXuwAHlEE53r46Nc4Isw5XhttHl1HBhODzDMB
zutopWCzz73T/T7E+mY5xqQQp/9+3aHeuYuyzS8PDCwMzzyS53eIrT/7Db5Dso3W2yng9+V9PQEL
AyvglS8J9rFk7SGX1hJ6qbU/l1DfxfLMZA3xJB97C6zJyQCWRVHm/bs3/vltsYaXbJQP7Zr8uCGw
XgJYD7MQAUqkSRLKTZ/zuOkSMAhhocnhmzIjW5WBCQN++jEGE6WSw6JC5sGneH38m/etdfS6fBzo
bd9835KlFJHO1XPg0ArUy2dV42l4SUIn/+gNCde20e9tq9pgNsGTnUjphA6xcsUpLV3y3b1INNd0
+ARi3aulGD5TjM4uEXZG8iHw7dQrbQbMdwdDgnatsIhFY7Bpy1Uxe48GyFmOz6xT08qwfIgN5uMk
/4HB8u+5J1V2s/yOA3+7iL4LX37eZZieNAGC0eos1TGS5EGQO7+TtWOZWBN3k0X9AmH6QPS4bs55
lrOaLawXoEhIQ7k0C70MiwbdUHbF1hpFmbhZcKR6a18P3ET0zPW0zMMNIWrc3FdO7PuVVtVZFutx
ljNZ0e2qFomlNzX8NqWGv4COAoSX6shYD8EMGWHY9+yI2X+SA8+5NJumS9hRsUwxWgU2+8UgsvPn
hTs6x+dJur/KszmEom9uspXmbVYOT3cT+MJalUsiQ4+H9Qk3NUcu2+5EXqGPWADcg1pwS/++oVXg
kaTWdfV6pgTTrz9/wEGunefFP9dX6n3PSzU0YEdt+8MftAHzmf4xia0fYNIXgIBd7ytbYsb9uix2
x1RXhfW6C/2ISs7KCatz0pZ/xXZKrWtUxfxe0Hf6VvW+7UmGTP7nCjgpkCO9KYwZV3EkWmOpETQp
xuDIN4I0coNscqmXBR30Tm1BNAecyM6RTm7IN6+UEpNKcAgjbcUfbRs2ABVbMWMH2QSCdhcsrS88
qhFaXXrthhystIC3O7KzKK6JiPJ379zDTdLac7xOOHyeOX8iH6RjtuIqUuPefCPAVa7vE0gIxAki
Qcd3Yh4cNGjwGsOBZOSNcnuSrpaiPaQpPRTX7JQd4Kj9xC92BKDBY2SA0TgSlQUg4QZLkNAtdGQG
rfFfDuSoMHOzfoS6YT5JRM5tW2Pwq4iGDDWENsaS3bRGYwUG8ht+1cujBtsvs16spl8BJOoKoOfu
5GA4fiBeon4/+whSs800Ix//BN1sfpNag+dhRdqN8ol27oXbm50BAD2pYslqmXxuMCivxLRys5bk
GR2xjb0rnwqWPR2bvDo7yPqEz/hs0TThB7W4Cmr5Q1oe8DTtcWXF+aOeun7jUcaeCcE+wWhwEvQl
hDmNmVPF1wLwRVg6xwab0sI7RAUsLx+A3ilcPQJupM9KHzidFmxHT6dgWCbZ2fGysG934ROmpZ5S
KOavJFsQBW/mhCZYv8pSWpVI8/HF7CR4HxRkIhVOToazl1DM1aYWT5RHnGW9zQGBzjW2N5WOVbAD
hmmFV8FwU0imRiMvtFvfW058WQfGvlC/7FcME5qn42CwXH7UMikoa8lTxM12cNXwXF9QSbpMZFOt
9yLkWlfmVqpuDOFL3xZgp189p1H68dbx/5gzwJazAH+Es7mMwGft3mn/HEl4Aa7+Shd9UAR0c3MJ
oFhD1BoeOrZl90BRO9mN6Cna4dhlIdcrntjPcw8epbNfEks4EvtdY7/gq8ay35TotHQoeFpUqhTN
iHnOVzw9I7RxWaMcNc3vTGBsZx86W5hi96ojE9ZDa9K6OOb4N6g6kyl+TmgtQmIVpxtDd7YXY4Bq
ngIbeXCdRWCdU5h6BsnA5F3EzB9aj2mr2Crm5dw1CLxy9KtuLJdGB2XzO9XHUKDShD+gVcbBtYLf
wjFEQfW522CSpQhgm92B3+4urE7V0TQbvh8jUvoRt95Frfc9tN5h6aeorJDShOMOSiFW+tFmBoLh
yv6Ygy3HJUbJcXTUASoBDTY0BRwTIZcjYZwbvWIqPaj/8MtzS7WFeLbdQNrYQDLPpA7Af3Yx11co
bDuCdSEPNh/x4460pLUiJSFVY7lo3sAQ0WMjxrfTZZDO/RhKAGarXsDFL/6mysSjDDKCpAbpeZoL
H2XMNNF2bmvrzzJWBgrvcYTKgxvVURLNwQ/NKRNVOYuVAc40RSqL7HnMd9JpYkbqPHmZ30BfNrHX
SghG7R9h65GA2OrF1QHPhga8JD/Og83USrzJM0E41xyDHU0gZ98QEJoUkOuHgTC/Paf15+Dx8Hmz
F/uzmMTvfrD8hCwuJ5bQ1uMXJV7Upu+9Q7x+6mUleyXxrds0bF2bRD3nJ0zZjQwY+7LapY0+qose
yRyEejZIqhTOQ/SSswgZrvOBHHWJe243MH6iFwTIaiK/LtSteunhdsrRUGoGpbUxsFGEMJsqn+ZM
KJB/ZjfT/PtRm3mbCRDqQ2SDekRdBlyJPrB+wcI2qZhJ8hvPtx6A3sC6S1M4uDv7buv1M/5KOBsN
gooV4S7R8byTgmPrB7oS4mTpZxZTHZrMZfFJm25CID/gY8lBFiKrSii4BR+4Dt2MaWiUSuTJHrWu
aocNRJiHWUl1ce5/5SZxV5RdXZiumTP/IPtqIjs1+/1zeNVsuj0GOShqvloeUgD28NFhidLNGQL6
gnlJKDs9AEqSsx5RM0JLL60uGKkkf8yCwjWUelvK1ExUmSai4NH6+55OZFqSHscrJFZ+0EBiWwTO
xeoDJmY1e2e8WbwmRhu/px9/dDM+BrZkN7U6wHhfzLUeU/X/vNW03tcMnm1t7253VP2aDrxAy1XY
UA6fu/Ky/t0s4c63QeYdMiBLx7AxiraR9XvaAx180pJdzJWPfziPpXDIHJ+WRvfWFT0qo2+bX6E8
+RTH2+HINzLMlwLZdZAK7XO4mNByUtSBh+gk6sObCiVsIktgSW2J78cqHbgMlhy20e0w9XkDLQjc
IbPAPwYVu2nco48k5xCbPsNfdJezwk61O0GmJ4mgFd373JNNdUT+wQ+FqXOTyTOn7GcU0PUcxpDg
OnnT0APZ1NtPd9NbPY0Mt45OCkMLljF2szEi0+6THF+QD81ZXVCGszCeVGlJKevbotc4VCQH7of2
ZphzN1AjjFhI4Q22xzCHJc0vkVegOaLXzxRhdkRt0+fTLM/98ds06gA/p2h7NkCcnBZeP0bNwxES
cYNPO/FpNnMT3Ks/Z1b3LkHX5cbCxmnQ812Hbin3XgX/0JZ+cN9JGmuIEZVKrxtU0cuiB+Z0r68Q
uqo4TrJH7B6x/+276gr/bNQDJ0yYJROM2cZsMMNnxgoSoOvIaei7T5amBcYyp2GZAriqVAozpl6k
8VaXHXIDx/4EEaWePwCm2GNMdHq+Twh3tEbrp+P+6LPU20TLHSwboLGshFnRsdv6kBaQCJVa5Q8h
JeH1lAH6FMptYYICZ5tOcO0cqxu3fIQz8pAtGSgMAFHDorya0n6TG6ZM9qxEQjcy7g9jkf2XF4Ft
UHyGlE8/3XQuy/BbOpZ+H+m9t789yrU4/kgHNWzWmxS2KwA74xcqvzt7lLAfSfVJtqsLm3cM5kpH
CgZ7IYYYe4CtctVOU5aAy+Pn6RlviNnBZYkoAkPn4RvqAB8VH799G8AEQZhQBbTF/+CG0EczV7gb
PtzktCYkM/G4f6osn/HFNYkXlqdj5dgQTgbeOedFskG5nBFHOessCC6GGh0Lf5hgMtYcjJCFx70x
y3n0FhmlHfjx9DVaKViU3GGaH664XFwHz4Pfa7papCclQCPCU0zndc2AOUQi9aRWPGqA2OgbO3Ja
hanoYIA51Y0M8WjZ8ehwyM9GkaRdRxGS3iNb9/z56dTch/yJLeGvLse07yV9L5men8YlMBbP5OK4
dg6RFJxwK1HhuaeaPnde/AZ+simkJSx4Prs5uLz3bW1lGnTTox8tXeQj0xWPBktM0BWCgnSJ/IB7
DDg8JgAd8VKcem5VRXTsH8UROZ/sI3RLqjXOvrZ6QcP9mk/Xnd3XlOT60GEcTFHmKlMZCz60hJBw
mJRLh4tgylMQeL55tSmO16tlwtqYihsPJl2+9BI7urE3atKEvt28frMjg22qqKs4q8SsQe93WtjA
aNjw4FJrwpXZRNtkgwPxzeHwlsm70BLn0x6AFQHbxni6lfI5D39HMwSIqWVHvMwIoVKwviNL1ieJ
X1JdII1xcsDuLKNat5lBfLb708mx1E3ci5br94Z1okzmdoGkxtt4oZ0MD7r+ysjlayxLjG14OCIp
IKVcMQcGjTDrxzGxRrxwe43VJO/kI4hVlSCgAkQehTOjhh38+OaB4Si7fk40elQjmrR1Sm7PIBF2
09tr7v907gt2RraKYF5vAxAftwUV/XLPenQC1gR1yEARQDV+Apy/4qf/GbzbQn415h+BKapXUDvz
j7/1DlQhtF9241OWDSwMz09SaJgL4E0uATwfWNis//xEB4pI1omN+Je11AGl7B+ssJ4JZcWW5nti
PEdKW5FgGz9eaecwi+CXXX2b3AnHl9Dg2C90TlgpeJvGZeHx/tCUa9wc30g2ho5yufn/ETj+jYaO
8q4MsnihiXyGBgI4Yc6TSEwB0lb4OZY3gQvfdpzERnunLAbqBKDQY5Yz1m8INHfN529z/mHnvstx
bot2yAJcUVomEn78KzC7gPzgChXmxwRXfHAXFTvkXnuoOhOhZemYjNH+0b7m3pw0KiH54aIqG9q2
RSTN7lj12ujhfT8fTeuDNc2P6pu1LeXShZbZwpsZdvSmiGh9ioqvi8UxtD3o5hsWUFtjDz4cfAje
WnZocC91Vqs5pxD2vVt+oP/P6ty2651XFutX58KlhXFMLAYO7mOtrqKFGWxXgzfsjn7wG8XWqUvr
+gW7Ja/sjIl2gCO6zop1zz3d7Yj75yyJo/YQKdn2l4/RQAOd1nNbIIhuoL1t7s0I+gXmokYNIMRj
tTu3RKq5mDcP8tNLMD4vt2tinw9V7QLQIE+4DRR0VmA7btjMB8JP8vMIzzAhw9yKoqQi105vgzPN
vfIk8xR/9MyBZN4JqWLRTjRWhl5LvVc7478RFM8sC3SGBqYwCe36RbfoPjeQrn3cSS2WxX3wCrqA
uB4nlPr1822nXVbqrlQ7Sgb+nEh4+xFZzfAk49trjvY8E2oVHiikxydfYxBQ0U5C4C1nyVO7Cb6S
Zaszlk67Nvyet3lzoRdmo7SNtND3nonWxlElzJNx5yRUd1fnmhtmvLj+apjxMGbuWRdprtanw9ek
jHAPcVzfeU7cPWire6NArdWNarEurS4yI3/vQee4imErfT3pZV93BdC3F57m4/kEIeE8JWQ7NxIt
H0hb69/LSzkElNdFxNE3o1TJ4OsalUXheIRR2q44B9ud6A9c5N7KkwrIYTWmEm26rNTZVp/bGB5v
ol0g9BrEGSYs0ywvH1vZ10uJjIRMW5HFMMEPp4i3VVwgwF7iiA5VVNCp/4Zi9s8zm+gw/BuKqgAm
5BrkYZvpi+hGlZWeQkkOJ/Mr/cBDurhi/B24o2kLF5HE1axHOL3aSMb89pFPU2e+AqgyTZ8lfYzZ
LzJMUrBlJQDLSmvxGLJ+GwTG+8Fy+EpibFOqLGYzFPcd5qKiINYfh2LqdXFtCG3WpnIcS2Nr+jNH
ciuglnSG937YOYSZS+JdZmVtCsJHJXyksjzzo/bP68pvvMLG5GpB5nzQvw77IT4HJZNxFkqk4UH5
ecC88HJDLXwok2DQ3ZA4EAJeE2sKJED5Q4vekdDCRLHTLDyrZvSsYXrL01i5W/xs2FH+wXuuRX/e
PYbLFvR8ls1oKjcdjt1tAOQYaVmj7eUo8163KADndo0wx6MMLhryp9GQDo4YOOOnGo3Itde5Ihlq
ANvh2NSJgDcaBXlRRZhH10pKrP1WgEkor+P0f3J125PMh/kaDj6ehCHUC5kUgdFUJ9pSsAKh10bB
nGaub1JB8xS5ZyClZKmQUS3ysYXXdeSnNZEukWOm7swYr7pFVfzg15VZOUJTHaZW/yg9PRZlGHb2
Algk6Nr1Uh5GAWBVkD5/7cQAfxjFtS6xBGSXApzyAjUkXzUSwe6Q3Hk0PLub44UIUSME1akAG8UY
C5sNMUXFJp52uN2UTU68fNcfw/+o9p6JizVf1mous1ovOgTyPqNpnJk37yC0ow+OX5n1aMh/hkNz
vEix8slF+XvnXkg+xJQW2IiqCDr6pGmeT4ljPokaPDVpI3xpMqRYOSVPUdQwrRBLKgrvswNTcnRN
11B3KMVLVgK7y2wOYGya2BP04v6ex6A73Q42wJFnAn5lTG9C9XeNKkq5kmG4ZxRUtJnc7jVDByoE
9vBTDTS9Qf2Bc9a2jsjQBE5vwzthjJi88CM8009Y3Cy4umEejrgMss3aP3X6CjAJxF0pBqfsFfMW
a+LykorLn+sUN1icWCgG3kjcsGMLQuOtJOTU31zLiz+p7rSN9v0IiI32xcEqLZDGFZFZKPqES3Xa
RPZ375CObLx3KkWrhvGo/PUqYgDd3mGGfSLEu0/LRSzR4rIYkX9wx49Q5NiB3W9XoalVHg70evYZ
Qmm2tQkc/8UyTmKLWR810rvA9mIL3w4amoKPREeVuCe7t99dS+gfMQ9XvOrqmXD5zfDO+sYyzWx8
e+QwCMeLYDkde7R2+Jda5Jzr4/q4Kibb7vxA8XT4zTwj6l6hrl4c1+vljFvUbTzWGvLovCBVivCN
zqt+5Ldm7GdRVI7RfBCcUh8OLVtzWJ261gwzymI0bieQA70NxSk7gPFBJd2L5uAhazTE/wumL3Jx
zEFbZC1U0UNiJNuxvO2rkpGwMfmehgNyCfriXlv7GQJPBWMS7DcsPOARWP6MZQ0On5V8Cg+w2CMZ
9HdgviHGHRqieNPG2VPGO0lXszPAtUIy+Qh6iIgg0kgbhqcnu9GdkHvPBxE/xwTLl8Xu4B2/KR+I
WzRkJLm1mLzf9hTz1LR7kfF3zNQFFLBSeaz6mAnO2Gh7C5Q+2CLj/Bk7BQsUG+HNeYqMGUlBlLSO
zAoPZpKX4eacuh00rJs3Xhx9wR2ZbMzR8aIL21nbFp7eChWX9rZXf/NPBW2UtDaNE1r0Bf1NCaAj
ELkJhp+6rPNQHjNrWl/wV/3B8Pbolo+wZNnZ3ZJV1+FBfeJmS95KUF4an6kk5DIKKJbmgWhjNl+n
cGc2l9ifl3uja6JESz+S/BuvBH9FDsRH7lhTUrEyWk/+BMuXU/igpXekCBbF0lc6NxuvtoilwjUs
5zpvEfNrmjScfzIYiCDXsqbl8Bl1IONfPjBLwaMK5WxpYBD8ElHbbLNPfK/9Cyme7w0b53TNAfOL
YB1H54Gp+UCxCvRHAehBZqbiXHr2JL8H66+vy+cpFEsDmYY5W21vnLOZCIbZ0wpHHbnWWoBr+GjD
6p1aGcX/et/TmdoL2i4T7lvcC3UqXGg51wvxEQ+YDyoVl+OUliOsvenam0UFK9T31WqT49VVNTD1
+up+QcR0VntWVIuOXj8J+ksqCfyXgHF1SEK1XurORltub+NuZcKzb1Cc90jNS2E+x1EnEYFjZZAG
kq+ohYcMdd3gbCssFNg+/DclM8zRgUC2YFeK4PnyqFa9MjppPH0XV5V20gVjGrhZjuPFJY3B/2S/
MSwaDh3nrCBoSUS9+SLqvvmuvjQzwgG5Ds3p41CIRX2VBhpxnQJ1J0aUjl3WOqJyOCjxeOv5TXnn
28+lA00IAE/KW0pwMLb6dekxWtmXA1e7gwpJO15gz4/okZdRB7Swf4kTDaFTjJFUZu0vo8KrlwIK
k0TtqYd0JPyVUEFk0XiEpfyjYvd3mT/YMzUhAu5Td00Cv0FBvykPvPnLDxO90AdWaMy3o5+uq5j1
poSX1wuLvRofU+sXljZZ88JvQV9iYHPJ1abk5ddil8kuuUjzEFq5WTIazVYsSVyc7dA7NYbXOOgH
QgOXpMGLJRL075VE0o2tLOlMYbJjfjvY6e1HG0TyQoe/TMQjjzeeEWAKDZvGkh47umCfryuYuiGS
cXOhUW5V6I/nBReHXmxXrWuxM35bknSiZJwNpPB1EHQsOyIDanKXbJkSZ4t6AJDp5LnPL05QjUsn
aPxlkKjyse5M/3eSdyvFOKwNew3dBReEpGd2e/qePzDPC9XtM8iy40YyAVyNEnIlhjgW6qHE85+d
uXZhGntvMuJH6j7Wm0yjvlX9MxxjMelYoUW6KZyEz5QH5leosF77WwBXKsYK876XeK9Yrs2XBewW
cPFbK8q/K/5wwBqHMI4qJHbT6Sia4O7mvks7vtLfXC8ln/vDcWQTjdue2ioTcw+hRmCHEybnqsB2
IMXY+uD6DkI5BJh/EWxH7vZB04RinERNs3P/LFzZQE69cUwlzTOXPrYng/m9Scvh/RA+0HmCRFYd
slwPdmkG5fS26M9sf+9dhguX2VzNWQxNHZbEiUGnrgnnDzMCnvzTpULy8uUWP39DY6Mh4hXFU2d3
rGAy+GxUj/E18hpNIgFGkIYxRkqPZ/9wDrkVFj8uzqX6CKVoVH/TiKsma6g5RKarwTsi6zW06TO6
tVHbHSJDgw24r25OPiV68fxns7QSkeUMCe6euaeo8hqvedNFPqen+Fvuigh2Omhgk8vHU8zEYQjA
nU3WP2x+CUbYYOWXvJtWFUzWCLUYeAxPeCgNnsAs3YGncfjU7AWc4c/NLbyLlH5jsw1YbaZvK+3/
Trfyo8Dtou4bG+e2JVMaRg10j2Ba9gQ4FOFBdLRlVao/KIF76LMJ494R+KZKExL2URkWQO5rDUUT
IQHjf1+EDVJFBQs89rZy7HI9Zs77Z55j/1NOqy3M7YwVgBSXFmg2dCMD0j42T+0IIiftmXUaOFaM
Io1E8XICz0/3k6omjdjzZUXjWvLotGEVzB8ETEp8GgrjnfUr0KZbbjFh0bU2ZRDrKiWzDhWDYJbv
6ANX29gSVKL03JZJantQUZxmWD3v4UMxov8xd1DaAFHdIr8d/KMBzTkp2Ymwxxn5lWfysakIZ8x+
OK2KH3P4eY86WihtUjctqt8QG+e84scU0x28Lfm0UnYPOpIfGMHUIJHdp/GK8ci4RCHc3jcUxZvH
aNNlCxRDh8dhOndDw7F7l6PWF2lQ1Axv0+MIXle0vZnTdHDRnZ5o9woUpMqJ8X5jmFbhNuocFxzG
S/KINMG6VX3dqfFI1sJdnnynTcGACLlcx65vlTfjzU1pV/f71mibSYZ1K1eA6KY9bfxCLO9zaPE8
TiLp8cApFqm0nCTZvE0zHYRZS6M5BvoDYKetxKn6MxdFBdD36DTR7Nw25uUd2G77PeWq1aGGtKc5
w3Fh7izNLxH6PSE85+JMLKSgpfK8Nbp/v/tqu20/BgncRFx4GgEQoirwjrM6U5RzGFX5Vk4ctJMr
GxSHluwgCdPBtk+nNbbynvng5w1C0T87vpy5KulTHrjkbjQwiC3G0fMq4sioExNSSvSequsudVev
yuENVrj5bcQbvygLD+6YvzWgXgbIcBmCrHxYXz04U8JYZZZp2k8ITLgVCD8NcA7pDLkb0Cjb6SYz
k4Mk5L6+4NNMzwSGr2OlwYwc1YMB7u5kz6OcwGi17TWybg3FDd9+cwk3I59UPBAqfECt4fNEeES6
M0dw59RHVK5L2Iae/q9Aeklf1U21kxQeDrhfUbfgkFE7Q02Q0ZbJEI0d1yhGnA1k8tdg3fKKQ3sq
vF8WTcCzLBv+GrEBM26sSK/ftZM0oisO1W+fuWzChGX55AKzpPi51jmJqfH3OJ28caDkil+aA6oh
RbYoNO4HnYiQNJAsXUT2wsSVou0R7hxvPdvkMr4UchM0JFY4jCEo/8nJ3+9iTvMqIcyKkzFf6fkJ
evbHnIFKYhUfCEJXsAN2Fo3IynYitX4yymhiejySDQVcOMLO8+R0PvClyB3SuGlrUOvRBnzaI1zu
lP7cLlXAXPPxDCVzNKLjPp2KF5S4E6B2S4eUj7HBIFXd+LfDTKjv4fZpv9pxDjxMHRD9utKjM3HY
l8U52z/VJ5tcJcPpZmESFhezp+zB1NiXMDmCh8fHHEYs8Ci2o4Ve2a6yIQXJzMNo2AzhTGgcMAIq
5UUHWWGpfzoO1n6JaUn3BtjD1Nab4o7rezcGc0g0AvaR70F2aCRIlqOaGcBNzPbMhnaCQb3hxRRd
s3ITYTmCyoLqSG3uhGzYzfh6nvtYQ0G6iztRo5ocIKlccxKm+WYuxygiM0xqiGYHgRzm6JY3mbZt
Y88DFYB/FPFzwNtQixb135TiRmsH3l2WNeO2dswC6+aOEIVaGdTK80+lbCI7U1n5pG3+uRDd7a/g
1QV7y7BVT8bmGnS5rGR+ySEVN8X62TvGrS20VCigIHtEVuxE7l/2n9fxR7OYJNgZaELbWqYmLA3z
NbjtmdLa8GHuAT5j/b7qqdjH6FyHULsb1IisDoLWKVMTcEvvKh5XlRAUJGmBu/AGaCIDVAq4yQgE
q67I6Z3jCyOpRnXY+h5djw6cYrvX+Z4/TJNQoxgz61tvxBkA67UsNpOKtgXSL/4U/WFzzkFA2CAO
mQuLR5rvwKcuxjOWHXxWEqxWhGBWyxE4CZh1UyyAoms+jn18jZ6HvWmlDomWhtD9JLk0ctbN6Kqv
95gPeXks1AxKCNIFlTfopBBfWjx0L444mxd3/5tTBcYOGQFz30k4D6uqmEyIohMYnzV6/XB16qTB
XlqUowwbFzCJ8ZYd87EpIBmXxPQl1Dm+FSQRVAKCh61UbrvSwo9oUVeQ7uHE75ydpxvuLis9Yq5R
MWV9jNaNWDYsfog65gr9oS02pjHyM48Ow5HwVCCOQsX1deB08M1YYH35OfuhzWEbD1Xc4rBE5ahb
evdOpK+XS5ocsJ3DhsfB105qWHAzvy2ZMrqJkhSthKCrG4dynJa02Je7usJXJFTDYmanjqXtyjXN
2ia5ggiqo8lsSUSZ+UKWdLkPJ1bw6H0UrJhaPP/N3YSc4scJXkOySdMXRDLllXY8asqq5n/SY5v0
sZ27lIlBG04RUcftvCvc/IV6Mu5WHgyJ3h/4pllGn6AywcKEdUWVOP0Ca+1ivK72idMaltCJzZTR
7RNbQMmL6lMuBGzhfPWyKsvJgfMiT+YCM16K06rvH/efyaa5MwYJnxl+FjHsNtERYJiieibEarts
pH1CsGw3MB/M5y30zJw7I+EADAhIWt6Mcb96pVdV5v/H3GNL7XeHen0Ig4NlN/754QM0Ie4pfS7m
suQ3dbF/4QquXJIdubVBLp+wbrzqj7b8v1pll7FfaCsW36KOARiVMMr5fvLp2eV1IVAM3SToxJlQ
SJOtEfk7vlwAKvZtAJsUBaxDRq3aOFC6ZGEoffH6PB6spv5BuOodhSgi9C2dCZqundcHI9LoGQJk
bKQQiZ6BHUln3AGOo2OAQUHefMr93MCaVJ82Vj2YVk9+8UQ8jx5ip5/L3pXhPCxhLhzINR0RY0yq
lnPx2SeIId+ct8OUM8GFFstryK9M/H91GhT5ZvyF9P9fwa7qvDSBvuZ1dVzkDwOAP4G7UG/YM6Bf
/U/96dsTcLdjxSZ5uIS/f+0iBM6QtJV+HtZ+KwgAdPNwuGk1V9+qDv9hQpN0zPaM+RoKe583b7EE
Db3TNq4JHYbVYS3qJR/dKsjjaO617x77SinRogy01vj+NZkP25KJBaVR5QTY8dNFmUnfSnuRHLEE
xXJR87dsaVacvjROYP06wz0Sxi9nBQpRVL40TfKub6vHkNMfPtxKlDGZkUJj7HV+A3VzNGnwQwu7
nJr37mGJtWUGl8AEJUFcfax51s41ogUB0WvruvhZxMefJ3cGUPGR3PEVJDGLOcg6hYjjzY9iha8z
vpJr6lUml8zixNLvadaG/ZkEFgPAL6eZxqMUe7vJhtU3RHf9MjGV0+MV11D+iyGlZnnkhw9lBkOr
jxp4nNjZX4RkKCizQl276zboSb0+xgJ/5+YK2S5MaqP5DGaZ0sHNKzvfQO6zMKlhdKaR1+swaAXe
wyUo1JzXAaK9ApdPk73bzJ9RSyMf5a38oPOMQ1l4QhO1cvG6hFjHP8evcUal5uhpr9SEIMgMjz5l
bT0DcebOSLZkC60n8UkzioC8ItwY9OjYF0G5GXtFBOm/IQLKHySWYnv4za3jkB2dY1QOlDkjtucu
yufFHdMJ2Jw8I3H4hUIPPGP0HUq7Pz/xuw5gUcm5LdYtxDrKzDTmiIDnZAoxS9bOUA+lb0xgiAAn
Vww9HM92ldYAkLz/TiUu7zCdgkgkA3HtaEJpFcYWBkbXFsBE4BUb43J8dG/JDKvMGOW/szBqpHzA
SjfDCzCNGoQbvDyZ2150+mS2lxtzvEpCg7UBKcM54trBWWv6zSe2VLeMtYHkL8of8JAaBPwlLy4o
pUjolOswcBiSAOYmH4QaWNtGmOGnVNpiDGQ27eCCAFYvQxqe0V27QfZsRFeVzKiDmPzyrYinfX0G
+m6HxuRZHvSJluzh78c1uNpHnMAg97+5oj6pdFmlvrqSY8anXv6mNDaxEO2kd55DFqGO6nYFYhgt
R08N+Ris7HP97lBgXCHEZBbGCO6vmKbgB2keM+g+c7VTViZe6DxDKs+SS1wH3Ve5Awu6LJdY6zXR
s8Q3V8GR7Gj6CriwFQS1gBoS8k8wsfYYk4DDbefbhK3SWwJkqld/p/49e3kJoQABoDiiAyW2JU5l
SUWL5NYHajw7w6EBUEK2rWqPuWbdLde79yF2LWtqSXau+FfUAJrpfOM/y0/UJMvr7+I4ZnLXqTkX
La3OaBbDUHFQSQnxGyNHXPTSMV3yX5c2jpvs5Mrp9SbaKv2C2ViR7Tz0nqQHxPUxJQIi/6PqBOhF
KZ2bYxNX4Tv0dhNqy2FRJZnQLS02D2QfU/h9sy6hipZUnz3Ln2/9g24YA2DTVw4ebL+wbUQSHHos
Zrk2DOHrACx/SXgfJ7QIEEz8adLq05eKwvl8hwfMSOxmck5j4jqXU/wsDmFxT+GydT3bIWB8/RQw
Btc69OFCB+gpZt+EermpmPyLpNWKJVmgC4jvM7PAeXuLhgoZfQbItaR3Ti453/eLmcnj3sATEP2/
JmZZzyH78veWM12D4M+9YNaaBV+DkwLARRNOxpMHtW2U6nqXJDkpuMf25C+rm8RXvw2emk3N3b5I
yIrinhrSdJ6Et89oA+AP4ntkFC+lGPf/arYn+L8RyZLMEGgOlOczBZm1e8pVMYZ5/gPE1P9HpUsQ
0oBoui4BnWpnt9lvTW73uxTsoZ7CGc46S2eNKamf6yvtg99JkwstCN8iKBZQq7XjWJaeK+jhmXHW
SZcNg89ZwaUpXG3so7WaHk55cHZtH03T0oQExyD021B959V2Nlk3iA9pm19CSQM7UdQDQxEi7xsB
ZTsPscndAgVBT/WT6EHdiAxgQklsnLatD8ncaR5QYmYfA6q0eCuO0Shr016n4mGKEA7woMIN2/EQ
znUjknEfVmbVaTx076sbtcWz9AxDmFqUk9MEUpzRC2D5UcCQzVEkgCE/YT8FkkMP46rqXuBGDC9M
b76888un6u2Ro82IUqp4HtY66sCo+NGjrk+RVPvi2aOtut7anwZQ654/dwp7lC7662Y4I7x1zB+G
GOIBJmXEjmi+whxGHxICk1HedZmNiUtFpOVWbkYxrMmGfzbOYBuOlAq7WzMUGS6Ejx1GKnSBUAis
/vCQ1SqVROr8VMK8H4apf0Po9CZPJDl8FkSDpHiEjHPPbcAppE8ubk6XgtkvHyxT71cy/raY03sn
HAPxDYsXSf1y4YTEUGOXe/zN2UXxxR8Xw9hRs5+WpqCbXq9i4WloproJWLdi98iDIYz81ll44xT3
2uDPwBSGBeSmsqu1agNar4GxGnLvY+Jl43wKHRXIdUnrQUauh8CQkPL+Zvp/XOVVKMGR4KfDgtaZ
ENNWJkOQzR9KjiL67GfG2vr9/cKAFHhlkbT2iFDzu6RCpMJH0YSpgIfpag+FcYlcvqEzGv6vm9Te
KhhlhpPXuKBnZCHqWZApZvL4yFwEixY82N7rZs65nieiDPjogn83HFoCaL6nCzHv0L06fMnoH9Of
vv9VhcNuEx8KP1BlecXpVit37yAFSufS2sO1TBMp9XXZJWGEl71nSUsyMWteoqvEyLozPywZNBc6
HXcRwP81ce1792ArSAAReVsr5SwfhSVzucZCAwzy8Iu/p9nxhLUQ77pIy8JMTIZ7vHa82MGgXLsY
43X3Qi4tBORcTTMLHsFwypZfpiOXsrseZNmuvCeDFrFTKmo+noaMhiz68M6lj6cppb3gFjNTXm3t
emNwkIM6kTH6iPsAe4+TVvl80e2UsBYK1EmhcSGE8qU+/1myGO7A6oTSjNXwQ/K2lPeAgNV24MtM
9QNQtCjvtagluOQJx/EGlSzxQPkuOwQtNtP9x0BLhHt4fpqk+pjRAdoyrLOo1Lcz+qF8ct/26dk9
IVO/YsgumciCfkL6yPoolULMyOzSillgiC3SmV0UkjmqzLfPlpjNPE8Dyy1F7G634gC+7LS+h82c
EJGTXgOwYL2FjB1hMmTeCVIRlamcJkrIxpe0LBjdXHWg/M5qtpYxfFkWPYXvRf0JysJsn1UzGPb0
LyTLGwl8yFvvq8bRSF85jRJq4asGwmzG4kqa5NXdzFkOC2V4IQxeZ0Wy3yxi8IcJB/fABmgiQ4gL
k4497fvJ4Fxt6AhxPjKnkuO/OYdvr5OOe7rUgYp7enFTliYQSH+O5UEMuPOzdxu0ePb+gVyD9Chh
bSZjfHQI9PvDz6oCXIIKyV+OKAFJmgDQ2azvpATAW4iMQh79r8EJwl+Dy7KNkQ7jxZxjkKuYWesm
OIv4f/fGIE8cVInIp5DxcjKNZ4ZTcnamvo+XIQLtwTk9/wIOhWt/iQN3vNjWXsjdipiNnMRnRSst
FqaAanb7ttsTj70QH/B0iWHt7GlHoHSM6P/jn3AJs1dL8JFFLKemfAgdBPDFTP2882/w4/V9rwcl
MANu+08Y9breSWiLFiQTcXfYzJTqOKFh5BGQlKjKqv4VJ7g2bo9PH+uhylQb4VmuGmtRf+x6OT1N
isUp8UzCFSN5O07vtwEOq6snCsLIHaV6RNU3xXNMbBQ2eg3aY8farhCJKVJhPwtBHPqSgr7oZCLi
T8Be3r1kdP/MqfgZAxzPzAkPm5Mt8lCMzuDtFThosrcPTt20+eIR1sKfeGLX3riMc8aQ4U9T24Ll
isumkjo7vxU1Ktbs15UR+nnrw7RO+kbi2AzgjVonwHROp6uQeHHuYmL2nJF0v65vC5BBKiIXwKgi
mUZHhOqZlj0RA7vJI9J9NIuikzVNbpLOISgAUdqB9Hgu4sAXi+KRj8pO9u1uflsgkBMwtwi6LN5U
cTn6jkulX1iNWdABoCLaLAuH6rPcnJcC6+9MGyPhwhOlmGaoMTeOXmw37bkK9M6QoKW8JusXfPMO
+TbW19Ny2QpPb3Eo+/tihDpiDfiPLod3Y9fK7QVmAJLcbcs6BqN5MzQxJceW89JryQFWNP0ZagBy
yERq0ZwAAIw35KPjP81v+vz7NrFiu3G1lCsObC29cez+ez4D5DdtwcLcgoiGnd/5tSQzVXrNZgfI
Tm5ix0BYHTLZ3A4RFx8eBL3+LtvTjD+wixlYJBGM2hf8Ay/yNqZDQh9Upsl5KCAWrIwWQJBXWCWE
fxYG3BbjPaPN6TCLThVDlrrsa0BEamwX2rRjg3u6fDCL/OI/QE3BI95iSRXu39B/8yatuRIA5tgP
mEU6LCL9Yo78WwffuWYuftqE/373fBHrcwZqkcdR8J/047NwcgqH0oPY/krVmnqdXOtFHl1HJJyT
Cd8YVT33KUnTbJXBpUh1OEEcwgl7G3qYtPbfTMWwWiOY4/t9sVkfZpcSY4tTsHpeFZyp6XQ91Hz1
ZThliJDwrPgBhxKc3OZwjxA83f1wuerGoFwX/qN8aD//42bl6q60NWFYoePOE13PtSuoTIH+QFfq
FvgEIKQsjvy3NHjCTFB1TPYQb3fvsP1Os3eGOX2zLf1h5S9UwURwiwhAYvVfZstHAqVUy62fsN07
IShVH/obzsOtnNVD0XZVLmjI1aCfWMT34J+sBCtvUWJjm12/Cz+mo+6UDAz8m7Ew/7jZtIpg817T
96+3EHg6SznSYMR393XS8ULqyh1zVoyJKywg++zrcBD6GFPBSRrwWB8Oi7ARTONXf9/vKt4vib0J
6o1FseeR51J5LEWKmf8Ksd5B+S6TURVlAWlX6/hBuldUH7RHQ5VxpeaaYVi4ZDZ/6A6WkZyi+9Y2
p87/8vkT0ZnXxN2g67J9vyFKrkpIh/EKTUPADOHwdpAXVO/9rJVbLaB+gOXd7qkAv9B0DXUSuOBy
/DRgY6dqpjjLalr+JGXK8n411rMw8SwWWPi6UIil6plsjrBBOoII6nPhHr1JU2/rY0oazvSN0pw6
q8E8/U0kEwkVym+sxvvkV3grBkVfPhtD1paAHs1B4VRHdY1pUOeWCfEoEZK0ozjnhPRL0qWx0ji2
N+kf1PyAYkFi7HJyUK1j48kS2554d3ybLpGq+6yMgJq6+yk+dL9Ynr5TOZ9oRS/HvLfIfXDJs9T5
LfCuoaDq/qPcKSGbNoCLgI7stLYzvN+KwOwf/umfAhgw2miswtkOPEhkfapC+MGojr84mVXwgte7
Xj9d9nqmnCuCuX0m1GBdh9NxX63rcVw0HSr3rJ352B1hlQDswUU8W9fI3eNlqY9Ix4rjPbdxO70/
et4h/bE6fhp0PG1YQoT5ylfhmF9h8epbZmDB0wgNPiEGcf/cnhRKneXvy/KfiANnRUezQmKWpPGc
/w5fo7xRMYMgSDeY6lm5bFtEb680gX+9bFI1VWcJaVOJCDOA41yNOf5U17bnaX74GG1ZqMEEVTj0
uzWvm4oKa43dTAQeLLUEs67z2Au0AfDwiDifpX83lkVtl7+J3LCocpUiFYUQsN4JGIhr18Y9FmIB
LPIakBLiBA6a1RezCH0S2H4n80Zmc1kz+Jo3jKB4cBsaFhmaU6i2D7orr/af5du6uTiieVIy2QRR
AA+tO1322//4Jq4Wm+Vb4susV9+Sc5LpnCIH5ukx7K4WHFDpHkWPPoH6BsQrQL/gxNsvUW2qooi8
T4npgZH1qz+jYVqA0QzxS1+/Vbr58KblSGIk5qP+B6BAwYvVwUoa/1vPkYX0hfyv6vGJ2Lq+gHKr
VYmZD+j5bQDTojeutDo/oP5NZ7GVdapBIL48cbA5SpsZYZPvjtY+Hdu7vGeprWHXdh8zJCcb0T4f
cQnflw4KQEM1HgkztV7y107HSENIwkquR2YLu7txpD+gKcgEcRaa4EUsHmrcbauBfibWklukJkBY
MgBJgZjxiD7SERhbFBP7tBzSmX1rLXsIk4WKjQMOW5/FPZwOwcw705nSOYz5WluYTHhQrodApM1w
xHh8pKD6d8bq968kOTX7kbSEY1EAG5FK0f2CA/P3J0fkALcQY7bc0TGYTX/pGrZA/Yz74SnTtZ91
NnWW4bIxfDfJzD8aMqm/Itv3UJVufPUHdzUgxbgjctVLIQ9RjB9t52aXnj/L7WlpPcLDZU3c0j/0
iRwYhQO2R7Xd92srz/b+w4OEUtMi3ayPFCdqrpaGUkZtAH+883tjl1cpMjjQ3iRibcb3vjzbhnzJ
pptPmLj+uoNXeGY2cOxVz+GEnbdqr+EcZQp3jDRY6VGqFpUSQXN3lSXtejX/+5Y3f5EmudXamLtv
+jPsYfPqzwNa02Yi0zza0uzz+WeI/rFC29H+jKdSohtZsFmGPctpuLv/9vYsce2Nq3TIKpyQBDdc
vLXSLSHh9jUcN++SlzpMQfU2X4K2qUJVZzK2v1j678C0kWElmrgdbOoJ0t+nmF+THyI6N0wUkHm3
5QOMBEyBoxjDPoEu9sxWflBNP6EGmzV60ExouwRBZ+6Jd0ZCRk4NWzXGMEhHT6kQsYRNO1qTtqgi
nWiU7nDpeoDGNbswZpC+/PIU+ilqntBDiF9Ndc1iu4NU/lkYCS84oZJs0jxr9HHzluNuBrjM25zH
WDKRMfFzwtGhyHfAeoOdieyxTL9zEwnu31p6VzSR0PTKsCQMKt87DK8AiUxe9AEK3230ExIcTw23
RYTZUcg77TlegVp1Bcq0tGu7j0oSfppkYnIIKklIf6Nb/QMKaJ3EoiN4ugQQBjaw4Hycr9NuOmg/
nvjN1zbNPXRK3zCcL02+GmZIo3fWIOqiHlKbna4+hKd1XdoTvpYc+9TA/RQdq4fPZVPWwbOZCh4O
iM03n57fSb4BlTmsNXyPbY81VmWAnFsv40hRRFusw43NYB2XIIpZ+eCUnZyKdArs8bT1jdQRzOSQ
z7ZISWFXVuqztWr2cFoGnzc3RiLIObSeNqXCkJw+rb5R5S/cUOcawYlKDkSyWOBPhW/ECQKhXVSh
lHum8ZZZOd1VTq2lc4fsB7uSvhD2jBgZg0FPiWrAgJV3+KGynaEmP3fNn2/JizttV/NV7YcdZIG+
8TAwhHrte75a+cuEuy6VP3ZBKIqLOj3qGwOqCV7SwlBbIeUbTTDs2QE61gPBqmTsf5TXMD0UhvU/
dc1FXiIzhZNviMMwDCfX5UgoaryoJ3SRBPxuUrSkLoIJXrxwswEOIl5MJWRw7Gf1r7PhaSAJkwED
virNUAFx3VvMRyaeRsRSbtoGfISDOouWMZ2tNfOZ7VDnpT5C3nT9UUJrQPkJoQnv3fHY96T4vL85
aNGpWNkjHb+RHgrf3H+n7fJEmYCSu+e5y4qLxsIiEFlTlnEkpYXJty9YZGBM3mOWQeVoRsEf2r5K
vyJm+i2z0hnpSkJuix2qPwQ5G7VyVYTV/HWw9zI2Ipl5LOLJbnLbQOT4GG8gwJC+J3L10A9mHEhP
Zzmjy0wHcPoCMgK8gdfwHlF3DKrLhTDPgZxdlfdrra1zshhmLiuQXFTlqzjhZlOxQzQrET0qjQrt
pzRxVSBfpYJgg2A2xXfz97ijFzNcH7ISRRF7VCUaKP/nj6SjGYJZATp6d+MTPDthbHLzVyxKoxir
dn8xiYSlRut6gwm1OYbEy0XIBrlNXy0GMbr2XnydYBfaZNSciRJhSvlU1/fgh3mAb/y0smko9FxY
cQrlVt7c+4JwE11G4HUmAzQdE/UqGtFGvWIhzJcYedofydMGnmt9SqEUJ6Dul4JaAo6vUknTE5PZ
ajHFrJW0TFMEtYdh7K7Igvu6tGg0qOv0D2hqnVI/gJ8unsKYhtSCGDPBDbHVrnbJroOAjSG4rANo
lV8l1qXz/COM9vV3FqwgFMtmAubzjxay0ICWVGearulCdGTllXXJwoSvIC2BqOOAfvlbpANr+YIQ
UwbXMs4dlKcz5kR1AbRgqRFqdEI3uqU3uBYPbLHm+NrQskWWyy9UIaUH+gmbWQWHtGbYi95w+Qly
hQBh5hF4Ajp8Dj0U0LjViXVJbwW0JFJrFGE5xyRLLCihaR8xdMc4VEKMBBJ7Idm+eUGMeqXo4rlg
cbhEtxySWavIeZcsZfleknST1mTDL6brJ3JoHRI9uBzdHdKAZ1zeeNLbroI9ZwTO0VSa9Qy5KdTk
PuDIGwt6pijDyNqkhnvQUST/yFQVBz5OwmgNIQv3viHYvpJLCOl2KmHAwb++xVO5GxRm0S1EC/00
7JRi2JSfR6eP1b2GH+ojSUMlKVw4A/AxWZem4Slwe7CUimr8OKDEwJvFJL0Lt3sytK7KFYhqYSPW
wLjv9JgvfablWMgrrP2+IFMG6pSW0lOotjsxb471ppXRwX1SpAaOWwQyDOHACiHWdgPUP+fRWQP2
NuXRZbHcoXPmf/66z98N+3I3x7+4Q3h98ktWZ8tjBqe/GmzQbpTD9kJgmQ2TCnFr9HfqRoqbL3TY
tYSX7lKt7U0nVIDmkf8vPCqKOZvTf5d8cVQKDTXdkYNNuS0R6aDBFA3oJOC2HtdJYgOrMz0K2RW7
nr1/1+bsxUgMQnjdGxLwaADqMMbRtC81QsMXpkROGRXSoPBQVxGoEKdkiI8fp/HSzS34vXISPEdr
rHB1mCU3urjQQPPat1d3y9G0d44Bp68P6mr1zldzoNMrTHtHqMM8tth+3Av25j6jXRdBHnxWQ2Mw
15qaKKWjtUW4fQKNCbuQKH5RtHmO43x/S4SqF2cZMRmVVEkLAKdlVg1+NQjaRwHB6Dq19r4FzriR
Nj0QM4PdPPz7/Y8vUHJbRBGO1vYYRbpRN7YpajqSZPpO61jRj+pEJ1Uev7stOjR0MduSAkH1Y3a7
BV5BxtgB1kGF2PJpw+EUvw04lOuS6scLBWKVAdZBWGCUDdfs4yoWJczc4enuhATG9xvq9EUlCCoW
pvr4Kcr1KIUxQXyhtgTblLCr0I6cwJZxfFwDVFU4iW+2It5emLZfZ+V7xJ0kGUgGp3X+4oKzjHpT
OE51tdLdCJ2Ah/9mFa//LpUu+QjuKCqY8pOkkfxqGdl1QHj/zmqX8QBlJcmjFKd/f48mJCUNIAPD
xkdLlVAY7AoFlL2ZiddxgIunRiDGzInB3qSTQbNbvYV1qjWrwxWIBTEP9OhJPEibK1imT1uuwbYN
8fcwMbLIS7iI2bVErhxG5ee2fOZrIk0Xn6KXN5Co+iuL23ls2vPXd0kNR33yTM9jMtayWJczz3WF
kf+Pw7emUKByM+RcDY0hCMl6BLds9unmf0PR3reDH+msGn3I2b+DDVm7J7eMOf6DYhDlxghlVwVX
N4qJeDzY58J3Ki6Magvq4RuCOLVeuPx0FL53qCosNI+jE22c6z3HsU5/8iW/sYcTG4VU609kiegP
lkx+E4xFlY1dF+0soJabJOPpq5d1Kd0jK3xjm4Z3/zyZIfKb8A/2L8TiWE52VixDHwv3Cy3pSjE6
QefdAs0ockdeln4MqY9GF3iFFkYCoMtrK2NeVKOVhSxHuArLvwMh90GMO7iBvSUOnLj1S4/xnKLT
MvZJV8DFVtumNyWVL/lKFuXl22LtzaLtCMsSFhPEcMWv+1YA1fftKiMvGZd+JcPQl2sJuPEFHxgx
Dwmq4avBKVhal4zMHXZM3RWICz+TMWUtup4g6WrbWTTYQAEvb32ZHSH6tkXmUq5qbTs5sdg1KeXV
T/T35KFLN0g3xO32OAw2niz7tWFbM0QntfRwNdklasqmBfb0s5OOzzTIJtLgIe5i8wdHCA9LAD7S
972X75POQaQhZjNzbtZecepiqGRLi/jkp7ylEwUoTDmJFqijQobNcP903ny65mQ4EVgy/OAm22TP
MmPwc5Bzkvw/lIWYdEPbQMbkbpPM/HlYmskHYdWvnOx2FoPp3h2Q+8bD511ixUOWq/OEQ/EPv3/g
JUxlFLCY8RsPn6JFHwezFMcRxkXEnSkN+cOe8l4q3705TNnc0PoQR+0WZECLmtW6+TojFTNyVcHc
ozLaUpeKnavQFQ1RCFM0FIAt91PBunHcR/kH/7SwliFadffiyWf08u7MSlJnX9Zqn1ZAjslFjQt8
e81kADOgfTTyVACjGKdjcEWwWA0wcpZLBbe0fABGOuyOI6V496AxdhCCI2ROl9AZy/Tcr3sG9QGb
pECkkzPHJk5CelZpFN/PcIOxUeosajn0uJxJex+YSGuv2lj941/HX7tsJOpjV69G+Kcw3hZwc5vg
TZ8EWlr5V2yjkfreFESzFteRE5u6kJb0LhC6ZwpsD3QLDlqOO+Q4/sbefEkSyrqTGYPm3CbxawSG
f4/PjFDsW0TBx8Y0Dik7dQKt8a5+rtIXRSomdyJPxPBznLDaxCnMXeimYGdU/9bEhP75mTPsQeW1
73diyGqJpxXi7APkT1P1fBsvY7K4+v9XAExsN9NDv2aCYaYNofM9f+A/bkqv+pkWlBaUqYtD0PPg
kVW/5xNcS+9H2r+VhctoyqeDJBabs0Rv9ND/b/q0le4XcVse13oepHDI3evr/9Wl9PdSKAz97r6C
RtXV+dPBW9/NGUX6EbnEOZJf8canSzWpOyD26zjLkLAWDrA3gz3ZHB0sio9gV7ogMjE5wlnx7/Jp
gpaarrDcW8FoCr7/bvlABJM7wC01yiCe0Yp+R8Hdi2gbfjJ7li9S5K/8ZHb0lIjMCrJXgMHsDtZR
xTVoOg+iGjSwPItyBjr6EW+VgO43BmAHuYcR8BcXdIkCrcuu9NkVPK8+xnwwiuRl/iXFijaoELCR
28OZDFO5fYgwC4tX8WGyg4/KyD1Wpjg0QC1Nhlqd04BlVOG95r56s9BAI2WbA62hc23W4f6anf4M
eSAwAWbyTbwpvKKfnIaAhWwscpexn2yBAmHLFtM1VMts8JDtCiIyi2VDl68QMfRN8J1lsqsBzUtC
a/gvpjv9QW8WcauzjbQs3pqMylWWNkN+2WI8OoPAZPmfsjy3wvLR7R+Z8iWluS+T2dyajw7FQ2ge
ZbpsccoLIabeSlbd71mijkIqxNupfryOYUGUCTidS8hxJjl56kWxHeJnXy2zOJHQQuRQy40Cq992
0vVqOoswqgbF/Lb4IvNM+eISJKqkg3bkpBhPPgY4TtP8wwyitmSaXxS4jNZrosnJ/O3AQuZ9wHKt
w5SgiafIBUpE7wUQ89tfw9mgS/qRs0kz+IN7whBBersCQJ/KKLEH5ANxWji33v40DDhxBhA1kbeK
QBOO4r1tc0Uia8vhzMfgZyxOu0N62VyQvGzZ7bH7VP9G2OEGZ8foxknVXP03vwEx4XZMl9TDNUxm
tnqKv28CtnE0YBskDbp/UfmpXsejSu9RvwPl3d9kDUm92HZ8Iz0Q+YaaeOOxHlqdHfM4AbCDSGXR
RPgt2j6Bn2g4/fDRgj9sap3wU81ux3v97Y2Y2aO0mvtGxa1ltc1p+EBAt7xcoPQTL/Ye7w1U7CmR
GAdggzzJfZ3eUZqVd5aPwxzL0ZIBlFlmsdy4kQLmDyIhya09QiShcDuP2xZTS3EzcGc6/80DBDYU
8cJlyL9+V01YBWqGbKuGYAxRWH8F3/Cc/ph9Ae01nXk76rveyUlqpG05qll2YFW8CwbGJwWv09rk
FQ2GhekUO0z2MVkSGsvGXkJhAEOql5NnzefaSMtfu7c9m/X0MY5bt/gqV+MIaY+guYaNSaLbT5/d
s8csR+p+df8Pc7tiV9iEv/xlfo7R/7NIDFsU9YHDbY7SmhiHMPXXVp9H+0WbR4Zsz+Vlr5XbBl2Z
pLqb1siiYCnyQXqFFGHfODYgJH9QTwsmK7roJQVIqS2tw8Y1pdT/+l5zs1BU7kMEiscIVH/jQLNz
vj+oRLfgGXkzulRKwSVwWgyeXoakPDVDmH8xAxspIAl4Apu9ljEt0ZXjfjCEpOJc4lc4lu6PhMr4
nAsJfK5gDYdc7xDv3fo5wACLui21KIPe+nMO+xVbc3XFDXSKYH9uYWK+jka09r3EuRDm0mDvpuLu
Ia/wPerQsJjE9v09gE9nu8isOnvVXV1rvukU4KT5QqdXrSMDYRLH+w6ssJiGzN/N+HxFSWfOqD3L
HZmK0erMyXKnkWXTZWnrnivMIx68xG7pHUHCetZfh+QyacLw9t8lrnSvA4G3FoK7Hu4ZDHxxvzCJ
f5GiJGR4uoM09iSWr58ZHUONX1Aut1Bjw6ILIowfHh+J13y3XQX4rtDJOfFBrOq+ukiv3wHoo15a
vcL1FuDbem7CwEuww0Rh4h9T9SdiGjnc6Uz4WlkFNrU7Nz8Uz22KTbihhnBWGsHUzlNfyWSduquf
s5m3/eWX3dTnoAzCVZInRNqPD+F9ggS4GMYtNr9MujA5AKoI5us45hEhNl//PII7YtcvdrsWbsEm
p8m7eh3TYhZc26YU0v8hgwO7EFeG4+L41/zxUsKW5bIJH16qcvg7pQfFiTZDvR/L0Frj7aaWOVZ9
gJwgdL7H1i5TecXYSjzugOPc5gfbjOk+IREX2mzXn5xd+STlvzJMk7bXm2W/QpMJG+SrOfy5o4MT
OHz3A/0K4P4wTF71x5E8WW5UN5DLqgejW+TO0Na12rFf+WZEQUGKII9bhnbHLXra7RGyp3e26FMW
ny1qKW03b9xMksJOyiAbu6Bi42mU5T8vnLxhUndtxm5hovyBDyfTAAgynJc2RCWf2xzgIyr6PT8+
u3InstJ8l/zswXkxptD0+YJEIxRWZkt07CGL3Dm8k79sGP6m8nPi8njfQMG8y/pSDMHR8+nRdOBo
u8eeD7+oy6mVJHK9rErPIfvkD1Ag6W5fb4W62SGxc6WHLFI2zgNbfZlQ+u4gaslM2YEh+2XmwADM
9pFMzzZzVct3Kpz16Z6xCL5SRcGBY9jUzZtq+cjk171i/GplMPJYGdjdavpIvt/bv0bnXlg6/9RV
+2gKsGpYwKUIwwer8/yXakvzWhar0RMInSDd/KeBI5yUipQOdJcqqfZedbsgln0geOl3T4QMctMk
65rANAUpCqrAzHJb7key0MOYUkavm8Q5Yrjq5wu1euViFnCZljAu/I68owuJ52PLNKvJyTwnKiJT
2b6PXx+vp+BUr7GbEq54q55xTAv9u1cK6wCQDaZwieD8RlByTZYvOzS0FQY9bGkPont0/8sslHmF
kfkNsoMGKk7qQRRdnwyqQvj7MtHj2v6g++vyWblf7Zuw7bT+6FbPdwAoX9RpbPwtRGvYM6tIoGx5
125/jiGeohjvqAR0fHWUDYha3nA6OMZNvKAIdCSWRJX8ImLw5TN/j7T0FdtbRx6OzwTE2fjUVPH6
f7UQ8n6aeVMG2BUOwaCsgm/NgXljUtjoq1varkn8tSlF4u2ZuIjNLkFsIMxBOxEFXjztktv4oSes
r9FU/gdB0j1xnpRgliFwWgfSsRsJgNB02E+qMeXHNvNkwtFxvSWi6Tdj+6msa6da0OsMFyC14JHF
53KAPqp691GT4JZiVvpx21TkoeFNqePMhhoDZ41MQjsO+Fp2h205EC7NGAoBZ5eq7WeV7M3ZYX3N
VqjTdVi54fkN6f+xM08b5uXf03uPDS1zfoy7tnAgmafyvGpS0Co1M/4BsI2nZbXeVoE8LW8nKZrH
WkLrLsppqGTwvwese8hI+xKIcqGxlJmJQeqqH0kgGmQeL+dbh+AKz36lGZkvbAGUyN/6dupE/5Qh
s3Pk0/bHaPnwoR91Bus6ukwHnpbDNIpoRMAdD45JtQZ1ZQDDiFSSVPgcUrAW3qYC+YCEfwqeRz5i
KRm8cgEKZ0jWEM0oenHY9y4ok95fP+rKiigGWLxp9Ph6OKK5eWi2vy3uFNkIySpUke0j5HCqhnf9
yiqlT9jpLeD4AZXuJwN+bKASzY51joklMRQV6W/rUVr6rUcwGvo7/PPNw0YEikvjSaHqlV8367m4
TtyKf+PpF5tYAS8uXELYM8g64qFEwXeLW7rmR3REx36kWzd4XIOpru1XClr3Ese3Tarsbrq5nMMu
VugwrBrlZ/JansPZtCYVbmjv87qgdTk0MUC83p6IX24pWV+JKdFW0sZo7CFnLOyfyl57BsybN23b
GhWfUxDA8EP5uwb86LF30+gV+Yqgw+dw/eBlIVUVsp17ahXGp4qDf0e1XW/9oslB8O/Fmr0MVqvQ
LdSHfa6A7XKpzeztaYYhnOJylSyKrVXe2O4fm/URbC1SDyH0oIJL1ALj9n8XJuOretXD7FzCM7Lz
LU38KR5cWbfafbeBFYeusK9Exj3uYPN4QqTdoYBbtPsFGCQsR1Vmj9xWrPkdyruWTyyL4Bl49W6J
gw0NVG2Zo6HxjleL6c/wgfBHzK5n0pDWlz+GC1NKLQn8JpMeBk8r1X4zGqz71KUoroNHIo0e7Qkh
Hczc/hxLItrWsRsm7WA4fR89Y8HIvx1ttPZXcuAXphczrpNCriJPCgEmBGGJ93KzhDEKJwR5D5AQ
2k/ealu4ZaB4Pgu4rS07rOwTUnfkH5jGITPE3fYMvwIKNeAETQAcbtuFbyBGpXDsRDcHksHemByQ
6smnTV4TvjWRvY11+sdw1CwbKWaOAA73KRsXOMgEtZde5wt4WeP/2p3xGhfZ8csxBx3SIiPk4ddF
pkcCoyGwj3ClskvRzm+VM6x4ksdE0DQW8nKPOP8dwnMnTG0Yz8p2eNcDvAxeQADcz01GOPbeu0Zt
UooI0h6u15OmAdY12q/NZYbnoqebZgNsfBWrYTHyifuOz/8ub4h8z2coG+0BEuYlu//4gmpXFjGw
JPer7mSXZyj9zcRvJ2UaY+LZWtDlOHTUGpVGlHPH22IfvhAEGe4llZjRTYoXUNqSqVZwzvPYdCOc
uqBpwJRu4gulaEAlng1WWftT6qiOAjNgIC7OccUy8w8+tw0vYK8MSzwZEQActyYS2UF21M3UKjj4
AvBcsT1tZJxegmbcc8Yd46GLEftwcq0eBa7pT7KzuYYESleNk5Gg1oXcID/5wIlE2WgzpzQgHRsh
o4tPiBoymlPAYWUmOKFYGGJdjPDopj5k+EnsFuprUCvZnkDu3sKAmfkEw4NRSdSuAjgPtKCJdf5o
+PrdNGTt9XZ3cxKY7Pi0jG15gGzsAtn2SWLedpLXWYYPRVqmRqzRMxXDUmpibmeCsfCCD0BZV6MZ
roAl/zRxV/JMxsXKuIFGaj33S4oqGc9Ur3qjymoYfry7BwzJ4+os6uNbgSrdCreE3IVE4jDgTH6x
3erAdL+Navi+8hjzWfAKU3RuAzzKSmOG/nlyYe3MNd/asMaRySeZZXPiWqmYPEZZ5vRxO96Eof6z
isap3DWuWAhC7vZJP8NjeIZdFyFSYMMWhOEVkb1a36UzlTMA3ChCocWREXN9bVfrlqYqIQ/oC+nN
iPbsq7A/zQkd1pLPmMdcYe1LaViQv+5jF/8yvsXhPqKsVNwTMXwJrJ4H8uI1vyyCDl0dcfHUwrwo
l8QYj/w1JLzSuXoTvbe46Uk7YQia9u7OJu327PjWf07U9RuvITfg6/AxCOheFjAxcteRCBIpH1dH
aWjXkybO7b9k0xoqtvD4UStCg7WZTlRQuBNW/mlvqfJ4vWjLMnezOlAYnW7VsGUBfHLR1fpBY7Wq
RUmr7K08WyFhyeYqF26SK9xc5hPKBNYev5+7WwuiLWsJCmpqwts5+f9ZBDcyp/mRR4KcIF4BE5SO
1DdabnxBuIAAjyubyd8tY8sFojreuzPiwnE/Zk0QD6B22t335BzJiGI6mslLn70u+iGPMV5cy88j
+cszvxOE+q1gCfKsMU+G2jh1OlQLywosuqz7h5jr+g2A26ZLaWW0kP6++POJLGuKHSn7SGHQ+Dai
Mm/UWadefbfzuSz4N/pliuahpzl/uyJyhFBEVkzHacbbPNpa+ZtrZJ7EK/ikXfcATkU2zyxHiof2
1pvsQmtqqxBiSUUWmrx8CRbPaD0orfL0YlyYqNuMo9Oi7EVI1/OVzGtvnaTK1R6QsBwpykz4mT4Z
edR4Ty1731/oXlr5Qsn8jbcEMJzvwZzkIUCDxmhaij1EB4RynQr0O6JIMtai367yMea8j2rw3jPa
VURflvjIa30nrldSE/hW3pM9tHMHurJyWPzdq28pTcRi1vgJwi98i5r0R9xPz1fCyMEwNYfmZsj4
QdGvhu6MkjOTaGhJKYsm3wCBRLjFk/ds52E49wGA0zuUKubkR2E6LBcHhh7GWy+fwPUtuMYx8QB6
eJKXii0XVfRrl1MYGwAJCug4s512Nd622ovuCl5cZ8zMDjhjJfnidwd5t90L7qZ6dUMIbh77zX0L
xmXgpD1IH6VGRmQpA2A2S5AzYxcM34oQEFBGz6npI8JBmRbA+rtg/3RxzkeaW+9HEDKuUZFUlO5j
rOZO9Oc7k3i0XERXvRCffpVe9GUgkZaEDjeFhAiXWBJ0SDjSrFwokSgOrPNf+rfN2XHZfoDm7y3F
4Z3ezrFhH2ejTKyVQ2L4+H+GSA4XfjFb4v54I8lol17ZU8XsMkGi+CHXqcuyWL7/LPdcr9GRM+zr
NsPu8woHX58SDy2AZbz40lSQQ3L8R/WdjS8Q5bF0R+EWG+HIVSF0XyoNKmXn0MZnYFUGvvxDzxZP
vHiDT0oRWfAnCkZK283QKc8OgTHYs2pGcGFVJ9o3Tvx9LolPlGHburajZeIbpEtADby2gvWPdQYt
Eiq/ngQrQQjLgywlC1pw+fzGrQqKKw0TOwmG86lmKZxeB1zzGa5ggcFYEO9DFTvsJxuStsqjvWMu
trk2G6uJp8cVvh5UOsvVkg2maOHfPy1ZCcCvCuO9nhWLvNLMDirJH/5gWOz2RjtOifSA5hO+jiDY
utItB02MSl0XMUTNquEWKSmhLHRcnTKiDqD4vB9fZGur/N4HVIGsZ8nUTa3nknWkSnrulntG28Wo
VraFHHag5+B+Jq0sZJXe2JqQ65BpkZTb3YQPeu4woq9J1nOdMIeL8BLLoUzLiP5iv/W4Umx1Jk74
bN2FDg3twRnWJLcFxw9hKV1AifD6k+rkyhl5NrMOJ683BgH2vWksygHvl/dpyvu4IZIHqdcDdozb
qT2L61HUCLDCW2CwvB4+NJR5HLJtjMs503dnAQG7u6bmwZl1qGxcnV4/k696CtIjWIFg79wt303o
a7L5BBh/ISdSBYvKkLB3KJneNiTNS6ZuTthxTywFXanJDGCKKAzm/A89ATzRr4i80ZKkVuJV7bzm
b7F/anaqrH3gIIYzntBd240iRAUvcjdI4g/cefJC5Qrdl/CPijqUEPgBCefBmj+0MvJ1vU2lrVAR
viWjv8d7n5/dbzMJNFl4wt/dhRwyltAJbJUYN14qUrBErcMgtzug5PmaHZG069KmlGMBjXuTtALZ
uEQEWCpiPLmdA7NZqDM4mN3vP5t//vHzc0udQtNRnxjlGhoRlwn31cB9mM7mlC3BkkNFfIGmMMZ9
3ik6zoZjbkWKhiMiHdzdMacIr7e5zzmqJCJw1LCbJxB4YTpVMu1Lp3dPDXzf+rGN4V49dbDhasEf
7lPcnOAmZaCDtayWRO+a+ufimz+dTMCtJYIYlrnvbpQClMl5KCX8kspHhbQQWXGaVDxiZz8WYyfP
Vyn/COPlHoJjqQm2vFuK6M7JGOEZhmye5zXtPXlI75b6qoQwoKgA2FwepEhuG6gTYqBfeKZckxEb
1Oju1VzFFvAmbWuSBPZ21OW7d1xrvS2axXpDKoE75EX41ymYLkekQjCtZQjOEWLCwhkawOVibQAO
Eyd6fjcqtDo5yRqp1ht2bUrNYO0+pmPRntXWzBlx0PDOgAtJ2gN//jEF05ZB3dVt9KNEZgD+SuFW
S/CFsCypgo7/LVBz8Y1YSPsy6ZfjXFmGU14pk24HENmO5SM34htcD1WaUpvo0O2PBx0S+T94yK+r
Yod3GCVX/Xb6+P9ZurwGn8n0C+iMliY9S/HgZ4We/g+flhOuZAxrl613EL1SXLsDPXkPulsdlhmo
ApF889/GfDi3lVddoOT7x/004UIF0nntQy3vTK/HSqerJuSYngBSPOzWtXMNvZzWwsB+kAYE2Jkq
p5W/cU3Jdu23RxwW93JpeTUXfRwBRFRSU97azlpAu1LX++DZB79MQeMYAvQ868l1fXVDg94YKSdf
Ax+nU69MJaouJhkgE9QFi9Oc/VVVyLli3ay+5dCeq4aOHZfKQDPLCmUrflqh4JwPTtLtT1dbc7p8
QZBPPAIy6OUm9VhjXkJUDI+Ojtzd/SHBDuaoUmbFF3Ht9jK5df0Fs/dKbkjGIwZje2o9XiHf7PEX
zG1hUiMFJWiBcGJNdFcGfOm1/D9GTVfryfuCIU1/SdSr9H9mdUZdFCFbjAYEbckoVjXBwXx+0JIS
E3u2hqEC9JqkU0ziC1xzIGwWbw3YzspSfs1aC6RwQmDNST+Y3Wy7It3rt3hSUGIUkZizau0fiL5q
RmlAtSO/BSKR28wXc6rxJ6eG6Tu3RqDZJmL1P8Gnvpi98C9Kv9oEwrVMXXy9bhTrPWPRJrclozI8
14WUKnJsaWoK5+gyJmme79UFsA0HTmGb6X40VambKPIC3KE3LenEEUq+Yhi3tNq4cS2vzWRKzrmF
EGoBu25jfZc96s6MT2W3fBZkMgmSYVSab53+XWlWuBiZR2+UUGhxPGqQBo4tPYUBF5xVniO+8Lrf
6u3jXCkj3XbrSkYnSAY+U2Fr0wi3ppRypQEt7u33rKXhJXvZb+e/alabc5vPikfPikh2XgEoxPj4
LMsA5hdxQnH7GXw1tjzfewUJXfLgVlW0ZFKdvhx/6IDM1a2t4c6AmWIPeSuRREKVmlF5bbQGLGVP
slzL/VuQW/FY7BnVjVle2uA1iHVEW0DO9GYVUJFUbdxvZ6vSrHWflpNia3kkHnxBzBDUDsUX7nG6
tpnmnqNZdQa0ZEYXG07iu3ubkyPFVDhxJlD0MbI/f/TAABqQivsVyY7RaCqZ8Mc/M05Uv1gl9mPY
SFwZDtT3ODNe2rAk5X9S5JLFatgKyop/AOJQMnFtuTwIasJhYpkn5jt9Ql419lXKWViDy2Qrv13A
3lkqSauBJf29ZRPTkfp3hvnf+RFss+6f66fuJ5vOSdVHqoRg2I7XF8ihaYqfXOwwHUOBNMTXPzbe
ZlgPa/l6Zf5AH/kH/V2rhT4VecBwa9z7YGqGwQtJObOwHOJ9xT1UVWbKh0GqS7TWhB1ntxQ/G3n6
h9z6GTe9T2+mlfaybROnCoJimmpDZJD6I/ycS1apQyQALZvtCg3EWPiB208LmnOxgor5u02Jomco
MKcr5eSH7wHPUoewwReP3dUIuLCBMgRnOq1p1GNADIrZSVWwR57nE1Q4sDTmhYeyQ4xloyeKGSxa
VpySVcQSChet+o9RPkJCSPZ/ohv0cNryiRqlpXpUrQsk5C7iTC9uEjkpoes8LGiiVouvMgm0rmxS
qx3KddTSsKdcrCBECC8xzZDPsbWF4UxzP0PiTQFcpChAESqilzHZOifszTQTQ7VnsNlcDpqc3XQa
fy+VvrByxi/vmwCxET1edI+ZbWA8Hl2RSZ92OiBB6oS5BSkb+kCoUr4T5S6zR7l1L1RbBZo7rd8P
n10SygNNp5OKSne6qCprP1hXB0aTTPElJd6Gxq4WWAnPTy6fjqZ/Qn+U2fhNH/YCpFXUSZF/cYDB
6qoRf98ZCBTuzW3rIxR7Cli0EOo7FIn1op/WE6BjoQsDC6B5fiki9oXjtGicq0u1W4dkidtOT2+a
S3LO7Ctfn6MAZKKPVes0haE0eqKvrq2CkV4MqEIBvcPrEfaw7WA05I6Sq7Qm3bU2P8FqWagYwzoh
GRqGDcp7R+ckMGesLCOtEqSlK5l5udVyk49WMVCme8LCs0YjM6/69ktXCWzBhLeC5GRyM7dB3423
V9Dxlfy8zUKKEeyh3YvkxvovHQGqlXAn65v8OqLXTmpIP0C0mRBMjWbSAqCb3rjipMRtY1B/4oDU
Ew0wXAwJhEFcO1TxaX4mZN2lVGqSkkMZ6YPCV2Jiz02COSlGO+WIgfibedwLY2HATO4bg9hy3qzD
eis0+ZZkdJJR9IlWdsjrjtc1XxzOs83VCxBwtYErmQXLR46upBvh+q2420CVJwcsmPsemiewhKzq
211loe53OTlD4vLcPGQjPzmyPhE76x29w8tUffNhXDW2VQkRrZpg5yZgWrVlWVvhkpUpaxsrR0Tz
VOBMKLXgC/kQQtGabkXJfHtvpTuZBH2ZLMLcBwY6RLvk/myCDMOZhtj+mkYrlu7wEh7LiO/ee4Jj
Md6/nfcInwWyi2qgzcvewntSke2/f2D9igZDOrXx5xd2TOcbk6zzHL/j58ztuczGXjL7egeHMkyo
kIprwNlG9fGa67vYJFzOxXD6Xj+8c7YiNo3b1LsOoqsW3YLduj/tXmUgjOoUVCbo1VYYwoDL+tI3
RYqjgJ2k1Mnt2bCgjC6fmX0Ve5MYmVHwLDobPBIgMt2zoo+md9SSinQBBf5CjJAcMjMBARB33yIl
DZXiDfMFn2tJvNarWVAq8ZUr8ZXwBw3Wmumdu31fqxtt2+5jjGQzcsc81gdqeC2j1PFG5N2VtMdG
gPlGIqv6VR/zjqdUT1IkQqsew6dRd9mXxQJXqeIND8L1IWHZ/tFADE91qS+HuZlQFWeo9cFzmVRd
BmVsLlpJcISi4dBB8d6ady2hduUUqdoLwaJN7/zKqRy7eTeO01DVEcUoOsjAidaVO1M3rR7HhLXR
nkd9zs7GCZgNT+Lp2VhPj3FD0FOLFYGGQcpCSF6KTsXMIQxsDXS8zYdYNCFQQ6PjsLldx8aVIgAS
K5xnJ09oTl0Hqpp0mviSCRSd5qkEa7pplQE3tXDgJf/z1E/1MNJrkrMXzMG6dh9zJp2YP0EEHsBS
j6wm2DOrGnN7OSH4VuWSvmTJhPrhbMhsqUQb/NY1CFAJsHVRBlHOk+yaJDegPRfPTG16YXJho+Md
AOTQizH0elRpOWAat5Lw6uJGzK3WWi7/DGer/Thxfyp/fopS6/PdLDCRp42GjgCYjY8D/EcPVGgX
TkDBMFdxN9IS5vm6elkDJ+mmoFrOmv1tX0XZfo5pxYOEB2s8k21VkW2HV11Qw1rsj0aG13lGQMOx
rWCRHAvTIuq+8P4VjkQLuMCdzH5LG8gQNEk8IytSEshoEACdZrtYWwuyHqkYgrZeGIi8o/kZQaz9
BNfCfF8/ndnprWOOgzCAFrNxdL15b/oRfr/PRbgp8W/VFff6/cex6fUp2BftXBCgA0Tn156EhFp4
cKbmm3q2fdTw9rFwwLZm4QNR6+51qMZSgfXM4lvVgtmbCkfQ8UMYqKGGGVyHaIWR3G+h1yoghlkF
T+t3i1Mcm39e6dJsp6g8+YL3g7+BraK2/XVu6slcwvRPwsok0+ymRvLk+kO5Nu/cDUDpXfCHtfv5
ldqjZODsIQPMS0O9cpupl5SDY/b8CG1zCv6+vxKbaKzC+b7OHWIqml1RoPfuG9H2AUsiv+1GODlR
5dPWMsIPFV3vyqgreRZovR2QKbW5brO8GkGIU+aL7txpnscVKeoFDtEyGAkA4Fi0H9HB0i5lXCJR
QCZfrK/+sXdmVuCE8NxG4i5XRnaS0ikrDxMSFd0WoZRM8jITxLmD38p5X//JFV5UEsGWZmhLA0Om
huWwscjtnAEtvMMoY6J/sIPv+Pqk2+VSb/VSn0KHIrSvsnOtlbgm/ETFb9XxuE4tUKtR0Gh/GtJ3
FdReUUdrVdWE+/yDR/JRZ3ywDqyzwiGfD7h6vXfitvGWE/6r7uABGk1QPYbb5CeQpxpRFgwsk+3W
p5ytrkBEavV193A9DxR43kgf62cVe+5lMK2s8aObA252PELg/UnCNuaQB715fEUIvv8GthWK0lID
FEwlc6UehekykpbAJkerNnUDzFpNqxWypFD6pIBI0xTY9C+TfH5+8ntQ8r8vE8Ov9QzNGB4c9ePt
V4eoX0tcBNCNMJ0hJNyBPgI4zCZNGjlf/eMuQyL7q0tFehEkEQEPA+bW1isEIdb3+L+CmbXZUCT0
e+7hPkl8yaX/gYyE0Sjh6zW91L7Iewityawm6uUhmzoQv8Fr2l2lAgYQn3RAhrQr/dX78YrSvWhM
PPx2PSX/ArfccDpaiwP94sVarzd9DZiEK3yboLrQAbMZPS7saQ32zFfuJntJWbtLHZJYWVZ9KgwA
LrthF3baBxxpJq+IsYLB77cjX29ECKvmUN8g6cBmwjmB6GrRjAfeSjC3Jwqe6ejiywuUy4iwWAZy
ngYgIi1FNk4gHKPSN3Z9VzIpLxSTlLIxD4nc4xpNdP0ESYlklOyK43jOKcsxYE/vnyK7RfzUO8cW
56VBHpOfFrm9W89haXllBMCZEJmZE4HJ1YY77DVrZi+YrXrtc9AfN+6oVMhp7lku/5GGAAJR9Odm
K1vicSoa8vVIriCfdb6VWS8VJs0AdPm8gmLPSW7oIKGCI58GWQJgHg1X1GnsyxaNh75B3dHVFmhH
FiTz0/OxYnvYMp0j6/q8s6euxo6CG5kNn51JShSxeHvwAb/oaj2aFdix3ZdFleKkT4MSxIxQxNCS
636VJqKtX4NfBJiQ5JPfZ6nqnqiiBpH3ywbrFMYiQOnIJ2Xk3D0mNtdA/GsPJKc8BMm//tD0TLp0
u+vdpT0ioK3rPh0rJUX7Uwy4i3Ff9WmKTiF9orylxkJ3JEfJi0XysVtUPrZSyhVZ+Vgwu2rqtbHr
v2ZFJCGsto/Nxoava0tn8GAi39r/Xt2HdVSKNgtnqTIFL1gRG1y1Eh0iJjObcLW3z0mng8o0yP1o
qp93LSCU0AJ6BrI69DR2CbArA3p3ptiwgOkvUWCekHNmkIMdIGW/S57YK69ksIAGFNpG4ZhmX7v9
MIuKp4DDOWp9qlcigLhS13HLompfDO+nVx2BEufu4ueSmdfCetrZPFVSaBOOFIMnspZzR5MNYdoz
+PlF6ko4ZiL0pXGwlQxxg1WVfkrSVEi4boPzjm1NB6g1gpBdZyvPLYZdEDS5fW+pXfSCyGjn0lgM
FmPds8vWjV18TTZGrD7JFTKXgUa0bkJIEpFII+/PyNJkgE2KYTO8G67vMNOq8W/OwURR3VRMweBi
HXOxZ1hDdvrS1e/omME/h/0xgdV3ro8bvobWR17KPqrBvDD6XlYV48q3hLvaeHM4VU65pMX/e2tV
7EmAgxDJ3r3uJ99XFRQCAKpY9oe3XpODlunnkHVMaH5brqJHtdw8F2CF7OhLbcuPDzpYKSbx2COd
3Y96z+dydRPJTl8BywlugLbw9eyKOAv6OWA4U6j+6G8E7b251Q2I4iuhlruBKd5HEZ1wo3KfgNWP
nN5gOtPEYU86KTc01fEVGsR181bAfGmYmJSR/ErNuUfX8a7po0rxbktahZsb9zw61JLN/VnwSxGd
oCPV8yYZxdZAKivUxdcXy4X8BK1EZp210leUB6Lqh4udNarAJDweQlWa0/ROgdRwAA5B8yRnncWN
esU2AblMM8j9+I+PR8c+9a83ntQHfmgSLvXfqE4sFv61jKazhkC1pMCkNFcy2liEnWt1ZUTDUZui
P+bL28L7EUkS5LeqgASeyEozUrWyPsKnfQ+plXS/nLz7A2wGe4+OOd+JT4Qm1JpTVcqQP7EtLwhp
tn9S3onIh/rmQwE06UdfmepYolhB88gW+sKJa0bECA53UK2vaFD+4/pxZDmOLX3yKZSEaNDAAhoU
vbE6QfgVurSiyGJj7bY5bFfD7MKXj3xzM2lnZ5JU2P27C7ui7E+AUHxlLue1QTCd+T85mY/Oc9mj
yxYdIIs8JnfqxK8gZauEnra/S1TuBs+FwfkUHGaMVEtTNxcBX6u1LFVtFUgY9M0W20qXePKCJ3jW
ycnzTPXlOXGXXFFfoKaHK3pmzTZqE/7SAtjv1vP8XAH5g8iFiQY6MD4cNriiA79NDxyFbfeU8G8D
UvYMdCRH7ByoMqrN8/ijztKgomEtNB8UDoR1amXpL/w8ikjUJA7p6u5shuA0P9uqIqPaG6siGFeV
2bZqrcBoZeaV2DoKYEYKg72yTnB0YonQzj8E2uDt896yIp2GCTcdm9dPGKrXO7unbSN4vWIv65aF
x8adqfH2/4mMWjVcL7a4Sai/mYXYvzKN2HN6UqIpIJO5lBdzixK4mIHJPCLf2k8zuCNDSXDn6Tb1
fNjXKGI6cAIq4QT8Z7sh+ss+lcjNhpSnpC7oQNwMzfDjlMvS7de5im3XvtckRNII7qmJvRk3q8sx
47clmzLC3Q4vxlH2Aog+cPDbNRMarY70yDcJ4F00M3Na+q7YtDH0moKMxbKwAxU+gC53X9tthwcH
2PwFULI6l30k5VDbBBz467TaQrF78X9bUG3lPsM3KOPrNdqmrpbppTo7p7cO7GCZiFL/tOuaphZa
tCS5EHGfQLob9sFTTzaavSRYDUsbSyOdFyPu1IoY9kQZllZLfCw2Pa1EkbU0RflAWvrX9O1Cj3DE
aGMo4nmYrFM7fESCNVZqbhg2B/jIwwOni9AFV3ppi6i8LzK0ZwILgplM+X2DGfdkaF/vLoQAUN1N
j56IKB/igXnKBsdpeeOAKBoCXdCA5VslUxIX+RvdV2h1cifg8WhrkTtcmCU+LthgQP6rQOZ6Pjwq
0QbeentNOJMykPaBPIDRbv6Nmpe0vCabIGquXOQ846NLhQ4udHgsk7umKKa/9tTJaqjYzbDuNe94
BpPowC/fSYxsKypKIYkE91C4u2khrdgdwkfc9jW2p4zonS/Dikcoy20O+r8+mPSuKbijEN9K1/xK
yFwGHaNiP4yLOaAXZqUXdMwINirQ0uwRgv+chJmxDVuk5N+21M259f7AOcnpOpA98s27YCZp2Yqs
80cq5laCHudEOn9aLcFAgWNL4t8u2XDs/LwmiTnBFhfH0o7cEayA5FzD5g0/Z813uX91L2nGG6ux
3PP5stmNSOqSPIfYm1vURbPwlhSjb/vidHykNLdi4NYu5IzEJ1sp6uyrxlsx4H2AT/xU/45vS/lO
EjrY3vdGoVkX1+pBBSxB4HLlk2OmXkk0mYkL1W/eTQ+yd2sUWC3wATZ+SNWuXA4tV8r/jLS0L7EB
iJXNt5RN0p+z3xOyzQC3CdZNNczBNM+DNij5PTIgaHixASV6ng/5usGpK5wSPn6teR9rk7ycQbv0
xT2Ie59XcGjJu6h4bJGhUHHCaWFzd5VhqBlTDzXnpMSl1BpGwb2rf7+8SSFHCnHwHXMwODcAu1Tn
UlPRX87gJMFHuxiKzSAaikfomhusn1ay2jXtaBfuM54HVS6RnksXr5OANt97gTaL3YJjlUTxnWQN
pT13Y8Dgaao4eq6RYKmqh8o9ycT5wfljL5ueDPS03S9UUDaNEjZ0GoA68628oKuhN4eBGGyihIP9
MVo7YRzBrJ40L/L8kYMNt4/PJ1IqNYOq6PzzJKpfmWElYdiCNeV9slmomjUHTJrJ+p3pSR8Jdhiq
XKymOENZ48Ft7a83gwvqbXj/Jja3ULFc3LOLsv1zZmFfcAx5nuEvRDZbfDgpdZF8yQJ7AhQbzZDJ
hLshdfC1W1Scea6/NItBOUD/kHpVz8UXArWUbmjg9VQ66Ipy6AvI9fKQhIajh5oE1ld3eyo21tib
A6XrGrE8OccF8kLVzTGSk0kXkyjTyWxqJEVH39SwI82oipwU88wMbiVJmrnUtUfuOZaGW992xvT7
+WTZEt9QYip6OmtKVBqfmpX9QeHzwa+/9CNQM5KIK5Kmc2qL0v+i2H7XsTKx4dsJVB6frsX3iRCB
hzCfIgB86DjMDVm08b+KNxjqBDZt5UPTWLYeRltu0oPTbmUuzjiwfRarlVb9wt4S8Rw/wVT+Tc2I
zVIIX+Rbyf/tYTh5g8mm2kCiN2BwV4VF77csCLnhc3TByueLO/XvC38esX4iLYIMupYD5jhpAZ/k
LSbWOhouihNMDdUeyYaNOA7Y/1t3trTzOnnUdW3T8zb4Y6iocJshW9LWf8F75irt00jFgP+l5E0+
SW8Mjn5Mq+hJQiVKN54KHbebn3XeFqe0TMbuVRR+vVDChyRw4E83amUqaGMztIvoBLSXn8+0j4/j
zLDIMfXT9Oh19NWz2Te6HtwXG6rkEED+62zhbBqQnmpYObj+X/FgzDBcEcU8OveXoxPLEgpmzLY2
3+uTy64IEfN8RIgISmvma956VrH/b4edHRAJkzBwvguTLrQsImh7jJhG94d2Vd/kDZ2leuSrqrG4
xTVkDKsxHy4N6hmZR2uMQabJY6pN44AxXsDttzhm8awvM2DRK/7OXSvCHHMkuksrAbbPaNBVgVsD
8MJT0NSC3uLzU3f2DFbTq/gkXk/L+75MAB0L3g7GtIjAGRhin4t9nTojWZ9BNt4r6AYhj/poGg+0
yQpex3n/e7GT5vSGxaRI+uObzMr63+27WOywCeCwBH0/I2Ir0EzFmscvfEBua6ZauQPFj0lT7k0W
QJnVnL8ApBtrAaig1HZN9QQdRtv+2LjDO29ncbmq4hY/0JMZx9lCRImLbXv7lUpAs4ccCMlPCeaL
j0wD1Ydg19HS+b8xMOUVWhC7J6eFMiP9TeDtA1ZkcGv28ehORFYON7Dl+WtUMgaTiZWPR+iDkdjZ
F9VQSVzrIx0uTGEhKUgFcNyWft7155aK9jn8t3XMMGc4LJOZkCjU2qLOiCskCpNHLO/9bNj420m5
pNnXlTtbBCdb4033bDAMKkpZA6DCFSQH1PuyH7NDQaC5mebKRA1wxX9ooJwbZUAQ52g34UrYDhBz
poSvPQVeOuG0mXnutEMCy5IBx93SkCcLR7IxoLwuALU/UAEnY7QtM3j1d07Bg3ICCnHD3qwhKGLM
CVvEmo6vlMMoSKym422gBovPr8TsHt8YZ6CHUn6OcPywQ5YWdPgv6YdC/JCzYRX7Iz7FwHWoFgWm
dQrXpjBxIM7Ywinvc/vILgaXsHwFdSk3qrGhOvELFZwD/JnG/qXAc/nOEkUmHmN1QNwIf6MQ6tRx
ofJYbgniIkTaCpvivmdM3qyw7CrWV0M+g8cdvmEhLwPgBv8fwW2D0lbmx4JfM5YHcOAdpDX7hZZ+
0JkycIvpMX/+z2Luyxs5mcocDBFS5iLrZgbpv4PLSeFQ2iURJhFHxnmKClRwgLmfluJHP0mDNIIc
WmoZn1UIkfqO2xbc/Hri1LHlvQdvuTSm4NdG3q7V0ujsqTBY14AivUjcHOrY0z4MvrbpWSksjSBV
CNybbfZPzkNC7vElk1UBwIyVeeU1XMfDqQ+RJz85eDvdzEoWLedg5FHU11184p3pc2/d4CnmLG2V
dIEw5sBPJ1yEn3/RkANJlViqK1iSaTu8D+0/8udbFr+vdyQ+YT4QqEfYwa2gYCbvP0n74nFRxb0T
a3uSzd2uADr5Y8WUqFcoCcFhok2O2+3Ujmm5R8JEN1dOihlb9r8tE+0ybQPLhbw0Kb83lA34ZmG1
M6u+RXOOLwa97iuUTMcRPbSkufMyBuAOezw31tG9a7KAunjhB3j2vrvr/xw5Fl3KQme8hQBWy6At
csv0BtWh5oc9lziqhTbEzvSGW/+8iC+OXFlXinOdIyyqsAr+D4YhnCoS+c/h4+05KHbvDm662zK1
SUZZW9ZzCxhILmRL5xXgPHRSQbiEqdIKe0SCNFbmevP8SOaLH6ZqKT8WY2kOG0J+NPfcV7LkgGXk
674ad3T8CSGMrz65FxY8AV9BeyJikB9GbgEvZ1Sc6hNig/E/d8tJr4ckvNpr/KHUDKtfFlWbbcWF
1+gwTaW+cW2XizZjshOsCsmKoaftC+8LU5FMakUjsXjJvtEUgKm0WLegsQdijAZhjfgqCdue4wYd
vwAEK1i6ERixhxHYSO8iEyt9xYxm7pWJjiYTfA+VNzUiKca9YjbwuStHPJsmHPb6qBpH7IC4RN4F
M/4Sd9mbY9WpMxiAmnlOy9DZwJeneBAocDfuKv1mB6hFT93zIb26wzOsCvuh/Mpzhdh6IYalOAo9
Hs3bMZR+wrE1m17IWmE6O+5VnjUbQV4vOLlwqJt0U//isF62d9+iYpmT5n/ATYjDvwR1TNsR0o0c
M6HIirG1KgSQrZxk0TnxMcNP8XRuWsNXimBbBoYj/LLVgQivzmLZ4BfojmO1da3DQdbyXsBxy9zz
XTcFf4N1P5i/sfvpnkckBQ36MLJyOqv+stcXrUay0AwVhL8/6t0zTwAOTj/wVVjZHAgtRV7aii5j
dfq0iiPe2nIU8eJoW/yPogr64vdDQ2/tmDoUF7t6FHy8V2Y1AKJb27j7HgRmpWbUYWkpp5ym8Q/X
OxVRZKAN6xL7YYXxiZOo9vEn/kh08XYTRdXbNdG9gaJ6jalgneTgEGZa6+kl604JJQcEWuxn4OQF
EZDWAcq7OAcaONuOsoE5ck+x90dNJGv8iFDTXi+y7AEp3JlIFF26zxrrEs3aZpFEKIItiPrEAd+h
fggWTQzbQynXpc2Y3imQCP8xGXuXqZOzU/x/CIXad2toZD2XrGgBQMGNSMzBmTD9n3g2LlgAEl8M
UnuW03573Qlhmqxh0ovr/+7ufuHNFKIGEPDm81qB1xYKIZq6NJYEHDZj6XWzhqtoUqw4CzdepCoa
D6R/h3R2cBI7mutwPrlFp9nnINAWLsA/P3q9yDX28HT7EH3cPgykCDzLSSthGPIVnFAZJON/s9tc
OQx/uni/Z2JgcmsT+aCSVAL27v/qsy7Ed/Hb7Yuy856x+9Z6t0UwByw2lWweHeGV3fwlOvZi6/R1
ndYWDGA7jkCCeZLwWaQ7L+OOfcS/JnNwRGwI9l3PDGJelg6jBvmf504BaJqByaePB3dWPlOrPsOy
5tz+8+qYfRH06muml2F5G8/RzlesZbrp4OTYzRi1qOtq0zlm+vwFHCMbCRletJ7yvCMMbLZSh6Dt
XycocRC2o5ZT+86FQyGYFt0Cxh5qKlyHeWtYhBN/44JgHnMovAYJHr3WSgsQtwvxr+3u0M4S6eld
eOEoI0AmCx9mTbcRApxSVYAXnKm5tiWLHQhRlrxxbEbU4RaGY51yGQFyEhzisRgVfheetwEin3aN
brH0xCynhB78us05wFueR45zfXi+zGCZqgH07D5UHItO2/yh/PDeLXS4rPazSpg7JBatOH7oVNWv
ZutUd59oH1fPb+yMPfnSg8pun7hYAklISZBDi3owQKxFf4BBWmjgic/8PHTbb0gQqsZEY+EfIBXu
UE3gNXZoJHQOIwrHuIVcUvw6rOJHPc6iiD1DPMy/sudgTnbdZEJxOcPz/iIgFfk+o5YuiUu004T+
F1yvrODPFMtPbI0xSwKeJBcoUN2Q2nYRq4yuB0auoqWpk1J7M7wJBv3arpiSX4x3Ed0HaVWZu3dH
dK+b7+ZZDMFPwfDYaTFsMUobD7bVX9tDsoRxhtlQIHWG8Nw+64T9JYTyw2lQC9AEkj441Q1zkB4D
j31BF26iMWI7kIrULEd0tHfoqtUSgFRI/QMJsXcQe/2q8b/YP7965+RaOifanyriElXF9k6i4db8
5yogb+oUnM8rOwrvtA2kgE+RuoAmLlCqJ1lgFNLEAru5joMcInE+4aVrk6AhAkb6ffV+EcV6dKaL
GWY2SdvMUd34lI/p5JIPhOiTGo7JsNgZEGzlCYF+L+b6TcKLeYr33L1oj1YJOtV5CVPbO+ctP/In
m8OP08OTbUPiXM/61D5Z8Gt9dtfziY0zQJCGnubyxCrydcqyp2Mrvj3hVJREpREeVfGLmPSOW+2G
GKl6A9ci2OjR4vkkVdtD8L2h23XeuNuTvStel5cvDP/KaYiSO9NOeJiTnoSt2FrMJN1YPk7adnkp
EBSfy1Rk4NkfJqlXx/LrnMX9AY0bUh1WwlKUGVlqV5UCV/yXREmVbP/lHXW3MW2so//KvdOU0t0r
ro0q2lKWTOPjVLJGb9vx5L41fm1DT9zicS32G5jBbOwEpsUfLccqiCRF+RFEWn3scgkBaQdhLmm3
9wNRmDCcx6yxoUq/YFKjWBLWA9JAU956dI6qW75xKsZOUmXy+/d9s5ib5MPkMX7lyM83AF1PCLfZ
vNUJGRnFfdZX6zO08Vr7dnZgD/EJ5sh5uOun0EG+vYerrAujaXpewfx+m63TUaM9t+M79NeV7eOF
VgwvLFLsbklHBOuy/MTae0tGeduLjARX1J+1vmS9WEZFmtTDe91VQEe6DJ7xdbYeiplWLHeS4L8c
EExiT7ACJ1dxZ9WDjMNsTiVgBxEmXg7xoFxiSEA63e2XbNJNzp3vIiB8VKadRQuaDvLnCxn3DQ0o
ZViiBaGAvtyHbqEKttl6bt9RpqE1af8vCF/6uiB8kAxaWLWrWbtXUZGLoxF9jYKLa34oX1OEKJ2R
0zF8dM98AMrF2fB2RP5d7mlQzqXV3UlUbN0QVHSYOJHliwk4JrBAmJxyLQnSTN1PXd01oI+iKIRu
cTHBOQN8pGeG69LfvAzHXBLiJ9hTOgbKtFsnE+SaKcShvp59ZHSLVo7S6L5FckfrI7juGJf8/kN7
vFm7os4zs5acolSbpzvem6pnSDIPnQf3c2nky7hjM+Zw/YpV5sCv5UB4wxjB3EZW6DBJ7zddpxVC
2XAJmoC8O264/Ff9ScTglS95rKQsL8caEy8BejoM09Up9nQzwc/42BFvIuoFanf3xj7KmmxwOTH7
6wzYorsYJ+oTrg7Z1cdRJdB81/t5GFnXnWQrU31tTD4ldOlXhfeEmYMOB8dWDQru2xl87KM40AEd
S49i0+YLIwGu5C9/ZfZ1RV+AEKGwjv8uJhK5IXssKUEdIdtE3q+7v7n/8nVEbcJy1PcEArSeVBke
Gv6mZ8bG/xuiJU5cU1+sYRM3oEBBgruR60PZbYdIdp575szkZ8fyQcVG9Bx+OU2OONd8rHqkpeVX
mAqTJT20m5gxQDImKp1r5SLoUtGKzcuHvN/5CPhKRdpaOUQlJh8SxMTx2wlNJn/oVULQ8avh8QsG
naU43z1EnDNdPBTEYDgEj4SYUSZ7aOa9EfCyJW2b01rUyXlYkKikrUA/so1ei2tvAuLX19dZUT11
OKNUvJ5NSoDItrhqHW08cvPHSjP2zSkuNkMlzl0UYQdt6LyUdFPlHeN4DcgHTwnFQ8SR5B4cCW8c
awG81hstIKm47mKkc8iRggJUW2lvvAcHxOV4rqjsWGDFAdLB8bU/DTHffS1HsY7Q+vij8AJKxPnH
+ZofgzvI+6R9FQA+VAlE0Lhhtzdmu1s0jV6JX26C3JrhWpFQyiGSbPsjsCcCAnpkxRmsuQk/rDYg
v15WWwjs+zuwl++AaKu1LagSO/tHrfLTJqUddQlA6OUSAktQHPhko7jFnx3sbHcWhwWDZsm/r/T3
equtzoJ0UcV02k1mJIPGLWrceF0Yd6bqNM0e5YjgoX7xCFF2gH84Z8Ahwepsw+1V8wa5YKbr690Q
zIVJtYPu+WVmhvpbcJ1UXH83H5L2ToSl/eYCyiin+kd7nu63azmRmhkDJnmTughY1PP6hqPWV5VY
fILNK8Tfe6aihjiiqemu95ftrVhJ/U/Y4YIpFGash9pZwC0EKrE4hapqJpVKZVgW6s/Cpus8Nxec
11wqrTanru2LjzCRpiursx7xMTtIO8SNO15ClmOt5P6UqEOz9rcujs8RAPe0lVl/+HleELMT6XEy
FNTPNx7zoLPB1TIi8Sa9H4r0HFlFI/mKuQYP9Ezrdq9kTmSDZGEt8GjfPR92NwJA08HA7CUS5OGU
Ct++b2xQvm6P7X7b9ti0IUGBIrwGMkgccScFkrPItRZLJ7iEWnxXoqcf0ewbCL0+qcY/ffmfPU9I
tPbJuArweRF49SMuY2skZtceFh0svvZ6dlqyhGITZI0Jj52K0c3gRZjxjRKaUoYi2PMI4+BlIxf4
GzDeb9oxvPFOMWhkAwSqCvETNH8W3iFcGO7/feQ8fOH8v12HOT9pyCpZw3OmRUTxGdd+SCRxcaWW
Ua/7TVN+WWKHSZxcNYhCIGGLrnEs1enGz91RLeWush7yraZzqr8msP40DvbE4tDT6c0oWsZp/swZ
eOFcTZyQhYbrV8vDas/NUTQuJEywxOcOzE5Zv4CLOtbuReh6dVnnq6KTJEYQMeYrnXxjGqG8HVLj
iO/K90g3GuuJUeZ41KzuL+rnzDGCXUC8KjAFeLBHtnPzEqkrne4OpSspXGBHlCvusO1k3EAuv9xr
SgKR58uTuYJavKtO0YpagjFp/KIA3oaLgKj2xJBXnhxECIetV249/trna2uhE1fcYTwUxkUxHxq+
RxEolazeVaRKWet9BQl9yuQsug7NGgRSBmB57RqMstFKIvj78vruB3cgwfdNpvoe4PPtOV4Rp4LI
fKvuhN/tc0Q7MJB9MHj39gmi3o4Diu5kv35OCi1T/MsOfH2XtR/RqZxodtw2QdrjHC04vWIatVH6
Mc0lAJcHRqMy9cK6HN4MJL5oBz5uZWPdWbvdhRJ+bsPjd4V6H5O99xfQZQJM5fCjl0FiAXOxC+Qc
SRteMdQMIMDJfBpA994gNVSSdgvBNYsigQZalRRMQ25/bTUfSREiSggS01ttCZ6Woper4Covc+RS
WYlxEODUEk9QW6CPG9TFPoDMXNxC4bHZWBBKTqdkV+8hQtHoJQSljxtkCUsXF0iq6yzYbFvoFndy
svPtYMnyZqqmM4GjQ5gAwcz5zM2kSGRudH6RblozN0b0zHEq1ZVlJfYQZuxJ17RCKnPP95VymqjF
ttR1OzkCGnCtleDiYxYm+eDkRobohR2hW61+wgqc04xAHynwl/MiwnPpNLtk9kTvdS4Tmr4ODoa/
xwMVill5Jc9+htEVs14sTLGAn+6jH4FxStWbSJSSf3QyxJEDc/O/uP/QDwjhn70mdWLCyHHkucYo
1aPtsv1bqXQVfuFYFDEXmRk+STW4m6quhtpIYYOLJxmmUCQEl4vpVfuq5iyrflJFTd9cgGZVyHTn
K/VCkRYPR/JmWjvBiYbnQAzlV0Ey4NrJrPzAUHSagBNC7EZEkLYXefy29HNRvcOlsQR+d7Ud635i
s0KPFxE2RjnBQt9zdWu5FST3HS4CIm/pMlDp+EVp8ZxUMgFUi1D5OyifPdkZDDWv+Bpq1Sl+cRr/
LXPcWBiAuNla73uNwnpGmbZkumNRvFCk9R1qSsxWyaaRdETaQ2ncw9ZYfQvmUyn9PTmux7574SFG
p93AJ+5TqBP20/vWClycMgcSIqQxMsx6LWXWKIvcso50pfdTYb/4b4fd3nnsWd65CpAx/nRbQEkC
MtOEm7SSlJd/JWECSW1ujXaB4YFRYALD4Q7S8cER+w5reUMuIhO5trHIPBrZTLebuCZCVGY/69PE
kzwZDYHqrWxaQajRjV8HCUwBygBt2Vg3eBlTQoiViZCvt0AHuC4rPnRcOWGSJrlecYCrCYW8TiQp
u2jLD57OXlntlWKTJdMX9HfU6OTAtzqY9UJOahB9gA2Zqm0lJnZrg2DRjZA8D96VMMnpoLhugLXH
sQAfg31UcQIYOa3rbASsN8qKwz3mkDqwQUPBpO3400LdrGbvgzRg/5Ekp8e4/5+ikGg+lyJAowYd
ySHL5T8Oa81PAKCxVhhFhO1K7UMVOig1ahrxZSGDnu46G93v2mLJS577Min9A6t5vUFPQk7cbtec
Qe+sczxZtBJ/TFdn/djOF/W3njqFQgx1ftNRYGfl8u3Ls5sxtV80cmuW509tkEXbFo89JLWVAdcQ
8wNsid73DU9Vza6hq4YVXEZdbcQDLQ43mpEsSKLvJifh4e+0/NwS3ktlCz8ze+jI0/344PlUCdTf
mRCGOmCY6SstJT2GPHemIRf3r8f+A796svizHqB4PpenPjySvgnhUQGU0ZaABHwZQSNi5HZX2E0u
Z9mj5RDge/CGRiBFn8Ukg8s6EWHRz9EfL+FCXw4JN00SNkUOPG2kyymYzd9uHbbDF2qOJOYZSflg
Nr69HhR5lQtkvT9kgrb/3HKwsgeADyfUFKQMDjD3FkIRqLjGLdzo5m8f1FeaNP3/EkxI9cFknYve
UqJzdHCVnbp+XqJHr3QGQpC7d7PCzoREgU2uZp+8J9bzxt1afgigM+X48CSkWkAOl/3YBd87jeJk
LZnvP39Zc8mmSc3GH393WnP1OhBZob7h5SUxGt3eYh2W1YKoG16xr3+5DzoCiB2QwRccQwgo2+Qe
8BBXKXSeDdniStUuecPv9Na1eSzdepsWUMkdkeQEceDg4Sapm6B7GtEFJnkrk8Un2mTC5dFTSd71
BhtB3ONADxn/f2b4LrV1HroPtM0CSURA93TfsIk/jb3BUh/O68s4mH4G+UN1o65sNNMDsCcrZVah
l1nODQ5MLGLOnAJ0rMprTcRWc1fIa23cpF1bWG+P2Ov3dgRxEkJsDKDktM9A7NDQRD++WqoWwJz4
LfgrkhHH2PMWIDa/xdwsUkEMHwoWoVoGgKexM8izknrOU8yZhl+AxLHc4WG360ai5iUSeNDHqxkg
H6WV66UVP2DXqXLTD7BKzzrU4aBHBgR00sbTdWTedHeysRFl6w9ScueYPmGZHEzBrAtnCK+u2ewh
koMl8RXhg+UeMvuLhoXRQqhuA8g5wzBcZBHTJvfgk/VOk5i/hMJTh5kvpARrdEBxKtZMgFUGgOV+
YFclhnNalNGUGz8HY4r80WNe2iEQhh7O9PyVRmcMhRfMGQSI1BvN5S0SunpciIRnjKWkzNIKbctf
jnPs7ZlQdfhdXWPU4pkOmy/aFRYfpX7ul86KYMj20CgwZYJHmKJQc2q2epswbdSL17a/DbJQqvAy
V6YIhy435feaqFwUOwK+5pavT0rJ9ePgxnYQbXV2ffXVIJydlvyTjyFvYSq4XDW4bWiYwVDxPdPS
ldanF5PC8QpyEmXlP1EkdDgp19sxOeHN9Oooe3YNmvCI7Shts6+IP1KYA2kr7NUPfsektl5UoBzj
002s4tnFH+f5/aev+Ag0pVLy/Vra6dvHurMNVHaQ5UsTxjHZ+QegRhRVO2cdlN/+Ksvn5dA6Rz2L
vEtV4S3VZDhNJbvurlm1dOY7lc1DP1se+zRRkaZPr+50wbZM2yXhZnA12ahK/YdtmgcJZFap+10j
yz3IqRhA1WWOKmqFjizKmbHUkURe6ReSj11aUr6Tn3qKUxB1x4QTdZ2QmO46wW2nsUiKK5zXWr09
RsAYHoULAqPKarncl3hg1chGUwx+UzbAK50bGJPYIS6BLzsBlqR2eTFrGyW3XiI9M2Ep07OpZzSv
ZwfJTaOQH+eGBwvnzRnuhS+FsrRRf+iSyQDSK7A2MgpTkVb3vFHZB7c4Jd7+14/3hAMXVCweJLkx
MsmcUvQC5QMmAXA32woZjYaPsqiaxkZ9ZOYKJOovtzWPgfYzaDWWihDYYmD96GnDLY8cZGVPFPPP
ch2xzH2go6moPmll11PUo228iGVlFMC8fLvtQJvaz8bmaJ9n4PCkzDXI0327KOSAziRZcByPUR8K
nEyYiyDJ7f4eNlBfNScYgt9I2HbqfMzPMch00swpI1bX/IoDqG95dsEB4o3IdDCM5R7zDhiP8uWw
gvu9Ih5yQt6YUUObWNEj5IMtt3BiJUpH8BFs+G2ywadsRRYk9Fafz0pAgNTHyzR9xu4Bkp7yuIfr
4E8r3n8QAo1MwXkYXfrjjSY6dOUMqgxU1yhf9O4Xpw/tpZ1PJIrNj73zq/q61q0sv+WHb++xUved
z4O4VuIwLs+8ylhxE2shcMO8XfieGLIwjUQ4NZf/bxNVQpEKe3P1p19anbKr27maygiGQJ8S/RY+
HXS7WcfrKDcdsm7cZ6YS16Zwa15+tJ+CBZyQH9GLrx6d9ERlVL/sfkg3W1p/OsgUEqBco5DwCI8Y
0BhsSEChXA8iVAmDJVrkxpC07UAcNmbjSY2HA3quhkFm6dOSvlHB/3LwnCLe//brD56BJANTovML
u6vqUFDXGzrwDV1YPW0abnFAgNSVjkjW+KLUVB/lZ5u5hUToZzJ9zYFPIe99nLmyhm6rAj5fXa5j
BOx/JJv4qmdng+3h3aXYtNyGEuhK9KnnunUrJbCQ84RCPRHeFATvGPVOKIg7+Xe9tbhlEvvuL5Wl
d2RRqRz5HA4JZWB5IzcDseRQ/WVXcZUgouyCVb4sAYtwW5mcT1hD49L80mLHMRIz1bhELhycjZ3u
nCYfopBdwzmnn2A98zGo8XYMhmFn4kyO32rFX4FiG8QoVhrvV/GE5WztCEhU8IatOf1UE3YD3KMp
HK/SQ/4EGIK8bG6DpNQ/nBtDDD1xyNxjRBhdQzdBSKPP3CrEfHiqBVOAAdyR9T+uakc+AjLQALfu
2FPMPTsSHN5r0tP9cpGPnAh/m5hU4Uxeuoh1rm5vyVt9AfmXUJyB5eXWs9RpsngSIejHaKbw4vtJ
6xbYhe/N4XnCkxVIyKBu+nZiH7Tk7qjicIAv9zHamd5QlqRt1X1VNSdg/UaMQUdQNsHwbMdQzTTE
KAjUZoq///sXYSqxakXqi5F8CauUK0sWZQxbB/FY8nI5NlSZUO8yRreFla2618r8UbD/vITvI9mI
3RxRCjIO4BZJ+OUiKkG1MvIVyHWnT2TQnDFUyFVADXLIDPLkRZG2R0NY8bndq0AQ/Ds+jzgIu2Sp
AihLHzRInNb4MbN1d8Qjr4DjGRCq4awgVTBGfp34qN720x3BHdQSuDCZ6eluLjdV4LLwpl9XPtdZ
WZzXWP7DBIGCoSrmu1/5wZTu7TGE1OOBoDDllvZ7IZc87bKL4PPjml0hFK0RSDSU1YyyC9VEk9xr
yoS2m+OVzXQTl032d9mom9cnQA95XQx0R1Abv30C47MpOjOHenSlvyrKuD7XpONnT4pD5mdbFasN
OTp9CEdbDFrOiQnvgnQnATquKlJ7S9r7iHfYj4gRU4gmxSPPjZFNLPdiw3fZc4hrIgBp2fvivs5i
7AEMR+6f2UMhrF1P3MgOIycbk3v2fVjnyx6GWvuTW0dV2tdy/j+9wfGwiTleIgc3LALkdaky0ljC
xzftt+/OrjYw2Enx6ViocktHpXiCG/MfaPAhnDWyTjj4TiYkTZUuU5zfec3r4RjcPaweWjnjM42D
lUsrZjZqWS6ZTYgPYm0kZgGYDVDxhDZXzJgLwNrk2YN7P344CrgV7cnTwKTdYh3gJBkKWF6zAYKu
1j04L66KqRPR7ShBx+4dlrwD2xp+rOPJDbp/5sb0UYNSqtuYtIN032Rh+CCYrNx6dxn+m0Tp76iT
dwu7GiYwYVDf+muH89hZ7V3hQCq9uH/+wN7eTSzJKYaEX3S8qEpSqphAtixrdupTOS1ipyIFhDh6
UWsMskgqF7RT3aLUVBGPq9H1usg/hhJijLX3zsW8oGMFHxFIJdg8hEBSe8io+N6e4cXynMBfdBjz
M/SUnSQYQkIXiw8UblihaU8wiJX94cRbFNb8SxFp6/fJquYR2U2+6PyOoFVIQjR2ADe/4EXbmpfn
CkgjxPvmIYAaaqR1J4W6U9L19fj89LxDK2BtUutbiNrD1lwZl3jZi4Kyv5nAPFTztxQHwK8PmYme
Ff0ma9a4+km6TGi3kWA7qdDnjFqdsqA2w+vjrkdKmaJ4Un81Rnf7fsLM4Y9cfxaP+80xixS46BP2
Ki/nZTrUl3WficuIq3+mkcsnxWsHBK021typdptCzJTZlYHCMVFzcGWJI869ohzaKJVaWdsM6mEn
iyqKKEvM2LPZDE8hSCnoYrFsrKN8lrtZdaIv7Z4jRk0gwrlevdGC3Y7az8mbAPj3ciASX6902cr1
zPP2C6JfJNBlKcIGu6vZWIoauu1lOnMxlX3uNv0OJII1r2lubTM5rxQ1U/vwbR0vZKZ5s2XxyBuJ
AOJjoAFZ199mpPwqY9NTSifKJIRsEDbiDUAXfnwv9t61ivvYMo6rCjCpeCmjqr9GXQwHfVEL60lC
AdXNG5hPxAghLNVE4JQIHl9408/040xE30rU1zD+0f66Q+kgS0LMabg0uvuEB8CUcFDYe/lOVrhJ
GcK8B4VcDpUjyJxE5jPP2m0xVFCsdRdJYSKyxt2+nSQ3HjdMJpeNLiw60zLN3AgQIljquscMq7e8
sz0EzC5tGLm076+HT4TnC8sytMS8stJcU03EaA9Ax9EEPeAc6Cmym1YoyzNpQvSI6waozaboJ4mD
Y4+sv3i0OLPfBMI9J0BEuTZyGss9zQ9RIj7zYI0Qv/nVDQ6JLueRHulNcFKSAzT5KNOtJHXGu6u1
IDvz28MntJDSELRIvHBtcelH33ydUEXh8EixF2jN0BDEUW0pOqvpuLqC5xiHqrhAds9iCbJCm+YX
6T5Uy+6zPplzWdwq9WSXa4q7HOist8mb5pLs4ydzhon/SYF0IiGTdgakXwO7CK5KOG4RZSgXYbXE
yERJWMZ8OE4JTRqzQqEdXW8qOclAi11RTlSBRa6BbSZuOGNKBVENgU1UA3ELZXIehp3Xs/57gnXl
mIMe6JVXIZGfue9CWfvwD7wh3ZZnhHJz8Kd0zLhZRaOxSg0kk9QasukYgxwGslrRpFhFCG/nY6fw
TQx/7Tuq6CtrdwHBw/7+7Y6jkiv2/NoF7fIwLXn2Zvs1/hMeNm42sA8hNaaQaUU0NMnni4BYatqW
No4tGXqU1wzv55zPbftaBoSg1P8U2Dv8F+pR3C4vu+GAPXVbM2Hvxb5n503/epN+qwQns0mJOEC6
e7BPv5X/O601CjfHu+VDaxZ/1fxqbp2MP7WsFK+azppYpD7CcCBqu7oSVHhQQmAqndXMH0tFAbkf
70MyNAMRV12U/wWz0wn+moB//63cLFuYIvqCRXKbeXlWPG6nD4Uk0HRZpihNtT4LQtk+S8XiW7zk
y6D4O5XYYgzRi84+wl9lUGRwH1vgFEBuerxv0uc0jYvHsqDu1eaqPAw5eq/4+9KH3nmMq1rdc5di
7z014xA52hh58DueEiX2l3krBoVXySLWLfjmuSVsa5RxH+HNiid351X9slIitE8Xl4EMxnKSoUIq
F90lwqio/0NSql/D3m6P9YoItTgpQ6/ip+/uPlQ16D/3LMtP6r8HT29oK4laPakJOHajqS0U5+is
/3xcntxvKY4BvBOcTCSmGZ+20NbyWdOD82TiT3PxFTtzHTz0jqNe6nJ8ldQvNx9R/4CXMce+nC0V
zi3h2tfSaono/h1s3X2OYD62dxeP9XPCoZIISvF2afVOg5lN2sHEUNqiJU73QF6PWlgaH+YBasC2
RjIqxY+kkrScHs+ICdTcY/DZwY1PZTY3cuktEXbUu1HZPtDLzrt0PENwofePxocYbZwouaoQ4awS
D6y6PCWGMoECbS+qsvRHSCk9x4h3jsqP4rnFumzGhWDPcmbrOKAzNKFkH6M/1yeO1MbsFJ5T29Aw
RlplYsVFnFSOATNI5+re0fVSf1Y8s7DjrvskojpewWAn8KjYLeKnY5QJT3eWniF+ihmbjHjM5LN/
cQGX6m5tdY8otQ1dmPmRQETRccMNvGnGTx/UfywSIInkQy6E+A7HcJ09UO55zBscMW45wxbeweaB
4hRx0NnSmmSJrzCV7P8dOhtO9kd6Pujcd16MYR4EvhgejxJYrLTOAJJE9cxRAsPMMFNB+AeSBKTq
uFc7Bii6IhwjFqt/n9PbU7DhesXgHKtDTl5OFfPYSaMVCuRnl88nTnoIS/oc3DdAEL6JLpbHs8cL
CWrlA8c2YHU/wImH6iI63vqEWjVIm/gFjAWiiGgEl/14PPnNV8gn6gLCKDdSlfIWQKpunoAaHn5s
BPA3Ef9dnf6VrJoSDJL/u5IYMpSTsi/DV3WbyFAUI2UtEdiDfHDoD9bMcR9YI67Cav8WC2PGxdUz
guC4Me0iIAMh14F9no4WHuuxvSxcvV2j5hLQ31CS6xKUOezJAS7cE3hnWdJATP58XCCvX1s48n/D
N7VvCgSZCyq3RUwDOhKJKh/7PKAiFUIfjLDqURZQkRii2JSGYMtA9s2afFhR7kyO/dfy/jqOzTSc
AFQPfrrDSDmdbjYE3EpERfcciHKdoupPS5zRX88jzK8tlhPW8UEWB4Eb6PX82p9btNE0NOF5EobE
vTE0t/mUTKIXmowKSt8CjAb8UzohwHaB6qAgS13gaDC3JhpWk4IumRAC6W499XyGzjyHwYHTcB7B
x0OsilHns+0eSc1IrGhtyE96a9DMPomqdeMVgqRu+5R2UAX/JQ/JCrGEUbXuZbA+HD067fkSe9QK
+VtgbkrRS9pTzLqrS6Qy5iCM5DACK/vSOzvBeEkAtt10N6havsUbNkrolQzhBtVhfCCGXZg4j+eN
K7DRYWoW4mmdWO/Q8JMcjVyJSJ5XP00TGdry7TTHmYfDrGNynqbv01kS+LHfawgi7nGJFzBoxvvK
P/jsEcpvFyIJKDnG657eU/sD6O54K5JDVF+xkqrVfwv+vBLcYomHPEgF5tEOPTtdJewwQm6qYwC5
mOZ+f1cDnknsfK2hJUNCXZc4OHs6xm7pH+6altE5PFqBWbXrRDVl8NcGPgBHaAedi3FCsrIEAbUL
VtWBHODgNZoinps+lJQF6xJDSV9HQ3T2ClWlnM0xR8GuhVdH1tak0OYQ+w3PGFZZQoIr5dPQUT5N
SRZg79yER67I2sb9Y32At4d+oHNFnlUcRaUP4P+BK9getozbiq+8YKKXd2RZrwTj+yQIBETKIZYj
fpaSr956ZlJd+0Do6XPVI1rSM2ZdE+qpDg7LmkncVOwEplZbyWYBne1LvEirV3welJk+A7gUBEES
LBNkjQrWe4ZZiuNlWkda28TNBIpGFzvyXyXqxzFZ84ubuEXVna3C6ySKs3BMyeSrScdtGhqjz+DS
mzkboYFmBgrApboa0wfdLOZiZNxXo53Si1cZW+LNy1PggFcDbmdjSxW5Y/IdpPSH0nRM/IU4YjJv
q9A3CXTPWxEL4UX+sC285dyPCpsIcirRh8qii3/uzHdIrmc4zTKajX37VF4swsQtfX14RgYEFp5W
QVAuX1w/C6hQfNzveSbzNlNYDQUdioChlblW7R5tZNtwNLeWcP6iII6xecgohnMN9TAAXCyWbH4y
KmdmcMvqrEc6awtBNbVEO01R7qDZfOEzFqmpKX1yW8LDCBEQel6BF8Q9LglDh5Vp/IYm5busjWMu
Jx/1ESl6k5uxZnxQGO4VZzSqunOzFmbpIO01B/eGiygsAw8C1OFRQ5BxrTKAumTjrM8XBO6P+YSw
2DuMJu0xJZFVr8Vqt87ip1gXAzJd92SLOk+T1Kciwck3ZvU4XGe/yBtQolYZDjlKdjubrfkJzqKu
GilVHc6nAgUDNsDiToEE53IswXH7zG9WYsRpO8NgsS4j8cXme8Kf4/cUdBMhLA9BJwFf90svhoBH
rE1GmKDKdKytFP2m1eCsSneSnBiS/Uj5d6DAUwOlCv0/+MBm4dfMH6P0fMXAtAlQ3XDiqya23ssE
fLAaLI1NmDEGhFKeXDPSlPzy/WfPPjzGjdy7yMCzPSw6cZ+tiA9NXtuMchgDPQxb3jkLSTcbcvWV
c32K93VHbhH4hvhM8LkLDcBsRww/WsXYb6MdlPZ7ImgSflVgfxCjFBNZViPfL1kX3uxLFtczczER
hTKIjsIxkVYiiASS+C34OZ46UqhR1PHYdTwVzlYwGy9Elc2aU7fwZyyz0emfMlc0YOVv6ExTd8tB
5A64FFcifxqU2tuq5icy0YcjPugHPp2vvfPX1Qn+lR509oC1O0lMcct9+gjUn92sHQ6ZsFkZiajP
E1aBC44yfI4wHvlNCJNE/JHwaWckhxAwkAwDBrLz42KwQFv9tNpjVtT08ZVgyg5Hs6lwCpUgEbOB
FQVXCMKbZukTz4l4aYYKPY9S8U1ChzkxsdeONRECLKHXIDyIXcnwTqBEcIW3o5e3rz6AzOqpCwl9
gNJ+5Ikr4AeZPFeKz59NV3EIlUnL4cXsakM8G4MwrIYS4BEey2qcgp59raLZ9Wv3C4Z+uNm07M4i
VMUEovxY8AiNRgY3bmBYWejPasiCUvg48bUIFUjrKfA9G3ROfIoq/cUpKxSrEs4m8xw71Mp7LwXM
Wk6Secoc1ulw6OU+LvdQk0UflIMrwhszOtMGph5s0HaV/Xgh/JQcGlLLgnAg3okJ0UvcmoAtKW+t
iMQLTG17+21hMl70GpC3d8yJ8hiUEphFURploHALAL7M72oIa6BHM/5FdXYtij/qY/TZlmAfhCbN
5CyJLEegE5ePM/SzSbjOyMRxqh3mMNZ9Hlcfi47R0GQZM7RnAjkR15r1hkm6KiPgJTvyu30CQRoZ
P1VT7QBZmPvmLIgO0FlK+J33t0uBNBrOVQzOdjZLqnTQTmGs5GQlsfYqv6dnrbj9VuFhOIkj1S+u
T5kZy+VzMHUdb2YAbhkkgQOeSm6tKwi6oDpIvIN/tJ0vQzBCk06hHZFv3dX/Unuc+M12QCJzD2yu
YTR7AYj+1yb11y909glijLK2K/G0zufPApyix4pbKXu2WKX/cgtAWJ/7hY1nm117+62AT9S9QDKQ
aCyKiPMEo25kS7aHUTdWHAprAu0PlNkI7eemwcRTsMtcsSfSCmHj0/j5jN0Z5sdTua/Rq99/qaog
DxK4nhnqX69mNk9QFAjqx7CgnxA4z+PLMIkWFC/U8u0xPjBKakTEvwScQwD59RzFeGV8nEu8sWd7
TWXQv4jEM08mqcsnzqyoUOp/z3vMbRXuvf8cNqjyvAArhy/ONW9pb01zQS5fVrz86wWjgHoLUSHu
Y1Razq6w/lX/s5omFfsojc+tj6JursCh3513H7uEDjr4S40yfS3E45e5wJNs6BkCvbzq5POD0ZPo
xQzuVKaz8zcg/jDa4HO0LypKO//wECuzhLqRJJRBYNxdhJERG+hGnd4aQmtUk8dQVq3v7g3EzDMV
dm0K5AZFSz0aUhwLtqalmAgBZkYurSTF1wrVI1K+W4+JXSbmiXUJZUugotZEanJq22VnHbuPaZhO
ndMxmsXolV3wnGB8nCwV2txCaZnPKo7gBQtdL93iVVXet3nmvcfsIN2Ul+I7yQ2btK84PIpAq3MS
OCG7OvFQw/WgZOE0+OoaYiSDSqEoEo8NSC1mLJUexkm5EjSGe2b3jNSiyXAcG+5YZpH+xsWNFha5
jSl86V6BqL9LVfUcwwGclWdXOMukL3lF1quUJBxj/ePfM/yjk/v9JWzP/TgBI55mkJ7k9MNLjgOG
xSYWiDBGDrSboZg1Y6UEhnJZFpgzIrXrSqP62mBehjsIgfsuo2FTxKECzCw6peVRTC+9nNxfglcu
qcFqHM1naf1h+yBY/5qBU3m6ToEB5p4J+eI/hze6rsIaZQRykqfuF8Dj3cs1R4nX+4/TgRtyiyUb
LVoIfn8mEiDthLBTcmQebgdAZ5ZKmcRL08NHI3mEdo9XxJaVyYGnPuRFgpWsk/awObMiuVHIkq5t
lnkE13Hyit2uwX0yzV6S6YBZT6KOWdyqECxIvwa3iFjVg43ZGlIxrG4uGgCqn2dkbZU/WOHJfpm+
fLW9y3chHZCSP0auq3zfHreUxatuvnHPsQGT657K6/S4YFc5VqQJKZez4CRMaFKcB7dHuam8MUR8
oXLy5jsGHIpGxjwwOUgdKGbOtD2gD+qak+4iINuMDUSy6DP2pX9ziXp+iu9USxWy4wkwCjjzAGAp
hadcpqHKTxEsFIW/bWssHkN++v7QiKDmHYUF1pN9lv6kOMQukSOpKYGvQltvC6UwmnSnj1TSjDMR
BFfWbEhuJ/0Yxk2Xyju4vyNAlPAVwUFyAvJcCrSu5DpdgG7HRHEoxCoRnjiMZaPtwj6pibgsbCH3
883wk1UyTm1z2b6e2AY1q+6V2AZUyQTNykT3VzHumptzXTLLIuMy8FtMAV+yod6/OzfReAmRyzPW
AD4KnpRQK2U0ati0zs0QIvk8PHa7tCn/xFcgHyPzm3h+6EygKRoUl+eKXBN4Kc+TMkckI89GA/78
lV5ENBk0zbYBxTfS4nHm++ks02O3Twf97944rnPH4EraY1nRxG9vdz/Terj/RavImgb/dwKve75R
k/4ZRpMwpMyYqWG2ChQpd+X2VkUTUCLuoeaPDeIxn4hgHKxnfTeFJ5Q7Tpmp62Z+3qhHq3G2JHuk
3lwDArtR6AYJTGHiji+yRc1Ir/g58+k6vjl7a/2tNQuwXZ11wsJuolFu7WgJ2hAeatNoD1lFu1dT
Mxuw68QPW9r39TV6TMuEQ/eCHpXqRUyJj9x8qFcQ2NgSf3qZSA/5gJ3QA6Mphrmd1GJDQBRjX5rd
ShpJGwA137Ma19/LGbSlIJ7A5AX5IVwSytHy5MOm573+nYw9kXsDc/NNhsiX1Qsw+ReSW1XOldhw
LkRVeW2vnxagtLyLPzbt3XhDtB9LbJReTh2EHqrTc6LS305pYgV5OdmEN5tT/93OIf/SVxZ46vqM
tyBFeeqIL2Wd8SGwNG/mMf3VHONtIcvGN3SnBjb7hZgnNlKwITF2VfUKILlS+PNemHXQ5Y8RqR/2
hRHK1mA+fDlCoc63HTLFm63jAOTd8b/1m7uTaEHsEbDB9cYMjtclhb8bUZQFKACa5JPVaR9y8men
138uxt/r2hH83JHmi4+SMhbmXwvDGIg92UaWFpBCvx84aajK4XL2KG8q1WBUuFoAFS+jkZ2tSWgF
eLPgR5dhOVHXT3Hp1yf9RsK1C5UrgwEPP+oewviJtVyf12gP7JZUXQj5kRYJc/xRLzkltbM0L5W1
9jkYFRGNCvRKkx+1kaqjDL0YA5ytyB7nWZ1zuhJg1U3MRkTSf5Pewbv0e9TrbVyshyHeUoJ3zts8
WNl8u6Bk/sipxnain1VFGuZGUzp/eQ+SBshUAP5ucYBuBZRor561La+EHj8xRPcnrOAaIjYZayRN
wwAiEOp37LOWyTAwoIwpKLcXm5JHUGj0ieVWz4A7RldJIlZ0VTtuMUsDqpjLhoq8Emtybw+KjVRb
O8Ts44QcjV+wswIEoW4hPomDj+wv1Ji1E3hPuItbB7tynT6EGZm+2i5U7nsg1+bfS2i+gp7wcUBy
EiD4+2Athh94jpLjIdaSCxyHPoUpw2Eh9rzFSUkAY4kgkljAShzE52dcWMysrSWwQXArBonrBp+1
Re7fTEqIhY0U0ULrm3o2BVcA23e7vWbcLGHkp3SPvuxSd6dpltbIYm0gMjnFLHeG2EYMmH7T11ol
xhIqlYKZSHSwa5KpT1Pp9wtiAio2Afz4OxCxvSco6uQmwFeHyFeKhDteYsGnfCMXrmaEYCd6mbeI
GOuyLrntINDPaM1dVanD8qFAZaCUMdr9ZxPu+Hcq5lakzOhr3aDs1GYR1sjV3erxhHcyhHxpsTmo
lhVQ+3xEQMnvKSeGIFl9Kn4h3QQeMOxDGz2J94S5jn1Nm9NySHM1S0lP4bCAeP07JF2IsryAD5vA
f4L+uQ4DDGzdRWCUmuvrIG6CBEbpSB/MqCWBdfjCIEhJbRzLuV5EWwHkAmKug9e6I47lKbpRKZ5m
yiiT2AgtdbEpLcTv72gW2X9ssr8qh7ioIEpve/oMtAuy/biyWYkyOnR/JRmtBwMfhUKs/RnY1rm/
0X0c9sBQG6EzNwJsb4LxHhcneIlOfah/tsT0ePxgERJL8l3uf1YjmYSEvZHLtrhB/6kR5cgZ3ZCa
DrWGmwpgi+zh8UwkIJKSbXCxCzu7QmrFWgdxr+Ngj7iaYs6BQTxSTMA/26BGiB8oWCOW9kRo+R2o
/AAjAYmAk1Rv293H4QpvapsQcZT+VEQlONBlZ7WVMunhmeJAk3aWPNN9COjVLD3qtfYgDphHAUFs
P3ZL/Nvk7JcEdvFWYOF3qota5ptbzUj5c2xJtuVdKNDitvt0TBpaOtD4NcBN4Bc0HRFxv1Qc3cyt
rrlFHfFWN6TzM4HL64jyb71pEHv59OY3YOcE9McRW5QrsuqTrw8LMrf8iez/ofIio58bMVbKfED+
++BVwZ4wAG233nSOkhhwYay833rMX0R2c+Rxb/XHASSSE11gA04AOB3uCaHdnKA8I7yYvn6d7pt7
rzFNBEm1DmKsPNmGlTYF5iHIesIJEu+MHTNwheYgafRraNGvO0NOCAysrxlpFe/QfeGMTWm8qdMb
54BfFqs3gtR7LZB6Tl8HoayDGkH+DJa01Vza86cbdhp/qt3RyVMbbDVT8fXtxNNW4jdWh18Oq4N+
skOmDjn69HB0WaqEFApBswJW5xegL8tfbBo3g3I8q3BX6H1uZ3aNnz1b7t791TR9/HzOFSnhiOvd
I4RvPBWSzIlmnJ5Z4Xq+yXwC6afzCU5qj85uLxAlklgJE3fTuOkp3EZnnqR7OdLAtGumpZNm6DgW
3q/YImvOkRbNzPbndPQyGyfj9def1/UlEDJ1AMYTAn7fl3EP6KMlmCKMoJkCV/h5mraQV9H5+eEb
rHZE4ixHNQ8u0tJzE1dDCgxfmQLTnv/383AVju2Uvf7QIYtED5JHpdt/5+/WtO6uRdHSk7ii+F4T
J4s4wSUCJjkv8MbE52wlI7cR4O0sCz0UGE3N68GMiAotOIm+GDhAeAnlmB9BhGiR1iqFvLF5BW7D
ZyqOKqLF9otSkY0gSNa0XUWX+YScNv0Zhlc7aVj23j90P2LWi0ebEtQkKBs9vG9BMds0OHNXOljC
H76EQYc2ebD++DpIBF8/00b6EuIgwL3MPuNkRfgnCwajIS5cEUCHrZTeFICJ2WkXXuypsCbqWo3q
836gqH0YKtJ81RLzjLmGxW5qnHz1vpo13W2JvCVTHTDDMgKWs8INt3US1niahbhBtGgyoyEb40VB
t/tES5BhyprumN0AMoWA0qmA6BWpXOBlOGg+DJdMv4MfStCUqCP/61zU8p+oSzI8hvZ+RTrwrk/j
QJdbBdjPqb9PuJP5fAMMbXTuIKkF3WP1wpZo8f7bHCluKfyfI6XUT/mpNz9yigcepTA0wZJhATtQ
5JzUImZP/f+RZYVFBRXG9YGL5oo9TPzftTiV7eSy4HWqWbnJU1NaFHDmlQXkAGLmt2C5rInpeLum
g09G5f3EeayjYzduc05ZPB38eppqZysAhs5eFFRHXBS6qRHFlax35ccFkkjKHgFZdG9ODfaWxkDO
bUYMDILFS+XPxINCCn5dz1VCU0FGjNptNPUWlmgOWQUn/4Kp44DEumYV4UHRrcZMARcUO0XuTJEZ
CcBQBUXV/4bYDcq3cKBkd/gTaYrbWuXemauJQpi644Od4jEIuz2KkoeL4v27n+gn/D2AA/Pdcgz9
Ie6NN6lFgVcpGVQnEWNgiW2R8ZpKfo4Iv5jdoGkENMH3kIteSFmHL2U/ieUf54aEsduNrBTaLBa3
g+PmmkdVXhjChzhwU9SS5oAkNWmsNg+NbtelhERW2EDRPbxcD5cAbeRsveZJyEP0weBiqQ6+odYr
o61vWBVWxDIgZEtUkkRmB9Zh0JgAAh+x1zLv1f5TLwFDVTHB+b5y8AdhuQw0VQW7hU5BBqVxdEVL
+EkXg7DnolYTSsbfdlfhenbdcUvxuGDGGAxVU3F2ExdV6XzVT7ZV9koOZ3PeTilxGZ3rXSzry/pM
Hhw73gZbMBzlIuJQNuNX7230L0zj8uCBO65rxAJBz1QPDcqMJzEHwP76Tdt8x/5YZd/PV8Yr+aBg
Gzn7XXGP9KLM1RlOb4x/YknRb7Dbi/IPkVJ6hnhM8puRGoRQ+CKGZSdtAcJVJz2StA/CLnx4Jxkc
ct5wcpaI9xXX+GfOgvsYmZ7nqu2GRkX+NEw4/O0vc3d1cRHMbynR1LgHzRIDl2Q8oHZMA/p9b9W/
G7U4AaU3K1ZPIM0IC3U8gaaHs1yfViUXc0DiEYXRoTR6LQ2aKePoe5Q44nEyYs6ZrLWhQIULfG8K
4gO8dC+61c4plWyxeWqy0Tvx6YL3jJOVelVJJ3sZTD/I0/mgk70+v18M517ygYRiA3/HRicwwSws
Uz3QC4HH4SV7znS76V3KTUdQcF95JWJW8Gel0wjh0DQ+R/7EbXBs8ziac4O40gZdemb3IAcWMkKN
+ESsnCeW9JWJjzrlUY4otQZ2caWWs58Xb1giQYX8r/O1ApYiutzoYfIKd33eL6fB7yS4yCyWbcE+
B6xQQARmeIwn8EmGsN1NccMRzzo2EG35IYOY/KSaHFw169fzVFqo3qgbXJi0WS2Yee6mg2M49NnG
N812iNDgw1JfBxKoAECRMXy4F2c6heLl60JCwgp62/Ld1wFNCbQDDMJWTN0UKPH+Oqa1G38NZyMq
TCtGvthwY1vTmF4Gxa8gAaqxOltGyz0ZHy/Leqv3duRDbqlL7ceGQv9Cf/Zznyt/uiLwgqjxPX+S
BoALQVK9cNW/bvwjJXhHI9e7DWHfBZEuPY3OrWRodswrte0J4d/ENtDVJVklazw6C77ZIAej+Na3
0AUxVuEIoZuSugA5LDpp9KujDXKoP+xx6Kcev8dF0eOyeH7I3QlVBEntCY8Zbg/INys1LtSBBypf
MeSwOAYuz3EMhY3aK3G+1x9nuKQnLMJ8fOGlh+148LaCmA9FqRwTOAKv54gQwbZ40kinJQTo8sdq
ShPtH6TBlIFWL7CqUsbXRH3tH0S804HApVBsQE6g7fe9DSCL4j10Ca5k8fezXSn9fj+0axYPS82m
E4vJvQF192Rogww9oqa3sXhakBKlRKPxOeKhf8NvxkusHjjbYc60xkDVHyvI9o5yrBI/VEVZVb0k
ptzeXuVpeNdRpKiU6o8IEwM9OkkJFk+h4ZugZCQAd833baxslASjW/dMRbNNU6je+fikenEJwRe9
KdVR1WFWi+MT46TN3FdYues8h+ZPsavLn89ipHInOG6r2MbgpXwMDwjGAFResR7Ut3WsKk3ZkW0d
3/2sxtINfyFY6+Tl9XRB9CFyBKeiFn/0nzgImP1CzPKAULeDiiasNCZ4w7vK4DA83OKcy+W7N7kU
WkKAIfanQ/sj8gmXCI6pwPhwhsp0Kb5BDiL99b4Yc0k+xtILFGJyI3dPxauHDwEe+GjB9aoAMLGS
t2BEqm+Q7NkNFRFbE/6d0iya48oYJlMAvG8qpiqiY2qeQAqD+abEcnYvVVqD4pzTpgn+RKhLNMV0
4kXre16l6mD3MjGhJG8p0JCZ3z76J1W3LUArrDR/P1oUl9gPADOj4mXrZyQIXpAkqRZSjQkydhEk
V9lcExalu/NGKEfpo/4XEH12Vcn3RmiLkuTXHUySgHzOrcs0TE+93ezfEtKz3rhlbApoYM9qTx7r
frS8LMnvy/FbwhEvdm571LvhLRARX2CObqo9BJ2QzUAhxpSuDc/+dFL913/6AARDmY06/3zJA3tm
82nDPI61iucaWO3dcl+ZfjDeuEtD3vjQL5KqjASBgOyPzUWKmrP1pqFI1nBNdUUMnvkfZ9Ag1rNV
IVuYoWlC3PVMZqYjLnJid1j8Y5y+pCmTAn3HwDwKGl0JYBhZ4KmCVzy9eIQeBAYL+E8OAfG7hDCG
dIHIjTOi2xTNNzVzjvbvBoFBpyDpmIjw9/i60+7jGaNb2n0t3zqcm9ReghwfxV5bmNoz6YnIzwC/
DCdegqBcRdcDy9rCCnAmmFNi+aUOJyb5Nrg18rcFY0H63IpfGQH6tlcd8EboUCV+t4UEvsdJdpiW
YqMj9W2TltZ3eHuN9jRKbSjYNJu1g3H0FPDf57tR01IpgkHXc0oB6neVpCvtSCA+AhbVoN2w2WlV
WUaP+wPFQmwTLyNA5p4IuZ/l2ttEftZdOBFsuIXuVEq5pX2sUv2AtjsuM3hzoZfxCE4714ZCMkCi
PkR6yi7nqT+hJ4E50vGHW45bkLB6G1lX1nVHTp+HHq+CAaooGQimpKRATa/xPU+nSRKI7Jyq0njB
h/ijVuXI/YJVp8LNBB+jzYNkqERK4ykZ1lPUCiSyctdFCxvVWuwoxZ7jfhyOboR8kRknOBUPOj9D
i5+vVX55RMFVt8c6Zcn2LGsyoiV0VDF/Ih03YmQmGNk9q2OBeIK4W5pvBmvCgAwVW1iZ7Lkxcj/f
S8TzGDtm5RQ/hXhS8kPKklIoDiFD9fDpQFmvIVyHflvtjAFqnfA7Yfk3kzL2KbSxS+DqZs/b3ZT2
YmWyYK0WMf7fPzgvKVR8fybxedqmibPizI9e9U35LxE7G9+V9uBM00H1Cfk+rMF88yGckp9Vsi3M
TBdVwZaZk3nOx+NR6pF/amTKToOc4o6BWyxIv21Vsmn7JQyJFx0lEmHO+q16QVxnqMuwAvdyYJdt
o2hm1kfHkjg+Kc1zDmp80jdu+jzeRG+EeTRf8EGkSsK9JuZl/Gp6R04Rs9ZCCQ+F9+0RzeVuHekj
Nv2QKx3wCJeStFFOhMcZzGpKoRBR4xc9CSvGmjiW2q7xmf8vOxUrYPASCj7hBxUwWMnvOyeRMi2p
yINrwGruxDj9AI226hnrYB3mlmnmXxq0KnVVcKcZl3CyP9dBkfWSvebU+pa4JhNCBlb0ubpzz9IL
+TR1xuB8hE0JLA7trEVHA7tcaXsZ9Go7EojDufL6xDQz643SuyS4VXwaugQ6Y9vuQJe1WAODFIyN
vpL9EFtSuPHbB33fsn9wkKS0IPGJoPanVPrkZ1zSMvXiGIqvewwuDOyKKc3Th0Nw/zXyy8geS/wc
RExdIPBZlOkAeU0J8hh466hWuAT021rh6djyt1Ku6Rwhc96MkChouzl/IsjsNIJSVK59VKwYlsxG
9Cnp9sZKVi5/79n+ZxuB01vXzAegxVhHgtI49F1Ifeg1SLk6dd97orvePzrnq3UWE8Dhou2nZE6y
vzlwWGazHpawidMETf7lmORYH6Is5aXLk7jWB3/+zT2/8pH6U+FoyWjxo7XtyRHZuIukHXeucmKV
OJ955zQS/52lsBZcOY/Zg5P9r8Nf/hKn7Lc+jD2v8Jq/Zk4lLbkz4UsODuOWBFd14A3Nzc5rCvcu
04EfFIzpZ4gpgv40H0oGZiil97aMFRe5NdmSSyiY21zXJ9CRDN5/R8HE6grCvwmCmPzBTpCMthWh
d8khRS/It/nFjt4VXxbOZxr/lyiQ0Db90Xlbly4U25zcGN3EGAg3e9Xnlk9+1HDfc0FALAiLfp1N
BAljf35Kv3UqEBQVkZUYi9Zfi2GmakWWEzCajjgqsYrbjHS0CNb0ZQ0V5j7OzGSttawWPfh42CaH
Il5klGwfl79vUN4UWIrx4vf2Rmw3426cpGGAOf78ApOPI/YOAbXGqT2v17oQTk6F2mDlBnNH3MyC
7k6gYu9f1vP5W5Sp1dCkCJWSpQTShrlamgAkaKSGY3/U2NMz0dur9MTJli0nb3p2q9wBuAqbT2+y
UbwOM999uIWIFNAqqAAExscn0GJ00zc6dUdBHXW3uBeMRD08AmhnK+1kfFabhGvnTRQIGxM+Nluw
XAzgBpbslORpkgGMamrP1iCr8Wm7uXBOcQG6pd9L4EOKXhl9F28LkSkToY7qqVfxUYP20nV4+Bam
KULHZWg3d6pr8oPgm2NX/RKM+p1zxqWLogNIzSpmiXmxFaaHfL+6uEVqbDDOchwBJ9y1byiOl9TO
zcf6qREDEihgMTTB7w/kMbyjBcuOe2QT9FWZFVuonbJR5LvGGZNkBwnKTBi697lmzlRzlQ3wMtaY
dK+pvCtXrQ77HE6lriaiT+S6S54aOPt0lSLBTPddQeyvHjU26fiPlUoG7Zbu/wPq0Vu63YkALNMm
tDBA1x4VKHiX+5NB4Pn1RX3xGmfynjHzfHxr8Yh1ghtIqoBB0lYXaNpY+HLVTG19cSa4ZqeyyqrP
ADSPJ7+K2nmxCKbusuVFXXRxsnki7DT10xIXVNzVILWpS9dA/yh9gwI4o0oSZXMolKZQxl8chii2
2ETxM87Wm02Q5Wrye8CjfP71eVyJSUk5JLwFTGvvi6twlwCuc+oc4RJvjfXEfm83gbC1hIrM5iIp
k5/WyYcdaJ6gItnCd9t5rvE/PoVRiC9skYsyxiw7o/FANp1bXiUU8TXRNzdkiLk/S+8Xv6O4ZoDb
W7oEQ0FL6Yf/8royR71NFsy1NtxIq96LOyr5wQWE5ROfLxFpy78N+7LdOu1ZV0GJq3QO3eMyp1Bl
twxfJJPQ8VQ53QTNPif7mS3YTLKRMZDDV4K/G1UhxOuWV1o4nrJcxcmxn2yV8R0mqRDf1dVKYYbh
QiE+z1W8wRaoLUOSI6JkvzcLcfOeNS6vVdBCjQksOHeCC5bzJK0HBtCkz2aiCAT04EAuqU0O0L+b
vyRMFTmQUNwtnZY/awHA8PUfUtayGVtvoo5ONVOVbFRV1BDq/m+AiuZAD97FU4qN16kaStiqHzQB
fpF66bwy84i1Xm0VdaUXAfCYv860CuKhpBBtX/9wbs0kGwbE1uisGgFCLwmC8SlgxJVNqt/++5KD
RFplD0Wttat52yFleZArmQMIA59beBl1nOx+EirE7xLSiYPP4Z5TKmaW8OQVRWB/c/ZaLPEaVt+L
VFSEFVWPwRiBPbzriS94hDcNyQ5ATSH3IApe+B+MqhUrOoXPp0u6LOOexHQgqns+1xGVk4eNPI+o
IiSbmYP2I6zLHoSUvy83DrFLMsP5hGFFzHWcNEMi9A90NWjXaQM1bxwOUek9o2Vdpuj6anm0Dkhz
GHdBN+3ogw/HPYhSRVesESOmSe9GjuirR+zYjxGKNrJ/rOsSAg9LML2UKiBBIDi1jUq3jCpQ7/6Q
G5dBqaGlJqDRFOiIzQAb+dvm4Kg59eBv/3q7HYzAZeHZ2FkCDPSxRm080PvpuRCHRA4XGfbuYqe0
7+cEmfwgCdgmd/1tRxmCpEAx9wL79LCECe6EZMf7rEbh5dETfidb6utuFv3UjEYK78pScQ9S4zvQ
h1hFecjG0nXVOxPtfmh+ptuDrA9GB0ssZing3oZOrhJQEZWAdPtZMBrEnPHGWqV+TfmpbVr11Rva
JLLXth6bcnlV7dOgJmc0HWnJW6knE6ra47NjSSKOMgc0PJ8R8ousAZqqY3rIAQfSlxEeJzc+SI8B
k/iVHGhHL7yfUn/+Fv2Sf6O0Mc2sCDFKqaiLuW6+D7p19lvdyUleGBF0fxqs3nKflKhixay2NF08
gx6EVL+WejbOaKi3OwRCFkUDd78QSK4M93k+caXNjP7aAzXYIkrLbqKTxX0ppEXLqM5/ndvXZwuo
VND8oPhIrXnYW9Jtfxz87elN9sTPKxe2ujA3uzBwuzCa2kJpa3baMI1Six+xeVVJPH1st6dZ+Qz9
PCYyuwN6RSryX6bANMdk5EzblQoy/Ba0pHGh97UIIezlGYmg2QwLEHbp6eZHtYCHXL1iwZ4YUeL1
tILTaz+IU+HSUAFHxEHnX9IvBc+HL68rJmQYjyG05hM4gg8m2tT7pMmz9bDx7JnlqMEOXLSOlSfy
l142M2FtzG1NMVWY424WgWztYZh84Qcly/gbcxQGH3JqjaYfuqfqYBj2E2VIjjtkxiXyvhqdN01F
QDL4fKW/dVJ9gVaJyStYdZydnpBht68Xvj7ksEBeAPcGmRgzzVOl7EUKC+eGdwa3T5pmB6vRwLQT
d+RjJpDv4FYTjgsiAcH+oZ0r6Zvg+QFuAqq9XfkHHsc5CLxnZakiSV8jSbX19kL+dHHWGZXLxrys
l1Q5HPq6Z3avzqO4baAJYa2boO8cDqA3unxJ0lvVnzeRbeT6scVN/R0bMA0piGxtVQOega48ZlU/
13j/39UafrAnSwBS4flApowy0Vq+I2WeeIeavU7gtgJW+FQLJe6/nNapfEHNUcOi09zRoXX9bpi4
Pj+QpEN3+kd94QrWeorjfLuq7Zkr/9OrXFYgSLvaxR2r8Z8iEi9dNFlkEj/PVE9Ll+Wv5EBvQG0B
3IsKdNzhC+UjloPNijScD66R9bS802EjGnmHxFB2sCKHEsq0fHHT/T0o5UP/av/l2Ja93VbFJHPi
7xNvojzprl4uX8guz86ONg5s2K7a8t7tssu9RJEm9burSmCpxnUF0jVoRDVq90e4Opwiy35h+Y/g
pEQ7937BENFaGwce4/Wukz1GgMiiK6fOw4g8mI8QZN2LsSNRp4cjqlovabe2PgHDobItWTQbsHEG
eRPLuBbqaqXyWts5Z1Y4Un+Q4+KPaVVWO7kc7UhHQ0xARTzdlKiWbQNz3s1NwbHIxtZ4n7/ZHP5/
JMlgWT9J1nGTVmb2XNCU+cc7iKkItd9PuJjYogNM+KUAn1nUyDgsUCvWprWYaeahNuOOqI+EuRJJ
iStbeN+rt0wirCPIewh8WItjIgzoeg1QEihWv2P6xIcj5XKXe+i8GPI4/QgFYyFw12LSVPhJ1WC8
Gi6zsqeqkRWvIB5txcObbCHPE5Y99esA00r5hw2yn0cuDS5sM2P3TYytOVIu8V65gA7+m6BEHI3/
8DFYsz3k77Nx24Cc/kGqz72oxe0zbjPXVdSHgcR1kJrJa56UpVvWzDUyp/yQa0afoORruhyT//R2
gtw0B5LDyGTFET3x6AfvjUVMJ1iy5V0hrCbGVC/dmpAcIV1piVzEWlCvfP78b185w2vSwL7PxnIZ
tMwvR1FX7Zr3hvbohRXEstSn5gtgXGDwhKOlqgC6lsKs6evkiRpl7GIFTOVfKYWJVbNQNbYKvL3v
jBfqIXEISq8V3q2shEImw2dlAPLEV69bHWnUWQ0IR6V56UZZ3owm9ql97CHAwOLemAsQ4S4PiBnZ
6x90UVuhzwansMdCWBdRp+ug2B2k1ejyMHl4gdgAyY7CFZHbkjyGHqJyevN478oS1S/Lb9lMto/B
jEEa+vlJSVskRFnrPvEi4I/zSJHFI9iNN17kE6mArrVCagz9unuNLyiDOaBGGuzWD36F70TzxAK0
aALDQqs7127dyJvbb3wP2j40uGX7HxQ0Hw5/J47+pre5IFaJ9koFVkG3xKVXJTHjgMvSg5XJqiSm
QoVdnM7SmacZJF/KVyfDhO2zh6oEUmipkrNQ5JIVdRRvEcg/ZMnyreepa7SKIARQF8cHGRiGcU51
93syV4w831gZGwLddI6pb9n6BxKUQtZ3/mS3I95+zjlgAclceSxA9j2ITMzQl9YHxt/xF+Oj4a9u
5Z/WcGMsum3kqTszr4GjG894jW0d+Sf0ghGG41OqIypnUEDLrKO/KbNw6+5X1b9IG9UUela7EgIy
o3tWPFn8mvGANcLBVjd+In/wQXX9wAWn8WBjDW1jNsdfuhsTWu51lE8wrUfrodY+UGPR1hjsm2v7
lTxWHihXo/29pthJScXKpSK73uZPyXNxxROpv8Q9UCqUT2oDTjNsEsD8UZYh3ZIKt5vi4mbTsW/c
yzXhb/QvX60hVZDahwI5T6rwVuEi6Cy/Rbvjj5kgYUUHeQCyF4MGsmjL4Jo9Xg1yh/VXUIne+Rnm
QDZnFC7XqvBI7Tb/j4VUvpD6S8qx3FUr0js6RSIb+PYVgr7DHrJTyP4bBfLhZR5736UReyXIjlDF
XFCCdKvmHeFE0qjyhVWQMYutQoJNqhQbz9YCilBjuwOwyOD5PCbGDSTjhAyG8SfD2y36IJ9ZxyNM
aEKHR4H3L7pKTPF7c5GHykpDkQjEx6d2DVH4QUfi1e8o/qvWJTKejVEbEySdWC5sMrMOezmEoKFS
AU3lT/b7VfC9JVIJdJdTByqousB3IZaFM9T+p5zvVsvGJIMEqL2rFStcFiA6vpkn1/QdDKo0ANd4
Tofq614Km/piwHMqV1ASHQiWv7EZrkhud026mepxKOpkG3e+cT/bAnWpXe1NvhcwV5wkqT+eke8a
74oIIkGYDPxmRa5VRJU+/+K69NMgXah/Bi7DdgfoWXKNBEgc3PcqB+fAXTIVv16U1nGB5qYidWlE
i1yRTV4cqr1KXwywz5owo+1JaL05bnxuOoIJRSWOfCu7ZNrFQTYC/wR+vk693mlJd/3uEmYDW7Ps
VLroAXhD8XxZ3S0LD/UJ1vGDZPdEUp0aTZmCsxqCs7sQye04QkmQBUrctUSa+S7VYAGyaGES0JN2
1pBBTy4ds1AvCySfcNcWYDbhEQ+sKKeTORy4vAka1PNN5T1da+6qSCq/o8lc+FLq6OrncGpPb7d4
H/DOeKoaBcXyHN8nD5s7vAOg2+eiMg8RnjWlTvyzhKS7X1Z1L0QhuP1fFKpgwgz+dqryrxMIw+Uq
ThnlQf/NfOOM35exBh3ygVzcTlOQh6TN4MYREoJsIPGjDBQ3tEgbYRH6/Q5IVU1B48UpxLh4XELg
bd1sJP2FbllSAtxAH1RlmoxB2xx5/YolmWVuciK3IRadS4GH8kj4XRGGQt0g6ULSb/Ke+tXzJeYU
14Q9xz4br8Yzi4vyC7kcvm6jA/WAquAbjRorajALbaebX78jUDhJrYPf9gxxbRq3vm6cxD43SZIU
knJXNDJi/uCD6qAIiQ36SmVIFoqubONsooY/8Kd110gZAS3Q34A4mKK7ECQk11+zHNQaTVdzR0+d
L7/4OT5OKVWUfTir3qOTO0ZrcBPaIRDRhQr15j4uWCAUWkh1etWeuVzENxxzKRnl2lQG59LlFRzU
TU4RlEJu4Li2NlIaZyJmpI9T4TY9dQgtEQNjzJB/4uSECzJbJSmcJEtd8HKHv5dI7VArVk9bP5vN
WJ2dYwh1w9/lSnm6MV7FrNuBJXaw6sG4r80pIzWBzqe6wJJGoF/qhmXNKlrwl5iuTAxSSsJ8xvYA
a581PtKagrDNb63cxLDfXLFjjxj3Ykn1BcodF8eIYUqqKJWsP2xkIskrlLd9pe4iQtRdwhOCh94i
v3JND4KC+XPt+Hk0FJxRl6zVrG9pMwMf8oREERZoG3CtQVw5FYgy/RYelu6OGvuu5MyLXHHRe+ob
imujewxU/3EkkEc+9NiDrepiyEij34T7HJkq3oELV6s2gQ2gQ9IjtRkbsR+VcE1kjGCUVyDOmdQr
HP1UsTB3Lvixu64UUWhzTWMUKOaWYgFu1R9te9uuZz214uYnGB4CTPWStWNDUiRB/g3RYG2p+o5F
ansim7MltUdtJF5kVYSxty5ndmf97/22Y3X/RuUtr+huzXWfnAgg9JxCK/ruAZLCUAhw+9g3JkBk
eLcwU0Mux9RR2KLPguhAxKfOHpfMd5K2SLOcWWN5o27bY6TB6xRXBdYnq/KKD8Aat9Z4nKwZuFhl
qmvekq/lkkVlNX03nqbiFxKNlpZEBP9GpPI9SGQDFA4MX6AKWt40n5VkXYtkLaXKDOjk9977738i
jt9UxCmj10U41b7C5H898CbDpXqHpsYRM5Fp4A4g8B3vcncXWBSUb6wq9kEj6JW9EJoPFqce1MjI
SdWQbDUpzBuZr/lJa65aIy5ErGNDe+TTZ4kMJAIOLZ83uZ12+obeVNZPl2JHL9+HWxrYOBs9+b7t
II3Pc1Ve7C4wg+lw3lavz+JAD+gJZRuV5W2mg1CqlMe1qdDnHd9LL2ZhRVeVY06vqOv6v6Os5dQc
eZy9sc30XKZsRhbRc1vknMcs9Zcf+tvrr6EsU7GbBmXKhNgBgrbzdLQqzL8eDs/YU2OWdJ+GAFMu
KMH4nZ4ZZUACG59rluYV5N9Av9SdERJtztxhGF+a67hHlqpbbV2HMdZ3nILUdQJZmMSpNfk4Xd4K
sb0UuR0ovWmV54777ZVFib82EMrvDzbfyM7yf5e1U1LpVDtsHuODnRI/ndD7a6TWAhSsdwx2Uu4i
jZ47rK+4dy5Gh00s/5BGV9xJxDd5xqql66T2jUBvDZEAqm5Alxyy/4LE/mDi+7TgNt2of2kUUFsb
WdCXh3ZZanWIR/61DY0jLVV1E+7O2snHiNH3duBfzVro6G/34J2U8DGkfExMQ7mhSAVQDjv+E3ck
RpVqmIFDLUvNLHoxRYyS+/C84MtGBYl/4aK646jA0dHXhx8T6V0+C+eKEhJ2c43FvmA3dvMy2FJW
f9QAglKnapKwhctCNxN88vJGvyROoINpmqCLFdysVNj7Zm8e6xSbn86BsBL7s31THi512UqSH1BI
YzICDHH3MVnJs/A939pHXo/jixliPQY9/2D1uPZpCUoCV53Ny2C9Uul9xjizxB8+fNP7XBrGuTCU
mOQiHhhmxi+ORiHjcqpwessRcjWC7uoGaS/2xN3A7JsdhKBk8M994CvNem6IGpGJbKi2xlJcNtKp
TyayGPX6LKpJcKZ7X2C2Zc/oQ132H7cnIwUQyagEMfcDfNdUOdUt2N/4dGIulY7jYEGD1TNBVPAt
2vP2nHk2P6DzSWPrPBxRaawA2QGoruHzkHdcUx7j6tb5yJSuxOIcskiAsoyBhzL+e/60JTLMM+3f
2Rw5pMucWimDfV+2igInAeb5YpeL3BWqaYStACJ5TS2kFgvXLH90xx+2Ws0EpfoC3GiF+LXU2ilV
W1wDdNn7IEvJkdHQXOptO/cYfYr8uhwDGGDJOQ8W0qAX1plNN/FYtV9ij5d6ui98pqkaeogsOM+Y
6xckfqtaPwegXFasYtAnM+88E+mEpjMfVulLjX6qPiEQVjW38f3ZEf0LWfkwGsgs5Jl4woESg9tB
TXncPx0beC8xwExRBSwKuQs/ocR2evggHoQOEEAM+RSBKZI1GQ/ajwu+b66nyiHR3v2kmOmSDZ48
+sXUGUtD7Sm9wR/bQZZQXYcoR/KpajtHrGxmaVErFZ7AD5Xofux5KEfuZr782+w5tv2qzrDPbgHW
68JCbGq/yywHxIMSa6BmiH0IXaSYolNXMcfZKIzyJL9+4icWuR0a061uloMgueok0xSJt4UuKP3S
0u3k/Doncvhxj+Y/H4IjAlq+Pqat3NqUSkpnGgYJ7Z6jOrvis0uWWjWDW47WS6lWs6HcEmYXezPP
z7hKLOLKnDUfIN9hyQOO+i0zksN1FtLuey8xRO45T2E+F7V7cwQQXxO6CqiwujW664DXi6zu+6ax
MEdIFC8MeAUg0bYC+nl3BQ4tDjvOVrKdWoT6lc8e5Qf8o1MdkjRgNZnf2s1axYrvevK9uQ1V2A9G
5xCKMGX6Okc6qvJHNZ1fqWPOEoayE2HY4eGOObIKCjum5BrSg809E+LOM6WjY2n49KfeOPC967/j
LFDBX+4O5GcJPb8jL+KQEd5ioCCVJ7pO347C20eDUEz21Meg7+IHfIrCJ3EeV2QiX77RvtgPN3o0
a03JsGs6KqQLvODbgNPGScYPZuJAHElF/ZuoeGPtjV5/48KSQDbBC5g0LWxBVwYTJYtNmfY+zHIb
5hw7O9hAn+R58iXWeWsJImHGdyzR5eyCztyQxIhIpOZZiM1ESU6wEQCH+uFsFI1PGpUFsvjj6NVL
PC442mCzt0RE6aGtowPSIhv8YUPrRoMBdCqxIJB2K342PVuANYjEF7dzlHXfRz9vfwJngbXS18US
jez8vGSpaSAZwVvQSsis2D4HsoArg+3YRIrJrdb7Ww8tj0JeLkHHcv4i0rcJ7dNAKvjeWVQxeoKJ
JWguF9qo0VJP49Rjc61v9S9JFkG3+bv8Z/S1xks8OVhEo/WrWfVQLt4HwtoO8PNoxe+FKsfuCq2/
OYwRE8rdUfaXkD7/OK6eCZpRMTZa5TqYyVGsiZSYarrgCadM3CPp5I28QfXnIQHVIqvIWSxqJLVo
SSaPI2BokRTYBGrIJCxy721qeDGmEmM/s+R4Sld+z684AASr34eE1UcKGaQW6t13IVg6Azuxhn4H
gbqcN1ml8UU9SvdFwXBi0e4pRUOSinmSuIM27UKMSCYtMySvtXOoUHPBIGp6VA94CX70K9NpApBE
dGl1nMnXDTby0e5DKaFBM69aawftrk9ePFuxczTwGjC9ia6HrPFYaXlLUAtP8Kw71YmXg9yympQR
gxe0reb1T08Q8DkRFS6Qr3Pw769e5wUNbBZ0sVB7LfcvpSU4gOyiUxSSSxYvvkUf7CTEr6XJBwk9
oi/asOOE8Z2oz4i24apzLffhbT2vlJ6NfhYEtaiY7Lnfe/+eOSE9Loqpb5wLZB5o1SWKI9Y7zwZA
siliSlvELYGOV+75hWdXsqVuyylW4R4+zWpT5o+M7jXGMqyk39YbShSEGHsWvbicZlvw+mMY9I9m
ueQJlUr3agDBWC8IhuxghMYBSgrA0SkjZ+d6RebInG8a+aKJ/yc4WJ6SViVCn6IJRTX5yYFZcL49
0mY/zciv4nEOcVsHsLzWeXBnQ2/E7Kl1ZaE7rXJ+a8l+ZXDvJXCaP64yE1PIsdD1VqP4lUkRH36O
j7hJH5VJU5InCttt9Y20fqPVUMZbGD9Oa0Csno0iEQMs74iP5sEfcwOvOJfCZY5z4qDx/7SLoWN/
66sCsVO3QLA8GiyND2DbQKyaR2scJv4KPek25Re0gAyxQtcloEk4zrzjL50WTbjQ89Sxlx9rJg5I
FpyZhFZ5Yk1DYAWsHcBM9PMgmfwMeAscAZqv/Ez+OFLqCrTSDJBqdnsMqVD5yoV19+LN/v2ufs8N
zpR5vfZj/ZsUxrtVPNFsnFYumAimUsMyLZscy9dKRO0CgqTZOpBKuL4tmnokOnp2i00hbRytEQ98
Tpf3AcYm9+2J4evKdnOWYfdnhPhuHxLVV6H/wkRuewc38dIVaWPNLfZwp5q3cgx0NVHtfWy1JwjO
XJAh8LT1I878WQgXEPVyumPDyD+Mw+E21qAXoBE0JMDncCvkxK3jpHv4S8PqlzO3PK//RXdMwyAN
pBbkWBk9XxvhyZjHooUyqnaDRGcegahyqrEfn1gD2qGMq+k4J0hGdAbZwwtg8RvTTW94Gqq2T3ow
XKjm10hB5mCJ1IyRjxcs1Djms9qrpreXydfPS01lpXdSRxn8rjX1WETEOX3Uw+9zuua59hV/J6/l
yYeJogL3IR3qVhNVzyKxdqu4abrpzx2BOpSf+1HBoooCc1R7tW/k9ulym/5Rn6aQnmHWa3mt4zby
FjfMHDpxq23AvkQE9UQrbtssa6PsL0OucAWzfUSjV/EM+NWap71m3bZT3CUEWoCxbtZoUPTKSene
zDNkb3KXUZelwGkoSHaBVYj7QNOx3xEbKnFHUJc4/SUD0yDrNsjuJf1BnQNSvA0QM+KomD5RS0UD
ZAG5IXBn16wML4LXVjQfRyDWoCC5NVZx/PwVq//1xiaBh2NlxecUuyHrK2Td1t0mDyOdES0rq40S
RCqRLzV3ZpP4XVcswU5xPHkEZRLHySvc9meS0MRcPbVfiNxQQZMgM9qjHEa4AbIEKCwRgQtbxBXB
cpEFR2aNalTcNjxW0Iyc+yCPe4PqW4gwL/+MsajB7S6GPfrKffRdqh2cxdaWtqZWSB4Xap7FwkTk
up7wG59F4ZJYMb/7Lrr4J/5CHs58OSskpUPwpRxak5APcSvvxrkdJPPfQHH7qAmHkq4kOhxdYPFN
r2PJL7LIaRiKRcph0ZyWI8wdElWUmxkHOqrzZQoJ8GYkn3/6txtBd33qelc5XMA3wKT03T1hyTvn
ABpxpMF6q3WvU1tGshfsKiCMHU28iAZVOTJ19LgCTxXO6dTaocqwWeuC2nbnI/clGlHdtT/L7LWi
7SzCyQ/ZA34V1L6aVLBmOMyFaRd1rdJ8piPBgWGM9391udjgsj/DI+kTNmJHMAmfT5Zbr00i0mkJ
oxeq3T4MYH+Z15G4hj9gSNBb1RDj2wwBDcxF2bxIJk6qQEg5+NcoENQohNwoNlTRPws4hqLdqJV5
PdahF6qxFk+85rH8ShaUVWweV16g5Xrov/qS3JE+1W92XNFbYLEv/pyiHGzlHhWDwYNvG7WZtR9D
pg+DqtD2gzopidqlB3GqhtZ7xjLCKrkjAu/s1fDEQiJAtFXz91SjhH+a3pnCFnbY8VvyzZzl48MZ
F/MKfX35CjFS/x6s1MFvQyNNHaMevMuxoxtOkw/lGfgQ9rbw20kEjngcQCI5rNmdJfaYnGbJ6Imk
fzEyxtTvvNUVM6mfa5QnRS7OYrdQWgWEswG2180C2D/uk8+nWNZ4BiR2DNpoJlFCG9e2YuQDAizB
OrPa5BgLwHb7lIiMhJS8YjUWu9o2jIeRcEb+Jglakz3AQc8XbIyC2zsF/D06+vcfvzATOI8bAapt
ZYxC0N0VuS4JWKwGnqnvSPGaFdkK01rA+cimrbI23R+dnHyV3InMJiBlkMQOAiViJP9khL+9vIeV
AGRBpqpUW72UmymMkPsLmJMfLuhCXWEU/KOeJdyPi3p321lqF2UyKQqzWq7mEwgQpFLEbUpB34lo
VdbAr9BE8qR8I4GrsPeTdT6Qp3rA66HFlh4S2PKSNYKbDr0pmhs5mlM546hH3mzk+Tw73YVpqT0K
GFOzgIWLbO+aefDXoWa47ldpNZgeoAnzOfrsY3u7jeOM4RaNKW/BXcRQFkejjFzW+88cWwDv0s6C
/xFPttk2gYGHstVhT7V7Z8iBujxvMo6CJBTp11z5VHLScA9KxdhvGhq9WdhRxEH4Skqdw2mjlfL6
en9E66fqnRGZmC3nbk1wvFCuZhGvQtHUmC5734xLFLgg4nSqWpyUaIx8/889oPicOGEWxNxTVZAb
Oa82k9U/HqYc5GM1y0ou2pESV213IccFSsLojKPqC1+U9+NDFcQjQHNayn7HxVxFxDE4EirQbq/g
djC3DnBImMXsOb0pIoGSz0MmWaOuDcHV7j7bBXHDhQBLsLfmV07KHwrMRHgEfHZCdIDrAdnADBKA
OsmikqTJbPDN96sVAaOKfAxUIi9gWSiaFSCbVjLxB4ixU/IcRcesoVSDfza6Q6bZjO+9MA20jvmf
CnPhoEKgoS+Tf77Jct8VWncinV/hAP4ui01uHTfFfMVzBXXDpedzoS0aBxSWe67ZekgYyI0s96XY
JC1Or2LSKv3Z/dfOBHJsfjYVNrWRByhq4ELdzmzHMRMmQ6h/oc4UoeBHshxssy1qDC+w4RLWdjcM
o0D/Ei3J6SQdoIhvN79LMtHJFGxYcpnjADYKBegQF4bXQExZmmPrXMsK8V7/hWYKvcjvxOY4AJY6
GFLMERUUsTx3wwAMG4uH4b1BU8lUyhr4f8OnUTR7r11IjtH1RwnRs+BmOy039YXmHJpPT/+Z4g1I
Ux1Sc1+BZ+HNfSyVNELgBNnL5CL+jiSQDHxvaQZY72qTpMHxE0pTGA3nzA9HPIs/AyYqaNElK/Kr
ELorQaswemvpM/mJyC2O2NyZGGUAPOJHcGqVYg5ccJD6Tn1NnnajHyGwl7iRmtQva2/XHTA0kcez
xm9FCu4latat1iqt8KLDMGDJe6/oAeA5gxOjC1P9f1Y2ao2llmRhuEXrv5o3fp0BlrP6jItfLj94
h6/Dh8Cpf39TeV4BwfyFgjILzMyjtTipruPlfn/30YFdDiXVWBZZke3gqvUkzUwVYnoUZwCBuKzu
72SDaBnTsdGczx/nDkdrUB2fUcmjaGzIb3EgIeRxpHMiXubVeR8iwE2MDcXZw4rwiQw8BFZzU73C
TkkWfAMUt68edqSK4AP7KhjyC4WBjQuqTKU0HQOB1sHAK2BhxRc5gu/5s+S41Cg94JnOpHLRQscL
ZQD8cZWkYlIFctzzafiwbCpjjpx/I4iGa1HujncsBR/yUAHzGfDdf1Dk46F+aS6C02l1Jf+y5W72
kQ20QOxvT7b0NPsb+X9BYO4pGUcdMohOIB/1A1maHo0RicGsGUwn5rpvQCvDQmesc+ASWQpwrE6q
TeMdmdk/dPDmY9AvTEcIEcXRBQkjL1LWBYGW8P7iErHB10M/pHgPMQ9Tw0ji8k3guAhNNXVx7A5K
9xzODTj20GBplyhR/x4R0NQCTet4IHqLFP1TaEThwAt2+1LqpgdAQWfB9tO10SX+oA0ohi7IxTSy
WAebBd0lH0njO9MJkenNWhY4CjcJufB5VfMKElSWFLLEB4TISzugax2GMRgX8Rpyf8HKgoVd4JuA
RPxa9o7sOnaX6hnbx6/SXLM4O1AGNkMbcTPrB3X6uZgFynMGsW7czwpLLaq3QYbOnnm/hq5H5IDk
ObJ0O1+w22wXAIOKq5erktbcrfX84BZn9hPyK7SSCGB9s6GIHcp83OHg9T2QIGP1+ig3ZIinN8r2
/nLetFWa+27chiQT3JlWpbeiDLiRbW9bIpspfXMEOOTM2ykfeoeRBozI7otWUytwRU+tN1JHydj6
QE9BCPhLFAEWyrVW6CSqKQ4fM+mP6oO5Pf0RAV7fW//5lBKPCYS9qoh/9Cxo+8WZ/Zgo1oo3xV2i
kNPZYVWddSiwMlw/2ezOKaJ9o5P4+tzbR01rbRCwz7jPJ/CKMWxVIKTyY2IKCYiFDvEZPfWHvpMk
8ImF/BU9/OOYmNwz68cFSQ1cVpCZzJ2BBSDTE1pzQYcmEkq3rRkT7C7+7ZvTL3DhC4cZOXn4YeVA
EfJyy0T8n0LPN4LpqJLdB3BCSR9IEIgGlAmK1wE45zNbZiQGeFJzS3ZBGQthaDkObUHqRiX/UwmE
zGnaXXD4sUg5Me9l+hoNjelXqKuhpe+tmL2fHzeCfn1eiGPGzft9oYeprPwsvtYmriieSQ5ic80r
O3gnRr1K26IW4sUxlM8Jly9UYCDuoUpuZnFC35m3nvqrBEPNwkSs7eOFyRifEClaHIXDKp/U/dFs
QGDLXJGJ8sl/8kSZAhWfvaZTaqtcvRxxOrdT3+/Af7jE4PMQebHXaUCziNewa+kr50KSEzQsPVa4
NMC6uvMPrlF4Oa9IcHnteFed+KaqkpKnrkoa07rZf6Maa6oC3YXND4+VdQcFXJ9EI52OSp1a1jnd
QigGWNWrqBSUsYfCBdsc/kLHvDh4wI8K29lQlxbA+o+o+dMI89uqOw6ZBuTREVSCDRlpkNa/Wf7O
ajzq3cph8+QcJ7egX683JdzeiqEk92n/hretLMtvq6gsbtpWds/xJ7Zzb0ZyfZkvawYaVt7O//mh
qLlYCyMqUkWm46eNg8UWFWqJbbLcYPvUSafYaUgX52wjoWt7GIIeErclHtccJ6FXJfa4+Unuo6Y6
uQ25gE1236OJoSQIjzYeKKZsckDYOOVkmwPzbGsWvGqzJQ5ELIwYWgNQlXFAms96ZSN/84JxYUfg
FRBKaWLbFFJKf9l4iZUhkvkDBEDg2VVxNqMmV/Ox0KJOIRw7Ey4DGqkc23BxSdjbbrw3ZLaPoCAe
fXVNPzazt7jmnZ0JxbZ5LvMnAxVW8VXQFvt4mrfUBVfi/PENGScB8wz2Le4EQ96muQikbci2qeI/
vNRPC/1ccFj/srXQKWGxi+U/qV7jFz+d83uq5d6bfd8gs0JcBqnKeaI3MSbZRRSV4amvvX6f9Z/w
pPXQa4hwJPZ+Ga9t6KhKHjyt3LYte6SaWT6+7/HGtJ8RcVtQuuk3K1mxjZPw2EXNWN1P7ZJLmmh2
hu5aIIx9zmcsGZTgQNltoTYnTz2UGUBTAoi9zTUpi58szn7xJOOeMYKUT59VFMRzvH6ZIzr0b6oX
lxcMHjKf74RWq+2EGaykkJdZ54TsxxIUVU1F00C4Fho52ftl6aJIuKEiNTboSPos9KA3/RonUbhv
hcJxlG/gOHlKVy0CvxleZp3dCwV6qME3Pzo7XF0ZWv7AHnzfr91/oBToRIMsSc52h7OgxxqMpyji
qItoYXp+x0t0dttXhYkzNgj4f80u8r93kkXwfIdhguaDzCVx4XM0IszWz4Q6GJqZwiBxYoStYXnH
8b5+dcoRMvL6vtf/XdfJNLYriRn9rlQ3FARgmUs4A3IGDNqqSov2L/K8wolpYFfkr2qKsSTkAckc
qGBkHXliCjD83kHsBfbbUTtbNK4muP0NcWFykILYrKgxCMnpHuVrb8ir/NIfUulhbPxmub6Qlnp/
gK3C54S2v1xwNjxiYWGEZ5zaZWj5xq0iiaIYZwCoFiSstd7jaannfk3O4W9LNyow1yHUo2S6S/Jz
ogF1i52Mp+Vno+Oma2ZqnSwKffeZBcQrjppuT3s34Dr3ufeDGElAXNn+tXuo0Gs0vGVcGocI3SVs
kBLFd6vvzgy99DoHs1JW7PBBbVIZ/LzYUoszfWtXiUnTaCLmEW3GIyIX28KNJYpBwgtO2AHIpVxg
zec6+38FHmWFykc9hu3+3HRDYh9kdGGx/RytbB+dTp4gd6ajiEhXgyzLT0GXxRDWW++atg/RUzZE
01noZm0LQLbimZw4VYwOyaF3aqgU4kkVuahDpYfgY6vn2owmvMQEpmiMoLe169WHXlLaQgoviMC5
CXTSSvI9FcqIQw3q7J3uGtfkFUXhhIJHLmPr7m1skCglIs8Cv0wRogC3Pu6EM0caA82ZO7qgRh0c
dmXU48VrWPosOl5puO2c+5caD+PqWVsDbXXJshs3lSaEjX+iFWupHiNtrOnTCvchHfW5CTG7G3HE
/oU3dit6ghbjH41ZNslcArRl1V13IoIRAafZ751w5LigOjPPlAlDLqJ1E4anuncpWVYHGgzDQVtD
J1RDQZWajO+58hPmou/2wriDnCXcjW99cgOlnAztLgBi4pv9PQ6PT+z6a7YPNNpqgzIBN8ED7XSE
xq8lgTOaReyYXTnTb9u/a9psG6HjCUNcQL2zk7CMuyHI7qr6GMIsrk+7z8NfIU3vyMez0YRXMfhf
fORXgcVRR7LiwbAbdiyu0Ii757Bonl1aY/uRHBTDtoB8cHpqOVO4kjTtNNmzc/2rbrLY4YG8VWon
PqCIP/tHOOAkcDk2lz1INTHmyxe2CPPYEVqb5p84EzQ5oX3jC/rIUuqp332jGen4TZWaunHe77Gr
5EBDAqgMXCjwVfPxvWtROgaiD0HsE8iJLl130M4beQBCGdArr1bNIa/7f6xlC5A6lP/xe3rVjFlu
l7vLl0/16xktW7W31yExWHHE8cMXVxjJg+XBEXugE3mDfG43mlYBhKGbl+7IVMwpeV2+FdTq43S3
tj9Tck6mMZX8bye2NIMsy1ZfveNW8AGZ6XZ9YAfxzBTdLQRY5y1yN+8uIar693zt9W6nOSYa+wSz
dis2oQSo0JBsaImxaANEYEwjoThOVAtpVwmYJMiEdaURvmIY7Cw2FS8BTg5j3c5UxDKD5jgvIoma
Y7Iap4fFpDtZl1c6NYgwCVKvz2i7r5z8VRZeDsm2P3thcMWw0yaGxr4qjtMt6MLZ96qr1Qi9Aak4
0WBME9l7bBtze/OZtLZN1T+GHBM29p6K2OHarGxkfXR/LatUMNME7HPL6qJfKPlv00/5gblMOi/+
T4IQpRsKDwr0KXKrWQZhLN1vZz+g9VBxBnTbQ5ILFgO+P4lABPZP9hDxBWtjMoQ7kHDd9Y4AxWag
8x5+fxPX/x70xxQs/nNUS6nRYfU/X0a4qZmyDo0imjup2s+xykqDxmIM8UeZ001YMi7wsxSchK1J
QfV+Ct2Q4xkX0VNFUJEVwA0lbL9zobrN8Q17SjhHEm39adXhPtB8uA+X21fCsZHz2j6KJjrdhGph
DW5OR1wCsP/p5cE7SAsnNysijxqd31+7aUsjdkv5Gpig1wT1GAdpK/fPtMuzzfIh7mlm9+tSjjwy
Uha3S3paUSeaY5peIqNOSvMBMTXu2UsC+LgAWW9RKwkU2H7LiE/GSEYycYDQsuhiRBBUhe15dJJc
BlmOCJIA9nC7rr2VPSOp+YC8dL4xU9SPoyiG5DXXmsktT8GwSDnneW0Wurt6mkvxW7IHnpajm+yu
N4wa1DS0k1WJdhvjzG/lIqfIIjYLfwagvQt59xuBgvsX9U1vTQWTsPtrK2nzW7Wg3wS0J2wOJh9R
NFvi8cAZL/MyVmF9IDoxHYISdv6FMyqjqDCyis9dl/HwiCzR3cNEV0qxMCBB9CbQABQEYW2YKNWc
0KKm4EFmJpPa/SAeb86475KR01c+sfWf+agmJ8ZaTy2nBjKsT54FMLsgimeU0H/UMrFeHz2IdF0a
naRYdX1umlLaRO1Gt1r7wyLNsFKtByqJvsHQvifVvH2ibKMAYvAw7d5yJhNutByoQf7HCVvm81qr
7LTtQ0LYKUXZiczH643A/k0kqKrUv4d3Wl0cNoEPpuaIPcoLC1DYXM+h8p9q87vw6ohjgfrVB5pf
KwC8VqUwQREYfVsEB+vRXXA0xjVFfW0/X8WHUAbqpgr1AO/0CgagDnDNmUSqcFQ1eYCrSkB0viZs
nAZ7FurVD3Mzt/V/xAoR79jq/7XYe9eilGc0afboIqu3FIpXiAvx6TOqDI/nuCWIANXhfth1+j0F
FLb9a99lm9IHkXSSjFEydpUt5xUCWYLFyMP2gL/txFQQIUPPs5c255tVlL5FYYzslpyh8EJ13veR
i84feVJw3ezIa8epuiFJ5XioM4e+KnpcEIg1UUQsf+XmjjDjBXGkDX4ipobkK4O8i2F419d+znXx
kenyZTANpvTXO9wdynFnzlLUE0y3L2+DZCU4SDTeyqB1SZMLt3QtP2+PpxcdTZjBGg1ySoG3hSEx
JjwJbBX0u7cilGDLDZlnyZe8zx1kdjH8lkJfLVxe3FixcnCWwH4G0NrcMg8pcg80x6ZELSOY/FEX
h5achcsZrpnq2DvNfDg+Egrp21Z0xpvAADJrOQ3Njw5HdtmZ7VLNjzt2TbjyilKGA4E/uHg9kClZ
DgGTzlvlcMs+K60P7KtaL5mVa8vH6CECEodVYVBC0ziNCj81FezEuyrgp1JdDde+Xt26llkBLMaJ
8J82LgAgV7jXw5amjgr1zTm/OcO4XwiicwhXjUt7JJ5jJgM0Tk4GxjVY9NWLrrJ3cL/TjT3sUHAq
gQ/bzfdsF+vUs7w1WpfTC3QV8t+Bi9HwaK6ZpOIq2t6hgYedVjNEjNMw+OlOV8gZzMSLVFNlZo3x
5ticNhduzlyDN+d0vbTJbEmNixIkdrbgvbuAOZnorSQK3/RMHOSGh+OOsfdqBPvoDEBX7sdcbCvQ
6hxpyX7LUx6MtLYvuNAfNZz7xdccBhHPwZtTHCVCs0voWzp+nKOor8d8cz291J+eCmuPX68VFz5C
EmOfTd+PYBzQB605314JeYKuGITMlwgp7DSyGeWb7DK+yr8lNslbdRNDFDi5VXaacSwYkEPdjagt
6KG2iTucPnslEAuC9Y+PCughIb/57ibIXk2BNwUtbHb0vw5CSWCTPp/5rJeFzmhlgOvyTT33rT/B
35iVdz/bZ6mbaXsuQnj/GXtwg6QdAhIzBUYZ66QQXdH/ggsiJS3WdU5lVV2WT00u+g/p/++mqM+i
I4553Au77WW6mlKgGOdZPlvTfF1BZXFoa1yHKWJoIAOLn4r/9xYxkW5fRMePgMNq6Gs1zkWru43k
HsQY9kEKmljbL60P1veI5HjsZL48MoCxirtczbIt1/CkwZS/CDEJoo73rwNTefN/RSwcTR2qbfoJ
9t2N2oOgn/rlXGjq6tHV5D7pwe7X7zNM4JTH/0T+IZwUMBDTaLXpJIbuvm3TvdMA4OcoDbybi6KX
AoouezW3aYgcOlcm3f+P1ucg68LPOJE6qM3mh8Yd3tv8FeJ/rVteQROIeQlkGvKhAGSS0QF+XcMf
l5b1/cnLVA7RD6Wu8El/B6/guDZKqwEtb2sr+Dg8HOY5XDnU919s0jKpdejUaasezE3FQXBTlDhY
iEs4LmCSR1W4Xun0HdHaxHAZptM8Uc6p/CmhzAyUH8usMgcnSBtY9mhkv+nkgfJ11OtHdSfjYzU8
1t6VqeJxprVR0t/j3RaQPDKUqidXGocvLJ4ludG50kO6n0Z0lMT6FJ7/4Ab5tmpY59S3XPRx7deC
m4UwAdCvFO7pOLnomWCia+Ng1ErUulV07HxizTN18Pw7I/EzA04M45QuOFZtBWfI/QwEhhYxEB5E
jVy9dxInY24Dw31T3KAKaD1DvyhTTUMJfsFIAMXMRkMwAmw8iOd0A2uF4lE6l3U7FRZiPtwMkgA4
BvY1t/fgJ4qZIxwVGTWKAFNxj22ZE5cHeaG5DALiIYpiW3BaPyJBzCt4TRsx/bQP3/nYm/sm9xnC
eZob6RMeodqe9hUex+FdKLOru3NfbT7GeQc4NrIeLj4e8fElD9cznDFSd1h2Rr6p60+SNsORaBQP
KqyrdJG0Q4i8GDLKLdpSFzh1K5f/edM9Gyk3JkCBKS6aYLrK1oM1h9DfEhQ+pLUPOqcTYgInGnJM
0sLCJOz8Hy8HYgXmTBpqyctMg8tbeZigZjYh+fGgKtiNZtfoX+tNWayE5fcVVfz85EeCRRNQ83pM
YTgKvWgBW+DTfvyN7FD5vT1epD55o2tUKAK85ajko0o+mbge2YJHeBzzTMjbELelT94IeK+fqBKw
3lMn5YBvCgd/i58dDmqgFyLS5CYq1SLOSv8C0uy8T77ROrHchLH4HB12l1WekPf/scGovIILWusF
MpaC9oCL+yFo6ZOepS9k9m/p44/D+IVBcnZxl74a+Q8AYGiN/ipfbOV74/pRU3P2E68UNFtPUSbT
FHhiOMdKU8xL15bREr1f5Bq9cawXJmmP+Eh99cT5AqmkQBxrfF0O3imeMo9TK7iM+EBuIzS5TJ+L
XiLW3z1fE4LQEZbiKaY50PlAoSl9RWhGbSD5EUubJdobC+r9n4JyrRlxbHMMqUQ63+QOWOrVes09
i9GZY3gi8bG7kR9seSQDkq280q2lhmIoDH1DOtGKI9DaSl8jeInMzbu9vgHSdb/GuK3EQTKeMk1d
K4TfkcwL3vpcoIVK1csMF8SPoPaY5ZoGd7fpcZhTJX7mDvXAaVecaFV42PpHr5723IfaahqEjtqz
uP7N2fCpVFa3Ur6eInS9GIoUnKYCLm8TfIBYQJu5MhL7787GRXEYxcTbvrILNhfRaCPtVmsusf0w
4jxnQiPdyGz6IRQLSVf9T+kFWMLSCaZXW1rj+LiAv7rES4nwCIhZZIgQM/BuUznng6zCUhOCwREu
PdbWZ8cHIPK+xadWrvROClPK9j7erSWFokqGcZ0KNFcKdgK5Rd+Ke5jsllL/KA739wuFbtAhNCvI
3uWIj/0HTQFN3kj50Y/zoY1f5Zu/5EmzZ8Sjo4hwG57NLljRr30FP/FGVl9q5m1z4HHDPSScyNJD
n3mzPLgV8YcC4jCgWgv9LjXBgFRn5OuM9CO/YGf2nUVyb3RD3YiEJ5VpMfZ4nGNCQg7ZntFcvZYP
/uiZuuXgdFwj2hYrN0nvN9PeWftn3c5mMfThhRfrM5Aolmq9ismvzvXS3sAG2yAhMEgN5R8BqCl3
xz/3LaV9c4tp6ZeJ3D3OQBT6b1K1pRJHuVK8Gb1KI0GxD5TI2cyuPVYJgAoW3BXVxzeRYnxl4Fon
iPAovlxf7TJ2d1yvd/MvElCiDNrzluCmI5FytKXRWa6g06vcVFt9lC/HScl/bTX694k1PTJCmqH6
s7X0xqfcQYlftL4guYad3ZbIbGMourOCZkmQQ+2/QyxTCG1wNCkRfF5BSXXsywlLyJCnQnR3teB5
K1oXe6bxRZIJHhr2DjCFNkLDV0l7hQXukl6RschNgphz4Y9wqjOPecS2X+itpEzKwtHqQ2ee1hgN
Ov2/wCc+wkBtWl5c0BWd813p4qaPLCGr+QOxqZYisJ3xz5qHZymcMP5k5A1tmiAr40yGFlX1BXLu
qCibYf9+RONwyanhtdH8iMC5hpmvuk2c5h49cwhvxTw0mEgynx461QzgzSL89j1uXFrtxHW3Jqzk
/Vrd1cm5TupUPqRkIazf1whZxk574bMkZSUYoBd0TYQAJZFPRvIGsNbdhqjoOT9ystQghz8SikLQ
zEW1/ccHGLydTphaf5FcTUKRH1l91J3KV2VJKSs+/D71+Hm6U0uCQyT5CGgY/JxJHkwHc7QMnLeo
wq0Wony54cx+cSd8jZBMIJ1g3IyOshtokfEZ6nEUjqrIsFDAaQ5oeciVpRzOFhKeXUsn2TV/4wcz
eD1FXT6u4RtHwtrR0PZOhoHsx3hB0igekvp9pSqEtCZt8h7ofv0A3BnTgNcPDowEurLc8JR6lRaF
zUiK+u+uHO41PI9632P7Jx+Merb6bWRJu3zBP8JCIYfar2sf1f6VAwICevDn+mhyc4pvdkSA+fZW
8zwFZhv+fqF6aLJQKLLQFQZ5/mKp71WHQYbE69EYPgO8HP/iHp4it7N+X9PXQq0Lqg7W2/ikXXGl
JaKJDy7HjI7Fx4d5Dcdkf5QXuMoOzb+B4cRExyJxOkrWrI2SaGpiBBIvZDyMZLaoI2eYL9bSX4Fa
70MmF+A271S+BuM1RINCaH6g8wXOjJ+wRkhw62HW5Nw1tI7Tc8NAGFUuKYeTYCx7HfrTMlTHQbGU
achfjI3lQJSrGcXPy+gRsYDTbQxTIMRTtB5EDsOXaJBf9it6H4su+hjVBA+G7lCYKplNE7UgvghQ
KmUkLf/Hi7D3Dhpg3mi8FYgAhQ+RWUD+BoaHnOigolUxuz8UGSRx1ldak0KnvWAS/Pk4ojyW0KxQ
j7r+xDhgccVgE9WxvHpeyLbHSgmUwC+3QE6l4yMLqOyWh+byaTfDIlv0L956vW0+I3eXr3sUBQrx
VBBLA31t98j66Mb1HnIunx4S1Ma9yLD8ch4qWpICnoNA4InSPvIb6WtFiAo7WbuUyvdUa/EPskCY
KfKma5+QbAyItTvkQYWFsHtxqqQQqGgiyk1dhIygmNPqrWZSOKV328tS8G9hG5vwoPOdGBkTA4zP
2dQNa4R+DavoPzSRITRVPoIAbKIKBoEv6wY0GYK/tN4ziImdiqcKrgnlLuM/t6bSihb7z+xT78TD
9+hWUklval2hvHDtsOn7docWdUwhi3HkY9222Kp/7VK16DrTo5qWDyuNkjwDCmwjOYU0YklOLQkz
PUuA4beNQ95HhsCR/UJsPowKBlYWy7leGwxG3nHMxZdOLWma4VvpwN3Rdy6p5swdSVx0BK/HXtQP
wGoOVN4FnAckeFfoft0+fFk0u3lpO2TPWDkr99jIF15f/JvD3IcbKtOmqTZk7Zigst/vuP6sYyLt
9x5UInscUHhLfw++wzW6b376AxTdl/3kYlNKszpQJ4fKVjV1uhVE3XMUk0KxqTa7NXcOMb7N9r5R
BSEqqpTe4MG5NDOH8lSKoPL6cur4qUkecEztsFxtM9J5KPQyVRM1HJrkMEU3rhCtQvQRCgMxs5bx
beKyLcjjA6rYe+zcCRWEwuMF56xItgDTFj3N/KLPhLTskS8P1qqal9UIynqOsOkqqhL44cHcNo83
RIEgSoNEteSjNwUn6/T/lIyT80O800VzMdEWjFRRhW4dG62aRB7PwF5FiPBugycRV5U1LtBx8s3Z
hqvBMtekw/dwLXcmE28nw/3oMRIUZa0bjK13cCtfcTaWy1xuWVROHyt0KLLoq6p0Pw1huNWPYLhy
7fhYjvZWJw4hW/wfzFroBYk0x8H/wHVQVcyloMPEpB4QLklslAJB7JczfdaEUiySgW/3EXPZAJw+
9hqPWEwrZMBHDMWfJjt2U/JRq2535TvBYXG8OeErr6B6TvzdmBe2jNHyvJTqzbWhU+rOoorvJu03
EHj2h0+x3bEkx9vLJWrtAsLiARXssKO0i5yNQVUvJAOJyoZzI2mlgkz6ZP44tn3cr1HflR5hEgep
fsOewD/L6+2uPBHf2fNFKZh2a/Xaeu+ks248XBtwiQG3mgYtS/ODV/SUx2tS+uTNmhX2mMlOSJk+
tV2OkcPFzKq8anCeQpazr/9RCZkplhJ4kIhSPpNUHIdzn3VPoT0XlQjnZQoUjwqqRmzAMkSa+gRT
9K2VHV5HvWI6xFvFRCEwakD2tW5V4AxGFhsNnHWJlUFSAvDK+ngRLkh3fGLdpvbSZiL0li/Y01kE
zkTT5szNRnQt/DPbTkJHqGNAMoJ3Aa/rjPXlZHQveh1Qp/TMo2SIxpwm+Zcjez5unvnKtneDzyM/
PkPV+HTL/HdUm+FAp3v7w3DVkNbBGWQJVomPiG+pbe4EMpTh9ZppuZfi3vxXnVjBu6JntdVn/i5s
lJej7K5NWwql66V0maw8sXwjMG2U4nJL7ejzckiJJiltefdhV4xrc3sKQe/hAFnfIuYhX0rnli5p
SBofpLvJzy2j5CIRn+GG0I5Ede3uoPK7or8tbR7wOW1ILpWHSN4k8xh13CxlNRl6nEEO+uVHvWX0
kXFuU8xwO+d4pibLlGwddcqKN0NkDEhyTRCQ3eomTirjmZTyxXZfs90LszuhsSLJjVVZjOpgSHuq
jRlDulYb/pF2XTXGQR2b2m5P5ERkaJMBy8fWsu3k34IoWy1GSa422siGLyTHMIwfe4BDXPOCX2xT
UMTgW1/ngETs3CyY1zhqkMH2Q58nbO4EB2PzHRqQcUH5iG5/Cwlq1Sf2sSfzLiPIg0ywIvW9DIqm
opG16Rho1705VRaOV/39cnZ37lgu8vOnlj0YxsPxNdRWQZrXfWtsby2/8KelkB4JGgJc7TLdm+7e
6klrKba3zK+ZJ3IumiDapvznXUTFZCLICdBy/uKTfCSkwnC63GEyvFtSL6E8nweIz5hqGEeMyKrh
Kc+OL3CnB6hfCpWxJAkTwOf15BHIRLo8oNiXa05hFQ7pdLiVpAWXl7d4jk/0I1EDYseXdBpHginV
/yu49UN+Wv05W/G8Ll8OetftHgoxmpItjrCjgPGzeioq73JDasuGw5tWlW/V/62DEV4EoOXPIrmv
/zezFBhP8a6CcjZowN/lBt9c8g1Ww9MUx7txthtKjey+vzCIUAbo6z1LNxuU0e1MRkQWrpMmCnuE
coqZ4VZvdNZ6dqDhBOYdEobqy27kFuFaHTCu7s7PwP4j6eRKmxuShd61ofl5Yr3Gq5aPshmCZTuB
5ELl3fNobBEzJ7WM2LVaDmFu8ukVPee3XvQmcDfTu3GmTYnvPuSZilmLVKZZ0LpZG/eYJ6s/WEuH
ti0/wK24Iz/XQkYJOMOy7dPozgioK9ZI0yPTUVNuXPdRbftUJ7RutxTOSRzNWKvUyhcBWAa8s9Sa
Wb9D2Jfps983bqBqGHW8xVsN6TuamJzoI7FuAjtU7flt39FSV3DTzYrMJsHaXpyskMuafUw++0gE
vmosiyyl/XhKmzUkCV9/ffEmRAmOIG8SclwFNimzkXKJ4kzB6MOMBk9Fgc6QsHIK55unPfsgM6ZB
EntLAe5EP/JZm5s0FoSl3LZj3iKqQMSVF+UoHGN2soKX2vUUyKRQp6AH0/VC9RMuEhc6Vm+OJ7kQ
8QSUv+PSASzhj9FCoIIyqBFHut04q/sx44f3B58Y+2wBMkMZh/EobFtc0b6OqA1ozCzipdRg/AaW
K3+m1jbme7fSbt7MKd60/k10tzu3Gqq+7SN+6DvT/7qmrXn77OkXwQx4lb/ZmS1fVNoUi34oTuzB
aJpsixMltS5Cvg9Bzn3tJStpMq4Jo1Rrcd8eOwgnk9Ydo9onE2DcUhKPWN/X5O9vFvoRCJHeRNCu
lUW9Gp00t7fs46xN6a31BS//y8tbnkLTL9rFMH2Z0+/wLiUSACEC9acHTuxUgM6+mb2TYRyobkMC
IJVNdyLC0yUn1XbSuoVR3DiMyP+MHyAY6Dd1TJul/tBsMx4B1NTfeVw5pMbZYKHmFzxaFbdTTkY0
uN3UJOz96BrLwDoku3uUbnjdqs7F5fdahB9HwSF29FbwV1jeCTNunGuNraPEVMoKpW+HOqVVPdgC
r3gGRy+HeI+be4r02QFvi6jUpejb9mhM3VIeey2hCRegMwz8TyP/L3y3IvWgBtX5pkj4Qw1E6GuS
zb3fR66FbvWrXDDxKy3XwWujQm/kktjK9hN05OWJSXtYrbhFhw6HPsFGr+wEPd4mSJ7+rECrNJsu
Hyjm10y7yikecRKTbmZSAxURRH3B+LmVABedoHthh66CWGv0duZv9zaKxSR/W1FZFNdysfvT5MbZ
7KzNojEhQu9/1DdoLTVohxwwnvkyDv02LFQETC1COQMRjw5bDF7ocoZxn10/q7CTX2gt9ptVx6uo
q6PCsyLmij/X4PYXOAoP1wf79+xNqSH0GmPA6cOhXaElCXNlEn4XaqEG/pADsfUeYw+GskqBDALZ
OHHFQs6fVGy25R1Wap0cUkndH20gDUtNThUR7kLVSETtPzjB3bgVrV1efwRGVVtBbgyU9zO5oVYR
M54dI/vUAD/ZTNGvI+dt2oeofRM5qIUBaMeQGFcqBCj7mSPSZl1/+BlOIECoEmYmHFNvDBvJb/nW
3CMgezjTgDO8frJw3v37sQ0iiiFIekwcV81MfITq8Fv98tmAd8fMaJo78QNpDCqMTDsaBFxiACgA
zvup11+WSIsPfKhjgK3qyc9vsnKwlOY0f2BhbYYqFd2g5zqMZ05TjMu2LV7lGW21ydH1KkKJVxyA
8nKK9waO+Ivyf3GGoE+IupPfg6hjqE5pGCd5iiQ1QcrAy1nTwMAF1S1wjc01zkgI3g1pKj3qe/Sr
q8DV9kcsEQINEqRH+6WTJYOsFJkIhfDhKF/D/ElwF4pIR6VyE6AvnBJvlCHfj0tibTh7IvYiJGWw
RUcRM5Rc3dTnamQeX8MX3PAT8QvkgZ4X2s4jC52vI9Rdma18tsQUWOum8mTHP90/xVO2DwRcSCqX
2ZyVV5ycnJzDAtjOvKaKN08efla2te/BfGHoXCYGQrajmr5LAsxedYJUHdCD2RsQ47bNtzh7vFIx
sY9yXmhHAAQfSOiwds6NVS+CL16CF24RuQ2fVvhHTzx2SHhWSYhiBM5vTKN0xd9YZAwfR4ZkyJzD
pdhOYisouQYTmFuwyJg3S9zAeQZ4fbQB//YxqHRZUJ2LdJLOGaM+YH8070iNRpUaKOGZ4F9LSkXM
6oxYbe+TQJzuB3Oi+eoJgyUn5726vK+7XxzReMYxsICMi8Xr13j16OZh3zujMhVOPcN9gtlv+QO9
5xD8viEjdCANHygGh6KSNw4woGASE8J5rnRJ28nnRlm/Rg01nCIMK+R1MyKgubelBMc3y89vjZTj
D3F6PUVTxx9D8iAmR5YEGL0+9WR8iwkUDObHtQEWiAS2jeBCx0/p95lfM1Q38UkCjQx5W+nRGlS/
bfpuSEkN2fp7IAoRnXdIQvV16SpLbi+WRN+w6uFM+JtRpLHclBL9PBIMbqM3MYCzjMWH3soT+8h+
u2QfLozkkNsJ/xbjNJn9YjWTumFBgiuOH5EggvJb3qRwayHWNidT6FeFuxsYwg2F1pSAs88LOKwc
+B/gAHPNH5NofaD+gmI+uQj75ya3X3rDG2qSvqibdRs8bCBHuHD4WiItlcfxXQWJkn4oYwhffrq3
kbNvJ0w9USmQ6u2BiyWd51ElQunUod18HzPimX1EtVSNncmy7CAQ48o9Z1RZ5UciI1yGgklyPks8
WcHLaZmI62x0VM0ZZ03gl2DCZVK8SM88Jv4b9wqseBaJnqflQgLl1rzsDXXuS4Z+1QVwOVr/ysxR
7Ftn8fyqfd7CoZLSuv6Ij1F3nLxiXSCvjj+8AYrN32oss6Vf/YMtIEeu0yMEabtRKs3l6ZhpUkWe
ktcN4Jn8YyJrfzlFfaFS852ztoVnN8tMbMHP8Bw4DxnbYSTh58ysUvAJATxYy2QUnDcjUIZaULGG
kD8ngT0oyVJtgcIQU9EPZLP5GtEjDX6qGxIU7i41OyT6cuP7OMufhRFpSYiJ0I2VoSUMthKRFj+z
HRktqhG8DKsmpA49x5pAwkI4Ylafrblk52PqTzbvtj7Ou7rtHkC8nY149WzazF05keqya2ri5hSJ
WwWbI7IgEuaEVGdMJo1Y+u4FP17vhYsh75bZvfS2dP410mMjHDsvRGeWgToau7JiLYSUizS32JQX
lI0J3fBO6mridxuWZoF8PGWJ9x7n/t+Xu3CQ3nKuzOfDi6gzwfX1YxDOGkfvTTpzYHPSPW1Pa1Ma
Ui/GHogO8aLCWsGHlGCeY1zRnkGZ1h8wlvv5bCOAWh/FxP1HxIinXoieM0BIomCZEXLyY8AmUJWE
FVuw5ulP5mGPr8IZCzxT4nQ1NSmumdsOGhd5/bkG/LgtreypsqvT4FbDHAnRVnAebpwCkPrXvLmO
+QlKEka20KqSBCS8ZrbXXzraTnDuvomXylgq6SphiQpx1F12GDOyWcWFDc/uLoXIYEnvIVlJ9i0p
b9iYi7WQfZLn0/BJh5a1s1Ly27Qg8axcilVRxXjEiaV1wx0nsvQH4PVYaHwsRx7Gm/QuoLJ5kkWY
W1wAF3PaUCRXsImFat18Et6jmAK1qs+s/VR3TKo3h0X7ji97eWgel3FCyKWzG+yU60bp8Ip/UC31
TkGp+dPzoVFHPfegyJgDd8XnRChzV+9WdfLcw07cua5jmFqLFEj/QuNpZHWUbWfH9eD4zpJ+oXZY
yTmu7MOK3co1HBiq8E5HdfNVO4nLFfz4L/V501AxcCMp+4OGEMhqMFu4zbCvGtRALeVxWWh5PJOZ
bxjOUjGXWmyxv5wQooiJSfaI6qjZPVKp6DPv2r3nlhck8rh0XyIamueLCfM2TgCvQUhR1436+TiP
xcfIa7/2QAKF3OLyDteQGc4s2QhC3H9WWkYD7epiNKAFjc5jpr7VapFnEwa7pWHA7wmOs2oTT9Sk
qDIaGZow43Eyam2e9rjfSm8bMfIHuf+fCgNaZVLIGlvqKqCJV9O02OBIqwJe+OgYNNgIvkboVtI9
6LixhtPx4q7wN1Osv80Rd/MjgD2QnP3rEhU5qLZsOogQNXUoUWEoLhnLIJpnEegP12rI5UKhXT0t
EDgZI8XBY6A7mLwhedvHfYxOs0M+M9kfGMqyHsg/7thlgzSnN1v6tK+tMPJpb7ImiVxDeAGIwGZE
W/VL6zyaisNIUrw7aHZItE3mxxO/R97Y52youoWZLTtXz5u4ARCT+X+MoCoOZmg/GcvpW7aJgWa7
x6QyI2F2citdH95ykz6fXsQehiizJI7Qc4XmqN1Q/TMFisMv2qyRfbrxabIO30EXeBfUXaObQI3Y
p82tkn1gJgV3A8nHkUroz/jV8+x0y1b9/50Ms7uTP3iZ5/UZfADURTCPjE0kGt7S5bg2gS4CFt+i
U0aCvnTJllUowIyVXmUxtUUFERxp2pPMxq8vZQXUEFRe9d+YMYikNQsY0h8u7p+6TyQEPuAW8U/t
z8c+IVoW49iNveMrgVsp5DvHLpUHxO7QRcG954XjEltsO25nITd/nRADd5uDhIuW+9wgqRYNdNJS
xwFdmyze0IvR6UqI8EgRQcp2j95j8SS6PpG/nFPe+fnOn8CSp5TGe7F3+vYdupBjAFkCr/kHRj7p
/R0oe+U815WW+xxBXviff8l8v6Wn3gJU0IG1+VqnotPHWnPkKiIGuK9tza8CECJYKJVLrAKNxw7V
ba+prwD5aIcKWdLaKUM48ttg7Vi9YWUjpNc7nC14q6lUe15VkhUPYrMnGaIB2BEe2RPpM+3pQswA
FsgSPrCGJLqB+3KOhxRZof5x5vga5TKp0WjcZ0TQpscyR2/PO+EmObfidZwgzEeySU6Qibr2O1LP
C/fK7rZY9iEDGOaRePMeDF5AsNuHphaGKD38dWx5dFnJPKhNWIzdX7XeOfub1pUuYXJA8RHcVS3/
VW/KkOFB4GNeIgxqyV4E+/NDmm/Ic7V31cKbg0F/XNkzcBCabMvE4LRLKtuIaDWoPsNG9Dw0PDcJ
6aTnzo4WMYpUa9ZMtKrM5cdnJfE0XQEgjVSzl2BCaMO8Ze9qvPfyhLaj9t2rkLjdilTtMf6laHPf
ThB/miOvI+pCacdw8/qxCzINo9IHd8WX9TLY5UPctUVhM7qLpPWIB65tReCnjfAtLPnEgvt0BfzH
d5qLbJJUFjO70G2S8ci9fhhZhxk7MG3CQyt1aLrnHB6qjTCq19eibuEGJeVGtpjUwlZOfCzoUezX
3j7WHn/jULReGS2HYtNCRdvZxAHBH+JSDNB93ew3GSxre4asz0DM5IJE8qzGkts/Zuk6GKfdtC2l
x2Pp5WnjIHql9wBXht9zvvzfCT31OcoIlo7Ys+fFoRSnraysU800DG/zj4jLcwm/B9oWXultdR2k
Uk1UzAjlQ5/m4WORKG36vpBCADwMAIAESQuycaeFQMGsrTdMKyrSAYBE/GpF5vStbRYfn9/bMfU9
OY+RBNXHMYY8Oh0YayW4o6UOCtefASlbozv7cbaD0auYX5UP35ee40udJRtmRkOcLJtDZshdsT/k
HHi4DFmATy+HdEYPdWwr6lzUBnoGKDLqhQ6usfaMY1i6jba9cCItrpg1t/xkoG9FFOLxkViSLHAU
Eq/iy1za08zsZPzNQe95pw/gIkvCXkq6WqSC/yyelkzCDhRSEH0m35uSePTpnHStlMX38DCpHMmc
4aX+Gaga0KmbRm9GPoMAxRg/Raldrq1rmUSTKQKsnGEDPlpp6P77y7qrR2d027oqJJMhw6LNWphv
Jm56QOCrbqq081iQt4c8KSG1cpnRaMAg0/AEuvSNfPsQVLF2nTeS3hbXAp0wY7HTH4r7VSYz2vID
3uKk00DTb5tQ72eTLlMev0H9nSoCEfK0z0wlicntBjvoqMKpXc8jgUfE2/+XPEj53PQSAOW3AQrx
5NJB7AeVfAOtZKC9LGKsbWE337Z7ifG56+/382v4O1Oad3bqXMMoAsMHRff9os9sBE1bgQAMTcQE
ZF8XnR6KxxlvTSby8gkTAzP6WoztU0rmnS8gpkYEzk80bJwHNKFYtKQwViIQiUgf/c4q8Y2MKEiF
p/BNdWv+eSdhFWeC5xoGtTLdWKT4681rIKBgTSumOD/QltuoDCv7CwXu84K8OnE26zHPZ5v45GL/
JQUGpFnl7mwdWL3Pf9A1/i426lRkUhuBM/U2cRdEN7u7smb3NZ+1f0Dv4r0z6mczzMCYesnTtMpO
CLl208vyx0XI1IeypHnEvxuzQ9csYi8eqneiI0/d8q2/2OPQMno/2dDlmKOSxaOMC0zDPKFzPkDV
mJDivCOCrfne6+37NbN4OaYhmcz7wm5VGAqzEls27aLFZQTMnMc2rl7+jF+hP80USwlSTnTakdjI
ca6H61/2zoJT2EGhD+hC4qeXJiTNLY24Ee6/D04c3p4PGnSoP/uSr9MSJKGHjlkEb9HuJhQNh7US
iWCIT78dzYugHII5kdQ1qPRFhBlRJi7ni4WFT9sq+QfSnzv9176uM8kz2KJ8TFjQFxZyPLP0te4H
8GVlA1cbHf+gEP7lsv8sY/1aTB8sSQ74EEKitJoWTFlIiWt6RfLyn17d2y3HSp26tQ9ygJl6prsb
cCotT1xBQmbKAks5tnHOdno5KGURYThaBxs53SFD/QpyHj/EaScsGwxGLi9gTppsMLwNwvxJWYbT
+bQbpo3ubZPFn6tWHBdAG3USlWQ5HGMic2J383joeksGtKDDk7Kupe8MSaQxy50pvzgFzM3GgoGv
bLfL70pH1cnvHEQwoZBIWumTU1wX5CWJRD1DbifffxCCv9KuMr5I3XQm6ePL+bqLahNWDwLww+p6
jZOl8DSpcDphfXE7DrNjwUMfZyxuVvUjjmuTqt5Fh/4K2DkcYMcPhwGkkCLVDepGLjcr9vuy7Jor
phGCj/BmKaPiynPAG8jApeBB48rrg6vjCSqtP4+MWTJNA/c3jGKkJWe1Ozk4TNB9SV/7osuQir7s
osDmHFDrKVdyVE84RWGSPz9V3ieHgb3tUvvUhf1jGqo4QF7FX5Ca5puDNwQD6VSfcjK5kJOYp7iE
FFniY9rK2VDDIlvtfSyOPps8Z2uv9MVqkcgCwOgyUcexhVKzNHBV5AqXGMSgIC/fHAQKHqMqwXf8
kWncWB/J+JMGfPgPXq1t1vybha0Jq10hMmoxTSAum6TpRe1q8bAuIW6Rk8LwoEVxnwOX/Hd1CAz6
Cxg6o2wbg6ytn37qfkBagBsaGQT2qwUrhzWqpE0p6pBMvFu4yKmIJczoqXOJX/ILlNbN5qQeQTAC
PKoomXJagRL5WOLdKnRIWom4SL8FtZ0KxwCZaiTwr8VxcOAg+s54rUgomGYwW3jlJMjTyGEcXNq4
Caf9buJHczm7Vov8K67LAok4YuTlR2tepF+/nlZpSm3vDNwhNSW3C0gjiNs4ezSLvyFkN0Y4mDNW
sKGDmCHczHdiK8FvjDurR919krNp6utOAQ42KajhPerNMK7QzT+rXEA/v/XFitjeC7Qq4MbhbgF7
lRgVP8mS44/jfaonO2hc0cM/TTr0jI3Z+nv4JTeNtc1v84ypi5ql9KtB1mKUXnxzviFvsVlJjDeN
37RUkJp1XfskFKIsOeLWxZZXcVF7UJ8bnVuVnUfH1s5SXexPUnRdbcK7qEbN7WsnX6wKM5JmuzyA
qxg8FYpL7rvgtnrOireD04o0jF9eb7j4MKsVbptzS5ccXGL6UWdAUouxi0kL9D4kO2Fe7Z9B0zHh
OgEemr0w5+n3/d12xBxNovzyPILUnRwf6nutKsNj1JOY9l0CHFycAP/KLo4qiJYF1aFelDgIXWWU
ZIh+ncLJX8X0C5FyRJtvGk65ie1n3tUAUjtTNZJbizADn3Rh0MSAG2cimvc+yZp/sE39m5049vFr
dv20kZtw38mAU9XEzSA/Oblpn1MyR+PYxodf3Ctq2hyTWNXv8h1bfvxO/nRUPTWnWcSeDMMgYNFb
wEJSAGvWnpjFBO9nLcau3qguQjedyUjN2o2q2KrEYr+i3NsGUuBic/IGmoX7DCPeblikRAf56hA4
nuaw1e2d+a2xxBjvkV05vhe3ufaNbFghgDZbPKvsBTQ67maDej4ihWx5Y69WYyFcz9s0WReCvo2h
LOIGaXAcz1YPxQ9GLrdx+yXvBJNGVjuXbD4QK0zgNHrUhjhwHuMKI6LTA7Ah31e1t1BvEvjxkdJ4
EZaxa8utprnXHjJfKVYdsHwNLkDmEfAnEf8hjaw9dgOxWIyEcsOVXzzpgZXaTOSBFRP3aPfWMjRy
ziYkr2AFtiXxf0KdY+pu6mOt4v/ellh/lHOlgraXDSrXjgsi1IbTm9uXuTYtE2mfB22+NOcwOmUw
S++wt+ypwRrFh6iCsRdVswhg/dab3xtu2SNZWvNfnfs7DnMoN6QzBGpLSwiOD68zBRbl/sNzJwSv
qkbTDzAp8KT0NMBbg2tuhyObQUyfxb+z0DBB4QriIeHM36zq/dL5n+cwzP79jtGs1+sZvvlU1P6c
c3N7KIxHV1hyYm8cXvVAUX6GZc2EhYRGkamNq0k/q7w8u6Y1q/1iA07q4rGpDr7YN7XgNS6a0CBj
MQ9S+RWfaeb4A/HR7p6qX+Qvu1LGfCtIVQOUhgOtMiH0CWVr0K/saLQ472sITeuJI/XrD/97T7RS
WDHOtTPd7FNwqaXPzvMk6O1h8z80kaZV72MREjeecDF6kARTcgn0PEKgy1VxPHoQgoaNl9FnP/Wh
mIAuCjll0vvZ+25KhsSFB2ycajouHBDdQJOLvLGtnEuVUGvXOY3fWvajoX//GBuXWN932qOaK9Ji
olQYCxdaiVVY/Itdvfr+2QvdKgpyCaoHKPTnDlZuEBTqigcsfsu30wol6qy9ysYALsDDAs7/i1eo
hjBG81guh2j0SAPlciitz92ia9YQVZiYQoqgU9VmoOJpi9XTvZhhCJLSpTQnia04r/ky50KPfPop
Z2nV3DXqx/ctT7ETg95sb5bAQiizBpAmgWYyrW38n5Tt18SGWGkA+Y9Oe+MMZo1NYQ0+6Cl0268K
q6uFDoEZX7hPHumEcd7f3t0oMzVwM7Dsqf/Ki72EkoS4iVmPAKKZfvT5oMGcvl8bTZxH2pvMOuz1
5Vdm4XrpcdKlvTvI3y6rmSpKGc4I3FpTsm+i1NoDMeGIhN/d/J04Tsz1UOG4/dwJ01MPKx6+W3pr
8/7ug8kJkeaHm0Rurs5bnLdG8YjF0v9nmQ3DulZxIukTvNehbGFBsdHYli5fxRn73UFbLjXndMFZ
rNTP7kK/nGQAIwehQIrr1bqTdsk+n7AYX089XPu+um2DhrN3QLutakTo3qiXcQIyAKydrkR+cS7f
9kNjkuxM0Mo/LoyE2TB9d7Iz8G7CGJOnMPOkGtYBFCr0EMI9aAg90j6neMmeXVPcbcPDgWAjifnj
90+EaJWv0vBkQiUZWJftuqLDtWXxu2usXnDSOIRx0UGAueze1M6dEVp3IRaqvo+pbMN6/Eej38OA
sYnMko2hrQ1VqKh5/ZE+cpguFjokmpVx2ymiFD2vTcsu8y5Ze+8AqoU97ovuxiExqtJXDFZAXoKz
9qMkHkl4prwE9pNw8SWmpK+WDS9pUBjLQ/Wddq1SwbrPrA4uAQ3tfuw0KCVUCMrS2fK0Th4pzXK7
HqPcfS0d4Hq8twA2gQknRRPFNUeXqY2pirDguNIqKW/sZZPy7qnn9BnqOA25kK3CFTQnuP61Vkeg
YoenebZuJxN2bZm9AYBtJt/Uy4RisQ+PSTYn+/g4uVcPtBXASGSra8QulBazEc+v+m6M7Xf2AhRh
Mnt2Co47mqv6228H1sJBd+xrdfJdJjxj60+qKK4vC6YYyCgcDNShbnhlXA37nplGhZtRDLUnKoPt
OC8OR7Pppd1CZ1nS0pdq7Z+8w4HvLpvV//S5MYVj/mGsC6DVUVmD0KxX1qLGlKPBUIP1m9RxjX4f
FQyHr/ABjB5O53+utwUGI2VAVo6cvxzqL1vmWHLM0WfamphLl6jkfK46WRUShyLnqBJZ7At2wV8L
KBMPINzx8WJ5GWCEFKIXyKjX+bUJBjUxV5jubXsP7N7S+yxYsQCBFb9Rn5QJgFuj4CzIDOtVukoH
MtmJ71fplnIwA1J7CgAGPDRpF86DNcEGY+zYel4eiZSzQsd7hKRR/DH0cLfW/aI5RRAX+1zQ6F06
AtIXGHkxIR2myi6hMd+rhVqg7bMvHfh8MH+J218pRQx4zcoYyxbxroB0a9MwKuu0nKl4dTyAr24Y
/fzZ6CEpX3iJVQbZyE59JmNkIXzT1xV4hBkLN88LY39zfQCMT7RPBaUaHhHWQYoxzBaG+skF3S/S
MajfCT5m8H8GgvZSkHamHtKzmDHkta8dpkk341cIYa/ZL4zyVJieyyrBjfDCtmZMg+ps8IaMFlD/
jB1kSmepKph9Q9IQW1K+PbPgWzlc2U/JPRw5wMHNN3x24B2fluFnzc5EZbKNvyb4xN/OnPy3HxhM
XMT+l6sQAfUJHtAfh4DZakXWBY2mV5EaEWqs0ujodaoP+fWeQ7K+EGJA3aoRUImueOyHQINwD/rA
LYH89obnNSTi3FNXnhtaKRWxh5oIgvXnSXEfB9Lhk18A7PNb+IZEmMq9su96nFTia8y/JGGE6k+U
Pd3nYyThxrQarkAQvY7ql23tUd+u3zPVyaHUzSJzvSBBFexLJlTAg9DvEQ9mQKByf1++ZH3vvB8q
2HC8EHPfGtx0s2sshnJ1xoTDdFckfH3awtiQV9ahbhRg5Kh0mhJjRX/k0tCpLdlONYishyghbIiK
L50D+omcnWoGOn6t8H7+p2b7qPnNzJV1rcr/+IeLEl9s0VeS1wY8DJKOhB/n2LCrQpXOGjbNRzH9
Z9a/iZCFVHsqroTj7Z6AckMj7WXeP8/wqRvk9TlnrEXSHN+g89WucPaEZfetYS0hbDYfNiNTFyJX
WaVKzZwS7wureu6x2YLER6x+Ej0V6IG08joFTXnGxGGJ7vw9dejPSaSWP0q8nYiJTpqbQj50ZKeC
iLC3teoqNeUC3MgqS7PueE8EWJbnihwqv/ydDKho4duLCsngoNx/aYcM81DEhWa8oJg6VRO6BANq
IJLFtxX4JCjpfts7ZnpIzneYiZbLqqio3o5DQjh113fI194pCU7DzG8mXuJPW8cCmsCAtHonihQq
2q+7x2UGLLPCdLitEOGA0AbzonDotSEPnXE9KVOx4AhXngX8uBkF+GYNm+7hhQtPsHQlhPv7Nt4S
jpjXlDGKpvpd1wDy1d68dp6WMtTP5ZNevFl59f5fjeSTpv3nFv8pPb+uGufvUanwFHxmqCb/ZPgs
WwqdxHEmmFsGAgfOAnWGnfRaQ2TSLjhSZtXxHJO4RvISPJ41XPRrfpHrABmXIW5tNWnqMNyVLZcK
HXbHyWupy1SU0/XxHbCM7GempivKkUn42OR530UT++H/nOKJWxCJnZ+N8YJutq9Ohc9CkI2bBLK9
H7bDxcf5YpUG7jhUKHMbRevvQyszMKD9sxmdA9wGSkSSqdK0kJD7E9ikQatElxc9knzR8Gj1LU3o
cqruzgq8h+XbpOwv0ZbKlY+Fk4O0Z/lSsrRMJoooFfhwyHqT66ky5l5DnNMfR5mbOM1ezGrXdDG3
qM8iaCaEDOQQ8FJ1DOYxBAM+wQrsWM1ePRbt2rO2dx/coELDNS5H1sUqXzuAkgSZtcNoJz4OgcMT
dvjppb26kDIi4BxLd8u02jGiacPwPpBBYbfdrP6S7oRGAsLm2BY0QuVCT5CqkA9kKs1MxZCdPhr+
hkosus1FPx56VMMIqva26xNzpaF1YnO+CWXCib5ARIBt9CILpJhE0zZ/Qn6Zpf3WOzAfFwk33LSH
P0I6YkN8OT8Rl+a34iYtqCr3N8Tw7NwzVshTQeyENWkHzYon3c9pjs81eSvrwgJQyUBpFXQA4Icd
Vvd6BuJpXfHCyFK36kv0sijxEX5YEgXiePyrej/oZttm0aepbQPkPTUxQxx8G231vHZCbyJkTBum
Oq+xXBWM/u7GH0rfWeUl6gKsEPVrNuXG2havfoDkUC2LZKWDBjgQO/anCQDfzE2G/kiIpNGxWEJh
8KJPk2wVM79eVqYJJXkALaAjMkyTmMrjNDhDIMGT5Jpq4F40oiH/Yqwemh9r0N3/6673CJDnBSK5
ns+laJy7l0sxVsiW183ZpUrr7GptEq/i+7XR2+UaJdCoZ6MtSM1yRZaEOGCRwpXKLU6UDiqGt/5h
8CgJFqyD2XnTAmE7zlbm1gVyekegaJHipCdr1O4eJGVczdXKsAFZHBKgYXIV/LDPTSiiu/ZXvB/Z
ZlMxxWIIICk+XRY9+nAtcEoxLBlk+kf3jfoCNeM78gm3CBqfW2WMXMpV9yE1DtYYlpJ7PT9qSMVO
mq6/PuqPE8ASp2hhfbxG97/hw99fFe72p/JJOtypqCJZidPZJeSiZgaWT8t/icd/YdvvtJjDhZJe
mG94lyCDUJe71kk5wNAe/RjnfqH2UhlTeT2tdz0vMvXKbi49fhBVDsawIAtN+bGZtYpP9hdYQ0lL
jv65aqEdDEUndqHT1TCs1Og5HEOrMtjIxCTNon7ZQucbhYdC3+el4zRVG8/yp1YPByOm0RvUTaPg
da21S+C6ZXr5XGqJTzd4sUVdXeIusEbVDOr+5M0v0AhYcIYdx8N2RuLjTWjrB/eNYImh3nk02xEC
bN5o7lKUNGOrMJeeXMwfH8sUNUsg4ElfPpjUDG8aiQxdokqCosWcshT2nbSfBcjSeSJY7nEegReB
e2MKoudCBqgyFGn5BbIRSsHSzW+gBBn49dHMtjUhsvrRZnBbS04lech7uENpF1vnmQ4t3FRKVv02
mmg8X9WvVqUjAjndveYTPc8j2bjUrHJr8IYuH8e3Ay87keKlDFQg8+CkXhLvUGuwkBrdO8SNbFP+
T3x+dVY2eWa4Rz969uoPCRDD9qk62MtC6szuLs+q/bhvYHzqQGvrE+aj2OqrEcHtrRPxTfKuGxTB
nzBmGXyjYFu1fGhMANmtBGvgXvhIJBBGCN9QiixmNeQME8YjBkITR+Y37l5wPsWbqz9soIPlXQJ+
slqCM13MwmWh48dxet5PThV9dAlbaQ65akltc7Ekc/pE/3hqmh4ZyWKsEY/lIb8iRlyev5RuOORh
TY3LMg5XjQmdO0vBgdI9btzRXUnBlPC8bdsSkEzzjGrHnepJv6xQz3r4Q+AyxGG+Pj+DolTZpfrx
FDcqzvJaP+2Epto7QIRtG+BQFPJj+cT6FuGgH/SyTv9ov/jA/M2qoLT1XH2ntj02vOYkgyk8y0Ot
OAsZ8j2PzTHfd9gaJHex7NjfsTNVQ0yfwzlWSmX3YTga2b+RwsFB8encXhOppQZib9Ird9fwrame
GNjFY7UeOsnttaDJA4TQnHfzjqvZY5oclbpd0YN2uheFrulAinV1AgED9n0NK4S1OPw1aVRVutWR
I8IZsDPvz8xEVn7fiL/EIiG+QgAMuwPHHqAMMz8UHkWLcuPt1ZDqMALwFkbNCuH3M5aKN0bdJtLp
xDYSChlHTA1K3BsKKEIeucsm3sEBar8fDkjH5qzYy1Rs3yow554wlrEzH5l6X4pBevvLMrhlTu0L
V+OG7z/Q7caBIY41Q8K0VYCaLH+cNCF81xLjbpWaQkA5QXNxHWuP7OLRmqzxGkLs99nU63HW2aOs
t5Fiqnyw5fk9qi7CzfV1wu4ejknDkPh6f3laB+HQXkF6yj1RSF5O94l7FsaUz9eLcEN+OlpX6KBL
8Iu1U7ThayhSgiryAeqLiPCoY+fcAXXMwRxM5WqXvobTGve1eba//zlhlta1CAOei79XZ0r9Fimg
J7grOhwyRNvc7xcE97/ULcW/m7+hy776Bwa+/xQiK6FhWqDgwZhFcHdsUjkFyqKkO2VR61gk+FOX
SySf+N3/YTlEOv5gApKvmwRJYzjRHbXswbNaKq8LWGBDT7LbBB8GUOfjiISRbZr6Y26bhBnhfYB+
Tky1N9POXu9AYGdcVmwdwoIklDvkNCVCIzO9Q/h1cgGNH8unraJOnj9S+vvtCTrYm4/7B1SZC9mr
rhSjgs+DIlxLVhpD9qfGuFl5IFX/60PHvY3QxImEXfNlG2aVPz1FhIbFxoUJvQu45xP8rcnwiO4o
UiZlzvELMVsnREleC6Op1qli/BY8m8dmdj01tR5WPtV82hxlIA/f2lEry2K8prHNDdBpdSZ+9wGb
jaisekwDtjdGERhvHho3m5J47ibKSjIBbbLNVGXPzRUEE98Nn4BjZVe9sxzl2KDhrQCpY8qv9Fui
lHSQn9lX3EISXM/K25lz3sU5XulYvUi+kxuhVXQ+Z9rXQePR4eTxBAUCYSkUzx/35VEZsPrtbilb
C4hvSpJye0mt44xZKJHHgEqI0wS1OiWv5nsMN5JhJ2/fTXWJOnow+at+BPEFcDYntnOGjgd6rIeh
b/DP2oDSeMCN18Ac/W7qqB6dYRogHlcyvkhyAqmcazidDUHPPyXm7q3Q4hltFd+z6NYIQ+yA8wXS
QUnJiOEUJjju6yc+h0N83VX4vF1aJbM/wYLU48xigIFKvMnimOfkHJUMsvM1MghA/OrYko1rFyEP
CtuAgusqnbN9rWFKJ5bCSS24vU/90qD9Cihtyf9zaYrZP9lPbnH9SsjxeM+JT008Z19vldbZmfUt
Ew8dJJooetKZNfrWOXyUInwy5bg6y4KU7V4W+lsnwUv24juth5qLetIzAO8FXWee9hOj/lpKijXi
pxJKvHIbV/4d95LWNDn8U7ZXJq516Xq/dBF3CV2otsSbHIerWgKqoHobXGgd1yAK8MpxZtLFwJRH
ENjW/vtrHvx60kFodr2eIW0EltFP20f22jr+SPsYntMQSCyNeQKJQabI49M61tSdtU2PaAwoCnJQ
T46RPBlUzlB2/LkW1cUQfswbSNDSZ+kDGA8FZBTxE2lPNSCVVZwhGHHpLxwBVKynLVpGVFBt4zK4
hYfEZfhIWQyVbuvAOLXRkGHlic9kTpzauRuewpZXlFJ3vWQ4Zh2tPnQaGszJLauQcZUU39HWma4Z
cxj6lKpRScMDrXPPCNlZEeX7uKLBM5deZcK7vDOGJtyOm4JsmR1WS2+W+NXNftGDMsWH+mm0mJ5s
Kr4iwFujnQ5RkQDH6DB2Y69qw5ng4dCYm7f+xBd1x2b6fqexoen27JOqB5rB/cU7F++cB/S6ZrFY
WzhqlZjZw9RI3rDUPJFM7b6qJr610Ysanqr0TgWHRB4jZhY/LSvDifpC+xFJSOJTKRpsA1Lq0RiO
8Qsh2f0PO2vheEDXqIkp4flpcPnDWe6ZFtu0gfilCGBVFLungyVj2B5UcpUzzUMEeOInkHSSmM9v
QgXGDY8JaMgvEXk9dEA4JDHSnfJ4p+bbduu/v03RqYQk7hkWdabPUTuh7plCHmQf+fxTGch/mCWj
KzNGwVtAN51BaegeFf0umNabtxUkFhXAO9pQ0gVphF/p9MsOahFMS8HqWQPmBvTxlLSrI7n1lcAR
L2d5kRv5kkYOA0Ul4Qxx8rr7bC8MKty+iHByook7V9xPLadhOxjhuvsnlRBvIvFYv+cBLK8RdSDo
ioHvPeisA4kbuXBE9QV7ieaMen3S3hC4dqtmVdDnc42hwaA8P3/jRKV7PjS05zTQ7xoE01PkpV7S
Axp164KwS+4FOBhc0pDUwJ3+944gVSDh2lvwjGM0G9RURI6Rbrr53Db6NSkbBB3egfHMvVMi+6Uy
ZpAJ+/vTi5jrLr+057ArYnT1ALh1E+2ypzikNVB+NE3vzC6omtUWfCc8Qw04wdsED7WOMJV/4Czh
GjUyszlLLBHIktL+QX44F+aeqPE/IZaib96nPISbqLJgqUMQVZx3g+NmRtw6qll6kHsYuOeBY4oJ
kOOizFn7Mlaj0GRLgg40JzvOBWATZWTCfpxqCRTb+SLYQVGi4AjslSni4exThbLZMdiA79R9oOtj
tYu3v0MlL+IFxZ6F/37KVyUcDapiIEWy9FFeo90LvDW7wKeSmEs7C2KtckU3dXVxb9u8632PuuL8
XX8ftNGZjgDu5uds30Wb3AttjnojyyebFkymxJj44om5mqS6ZnBYT5PXSL9JsL4Fz0A29Bnu3SrU
YKRMo/3lFvL4lD8cHECGQZ/mBYJVqtTwvRDQbI9cUjMasEpjUJlcespiBUWKSXR+BMGp2Q10UsV3
HTTUBc0XzFmVyZghnWUyj3l4jpHwVni+Sp+ZkJTC2Bf6xrUwXZqjvNkbiIoNh7yW/qIueNqf3vsQ
qzDT6VzAnVH1mIVh1CBWeSdAcngVXn90X4dqu1ws3LkkDMV34tuqqkaz/w+EwogwyL66Ms25yUyQ
wowVsK/DTdnJfefhNcYnsrT23OUUlLrh3AcyJq6uLUmyF0WgK8HQGKotWC64g64T4581W3ENJG3m
l4PBI3ZHfBUkgUJMWbdDsPFaPTpw0SOrHY8iP7UYKgMUJJCLRzO7B1MaRVhCF9BxXrOZdGvh5i23
08SGkVafCzy3y8bz/SKN+iD/epfbcKvaPafPsC+XQkWB4+wKvidxIlwuXUraniLLVPLPMHmDv/xu
RrIMcWsE0wBuKfWjN8BgGqIu09PrNNgqEboTw0gh94LDdmKomU0Hn41c1Vi+LNb6vABGvoD75dzN
ChWf98O8uDVOWaFQ890dw8nPN4vtiUazbBganBwZLw8S2+PiQ9eZYKtTMEmbbsH+IRbzJuXKZDiU
aDqcuGw0qssgbn84pQjP+nNYHbNT+DIFgbUlph2ucYAamgVzpzWxC4bn3LgeSWa5s5PU6UDoT5Xy
xhabVvHYw01tiii4YLWaPN8ez0MqkuvoGTELNr4ok9AXDvZ1oO1pxqq7gpvq+Ib86Kc50nHEmVFq
qOXhRJpa7020jR+nvkDJB5BtqsSlgsylRVYZskmtET8poAJU8O/933gXjcAId5k1h9PJpWxYX/lZ
yPeSGc9u9Jr30Rp8fQcDOQBQRQ5F9IufAO0xkt8MzFOh/ptJkIEJyOajlzDvRFQQ3CEDXjPMHl0D
AmVOgze0izv9kdiC5jgOSW3Q/inzplVCgF58mDfkOefBqtyMORcjYW9XU/8b3+NzCdIScqYqbIJm
IEw9BPleD/CkMpVrOmn1lvdIfOq/K6DGscf/+fK6ip9tuRzl961hwHA/ftmz94ckvqpC0qtT/rdj
bsy0CJkHPdatXKtGAY7Zfc3hxNZn5qQ7h/1yPYXi3nykPp7jfWWkeAc5voAJJoMQuiMTucX1jC5I
wxzMR+UAp8eYL76J36cLNX/Fn5W/WTGCMtlOP7YTQIe+s3G/RJVutK7WJiNGq+lO8EMDCyTkJaaO
l8u0BHnO9UHva0wSgBMZxSooUorgbrYYsQy506YrK9Zjunpuz15MaskTH2KJQDgZUQGfZlUvnauq
Z8SIAx7Qqp7oDYak3Mz9tapxH+D+dr1QCChZf9FV/lE1H/OUMZX5FZHMAWmcdHZxWQ3MfNlxX2B4
CfFPRuaOJ7L4XMl8x8sDGbJ3nzaSRp+Q9ScQsMqIUcgtYmptYX3wZFzP1iWaqJMMNQCKua3BbOpz
jBJGBh9YDHMyavLxUJudqHmfQRgnAMroiy3U2t8JoFjoqEjnI6lHteZKKrxgMF9FjjyFSK7WLiSM
u7lrI0fHzv5XhullyonNekhEV8AzQJoYL49nVmc0IISU9sHX+/dgf3L/KhbQ2nopRPVhzkRN8NUr
xgQK4lcHQTyjevYjjWVP5p41Ea5GFdQToc/r0IqLcfiAhGVdZQ7mjKWtJ9i3ONLMkiitZavPCvOA
UKHTHgMKMtD7xo9Vu0nURETL9/RBuW1tsBAe/UiPYxHoU+rsaNr6NbIYTEgqLbVtj3Z/mhJuy47/
tfQQ5MJ8+iHg02vfnJfhw+zKXZc8IEAc5UrShZZdK+teolQEqUEG0mEAPLxfaEsLlL+5fcJ10q8W
Hgsrpe4LuckdHvz285X6KlXeTKvA5GhKG9UWMXepTZUgoNOY2ThXzRoELtR8B2h9/xh3lzzlQ3hU
A1mYh2ru55x+fwdRZnklX7fvZ3qYJP5lHU79C2cYEDL8J1JD73XVPX/Ps1NoQcFa3oL8iCXqE5mv
Aik03Q66y9HPqeiCCej7OWGfALLRQqfIPyrdya3PehDFZ09CQLCsj4CG0bQTtZtz18wP5/vmOLZ+
C/C2YTI0a5dMQkOS9/h7RhyJUyx5z8tJiBv48+zLJmHN+N3H3n8X+WsnJi2lsJ8Ivz/iehCsbkRZ
MuXbi4G7ulrRTglw/caZhNDgGLYy7MjtIBk9H+s6oyuRU7MRv8YAfskvQF9c0lm8Dqz1v8/VQeLB
/1Ffpq1jwTTC7LWeqIo77+lH8IxzQor2LC6l0djxsFAKeZX/0lRGTEeoYJmODdKH1Idi5yrkxlQx
ZN9JxW68wOechbmc0y149/qmSbH8L8DIgtFqXO02QxGI9ULUXL3MyGV8Mw5o68wKQwk2PxV6jdK0
aTMMf9Cc7FLXb3I9cdP+MPXKRn1dYYDHPOZ0aOvCg+76TRjmEK3EjpueYJIf4UjDd0dTgGbgA2XJ
joGSw7QhFpqASK3QeO6qhv7GtUOvgmAuZE/SDkMkDbPezlKwWyZjoUzBEHtz30ESlmMyg74mQJCQ
qn5qXz/vSdJ++yXcerOfSdhneAOzbweyx0vT+AR2frgRcSsnQ2souDTY0G8KNv9QdC/Sr/5xKUaT
zbBY8cUnaJLKU1Q5VyqZg4O3oKmFiYrOQ4ZD7135kFldI5ZgIBak4JughxcSct0/R4XhuUPjW/In
rp1CtQiaFYlXK1eDMWXHrEOJAJO53ZR/KfKSUc+af7ccrMUsfI5BdfOOsL83E2rg7j925VEdxX33
iwTrCf+a7/TNBZBmhXe6GcI2DpsM7W7Ae8Etu8/rCZWR4OPQsvHILPWtB0cW7hHPhCNSRWx7nm7g
pNCQpcDPZxiZnw0FAvZT5Emm5DkkoUgwu8qsKq/EPnfdz3h8U02T/FUqKXUvitneVjBPocrGV2PO
oB/JUao93FKyqWhvqft0slAnD9LwUAt2EeKgdSskXFZcvdizEvVCvQjN14IFO+4hoYBacB/9VMcT
eoFCtRgExlHO3xftAHIozYBLCRoGgDEGYgyvzhJ2KNZQROOkahTbeQtYE67FBI24OB83mOL2z4cd
djy2OTzTrXD8sKNvA8ReWsry4tp96iPi0JIu3H3O6hVqIyAQVexUPFjj5O3CV+zaSxi82zE2lvSR
PaGXmQkO1Qr+wvgj8bvZRxCALBi/Vct60/3XyKHg7YRuEfK2QVT6VkgLa5YFYQYeIWDFMQclJSay
ZxvBKyIv7Pya16lbhkuaDtkWnSNADXI2nSoPKISeEADSEabByB6H3sC+gycuVB3dMX6QpWOXnfmv
sx8olUhtkL2ZxY2DyTDtaQXstakQxBATp5umsUkf8O8Fp9vN75hkSDlQeHUyXmUsJxMTpcqyTBQ9
TXP9l30wRwNVqS/RRuBrh1cl6fe02vsgz5ZcpYvi+JllsUET88N8w+dJHVnQ5SX4vaX+GdZY16wJ
J0nuC+wxchbJGbus0uPGAe3PZNcH8BGH/89Ingbqnvi79p1ayZ7zwlFOhD/37UjtXRXWXrLkw5sK
qHTw3F2nz094omRMCwSQQauI/hqlB54fooK5jugJyVBGonBHJmbSz94NHFwjH+xoL48P4uLh5sHW
4dqtsqsV8UQyNKaeuCbkKE9zx2ToczMziCVFfRbx9JyrlmhO5YKkz9EvbDHsSekiU9kCtVqa72mw
ncuiFG1m4A7ydUhwAh35riO6eKixw0JCziZdrz8LBf+0KJQf7F6M4d85sBXVTZysIPMayCLhkoss
/VFPpiUrcGaG4/Efioqvv7Gl6XX78+uHqhvwSt7QfhIMlFAOnbzfY0AHAK1OGfrb4MVEDcGzMWx0
2nakdRq3CTN8LQlGH0pDpUnEws2nhXrYTGr2YI7telzWWJ5tZc/KT1NTLO/AqKO09fOQFO3ZOUtT
RTuvvMXU/fzr19kMrgtxgDLoaQLWlgWU0n8AD8yAUCH8xB8CMoKJobe75hUSairUC+YnBHCHJRyi
3vyfbVSSqCFwfQfdwH0GGJKAhG8wq+gz6v+2OD+CHCD4J3ER7L3Bo7CIRXnS0CPndmQ+cO1h2ZAk
LpjfehylIBlhsjhYpkZ68LNVMNT6KoukqyDBKbJzB5Fessnz+n+8zAztMCzAiS/SDqVl+9psAnFO
mfwKYFbCkdIZYKxhWqmsdboXRk91rimZ8faKkhxd14T+B7mZ5ZSMBMxqt3QS9npA1PvanoPr17uI
NysL7u3jhjlE5vOfpMtHhbhV4JHeeTy5/Ns7zGZq2YJmDSYL3JgQ5cxlK7uLzn0nfbnVsiNSsrBC
dkcCJAdWghFtn/z5vVnUez8RWeVinFkfsoRHPshbdvwnGouKPTihF3PjQAK9BETT4FRpQjBvCkT4
uQxCDPKnl4JdhLu3GnUjQid4Wi73M9EGloeXEIei+wzCYson8WbqmgKT0nEKDqxFO2lhXWrl4vjH
dj9WtgFJyn85dztFw/tBiR8/vdfQiK5DLQjfSjt6ybXBwFfzpnamsZ2UMovfGURRzn6SJbh52J0T
dDtaWCdP6g49wkYg4BCFxhZmaJ1QYCV/rIuwCOPWSiq/87TfvVGsQHx7iKhrTGs433fR9AM3ZWtV
WsEAQiRvtFIO3o2qR6JUg5cjiPHKHVV+0LWkVT0m5j8y96FR2279Hb/es5c4P25RdnZ6V8ZO82Eu
77ZzVhFQlihR0cqntCeICoNg7RUJfde3d7q3NHY2AiBX7FTopOXx7VPjtSvjiwsVYzwsrFH/Nb2G
HRAFYle1UPnknv3pvoi7h2TDuNAeC4/m7710iCjK95nPLaKreJSir8qVdkSCYlPCICsL/sSX38/x
KsuT+yYUDQ/uyC3/YyDr3hMqTJa+PQtJ0PgL35BStZsBRX0Xol3zGo9+JMunvHLCU0jnoBp6DpaW
KxRZzw231WF8MAOagMvJGBn2Q2pB7bRJbiXhgXXtH6H6B2SV6RVvDD5iEJ3RlOKMtdtwUFeR9duu
JS+qB0N7Qr5bdzudJz2e1K4LX3tv3rLNGgPrQb6Ey1YLKUh6k4F9UftpnZRiLZPABIev1u0yGMPn
r233GCD8k9tof/AkVUxomPDdwhI7fCf0eKPYr76sFeUnRgX7oJt3VUBoJuUjKgzLZd41K6B8YHFl
ZpKIXACcyZ83xOIZ8631lao6U5jdA8XDx618AZO4Z/0qGRMpr7SGXWswy5ljIsYZsWdKiKPBnv0i
yLjLnbr2ZvM29LIR0gNsbckUIV8Wbr+id0NKjj8dbYsTKLVqpYWNY9reORmokJ9Lzb7B0YJTT4Zv
G00JDOGoOE2kcdyIBXvx90Qrjb+Ej57+7hIn2WaA7BtWwk97sQFDhEpqaqBFugGTWVhvbCa9+LLT
n+bWW4RK6luzhyNRehJvaCajwpDhm0/3xckD3pm1SRW0NJqOHjlNrn9YqZVDt2W61RyuMw0DdL8+
XntbfARzZVLnCKBwsaSnIYLodWG0kU/x3SPAmrsMjz3gDqKuqjst/ygDsunt7zEYWam8KY0xsec6
7L4W0X0ACwu6IZHCWOJefRJ4IuZM1b5wgTIk5IqErsfYj9Eq/AaORWjvouPL5Vkaaq3SmwKjIFwU
fzwwcXtSK6PhpdAdEECjnOul1J9quhiyDSKxHx+SbiP7Mst4vn/BVz02yy+tAMSITkugTBdcFoSV
h/wEfV5nXQp2ZeXYhsxpt0esJIHprscEkzCbwg5+8OiDo/iU7NQYq2e2n0WPKu0lQoxuyRg9A1DY
zJ13bkX5Sp94XQjiMeUeYfH+jQ2BKCaP3lVfDwolj0YFHKUAWVvc6nEncH9ajFNMyt4VPF1R97ss
LgJHZWQCoT9kkIcKO4opd3QQeedhWNtm/kWbUphj/Rr3Uzo9l1j94x3spslbcbVCHq6IG8I98T3n
BeWbUauckg254BDTBuXB2KviV31y5A0Q35KuSSIOZylo/SCIqE5YgDvm4qEKePYVw02vhP2tV6cd
G/mYYaxmucY+oVJFOUv0Wm3kDQDYtHbNoXmWeWdvQqNrAGz7LsHk9r/GOfY9r85M2xtxE5xertem
GpdbS39Bh3rzcFYN7WTLgK1YrnRwy/WLD/xKQ+qtfLGbuTzzQ2684ajEnvRpkQeLhC/XjDZ03EPY
PyfqcsT/5hBQsKFkDTHpKlX+dZJ6zGTN5AWMkpZp4lQ4HVcOIK+wuOyDGL3/An7XsU5obSDPoGVk
J0XEM1XuMLPYyUxDeyoO/kbK3TqCOuUqeZqhBSCwFfioVdy9/ti9P7h7o5DAFOTWqaSJsuuej++n
nHofEEJn23uncQNmKdsgKVuSqNYoPdrZbppaV7S4dLtZdN4VQlnJ+MGdYWR7nQOb3/7FpTWkBHiu
tYu+IMKEjTiIYsBo5Uyt4RFoyohQACI4ywXSVjstFqg9r0tQx21cqDNw/tNzuaNJ/Bkbw35XxxFU
YbMkeLOJu7peIuoTxAtWBC+hovvJ+XLxj5lUdoO7gzVoO8T6px1DH+tVJEx5Al+gQ1oBJZYpVyd+
CRArKJfI2fn402FO+9sfVLV9iaoSWUBMHW4zbNLgYfxjt9qL39AIKUGGHaiAp7YbJNSGbFeZ+1xZ
FjdmdH2GYHjlYUt+3R+E1H3pT4DanKoXPKTBOFDwWeb/MPZYyv0dugdxD929yw1BITWzR9efUgga
Dpz7U4LQ1YUtAfZ3ZGitTt9PE9i8yW0f3meWic9YSPXmDRmYhc37z60RNb2I610ipjDLlvrC8hBO
IMTOXIEsWPikW5LCiaPRuCu1nsWeiOOVoaaP44CIgXx1SjNKY6lHhOii9vOV3B+YUszoNpYbEApy
rEzdmtz3NnBv8t5HY3T8nZRnwSzX8QDW7jIaLL18sDfpEqIkvcOsY8dH7UYoocl3QhYVXd/qxzVe
h5mqgNfMDsdiuIkxASjObXQLrjhQIhbMIrJz5VXU7j6DKbZFh+/kGfE1PAd7q75Mm8FHRCODixOs
5mWJwVvbM7Gczwv5X6Dyxy+F2HkoMI14086A/n5CGsdqR0dkEOdsmrQfZPHm1EJ1ZLOuPAw+sv27
oCFjXG0SuF/MnpgryewUl+BTjWPTL/uZ/17Atyvp/Dkv9C8Hq8PiLkaKgZcI5q7qQa7q65Ymxbeg
EYotIvM1voE4OtMqa4lgfedVKueCx6lb4JDP5h4aPGaL6quaIr4vFO49rozjjDeRzqPbObvxkWD8
m/ZEGmHBnChKXp0HBocGfJEzfdMmvW7oiJ81guw9DwtS66aJBjdXGpoI1Tw+irsz1/y8QUP4X5uz
9MkCtv6OI6QdtoOyxq1HjR2Qm63xIz+Pt88gIeU8y24h0zZ+u7IlpcPoi1sYEroPkk96N+wOAih8
Sh/Z9zizzPu+EcuWESJMi+at4etHsTm6uKdZG7NP0Gw5zM79ldVJl9+j0Q9G+76j1JFtYACuAsEu
ms/ZI1LubvsVf0y7EU8xHamnlBkhoT6UDdRmw5y/cpwa7QmLnOnBETIoNMGmt9vt3IQyF/pBwySY
KAZjebHkK7n9DQPamKG36rTGBLfV8FI6688BsGOK+y5CLHbrOO5FZYOYCj33olyBanHVzHeGVQuW
6LbjIuBvNil/Djqc5I5eZHqsor01gWhfAgFPYWb4Bo8Y0xQeeIQtBG4SAPf+BIu+bUA/5FbgII9u
J6Snel2ookChmKs5cakacAqCBdoAYBOSeEGUbZTCv16Q3tiyoXnRRZLnJfwZKgPh1+ZSLQMfRJKt
Y3WYMM928RTZ3ENai4DQW2NITWAVZIlx7df+PV1e664yJTsJ0zx3LZG8IA/eayDsjV7Wl5JLtq1M
Y2dO6Oc7nCJPU6NJ3KYFV45TCIzcJxcus6+zl39I0PlApyJTXC6CRejog00qmqvarSCHzSk0apeM
sfGwsaPYynxi3636PbfPx7NfEpTHdZthFkzCjGay9TRI4ADHWo+Ba7qwC5HWOuyGMa4pFhiObHCj
VeEPGb8osDhYHCCsq9GqVgqknW981ky9Bsed/HX7dp4zn9iUekqvthdnJgYUxJq3BnfAAYsAekeK
MJYhN9WQnF77jb99jQv++cYcM+tNQIEdIP0cw7UvmPTlY3UFidmNH2hCHFb/iGTTWBhOjh6bmV2i
dE95jC5lHMPWRWtImtLBzQ4nQFlWijtur0DrUJDThyQrHOVqRSBWzUOsKORzI4Y9z2iFZOmrBtGt
XqUeDzzZSbmZTPzx3O+GwNRSoGJ5ubxUUtJEd5b8/sXF6FOJ4pzzdsAQaBpKBzV3JUmFH4hkR0kG
00YyGfz3imM4Khwz+9uDtzJXe9fHOChv7w+3yX/2olspPztFKD+6gyRQIp1j56CHZmExOLP/pI2q
+SAFgy9F4KyNhPRVBr39jA3DX/O4hDIDGKaxUVbAz8wvz2AP7Lr08GHzMb7i8tUxcz/X9X1/QFuj
1MAoWF4lm2FrIrcZ10xrABUG5UBwSbDCPiLEidGu4dDcJnPey+y6IhRhgD4DfAT9IS4olr7SuR3z
CcdwZ++hUzppO4x2Mb5VmueE3X5LCRRdSjHIn7RwhLag289gn4M9ajST0MH3ARzeeMtbY1qppEek
G4ew5MPDs8hU+1KngjKisk63bNpdmaxR7PEvvcwoR5kxEHtUJI6m2zSLDDf/MdO8ueNTNKAJ34N+
oDQslAxJW4ujsrsZtZq34v1nP269TomX+KXjWt8P3+0P4lrPj6P39wuC/ZGOxTkqa5AhabgSm1Ov
5+vhDOlgLPbMnBfOaGq4Dxc4C7bTFigwm0u/GBSyhCH3ZNs9kPlKGVoz645aMk5+z0C/5BUl9YLD
8KNretQWE20zVGny4LixuLZ8506jiS9MvensGDFeu63ArMBk9dUfyBvCrC3dYq3xgPpuTauVUEyW
HcxUryW3OtKXRf2FUt5kgo/1q/s5bQLdOGan5px3SFehazs6emg9QGqPXJWvlqfEfmEVOdk7efGO
p8x/CJx+703fDO12q7VlAaCjSGtvELD23n7PfOrMcXhfLT1PjQd/GK3FeZWlbZOrJ/8IDaa+Qy/9
CChINdd5vPAyg2sIrzCsxH9dvQdkYanckhUO0/l377wvwIQFoBjIesVdJWp5JcaYDjTtFJrWNd9c
3Auk4ew7VWJsISGUdbeF4+dW8hh/ldhKzLGAlP88gKor9JKdXQmTzXtRe0fjFvSZsCLGs5/mBHz5
LhV/wOMzCBQwaoq9h7suLyX/iEQ2EcYB6HhxHU8ASc+ritHpNDcMDLGqCVVCDoJONDe9YTawG1OL
MWKyzJNWa8NBFXWovfibrxyVPFU3W881AuL/rybLcOpHPHbR896WvLMptw6bz8iyddyxleD/y9wv
COmnr+iFPMbbUJOMEo5HhnHO7ftS9jlw/OscPH48DA+H9EXy8cTyMgMjhE/h3v95SNcEOQwagqhH
hc7FTbgHgiCJaNRw1lm+LhBngR+wBd8rwemkm9enf32bhSoUplVItV69vkEk7bsrSM7c36cRpcL1
/VQhtoqC8fFMcg3E2ZCBxUwvtxrBn19wxPZ7lITolmn8ZPUTBpXbFSpm/xLKdBXP+BIKZ7blKNhZ
XO9gSH0pOuP4QL7wFof7pHuy8jPtBOjI6MlESWtVVRe3KSinkJP6pMe/KbknucsYq42jcNY3XsCQ
1bejVILtUKpzoWK8AhuNDfqDD5PQuf0/uRT1rTCWbQjg3M+eXhKUG59COkj0zw7V8FXHqMT6jAGy
3BQEf1P7I4e9VXfBa0VAUEkLsc303ubmF13agAmc5MNY+X+xqqQesVDkgLjOghqhoJ6PcjIFeX8B
RQVCOviaqIH3u+wf6XRODr0UOFInxxLtVgQ+RWE+ugNUChgsVWtnLM4mCosg5XqRFnjtbzl5Thkp
P6jR1k7JF0hFo15Fq1SZVfjjXN1l12dqEppP1lO8IWUtYm2zMNEXn0eTHpKeNKhr0AR3Sk/rJb15
okQHpZy/EG2iAaq2iO+CRV8NBhGlbKrP6pRpWd6A2NmqkRrfcDC2MLsl3BMn7phnw0h5oEXHnAdM
rKmFp90Ivs9bNtgaEuN8wAfoEMINWQ1FwUWoLRpLo30bCIT1Y41FcAqQd8B3qMpQWd25nsfll/uu
LTKF3y3f6OqEpjRCbcnNCrp8897lNUKss1ZW/IqvevAQrzvvheR2qMy9I5nn31dMkG2UC0f/EqjD
koGJojdbfEbwJHy+wVCNqAkYeT40ejgF2eXom6BXBamvdyPYbZbR7FCQvY9sRgl99hThbINe1CTO
MMCjmgZ62H/CLS3XUoY2aKlE8xBJZkGvOnZt+JkFBRUpfmLldNYDHaeLVX2AwM9nJip7Fsh3uGa7
azDzUH83lumw6kSe6Vu0PtZID7t0Ap2MxNQgSkAVDHW9pUvCYHk0wsTqM8rbRJgU/brph8gVzuNW
5ZShWwfvBmzNDykVno4MZ4gkM4PjpaJFLLnxb9JnDEpVkgIH9SjIS4bXE/mP3gkEH7lnFILakNac
SaGZJsW8EunqIAN2/5jQA+Wfa7uG0L660ntoVl3q469xN7Jh9aslvfRRwKESbfuOzvMLfhekUUs/
cZRqfM3xFK3UiDvcCTN897tZXRKbhpkUIifyq0V05u6dleQKwSUTUrZ+mcWRlqgaJeMYNOBd/8ve
OHx/tIkDE8GUFPJDDSajwuOj9UkXeiooDWotKJjY44SLl61opvk17T9PZ7rpX+4pDS4ZMEC6EQGc
YyeYAmgmuniaiARRRh7gu/QbEXmsGVre/4EZ1tpcHsZA+TUo1pGEpYNviNZqJNxqA/ZPLHuJp3K6
OsCUY0wCC386FY44Iv78rQzq009mZohgsxuxgazCBF39eiMWgp4sodEusQcXbOo4QYqgPpttj0tx
S0EpazRSXXnYY3606CvOxbistNs2U1A85jOhaFt9TlBXqF+qo6o0N2YTtRzhTWlHqEdsRyNk8eIP
BhAeljpQs6Uhn1TADpdQYGb4mhZAvoLrJsI0Rv8YPVoeOITJ/yoLAoeoxFjnuf74/ExoqxRjhft4
F6swZ3+G9QRZS29swAvxwlkOsxKsJlTnERKBi6cEdRMXtE8dIlQ3UMd4dQPYt8r9TuesMCoJcZ6O
Y5ezx2lZ1XVxwmP/lxXgBQJQ0a8FfmFavjre4JeGQfOIqnz+dTQDmvWIAJ0l1kZx64Wf17Iy84IC
jIXIu0ST3yZNL1aowg2ZvdeJSukztbqBNng6lCxDhppZs9VJiR0VoxKDFReT/y0FUXIAkAT1iwv1
syDNKL3QmxYv7jBMJJNucmFs06n2zzHHhgU1ucANAAkPLK7V1TpBbjd0x45Y8NfihsC3nhO2daUj
fJheNmDZgcdIv16t+rXlmJQcbjhXL0lKB/5w5oJ6tzxtd7KihqZxk27rmQY5/TTnjLrxCfXNtn3b
UegJivZBwFf3c4fWWl07Lo7HRLFMRK8qfAtcQCLn1zBI3EdFQFn6y/at6vFftTS/L2X6Dule+/l8
XqKd7O02n2CA9BnWnrduJZjB3FAba1YJ30/aSzR/0E+zL536OjeHPIAMQl9tbJIfwOw7NAqfWaK6
sWG8E2tGCenx3psUrbLL11BHLXTYDMgpXRdmZOCib5iX2VFwtJraN6nNfC7p6+qZHFcd1cM8OopU
QqoctXsPcQ11P0ILEBcLMNehfXh3qKwgHx6q7Xxkhp9wmbxQoWtSGbR1kgjFBCwGFxYCGf4PKUhK
zD9fmxp5L8XJvo93yGgwDvavbAfot7ypl6aB0yY93GfcvBe8Etnt3X76l5NXvGnSZzALBhChK0YU
W4JT8wGv8Po1g73YldKVpOtzunWHHAlV1eXqb4eyamTI2aLQ5EqFp32oo/Gf22S5kWSq/ya0IC1v
pcJp6Flz4bccq/fHqHCMg6e1d4YgpY2LKv4LhQpheReB1BetiR4U0Ld+hJomHEsgwTPGrt4c+63n
GjABXdckdueLA1XPZujGKnVoZbTBi/FQ6dhEZSzh0oDdhinfO86eRZ66foT866Sszl1IceVXT0aa
WG13c60SzO2X6lIDFchZI6LF88dmifb2VznndLfk+ZLMztxfySUdz7p/ihCJfV4LtnY/XlJ+swOM
LlfsAjhJ2JC/eu6P5mz+FmECYjDurudmH/an6xMtji5kae9Wzlu/SGyfs4oQ5F9ypSSv9WxqQ6M+
J2TECN4BVsEjoj6z7xN6yhjuQQKgLayBxRPBFw94imTS96CzqLLkDw56smOyiVGSETfhLgrMxWUg
G9GttMaeMqDC4/WPcphVelTPJ9LyFskSb8UPjbEk440eyOU0yXW+XiVHG6rC6+2EOjH4XHcD0sCW
/wLMY0o83HMW8Lo/Y4Y/mcNu4rh1AZO6GTziaSIanDn/Ltg3XawmFXKfj6oawcNN+/K4CmNCg0sC
CP+nUkswU7PuEtaj3rdUK5fWGRHHRQsw/pWSUTZHCXFvRFVq361Mokf2DhiqF6nlANO5PKRuscNS
XflxEwwxJ0tFxpdlXPqNhb3qqQaKywGD/gWMWxvhYUWElmxnChPujtNN46IDEkKf4B7EI5uQBVfU
7hId5f8gYz2PkLkLXjOpzkArFJDEE6EbX2pVqjcNWiAjsVjFxWxyuL9Uy89ChXrEen4wse/jSh7T
RrsDfza5FIgdFaYRCs6aIN+8JNBTqiI/80NHhkJgxVMZdmSy/Oa2qHdaffKygQ9TqZoLBXUDJyVm
nrcFGKpRyg1ZghBjeliXNhH/YyRM0Fnhi7VmGzJ7LBzknyrswy4YPYTAyOhLeKFoKVmUBwaqCSe0
fZ2akfzuzhOikO1tlgQbmZnyEoZpZd5Bh6eiV/sLVQFNE07g0mu1jD9eDbxWlfgdu609Fyqop+pZ
C074kb2qBXyks8cfbqR0GIeqeoaV/Y2hRspCtyeF+mzvkYa4C45km9D5g8mgxaOByKJKJFJLU6Rk
IUYYdPhOZMgsbPKX1pevH9UExQo6zJ6LwYUGb9QEXcx46QWACfVWS/UA7sYF//0tdy6OgQiXdiGh
td/4d15apaI+QEKH56wwDjam/ox1shz9fWahl/B3JVagXXX5Our4hxhycCbLElEB3YJhvZPtnPy4
fnLnP55wmn7wCH+C4WGMqREJFPcjrbfEfCbPj4tuQ+t6E/Qwq4uSHoxCPgcxEaC5xQcOs9dfTILl
hTj0VIe3dJ+23HGE61UJyRxBv2yg8gZRbkMPOCaUfEWYUPg7kWnmX9Cd4Cp90P5rKVMmzc2V+2E9
8GlE5+mjRm/F6u69EMrcTDibg0rCQi/LiP+teQaveSMciivIsB9gi/3KgfZj5y9CbXTJW7q3eeXi
hLj3pPLvLKByjedeBV4ozEIvmMsOudviCA0vcLEP9XrBCWWiFUw8mcZO3xo0yrxPEIREINMR3p7T
P8Rm6/9s/H1wndBBix/WJQDqTQlxmx2M+bLgZsvY2ZLC1vh9mqPTtNIBHXtOWLbgR7XkAGhSIKvR
2VYqrmluu/RLFKhe/jOchMlAnjgew/bzD+8ofwZnvWpG+vnRvdQHkrx3/lLdVvACmGuZ74ZfbJiD
ztBtjtDmqbBrpPtXwB7KQBOZ2QqdjMtCIrkAfTc32GnOLPb6R36+bS5utt3/pvbjIOa9Y+AzId3x
MC64l9tuMIVdQjmslttaqpeNBnDV8yd1gm7E1Oy+2I+W0SN8VXKnaTmA2LbzpBFabYH2nXAItFTg
ukK8TCqMGyNuOPrPDcugU11RiQfntU+5ylWZvnKVXEVdB54Tcjscp/8gzO780ASlqGSFc+JUovQi
CITyEh4YZwjM3nNTBLXm1mNt0YikkUlX/vVFkgLrYDL1/PNNVXmQEw0EoCrsYXUsi/zgwg0joZGU
GggS820Q3v/HquCLcJ6W0fptJk/hA7WazMMhyEMd04oUXYZ1fGT62TTA7AnLKdyL66LhGSJlCQ7M
g59DKF6UNEc1tlxk1wyI4gLrBeCsXF5kMTwOz6XVIPhdDZPJ6y+x9LgUnd0sy1xAWLuGMMLf6ayL
fYlNNS/p1ZrwaEZFzICPIMbClK/OGN8D7Pz4FyzYrzHUQfLf16IYuw78UU4y6BRyTtTV2ZOLbiP/
mo6EeN5gftYcM8qAb9p4JzWEYMmVfxDIgGEDTxUGzaA3OJQKUIxrKyLrDEpuAR22vFdh/+p+nq8+
H+RsTKmpgiZNIJJ1UMF2dVBSgo0VSWUn+/0+VOtbitU1lp+ecu0A7hzOlf9ehhHzDBz8h3nQZSxy
OwBpom+3QgMX+2jYqfOOp5xdSXb9SyalPCoR4LKnSiobFA2rC556++42HHuKI1UUF6vwYWhgjfyF
q8P347nBnfhvmwzqtys4/SumT3xlLzgjqHWb1KNAoyy875ycaU8+GKy9CJ1kiCyWcPM96K6EYlhn
QfykS6Tp6nS4y1/8ArvSN769cPWPsD72wbMjOT0fmyQc9TW1oSGUdNVpYEBQP9B2TiECRU1DO2Yc
36GURu7npN60tlTlMq5LKuY8OFPzwuMpClW/dhgV5bFofkzy48udO3YSvelLBpCkuSbNaQskdTsn
BbN2V9pxAHYc1pk61MH+JqtXGE7HoQ/wqqpihvI8L3eFHmFBsxnaUSkjj3umPzUy06awECQ6xkz4
Pocr6z7ow026u48k2BtrcfioPE4TsWeisLw+yZJkTPgr5+uGcMGK9VkgRv35QlDOlIMEL3TRh4V7
DagJZK9WXcC944bPsEzNCnvXUGfkGltIPFr0AuvHsk6oLsSDLmCDlZt91vqQQ0ur8O5OKa1e6DEY
8NwUzD2DZl1RacMtjQgUh7Q6x2ONvJQSbBPwzZlPK+XVuvJMM7A1ZZJRVjJ/GHEiLDiBIz1Ka2tx
FtJ9PqZWeKKZNExiJLBSiECISM2M/Oa25Ih4iThPq3mv01lP1tw3qvyB6iWg4y+ImwNUPV/zKdu8
HwrMrIosQQxZ+fHUX7w7+eI3Uk91QYQ2K407UUnaW8ehaFuWRxuWSXPmfs+phAy+Dosdg0PUAwek
OvfL0fk79sfRikiGKxkBwLU+bxRxdmxyI2/hWDBAAwNu+ruMlTSRkmEZy6SZiso0+QuhywTSJBH9
Y0ftJxcVyks+fAEDcTJLRO7zAV1GHmKjUuADkDTfhhoGxW6hkzsXdvZk8Vs2boKIns33WMAUMFPv
jhEd77M2Ed5n4jhBY5tOc7y9wtimqeBbpKfMYdoYel/EEDJSOb0sE2nDoBnE83kccd+FVnlmNNax
Ur0wRN75r48zc+1l1ydX2Od2Pe5oU6i9a03rvX9716p6vayVFeixXQhbgoBpBBCSsJuoYXbRnm5S
Bk5yqLhVGp4Hk8LTiB1D2Ue7tyE7ybxJEauz+xJcA3Z5zP1mL60lAGcGsEFD0APVlCXyrKMBGa+r
sbTgBCDrTRo6IOyC5QgPSxKTWNVq0EkeflxbpuaGjA5VUE6KIG+qqdIQnIK3UuCRDwPakTG+tQA9
rtBwY+Criy9DTZYgL6Iv9SbbUQFVzujLDNGbmhdBDCChY+rwklqqJNmSiShGzb+n9vMtWP0v5e+l
/bqmiVSNHMJfzuVn7WAXp9WyXoUxFBu4XMl8pktYg+8T+mUFCjs3SgOcq/tKRBu6wKXOSFUcoG4e
LQUO+zMv9qoOwqIy+zebvY1wzmFapF7rNXgCbeQYX0YXgWi8+aglSmjgp8ynLEQBhINwVZyMb2Oz
OKEZWxt6hovXosTS6oYioDMSPCNMhL47s0WKfp7JJm1AfX6w/dDjdlOR1uNSBxVEjOvsviZIG1rC
h7WlNJLxMo2/Rl3c6ouKdK6T74xD/J6kufw11YytGFWqQt5T6KHSEcwGCIWetxJ4jYC7bZOShHAY
VY8B6QMSzvyx3OkbIVQUVrP3JXJfebPPq+pIMdQylB5ieh7mT3/AfRan+8b7JFhPSrdDtB39Kxqq
Sxpmt8rrRelPcq+aXEhD9O+SacZGXwftkVEOJeO8yXZfWIxrAKslgfOGJKJtpSfET5dPKMo/5FiY
pzbvBCdl4HbKYYm8ZSIxkrresrbkgmj1OZM4jSv/uJ+JhvgfZm9DafqgFbO6A1SEqVeN6qqe/GQt
KKSKY9f1rv/28p632MBhZl1g5Nt0dDMkfj9Ao+DDB7fUdbPELU10QWTL0CfbqoV90TNFrkzZd6In
tpgPzr+tvJVEpXLWCFLLgKGyohUMOfDKrigQCKwNarFCeTnwZe9jcmlBxU572auC62DlpP8Vdzd/
4TS9kBRNs++k/PUsa99SXXH06TEPIty8BduZyn3thVPpt+VY99gJwvlJ4Mwa0r+uW+3dctayN7hU
lQ24rS77VEGqhbJJIYpzKW0EJNNenCn/vmpwjOSZTQHHZIU16tvys8QFzNxdy1B1yJ2pAQ/uPrp8
ByDfQRIwbd3tb6XXPxfSzLtfxJUU0xbdpvZVtXj4mxHgSthSOGYiOuwwEiIm6zqwchCE/mw5bpoQ
8h1pjwbjjm0ssRErZnP2rVLaVu3n/m4/4ouykiNi06gsoCkWK6B75W2lu+RdGMD0AAvo9cDYmGuW
wRPlj2+mvEwUXxlgtuCqJfoBiGPaINCV43XzxWtCxmHlojN59yf0L1Z64jecrQCFBdcIP0ZoXDHN
qspxkCi9V3kT2JljXMlfzScuPLCw4U7FVrbN2It8EY/eB9iL1yEtEWHBycqQrFVrH+zPo6aZNyPC
4Wt6DhQOgGGI7VZ68BcRTJymVafFupA8b5vLPy3ISo49c/UQetHzoaRHXHtFlUHuNn5xrw9sayx8
y81tNzMmnxX0qdTz4kXdw8Yzx3y7oDUbsPZXgICk/5zDw4YYvjTAwCcrRsxKHwHyfKR811l4BkSI
3moWYFo33KlDtHOnVS1UCN2oeze6oMvb1MaIAyBRJY1sR9ZfcDARcVVU/JC9NP615qIfi8Kxv5oq
i3l535pM2UTZApRGKg8ACzMHOUKK5wkLIBtUpBZvn0mVkRx9KYbfbfoZyPbk8G8TPIyqcy72ap0W
mPp+7mZqh2tMWOYEF4BY1QSW/0weMsQEIGURpgrqZaTsuSkj9Anh6typsk/8tYccN9TTJ++r9Gg5
Fx/t+2pcHYjdWmvcIEMLT7SvBlCc496yxFSFaTezcmegkmvAVV9myoOyYBdl7HVzwJy26w55CnFE
Y3Tu5BrCZnaoxlaJ+QupMJEZr9j1znXnjjngiIDOk3e6IJUVQ+3KtPKhU6ISezLDoN5+5YFKFKPH
QovsVvePmnAvDQ6g4dmIkXGcai/tvXCCTXReEr0IhPIiAyZVbJFR0bQ+jFIQ4rpdSzoX6k67jE0m
HyHdsBe3u3+YZ3+D/ky+7QKhb3nY/8toOF+Dch7DzX4JE3rEdknc09pIeipYszj3VxxM274TscbC
XbNqnNYxrqseiPvYO/qlDGu0E6ElIrbEInFynVE+AWwdprdFudBYJEMbxLbxVEmONWEMubQ1wI2u
pDSeEwD0EICaBm4S1izCbR6pJnhNwCUsbVWv+IjRUkHI726RY9doMJvi1AbQwOtvUk68/Ab5cB/P
0VTsHi4Q3oAa00+pKnnMw7uxOhtA32Ev32zekgHXB7XtxTr6qS5aCk2K23nS38NeJS2zrQKngKLL
HxX/K/P2ehFZewQooRExABvteXFA7ieW9/m0eE+jvXCK39ByAwi6i6ZQmo5NFQLY3vlNAKuZb4dP
Zr6w8xQZ9UTJygH/P10st0kXsDU9P2wCg33GChTBIkdWHdSjgp5TyWYpBb7VDQoBz5R2INhrQlxh
MWuDbJws+JtfCnv9xH6RgJ+y8Bho7jbv4KzDjtuu6LjfphaB7cO/ccvsK54fS1zCMN2PsYNBTmy8
X8wnLqiUxwyjGZzu3xHrpiUFAHHV98Qv+5DpEdmYaq6o792T68WgOT407KUrDgibjuodn9N8A166
iyF8kM7bSID1v4xME+yoB3xCqc35MVaANazWIROv2ZR1fzfiG7yPTIc1WlWv2qvsLZnyQby+64Q9
cOiWdbhEaTaFwpTu8gPEhDJiliL4IADT84guhGtfAlE9NzqxNFtnpno11Ok7CzSmmxUsX8+hD6bN
zPZRO5DxoY1FBBIRhiKFPSp1GnnNC7TQbcMSYqwGD5zyo8wmdBE/4z2CWQ10CDeU+6UrnqQNF5hS
pyFpth2qsTJcS3spw+CqrY2OqlDU30SgokFrIJDbmSDC+SbWGuOv3V+NNjhhtNR9zIcFaVP+457z
ZdW4Jh/Z/0ih70/asAWfOQlxcteDpcD6NLw8SLDfwWBeWRhLwvYghdE0bFljz6Xl9QLPG5aDFLWl
/darZyfL03D+GGUriJoFsYsG7MwrTuyegNvdxNT4JIAs+W++eO6rJvVhXIecKvpZeGg4+39aJ+vj
wrvY/nNl+pGOaz+doG1WAk4eV5mlQdDbpT7lnYg3o/HGmlee5xojRDSHnKxf5lE+syMKlqqi8nyA
wbFxiZIvRDFmDn1yQK1xu1wI0ioXeGax/L+Eu0ZzVQCRCNFJ77mTbttfr/9OKJHhGOEijzrhRnAM
p+V2RU+WqJNQrCcIsq1/y7pKfp4V9/LDEjW6BIH8/8+eg2ym64YZBLJlos0MHvDxwzFMJgfaYHLh
oUgbBz87MbviTwh7MJT5JTAaMAjScB8WkR936x439ud95nXmZnn6osep8gA1Jn2SS8/mwNHZ8P5N
yhhU06/BWWgJ9knfcIlHrfvEFictL6pOfgfP7lEGmOQxDjdMT98Iy1mWN+G3H3/OWSBviY14NfFW
+ok8pyqDlnXxRnpztQbwqlOtf2BQGToiBr4LzspetolsGar7KUnSlsLvG4yPVbwRdm68WSsItKKS
QIIEIIM4RvAyTEYCs8jHdUVobj/Eo79YWhRvX3YCcMtkPEBvrd6aeIyt2OCJ/1Ezh/g2w6ntiDKe
V4OddLnLi4auoOczY5OSmLScPuDifolsPwxzSRnHR4HTrRfa8lqwgRtxhGs/htx50cHI5RvNiWqx
esaXVqRNSZ/+Zs6u74MPFfVIR46Zls9wtyufKkVKeXOsB2xpS0kmfmSeb2dfhbSu2zXO4GAB0sCm
aMmjs2gdc9YV2ufbUFpyL443Cb0gKzIsgKruHBO1f9O8CrRUVVqolhJqbkmdxCSkiIz/4W45hqUr
t5Nk4t0/FrD+5Wc4fbbpj6yhdAiF8qXGKq88WS++d9lLkGMpMcPOWY2O+rJsEdJaLs6T1qXRu8CW
8654ioyZCYdQpAlezRuVMX3AU1t+FnfCZ17sJ61RChZfLyzrvgZE4Q1/2o3qndoQcrFttjN+6JZR
Eg8pGH8ArmE4jf7nXZPZUgbkWgmCkF9dFPftc7dLKO13dPWU4xrPRDSf+8snxhTlCNxNc64GFaxl
CWDukA1UPH3a38s9vOXxHOixm4ZhyVzAj7fVx2UPuYXoyXz5gZHE54zFts1iHC/5ShOzKXu9efdW
9Unt9fYTa8KGo2q6cgrpPIjtGUM0IISBoDK6wD2+KlgvBVJdnbCJesDjYjaZOUTf/VPpPmUgzQpb
qTTZCAaqOnY/iEoFoq9qV22apBTiqFXnUEcWOgtRbuabcm4vGuUW+4f7E6vqc3vYlmkL/PxlXq+M
RH0HiKpmv67l+LyJL1/giaw+GAtn+KwsmaOUBlyzLjGkf/HltU7odY5dwnwJTbqAayXiXqCtwqrR
KnrLmlNLqiTypwkbbN/VcY28EaqY5k+v3XQbEUunMYgh5/ki0J7k+CI4JwKnpySftSB8Xarng/vn
MuSu+5A49pAZVbkdAfLHEthiZcvh2zg6QQXq2Fx6PaL5NijqiTvdeJPOJ1zLHZVSFLXPtG61OZF+
9cFDVoRuiPHPI46N3lOl/rK0FI/m6puhy0ypOTcXQW3Xq3ghym/HReoVAwGSc0sHdMmp1PQolphd
kC7ZOMBRyfvktUdotHTF004mVvEYkoHWCBTrBoPsBbOznIYxJOuQatcK9iHxFAq8ctj+uudvQ/3B
Qw9AL7MBAnXNu1+mLaId64pt7pIuYWPfTV8dstXBmywPIcdMf6Bs5ZfU8Z7sM4sbvbuj/+HvlnIi
10KNBgzVgVziYaqZSfsz39JkUusnXL0aJJqTCMoFWq5hb7e++dJLSLrDMDcz56zRpA6tIgYOaLdN
7M0rqfv0PaSysSH62v1b1b/BVDasDFkIskFuUWgEcKseoMRO3DoQn3qcCqISrkIindQ5S5qYfhmW
T5FTJQJw8enphwqwdD7hxzSmYy9n/+zXvGs4b69KTo7ViB03Zomg2L2qwrag5ry0yEAlLIOqsRlO
ebcYM5xEmgNd5kiMjX5+0Q6FTBkpApwnof1M3C32oHUWi7v/I3oIvOiG+q94GjOriZUS+5jMUapk
g7HUUofEboQGG6Kf+uTz0w0IPRmh9fIrHT2F8QeqcVIPMufcnKAg8XMCIi32CrJI1iuKtD/EsUzH
CNY2bj2Xg4ieLrDR+AKNVINFIKtdP5W51eZlk09rF021q9ONEd7fbmgQaAV3P1z6HRcUk5kxrbDd
OqG87/E/s7baYQDnsdGPqoGZ0cyrxM2VGzVLUPeOPhTRz4VZ1Z5Q+T8hc+3EVaTADviTlhpW2zBU
RcrBqfnIOS9duVuemM2qj1OBVQDA7UQqU22myOI9BemdGeoAaAk3uTJbFe0Sw/4ORLdnmkk92wer
KwlA3DAMCakrv3gDYKMbP+BIsYJL/ySxXtn6NVmq2hiWwtSlRxEc04tDEqcso40Yn7PyiTxtHAfN
WyuHpGDmtfp4LUyb805cQZdexSqLNNNxsB2tgUG9V0ZnfVW/o996SggkK/WdNwI/aAfj3ez8xyfR
0uMROYwzadN4wRvwbRFf1F1gTHqfGrzcUb2C04rYK4EFKlf3rBSB4Yo8/QSyV7Dg2bhUmVMeCAK+
1TmigqW3t6ijuatq4LZM56oF4HlALzoHUVj868onyAkn7ZrW7tZGkBGWiQhI/wWFna4QUZzNPAJA
QVM+S/lk6VEtITZalo4pxrsukK6u3LRs13fgSf+b6ziC1QrnW1WjhGmncqKpVoGJMCA1xBRZQn4q
R01vTLn+ykHcaJSmL9LRpkddyH9fnN2BxHPSu7gt+ESw4BlwhgkZhO3huv3KhCVfkQNzA3LNk4ol
vdOQBloIrcSBAx5f0r06+e7erEDJIBnbr/8k2++mSGHDLixes/Qws5k/ONZF7ivt4jBDUs5fhPBl
3BEBRA6di42pWDQdV13YudsbKMHPjUgu/PT+zxpEfaACQ5dq4Ne+ae0hU5sMNEmFBp2Q5ZYih78i
+PZ5ghC6ogxYGbj6YrgQayeeEoOzg7sL52FtYwYicVc9PL9U/gPD+nhVgflNkHUvHSbz3/kUDzGS
uXbUiqIA2XlyklFUlYPw9jQMX+AugB4BWWmKxfNfI39vXqRIp9Dmu06lsaLXNPKrPlm+c5nyznjc
/UcAaHW1tgaF5b0jzjkai8QDA72ui/JGxX1y6sem73wCVPRC58GpHbjxSKnuh7NXsWFIR0wvAntx
zfGJD966ZvCDJVQRTaNKEfKi9ufjWuXONMqAEO2edEf/Oj/huh8GrS8xzM5wxkBcB3CpgumCllJ+
XyAkb3iC55xLbmmrmSZBcaYQNMayz3DZDiQjkLucmYbr9Xlwan6L1yppy+TeZ8zbKrsXz0deJI62
fxG2ajPy8z+HdvSwH8FeICmXCfmCxgkl/i1tG6e7wfRm0zY1nKgL26AtRt8MXZj08pMbkiKdTpbT
cTX1Fzy07Pd9J0FsTtRKBPQM3LBD94vlLXKw/LOPEZkJ+P9REb6ZpHei14Jhaal6n6PqKMBUBkQJ
U0sDXXzoGonnwwAtT5zBW/4hArN8iOsOJw/jh1xcVAs25rDoNeehKo62GW3XxsXhdFu4t93P/srV
87CW/wKkkHaABidjcEdhZcwyJcC+B1KI9g1cE+1xmTWjo78ho9fy8vOhBAwvvYyhvbtm68lMfQr9
EUJQ2D+83twIb7xZrsMWVaYL+g9LfV4dOk+WKC6hvJQNKwDRbkkoImCbfgKmx+ffS4vHMYNZxUbR
IHHT5IfhFF7cR5AsID0SaarF1hIeMevwGPZDJBLmLEJLbFppWOMyVH1XM6ZAupUdqTBjQWgo4pNx
+GcOrS1xDT2yAzCGZNa9aZRqJ++ysN+ySJNM8RnGDcQwodre7ZThCs4dVHxjHv2HPuKLS0/p70Uw
mbfJY0yRu/owGlBvjJK6gJu2QGQT6e59JRaQEnX/z0w7TT69f/nN7jS7N/gZtVFNc97TWi4jHfC1
g1mXY5UMWcl3bABkiK9zp62brdJoeI5YpXvpTIwcGWzO1uVm3NopHH+RUHeb500YNhHlaBnphnQo
Bs3WygeFqbeEVbREotZIwfQZ7/knbex7zV9TIqPcasiIPy4JHH6v2abOV6Fgwm9OJBvGXAha1e+B
6fZpreVaFt8iXQHw2Q4OF6ESJuFnzw0VFdMPeANtZB7cUQs0QeA6khvN5v5reFuBRQY1F6ayfpa9
mDS9N6hE8dBAnNurZpsd1R5dd1aNfzYzoyndGG/DD7tjU1RTJg+B67KbqB03B5DoZZuYzvfh0rZr
/YuWpf+ndnA66tGTvUpEov85vU5+ktJd+7muXo3duoIKip25DgV6Md4iZ8UTxosfdJ89AjN0NJ9O
3y8iRY03LJ7ryXYbd/fw222Ap18Sq8d1tbtzKhG/mVJU5ZoRSA9YcwlkySiDm0jahAxeBX5lK7hf
eODRfosU9GIA2vcGZpNeDZYHcrhgdtj7h0adsE5Dpo92LvZ3ZVo2xwOLvM9bCPVwS95kLlJlsnid
MqBx3QWbEYxDc5kJz5MfqvM3mYQtmEK6C7cUF/lKH0wTMup8UqHmVkXk0cD1dF2zxuWReRFrSmMZ
BJcX6CiajwirKDpkyG7etg9k1CCkqts/UxRQabSxSVwRYDVS1WtrN7iMHjcSWycYioyczYFr+ir2
dDDnoaHHcBSn1g7E24KukxiFZ/fMWMw8wsN3xdXjBrgeZf4jQ1emZFhSXwrc0Ejdk2mPEeMFYZTf
PQ6xa49uP9AP020PheWB+gYdUna7ukrjcO5uagrO9dUCIgxpTe/MIbDwuphglGoYya3WibOJXGpf
enjrDsa5FpPseba6Iqo98vyqYzeLXZpMj+ws2UBVYz51BI60q03pRN+iAJs2KH8SLYyJIWsZ0WyV
6F7SzWX7jsSPAye7IcJJG5wzMp9Yv8VDyuB6m/CtwzKzwE+MsfGOE5f4+zfmHcFwAiJvpHIcpyCl
I4HDLfcoxr6H6uegPhVjk0KBISthXeF97kEoXHXqLEK9fq55uIVTb7OSAPEjL0m1ZYwVOapdyBbF
W/ZD2K/SQEsIZR6E+Io3vocpgDXN1DKqEiPWffQPVaRh8lD4gdfINwzNLiFlzvwRhMC9qNJvvPv+
2e5yZE/2L6HzH8vQqIkWXZYHpivfB3A7mI7wuDMtL9p4e++7Vl6pwVvqmAib9bwqxGTxqLHgmRcv
gluHc4UjWX+zq0tMcQvkhrLuLbZrDJ6y/QPxa8PBJbhsdZzNet3zXXw8e9uSwG9j6jZ/wW+naLBz
fhE9/EMC6C9a5gZ7QSV2HVqOcPBzeY4/OLCurE+oasUjlZmSMLvp+RNTEr+ovk+M7OQvaKygx986
mMA3JaQ+LxxdYcE4mk1dcswZL5PyKV5lpqZPQoBRs78ig/InAjlWJ1v2JlrqZI+F6KJW9jFrSBqT
J3qR8XksSAG3kmrRU0PdKeNx22dGoaz33ktoIAngZjGbUgtuA3jH1/hBdMrLvzIdUo5UNZKJ/7IX
jX2F+9eGhUG2keZfzIDI0OMFRKHlDI8OUiW/D4hbZ8V3iXs+JTKPvJEBXr3DCBpZYfUfBr0Oui9R
6keJLIlJu8z4rFuiqp/LJXeUctHvX68eBD04qyteLlOMx/QT51nqRE8BAkfc/eux+jK75G2VtDJZ
kmPa520pj8Zgg0A9Nc967JUGSkZAHHCX+DrHYUh2In32e2nBcHhyqfOnYa0EKB2vOqL+s3jfLnvq
jbzYSNETJgFFikoAEK2MNjv2acY78BxPQKA43dcB2ZZYybvAYAohEZlWEZhbgorRzOq88vwsA3Z0
9yeK8HN64/fX2LPOhnVzAt/LnUObS4FUHqJwsTbbUKI6yz+YVbkOKEj3QHpaBGSa1K/VDlN6dm//
tuvi7iz5e/1tUUFLt2voKPj47xHL7pIbaBrGSrNUC6mozVoa7XHj19XiP6PAiMwoRQk2+gCHLl4w
tCKreHj1LMlzMMFcTDqnWi0YtkApkc350gMyqWE7PSDyMrEjPbHo32nsP65jeUpcTJ8tgkwpod8z
ZBb6GYP3GF1yAwO2T5Tdizrpnq3SSU5beVd+SvpEZYHhBldcsSVDioNHFMfpdJAs8ubm+hlma9c2
mvltpio8OBPznx/kXEGXfgPk8RK4DYgJjdeTOG80f+w0vbfwnuln9hMG4uh31Z0DxbbtT20HvoZN
pDsUA5U5RF8UxNI+13bzFptlFMH2u6EI4Q02tIRPtcWTMisV5XG4Obm2p5GGm/XkWiwQNoDDXaJw
9zvGt961wDbtQl/zT+nbjtFSHKMZ7Y2nbuv/S+U3oCQI3L1ys1ZjVzzAd88OxqEQ6oquKCC6x4pa
XdbXK45B1nEJFMX7GLUULtKEbhVYRACVpn4q3a5uRBHBCWduUha/NU/XjqERbLEfkgh7JUvU7Du6
jogblMhXloAeVLGQRY/HlDzzWxtUNdU6IdA8Ldh1wbpKsQ4HEQunEMW7KLrIYsy0UBVSp1GByiRk
y+pFsGf/Ljp6uylrQUkWSSMKMi6Tunucrc+0vijT1q0/c2iCdU4D25AuJY2ZQsWM+h6UNc+8UpVz
6m+AJ6d/n59uD42K8lSlxsuYZIW10TZTdteHUiUFo9TaTe7BQlLH/6H16NapUJFkDOCrqsldYT26
VRWANTkDSXSBBtwBRfYkVSse8tgXgBpZCgLFO2pv4ieoPHGajXQ41dGdFt22ha5aklaGVLRwyGIW
JBSaGY9WftoP2J/92V963zMkd+v7vLGXTdum0aIRlL9zHXKLnf4j/9P6KprSQ42ktgwh1w0gQglD
si+YJs20729GyjCIp/sfWj6lXlgDZ9PCR0CMFgju8EnWMWbDYenrMVgQi1g3WKzRMb6E9PhKhcp1
sf0NfYebUlII9h0Kq0wvSAGdtD6ODnmY5FWnainzYaGKKDw0r6iWS2TzQxB1ocd6Mt4HOkm7B7Oe
LYmnSpWd7VKXTe2Y/jOVg6Krze0s+pOKG+EDEKz0ZBJFHl5t3nWlVT3zztHtEz/dbYTD/K4NjXG/
+cr82da4ouvqQRPXqHYxHKGghunD7XMe3BWVv++96rcflQDbaq76GOuHN/RMoys+nhP/sBM5k900
fT2AiasZKJvujSqY9pNkqYbfQ8nrbh3loCiUVwBhpeb/vuT7smu5bAp09BtzPJZMVRAsdFhIUYVQ
vTMm/z90fh/MFWY9nFROtq2X42rl1KiyKK9gpB10ck5918UOAPHZQ9yIH7DcHN6VrMLfIkilFaHX
4uATVcRQwlN9b2ITGdK1IOktoCm+5yU3lWV4QdIJ+yFvZVQWs2la6lRdW9anvfyTYETvTexKTSWP
04l3tEO6a6ADVbyPe0mbMJ+S91N86Tu8cEgSy2wvjcC96ZM95LYBMFGlk4xAM+PyTq9M9X7d0Qr2
ejvnqwljtdV0XD31Vn4PaU288k2oP6nRCIL59wwks2nLQCO1iIaX7L7ZMR3czOodXhtXvHoNR9Jl
4ciPYB+F78CIhFDoJCAa2JgNpK3G/0zc0T7gw0+YnqkYvayqPGaXvdhGRSVciKl3ZFtUidwLSt8y
o79tyh88/Gmbzh+C9FkoXlkDsN2k2JXrLrbe2X2WsO9/E9vtHv04Ksnav1pp7EdnvPNReAA1Cnij
lmGFbvSbscnKqVgcc9FnW5P2YAYNgtpKd9mttyZgEHiXJ/DSBr/ppDQ/FM8aP7P1UBwOId0hAc0M
RyyeO4C14qOC1Nrcyrhx/13AVoOvIpeohYYNRY5d0nD9iIBuTFrPUjfaaacJKV9G7r/Mrv+mYUJk
A9Ca0jrOg13A9kOdT7IYtifXYgutnban0VdGNd9xnyx51OlpajdTUUclznyoOt4jCNLfCcI652q9
QxtRnkvHHbhg2Zz+MOfIxm1GO/CWQ0F59ojgv26OW6TzTw0mDey8NloqwW/KQD0/iXtAgWOczN8N
08ec25W1xgaiPrt9TEmI+FE2YbAOFc9bOf2OQbW2Fg3NU7mbzB0KayJ2yxQoIhfqH3OjrMoG/ED+
hqylR9OzwFaxA0cfy1qBKw3E7TbezNQNtmYJQcNUMnrArS3hWf8U10t/BQ6wIYuS3C7OLP2Dvj8C
CebQ3yzrjXoe1rf4djCOGau9eDgtUUjf8Bfk62M8UEdThd//MZ5LDFLBWwZ9vpHQWoLBOy8gxl99
H2W8h4t8qam85xNYHPULiHXoTk4reKaJil+R3V4i5F5okB3RD/UPynnCB1pnFfaVsg3J4Y25rgc+
Zg03b0P9zz8NK77SNGKbIS9N3CCmKoVYF3wrEgBXjRjU+sMTfzJNLxI8L7L0Hm32c3db8OSVu7Rd
pI0IZvbOwdAyixv3WaN3kDT/JoQuZcWmaKWOWHrItcM4YiADu76P7LNYDF2op+ivpFP1U0TSrHAN
LHEXHZr0rEuxSHnKA6j1bNRSkuP7j2mhdiKAx1RRjioFvbpBmSp35Pmn4TNLfiCWR1mkFTvdScTB
+Fjc3a6ycKKS/tDPARfUYtER4xBLwlIbXdgRXWfUZUummNQqYAHJax41z05V8VGpVy9lMeHHIFAF
IpoT7PHt5gkjWm+T8+nKOHoFRUuVfpyXmZCE1xmY7vPNEL2VUE7Sv9YaVXPlWR9II1VL39Skt451
Z/daSFu4WtVkqvaQHHthRbBfh8V4HZ26yjVOftBsFFN0dEqMd88QK1dcZy0eyDZH+zYEz0le/RSe
CleyusWmaO3L1sWXICIiqdOG86UjBk83VJpQwYaHHxiUnoRaO1BtJPA/N8Lh49R651dp/CbITtp5
tHFinrvFfdECMl/VM/mSio0F3tLq7+sGOqaE6CrBGqHO0EqHqVcqtLuGiYLpOwggZF7Qwet0JQj2
JHIEsovih7EdEpsW8yjnLFiD0uFJzKJE85kkNpuf8VyIGm89bMJdKVFqPnd43WfRTcEoQWM+e+G1
kPZOJcTc1fPJT7wjbqGG+xx438etVcipEJfxptJ6Pt9/MtFOIe19VUxTCLvyg7TkGgjJb6huDKtr
MmfLeoVp7RG3//s+Aq/fRnH5ejo1+R0Jm2LAEmHQVLiFMhkDkjvHCSR4qQGJMN5h9F7uRSEj6GHS
/6BpDqWeqgRIkrN6xEtOIAr7sJcL+jLzvdihvN+78u8hgBTzWvHy1mXz5Lqd9cYzwXEuPSIF2wWm
cZLI9rcPNrN83QeHM4LYvGA8+yfnnZc1hv6VZ9DhRWoQZ2P/mVVL4byOB8JMpZizB76hjY3im4L1
3wDMLOIIG342ps1tKBFk6MhxvjgRChuTYC/i/Ca8fj7F25jKlCdVJzLzOBBdJEjk8MmyP3SbZ7Ie
RFtbcITRdL7qO96kyb+TfbBR8UTvIhc65X2UnCxOcLtLSjOH4laxTqw4RQoA7DZE/nBFMkQY33n9
KLPnLuy+5TquaJ8rXWCi12aV9Z54SWF1TurpwgN6xf8QkvrErw50eZ3uimsvqy7a3PsqpsUWi4kb
75s7fDs43tfk1ZD8w+QZWE7hjOQvIFG12DJesai6B0EwyFTkCbcsY6jxxx8olHXWxCxSrHiI8ojt
Znkm2eS0zoxuxVdQOkGpe0Guw38I2mvsfeifDQsV3FpKKVYf+Q4nkP6+D/rG5ztGTDZUC3VOhvJ2
sPPezdnok/C+QlGEt+crPC8p4qduDjeJIORney1rHwoB4ngPe0ZI9W6F5Vj26FSMC87X10c=
`protect end_protected

