

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
U7hExZJod/vUi3z5N4RSr1wa48P7uP/A8O0jgaKOZBD7WNfzo6GmQd7doggkH00XJgs7nLyNvPm0
0zWCfXninQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
k253ey4kkVql4FDzRxE0SZp0nnUl5fXV3ls/4mgbh/6ghGRjfZ71MsiTZ71s3tpy77tZHD0rpNoh
xUysBr1hFwWkTjAISVTsWyokKm82DELzMzaI0lqt04f7kevY+q4XugjttAECZCOOrrnUQb5ODPuL
TN/5/7rekkgE3das7WY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WoA52aV8kh0bkIXA7aISXPgNn7kpio3O4wNzPv7z4wZK/v9qsQ4Fa+1FXV0tZ0D+Si1URd5Yt8PQ
TB8Mp2LGBm7aAfzTAAqLpPZr3KRYlBsnuQptgQwkquHJi1BcDR3dhZHYw2oUKeYXBoZJ80Dg1iyE
mKNc2EAX8dBe7hH745fnWjhDqr0z4schwVFz8IHUPGI/WDdrXtDdyYzuiWdux2vjC9Gao0MkqalL
zCFAkEPTT0xtWcvaccmMU2ICHf+NVjiwhEmFT/vt1jXBw7quncqpEDMuzTHteQFztMFqsgBfXXAR
/Q4rfhaHiuQ7xUCcTEngpAsL2ypgKweMgL0LDw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Yb4xLqu3x9ghRLjHN7QkYl0tDMsZMeJQgGEQuxDwwPb+acIMCaRAm0LVh6gbF0arOSlfOKBs+X6I
1sCY01AUXvqPtXEUt+RvllN5odbTYkY9f5RujZ5aQ9olezUe3+JLEML7oIeJ23v82E3q5lEn2hpd
Yirga3+XXZGIeEC2Q5F3LdU1PK/hOr/QQAn7r3cfSPSRAYJBv2q0KFRrpHEdaRVBAVRTnMADnWqM
+83djfdVuwjO+GhXELQ+rhNH9dkL0cqvHYfgIcRG0rYfPORpbXH4Uiizi44H6tpqRpTeCgmUfW/1
kW3FxovGX7M2+iedny4BJan5eJXy8iA1/NmnQw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pj6m4D23BtF6RtOvVlnmIzux1ocpf3A3ahzdQxUHuwpW9nlstiQd0oSmGGaiF66UD31sHUT6dfQd
yKhb6vxivgHto8LAAEiyTiUmNTH/c41wB3zGzcZFasAPOJZMvUysBGURofn88ip4eLF52/qIKVON
l8AKPEa6atmUOWXPGRix1yyvpjUnvxZ+wFAbBvP0ZsReS6AW7b6zRE+vUOJaMz0EaWEMMRdw3vLT
W/hp9Ruis3IsgHsdn6M611ZJnxSa2tuwXuWdXURUJzFjnTsi2R7EoD0bDJINDuh7T6iiDjBFdO8L
a4ER9/C3EG6IOxU+oP2sYgSHnI7dLthCIjJ+rw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
B2bb9hbJCVaDRqGS393PhTqcBLIIS3eowUvDjLX1RVvD9vYwfdlG9rjfAUVzitJwz5TOhOabACyb
mMpxy7hxgVO56ex26Ce3uZlntRRrSfXZFQT0ENioLNV+BxEHrr7uipCant7HxRFrLFt9nR5wi4m9
ZZq5zS207DucLy0jTX0=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eqzUQVv3z3gvc1IAF6D1gFpnG3jJXG9SSewyb0B7YFlkq+2WoV55oUnb7Smo54ZcwqBR15BnF2xS
jlkL+wI6xvjzAFZaDFixez8MkTdRnrNZscyGLFWOHz7RNKwEpAxAm7RSsBEcZUaS6x+lEu8Fai/i
gBi8OQLkjYbSnKt8sfNmpRhCWxhkRR0QylraXCBqvJVR8s/2S9YSm3zj5TqvYxlJahDh9O3V0iE2
aVTZ//VjzAQrgKQboTMB5R+3O0GmOfi7O8vgrOvK/PiOq6kVyAYEvce5/1FU9VRi8AQk3Hi7BRZM
1pWTxx+bC6qDX+NQvgu8HPGpHmqeqS/CQlftQw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 506800)
`protect data_block
+VCObfFZx6npKHm4mI4bV8f3Lytq9qzugDOKrer/0p97xAby6q3a44M/YaiJM0Ob0gHXPp8xW9wf
WvON9ycw/XvAvxtDjb66FIHUJDWz/xj2ulEStzUJdDknC2AzgYBiVzVuHeKnQ89IDwmCCvDK7myY
ZLG3bVABPrsQ0GaupNUmK2JfEOGvUN/AN8o3vRqO01qzH6jER8ZORhE3mmCBfisrvk7y7DeapeVl
SSQ8X9tTd4so6GI91FIDxEynBu6uKay46rcDb/tFC63necVEVsL2y67B+h2s9cLd+2UoJaUCvfgK
OGHmInZWSXYaosSIIk5fLWrxsGrIn9AAxrQT+egwY69fBwcJoGUEAd3m3EDcalIPou/K4134a9pa
Gsdhrzb2X4+/kbaMkLPLLLPgUnWArEIRan8ObVP9PhPo9SWhNUsNEO3zP4ssPfP8P3gcJqtQdlK+
uQLcUTK0Bo4cFDq9nTbKs1QRDn3bFFuTtWzBpJka+HIZsCnE8bcCoZgwiCX+Ida4EtlXJ5kYd6/Y
CJ8zx9/U5ICGrjR8X+JIp9pGFVP/YjxyzicDv+1Oc0ZLepVs0zGBSGHlgFz3APJJxo0vHOAUe+Dh
cHrc5rX+RAcDm+xeh670O5ZOPRiPLEbmgyeFfPyeD3RfhmWqKAQXefvin37O/FZhIrFV+QX/xun2
7BszqfGTZmZ2IVdhY/bWq+hguzEy+us4WFsU4ijgpv6iGQTXV4DVqcg02jBkvwD0CHP9Vwp5+AWW
U8uNP40rEG0Qi8a0PmkO48KeNv5Lv2UD5kRmdadANa7yPPIeAN/a7GcxyXpM9KIv2mg6YVE1hQDm
SoW2JCKdpH8qyBu3sJuTlnWNIB1i4NOJtpDvIorY/EGLaHaxiYVoU+fq4X66HqfzVZxoBk5Bap2j
yIV34WOYuXT/4g0DYFmHK69ZV3yxLftQ8zVP7OCUdsh1vfJTSNpyKDr5ZgnUn40ynLAsjYpvWGHV
UMDe0CHgsfMf7EAsSRBde2apYqV+wXSVqUf+OR2b0NTzh6sWTBRUPrLHX9YD6vYtwazVGxK1XWuB
CAU2N+9PIAWYEnLQqtgqYCN1ddwIa/JnNEf0q/AtW0nxrd7lPwzbl7hl7WwSKGkSnFa9OTGgZOVI
bXxU3i2ckvB/8OSYkeX7oAycwUD8ovjByHC6ctKUT2S8hhf6hQV8b5qPPh/2tocDHzGIj3etA3sd
9vwnWFwAgB/2sDysh2CLqLzhzLBChSjajMN93I5YvlzyScqtk4FPcPVsGx9HHjuPELQXrawwgs5K
b13UyPzuf+wjeWPvFFrp1GSib7Ouh/4vq/yD6o7/Y7DJqIr9xgqRv+J/PPGQAhn9kXW49HAIv9Wv
ybugeQpeGBiWCTuot0cBUyVopky6lIJQ+Ju9UGnlKjX8G2d8NwVlDBqNulooT/crD1pBrNA9TrQH
H1CR2timXQJC2iJCGrEaN86YPBKCc4n7gAXsbqsCguPYkgY3e3bE0rmGT8NSCt34BoAc8qbhI0l2
AMcS7xIFOG41CuwpJofuIAszkKba3jpj9y64ATNMTGB4ECbfqB25/butK19TMNx0c6NBzuCpEAS6
WF8AOU/4pHOS69GHdtw9JeqFK07VGrACm8G085Axal19WxFfKJueo2HNwLg1B1vzxRaJpV9A5AiC
6tnm4Xf57g0KmPyN7+x6E7+nbr/DB5ojEh6oZIoPYgmqLL33/jaiYB8dlEOsG/o/5p+5hCJHf1/c
d9lKA/EvN6I11B0WU6Z/5oZfwJ31O+JIDvn8EcgnG9pawyJ4kP8eA2uuYK5geZXG9T0SuQmEEURH
AEvndOuc6EE9bkOa1VBpq/SgpqGF+XOGn7qJgLFG1WTsJfT9iTaeDSA4wB02hCyOsL3OXO3muCRV
IXpYK9OV6pN/1Me4QJfbhbSXClC0KsGkn2dnyDKQLRsX3Qvtq9hTkBslqlQrNrHN0BDz0fSNJPyD
ypxFfntyAgQN6CufSXdSS2dDn8nf77+sHErcVG0rGg9JOEa3onBZTh2AE8zJyKphLHxaU0U64c4o
CMHCxKW7oT7j24FlgRoHGu/DapDUKT9AE6oWF4NcCucthjTANGgp70JD1/1ujOqWQ8+jVPhsjevL
EQgDpwdZ34R6KeLiVhxCdv/gAPY7vhpTgxpEDfWSxU9y5WJClv3fMXsJWQRnuVA9RTN6JkZvIxoG
pd9gUdV/zrqWBRQJjXIhIxr3J1yniPbYFPMIdYAENiABUol/JoTyYPaCZtMN/EEY4NKDRgexdvt7
39U5WH7B1xKDFwft+x+IQ+RLiwBQHCGIx6t7M0V+yjwDH8krYiKYlL6QbYzwsM7I9j7DsRefsDtk
FyKsDGhwlSUn35BaAg1nwTJ0/xf/deIvNHjhuzYloQ6H0a067udkVRV2YQJhEKOrQdNMXMBJfKP/
jTQucWRf76JJCDpCrI6jZTpY4exw3VCUkeg8LFuldwDfi7w2T2I1aW4PX4uvSHE8LvE2DTIucguw
ImE8RjwFndS+nUgHX1TCuzMc7WWxCLAHQQwckfFCxsSiI4vVlEltUJjtRd9f4iNw6rp13D3EdO2W
zM6zTIGe/1zsdkZplXUEZGXH4BqKMGikJu9XPpXdG3QQPYv01KwbSe8BMnVkdrDF95bwZf5EOR3H
JI9VaQA7ebWJNMtzwzs0byLbcUNVSHaF4n0k7V52fP0lVXmRPHG/wriJq8M7EyIbejXr+wljXojc
jl7iiFsqea4Bqw61Ky2vi0ztvJ+RgDHNOGbtLFZGRHizVngBF+In7EWgF6Qs48ZgOIqe2BfN2NHa
03w05oDlQWGJRpjC6okbJD7mxxYMYntG1++KaCPjOL31WRggpXIXGT8LBCwxxa16iWyHQ/12Abn5
uYDRnzRQUgdV5iP6zkmDs3d/VXPBkYilU9r7GbiypS3xs5oIzp4bAn6tCVGdJF4QEOKZNNhrjKhm
5f4ZKGFYmc2JWMVdnkAm1GLzsuDiqpjbUe4ov0sw/KoDRoNgzutZh3fqioNHOcuRaxfDlcpAkDkp
xzNSTZu+LHaMtwByXgl3luyrM+fhjuxgOnXkWZ7ab6rkq8RegSQFbeaHX/oAmaChFgaKk0d6K5cF
DWjeyAeh5GMWWL2JqkjD7S72q4FHy6S6I2ayEb9lCmtKLiOPCOMOTul3vBEf3lGVi2QaMJvwvkDD
pfesuEFajZFS8yS7kXb99/07+57jjsAE6BM2L4Q9CWCB3cY254KRlDIIxW+TSBAFNFLxzc9utLRz
b2cBDYkij1szAyXgTv+7p9sHnJVt3D2PI0onPERXAc+PVlXl4kmyJr/JN0vBuqPPWxzUb7QdK7Bv
Lk5Eg4UdG8fidAOmK2Y/RtHjhg47wqjoySBItf0PoKqsX+qDNZsvoLSw4tsei6EQXMmbrW9JLBtb
eWcwyJQv96zSNlxM0sD4Y0He7OIyiWHgA+71nNQ9n8q5Ha3jCcC98S1vGG0rCQuZW5PlEc4cSKmn
jmwMpaL4R6at8Zfy3GTWG6ctOxiUIOohfSE7bz/1ufkY1684IAU299XNgtZGgdqeJxX1b1nKCKVX
rLRXS6H3p15UzX7fdA/WTh46XtyqfmUGHiuIWICvWlyN15efZqLyyEBK7uIxcuak7NqoeAWWZjgf
ii35gJV9e3B4K52GKsRc1ChD0tDN3egui8r6N2MVPeT3uxizGJVhtsrXWsv5tdR+0K6+p9DHU05e
wg9Bid2Yc4w3ACxT5DeLc73tLxwNnjc4M+yxHx+e/NRmOfMaiBm0rkwvnIdW55kzV+0gyxjg8/b2
GdgM8TZtHp+dEnbSItryYZ7vLH+sQ/ev7BAv+D7++Gn0ctGAT9bpnx/yp4DNb69jiGTTzZJppNJo
4Z3DA6Y6Fgrq3UUU8OZ2CDCCbTHbSJADN50OYt+XD77m+FGNuY07XaLC2DGw4uBYVO1srqx/PFsD
PxlucFZywOmhj6NK6qe+rTef2AmUr7/syaa4r68u6QHe5YpSwWmekovVNvtALjwRZl40YReOlF5H
R0ql+1LD4VQSLElxbnTOXdiaEuKHaMhpTWdlVyspFSLyUrwi/YUf/hM+HlzQNDB+IdZFpJc3vt8i
fqlISxlDyZvCJVSEu1SR99bCjYk4GobIP4tgHGdLT3xEz1948VqSb9yCMQ/54DC4giiTsE2Si7Xs
MTry52/czMA/InFAGfWei6KxGLGsNy72zYFSLNZyNOo7OWDBYZZr+RYTIXjsJCVAa2qh8Vh8FO60
SJe/Qo7V43gpK4cXCKWFVkAJSgLuLCPfK/y6DwjbgHq7BZTVfcNliw9DwTj5XxtitpWVFoHy46AF
u0pCIFMH5IKQ6k/G96QVUI1EkrROgdv/QmjowwgOCBatk03nrt9C8abyo+Jko54laIDlg1fYQjaZ
e9eFSQ4E4EyJmgYNBNxh0u+HgsrWoGiMKIS+c2o1GgbNDlxMmKZgKxZ/Qj7TGyKl4Rvo12pniL59
KDnipmMtFjZDMbo0YGOYWDxx5IwaFACdCJyiVO23hDIEyu2faw8a0eJ5D3n6/5T6sPXRsisiE9OO
1BISSOdP0B5jLdz0veiRTzXE2v8f7l7ZY78sPocnf5miuUzHGeRCmPDuYl6IlhN/BZ1m9lt/M1Ij
v9YLEsmWIdx5misARBuxc+uHv++8Ggma6QRfPXEcJvztFrjzS8iMM2IGROPqNMO2js4oSvUHTGao
SkwazHhYl+mz+iwVQF9eO3CyNi2zmNnhsxL339KhW8dcwGhmIiQ7rrZKMd3Mhyoy99Xpk5snXvWb
yhnG9ddk+oglNA6b1V9RLK8ubzOm9WFh7HqMJIZlYJCqI9zCbXTWF9UjFlzuaHEJcfuTTZZOOjrk
XOxndK1sekh6Zaemr1VeUVJlUQ4cXDWVxv0k5ClGeu2Dne33qTAc+CmrwFcXjgYkMkNZwDzdmjY6
qm3p1aRqRKkmgveZvwFqOOGsQVaxTxqyPS62Eua0qZpHYztrMeAjoV+KAptKvvZncwVHCmPa80WS
wP5M3s3rk5ImDucJpW1z0REZGqnaVa4AnxD6H3VHpHOXQjv+JNoL1FCUrTOOvTBiFJs6KSNbxuJX
KzEUhQCmb2Y8+MEZCqbL0QYrY4xF/dtMpZcAErm95M3rSZ923yxc+ylveONERqT8HJ1lWDj980R0
3ciaauB3bPOSRRvE8DTPsFU22knGRW3eq9neduA4hb9pbtdsdTXc3TwJhl+3aU+RRSn6OtKg9h2c
x5uZiWnN2ffn25RfCUg2rPkRceZ3nVWuOT7mn+Z+Rfy+48ekM0mQRd0InxRxSkUCqrSM5ijOlz67
7gRt0FzmcOb0aIMCVWuhy+SdMeUK42EFryDyqoltzx8fSb1M0hI+A+bOi1ordMwvB/4KTzsj6EaN
BxxRdqvPr5T55oQBmUBww6Svb0dTfiQfgdYYynIZ08dFQFCIHxbctCOrqObR/zTgq886gO2R83gL
n1hb9wTC0MTqrlxilGzBVm13w7EzdDjvVQU51dxqcSHVF3eowngqeBJxzPZgfPoHB/evzx77No6X
JASs4RWT7t4dt4gAt2ylF9EdcTL/bsjRZFCb1AWHbVHQM3YONNv8c0s7SXwJtIFZvEpoD/zxA1Ky
W+lgkwoZcf0Ara6qbwC01RxdQONp4pUbkHyON2FNdHXkZvTyUJ9GFppduJwHVqyQJ8JmS2YkukZ7
XvirzPSkrK5Ml+1MJZ3WyAc266vjnC6O3EFEJDvmEr1eguvtHPx2SXw9Z3d4j3JpmzdhBsDByxbU
Ogz0t5ipWSGbu2JT/K3aeG4JOaAQN7KGJMEjKkP96O6IkHbw3tUuO95ENCpFF2AGaStO0asgrnMX
bdgkQC85IAAhTaMKiBg+ce1XTmEdWJhbM7jk/m+UJpEpYfiMmLg2OmWQxln4vjar9tuvQMzjjzfJ
InglRfPxmWU6wF/rM+1HxI2Ba2flNpxWDwppdqFVXrkiTb8DtUyJ1GGnd/HnCiDceqcMPBSWg86o
f+xYtzpnon67xg4uwynUMj3rlFSzOaIE3gox9czqKQ0lwzOK9c8AvvHq4YM1aQOP8UqATskWpR91
AjUohpQdgr1onIw1fDNwfdmcuLxuhIsOSJI1AKw+xB79AXlaH6u85vqQAR4cQGG/VUpx6aRrPc9N
VNANokUCer21yARlScyk3xlWq7rukt673DDebQcstmo/qsx+T/0cwc234RC5KwmZTDFq+dP6u6/G
w9bhnBThf+o7AW7TBVCO8Do235vhqJi1NTPqJFG//tbKo7WyyaK9eOBogaEe68A6/f1CR+rqmL7o
gaQulYUWvHaBKLyrToUn1dMrnNMTRn/YUXg5MFfqGoTjSFvkugYFeQCn92NZaISlEr2SAwFFIvdb
zmQYPZ2EEKNzA+WCBYIafNjmBhvsWJCf2RDqeKagrAChNFeVLioYNWBzx1Kss+wni+qME0dcqIl8
AQiPJGPTjidcYZe28T966W7qmW4+HUk9j7NE4ZCPQ6Dcww0QLweuBryl1hZMvbXgInTdYBmshEDr
S6AIfyHLBD5nRVpyql/sIQHThlJHGTYPU4aGDJ0MU5TK+i5UBMEjLI5iFE4ZK2g+/SIaZimBxHOk
nmATU5I2DJJOLXXnQEwLcCNZxB21NNEIptRAUbMzr1g8GkfOYV0OwMkQiJt2D4Yv3rtPtirHAcCZ
VOW2gGEknEBXI9HHL+L8ZWd4JJ5YfnVhea6niv0PE5eOK7wjdFUCawpp2+ElL4bXeJxYRa7DBkLa
ccS6RfuOv+cW6s1ykqmU+taIeODoGXQL1RXSa2rjVRT7hSoCocNosGmOvvpEtnRfP6aEIccyW/bC
7l+LrH7usdqiXjDozj3uekyxGPmOX8MaEnO6ne5HYxh3GQ0udd8ecb7IRLNRR3GwLeMnVHsEcwQ9
g+tBPflXxUf0GEILh7FW+cAkxTflLkWNiIPXnZIf5xZEkKU4cbtFar7dSkdZMp9fkafjWv6PI4Yf
JUkk+CRM+ySHtVXqcPwhnJ5zpMnCwiqf9mEhQzvd2VYTzbJ47o+1phsWQWo1df2CcecvS/3VvV+0
XoR/ufoNLt9pkFe7x9qFYJTwnMCz0d6xBSQGF3hgspdS9A/YOO9CoKrjMgJnUTxUNryeUWolpwrn
jvEc3s5jcnNcw04mhb0eETOI8CoY8pYDzmiGve3d4Qq6uc8AewaoLNTMfXiLDUC3ACuLei5ZCySD
a43CL2wD94OdzG16aPwbKV7gjEMgRddnl2tNr7SBVD8eCEC/WYq+hrVntIe3RunvFdDCFXgOsise
8fd/loWqz/yDNVZUb0MR9CPh5rxhmDLqVwYmIoqWcKp5DRX/NW7ZedRX3BXS3oiNzsaZshv8ynJB
VdILh2KArbJZcak+2GFaqzUx7VjvzQok/nrgIGH+kyOjR0L6zNXjV/llUUS6K63C5M3eB4cQwt67
6LkLU5KlyqRXKWxp4pnvJZ0HtgGAOqaIezmb+mkfdRPIkfXaY4I3TfGhsuCFR9hE+M2686Y49e0e
3B8v7dwWiKwyMuWPTwEhWZcKtCpnDsjPM/ga6NLijVhkMRSdUjxX1zgctwerTLq5Bi1Mad3VLa6c
B1JCQokGenB6+VE+f1Hmm9to2otEDPRwg/sOLUS2P5W2qeRuLajM4UjhT1WeYRK+lBEU/MRyisFK
hyV+P+4ajLXgjZxjrKy7iOm7Ih8iHF5znLZIWu5l9KaI2UHrL5T9d4OS+KKpOsU3gg4zOUxAa3RA
Cr27U52Lrq3qQRIzs7i7C01klN8XZuEaEaSC9d+lwgpSU1+EOThRa5BCmp2LIBst669jLmeF/JzO
k3diwkblTflyPeFi47f0tEZKIGnvy8AYxKLdkzzLpsoVNSstLRuqDRTHH2+6zmCTkHwyKMeMPwhH
MuV3mwdX5qoFBgWWYfw4jq4USdYYF8BrmHD2Jw9npIW9LRVAmZ4uJBHKBxCy8Ykdo7Fiv2iJ4FE+
iUf4scLlb+WBlk+6RE1ZNEnnAaBXKnHPrl6ePwKeUS71V+AuLm/QhjV6fAHZvKeBtdvaS82Pii8Y
M1+uBcKpst4bfTdwaKe9J0MI8iZsuAW6fnmNpF5EAOnoEmOzPF5x7w8IXBJtHezpJcFH6Ok4a4Jo
kvodxXnuzNfsJ5PDPoSbLzbYuyQypaG6Ye9KNXYiQCBOSEnGlsGcp/aAiSsA/7rT34GBf2yCt/Gz
S7bzqKEggIY32xeXVh30X1e3GQ1/lrHqcZnU1a0F7w4XOTSweNiIgEavIrEyHIiVCzvcXyXq/3fr
LB+1tdfYnx+08+1hh3D8QWo7NVFOPmjA2O3AFh/o0soFxeVmwvq+XY/p2os6ngD4rV6KCuOYdqIC
kybHhzKogvgFLPjuHw95KI5TTsHnUUy1cmRJAf0XJnpH7Ppc4ERA/tStumCKsAhn2yL+QmSfqr/G
pAJ3QcKKhpsJWzgP7OZAfI/9VrTCUZCZ7FHvxOTyls4AiR/Hng+1q88+qL9a93d8PWQqLVzcrOaM
5H7MlRklusLYn63giR7STSUTxFhGu9KrdEy1GFctMBv3t7DIvv+ZyGQKZbRblbqC749nyYbUdw2j
Ef5CSw+r8j0hyLoVYhmVyZ5YADhnnD9dr9NTcEbxoPydpEa3UbQHHutBcT+8fU0kshQ4+iUK7yE5
wzEc5v4Z1lE8BX7QyOca7efhWkEHF6SByhPZnQwHkbCtE0pM6oUSs9LjikLy5tqCwaHmtuKCdOZ2
62XuBKCeePCA6wvk5FAI72wslvdyacsEwaYgU92/24gTz08nS4p3Na9/z7Mb86YGt52D4C7zLdXA
d5XPa7HrsiHWxh2F9Ou7hpQ08ls97FFKj+JlAMvBzOCNFJlHR45FsKe+p+SqZbBTa96kppyBTfpc
g9PmAniGvnBfF8X98R9sHY9xtVb+ZLgl2WyDET1l1kl18m1D9seM1NDJYLGjAD340gSN3wwLnlRZ
nR8xug1KdsJASaziLP86Db9N51dt3oqNe+BX9M0WuJ3vjGCRTWs3zeu/s2+hm1cOq17Pu7FknjwC
zjpC55JFcGZg5e+myjxSV+RO8QXM0oyo9F3L0Qa4Zak46a+R14wSgwnqcNnZvtfXtC6Fcz+uoSMj
GICHLC/mrIMl2xPPJ2fENNY9bBSmy6YgbWIuBYGbS9E4O1A33/F7+9GwvEtjfzeelu/9fFAPHTrG
3aOTtNs4s1yhbi2qK6Kjhbv42BdxmOwtMdDEXsNuyTGkcov6wyAeql1Qzdgux5KIl+dIG133lpUM
sfpkEml5fXfsqIiCGA0toSfpR1/iSRSHDJMgiY5vLg0gLuQ3t+geCacb2aERh/W5HuCNrO6H3rSh
KZcALYKJPs/K9nsmhbLvYF/D44kHClsku9ZYNcPli7UWJXXBOXpnuKmQrnNBECFiUm03MvYhjHRj
xUWY4dzx9R3CiCc5BYcdy4RZwrypLO1T6Y2gSpGVyA6zudBahVOod9yBrreqqwnWRLojlh9dWhp6
HtOfofkL/aGicZb4F4EWY83zz/54PX3Iw/bdw9SXRELk9EktaGETNQNr7AcJBsfyuV78wdxZMUwA
JBStNjY+fZn6+FEYm9bsRb+374M1Oj5nn2UVUKn27B1/00XVG4e060fNJGa+x4N6OB2NCtqkIkzQ
B5NIJYPbWplOk6YLneX/si0FyS9YMzgoDZNY0B+CXQFpkM5xNDnwlyWEsgFESRXRPHmY9KK82Vws
e8IeK60WP2OQ3GaKsyqcV3zTMESp26d1YDWYz4CpiMXV5m6D/sbQ4Cys+tgJNp3jm/J9t2acqq/7
lGLSyMrqv84AoiRgasamUCE4i7JQV5wDLcNG566imtQBBHhtpPw+nTQAV4m424a+7Here7ZLL0xU
w0Iw/CphSI6Hu6q+jw/VUd0VqL72shzPXccLW2+D1DjXe0Mc8ldyeolW9zSPUseYTKwln0R1VHDn
QKk6ar4tGaKm/J43WKU0MEevE1afih0pi/YvkCUT/Bg+i3fec3eeXc42zrnUg7FVHBGuyWfLyvJv
070GGrt8OuWdUGHF7YOSD/wXdmJ9a8uf6fu92uroq0OQjuge6edMG5V8S64dtLZc0q7btNrgpog4
n/A+lpauLfq/U3aiPan7UIW4y/mY1gbtoeChZFC1nd38mvLcmwTprTsdvOQeT/Cak4pjsqbCF1IO
s0OG1uhDoaeabIBoQvp/Pd6ZPoAUNp1BFRQEHdz8mW5537Qj+2A9QWC0RdhyIwqVIdB1wVAvwkiS
o4Pbp7o1pT91/dDFueJlxS0x71ectrdwdfcD7kSEUb310hPgh8Ky/Xjt6mfL6U58zqo8zLfjYs4L
BqilRySUUjMJhkeqKzxrhjYp8R7fQ43SLhlG37BiJu5auQ0M8ZJSzUtjdSd83wMS1lgoeAlddlBG
CIDh8JjxnVFVN029PHDIT+Bdu4xRhBgY50ajtFzJX/Dxu8twnnq26Z5yRc+6IZZUf+rUIeIolBrw
YFIVSxFPGtQecAw/0RrhYBJuRcD5IB2jwh8VTVX7ZqRrS7dWwK4chmqLAXC5Utf4l/QDvHiOZJAo
f0bClqW/zhmIb0mv30L4rVFvzcQz47SbRaX4PjvMQcfVWp0YzpuzBs2w8IAXaVNrOxEBiejI6Pgy
CryKCY9d+xADbFfu+YCSj8t7ad5duFZtMWcFokO5CApTaZ+x1BPCUOFLJHDk0+/3ztnbYFpnuyj1
H44YQuMKMJfEyRvXjbOI6Jcvm2GBmFcCIprJJbZeJKQkl1nUwGCkF2xF+X8HLLEwLJ3YnV3wIBPZ
nMZi610HilDmrOeze2SiFxX7XOjnayKMGasi5OIEVgFo0ask9NnsslnC77gABYaqoR5bfmb3ziU1
cZXxQVgJEw5WxU/BwGg1Ef5l2eDk5Xju958rsJw+Nr6cSEnAFXQ85ig8v1BOSssHpfWk9JQmsWag
aJHRv8NajvYcqmLwLJ7swziQq0lW0XzmKdMrCiybPCSrmS+bOihjTNUtZoF5i2359PL/UdazIDzM
mCoU4zbKZTlXhZVryFrqqcIrGHtl4H4qEhve5oN/PU5w0zewPskTywQPusQ2/UmGo5uaKiYbOkW7
T1NtHIKa+Lt+GxW5cy/ANNaNRFVmSurLrEmYoP8fHUkuonQ/Jp2+wecTwD4PE/BNRxl2gmGix9ld
IH9jcE8NTtRA4+GmeEOmslyua0j0/cUDXuLg9Jd4I0jevFiUiFyUK/DpFjb8WYUtwQrQvWA5dC/T
XfhF/+buMBFHiuvwnXin8kVQPcWdybEJ9aXGvotBaEjpFl4b01oOkKfYBRTcLxKeFQesQgnR4yMC
l5CULx3qOVMc2/H7SYQ/SzWVAm/c5hjJPTE6xZy6JsAZw/Lbz9o+U/bjbJKTOY8HJO9QFkmpE+73
14YIlD3e6rYHVdvJXHu5dfd6nwCRPicu/G+HbhPAcF+Rbxwf/T95hVtVbCXGAqHgSsY8L/bYYIID
NUP/DGrZQEn80Vyuzx8e1VzP/OgB+KKUIjrEr6wDtEWG2jAgfT5vrmQM8MCuIbankd47LFZiCRTA
EbVGu0pWxmNHn2mikRlQUxA4q8XoBqleC6DPoX2q54MCO/a/fh61KHQVZmx87ZS/W+vZwuBiO/w3
WXQbcLkQeGsqBhcQJvWXm+5BCiNGXZL5cZAHLuUprIMt6nj+n37U/R2CUDmvxPuJQlKJIr1+jQkt
nzju4NJR9p/CyhVCnXObywNQbkXiBgQLbM3RMOk84JqrDb3wDVzKSUnyegzWIteSHbpBLUpo+j5d
SUjErVzN9pZiice7eRNzZlb8U5lLFExk+J5uAGN1H8TNfctG7u19u4yZw5na7t2j9GaPGkJ92DIK
3EjRiv0idTdz/eY92yRLQl2OC5n6NZD9ZTf+laPn/pqHzzTS2ce6GcIcGPU9ok1vZ66RGJ5boq/m
D/MzltR+jWq8HSuEaF69mgEzyEFbiSFySG5w8ZsmtrTSeCcEwGEYCndjxcIezjdRtfg/+sLqcA8k
8BIWoVnSYlECVhtSoLmlk2taaEJ5aHirdmn7MhJxyP+HSHTKnkRiJDkJjDi794+FoKQAyVaqAxQI
hyTh858vKb43gG26P8QNpzP8RrN2bKWMCnxjJ4AJKI1ENvjUrhx8dmKucKdyi3oiZnmznmItcH5F
FSMa4tvM+bbu2h4Cnw+WTDK7dmYFtT+hqiZfL6sAaP5AxbTLU0Trxa7eitNkPsRTBXbcN41/XR4s
WjKjTPvnzZYGNK7IgdGEV88v92b6IY2O9YlHDpvnFFoKzIxLzUExAaTCzsZXzIahB9w1LTUFxk3t
jZvDpR7y8LigGWSBUsi9G/MarvfjsGBoM2/pHW7pccR0xbM919dT1hlGmNyXPFTJ6Jw7apQL7USc
dZEsD0uG58YNACUk7Q9tSsf2lSRu/nRG+EjtYxVM2TN2xpqyMhyAnQ6+NUs449w7ZtgFw7zwZLH6
pRSwYEbImwW1wWHKxOBBCmZ5ER3jhtM9sRBV7E0qIvL+VGAYCUD9WH1ojCSB428BbYo8BojWtovZ
MkY8Q0NIVDn4GwfICE90bNYN99MzUjUGDnrSwAI5/maqCizNMpSiZ1vMwJpegRwWV6HPIlK1Tvdj
n1lI+A3ekh6dMx6CQxhG/WJUoFkKDFPp/QF3KnWPcu8gQPbcfbajgM2WXWCk1FziTxISq6iHCeCe
BGhWHNM+lAOl4Zxw91T17jelcYilMA7mJGYxCwSs6uaD6xH1oQKg0OlLtK4LGcGe0thiZd5e+I9O
Y3Fbh/dOf3cj2yWvGi97cx+9wL34euiEA/57jIrMX7DLnkHkZQWv7u4d9PsHuOrKPJlDkR6CQiO1
9dE3EoFL+iMjboOaw8aNEX1Sd++1hbEqHyEKLxv/aynDAbScBfqhgLbeGvW/J4aauwyXtcVLgqsf
RaxXFLdKIbalSPbim5Efq44q/jq0L0rDutu+GMg3ccsIBm9GfEzMZJFBOsanRDC1nnpC1twjmOWz
gZMC/JTofun5T0RQztPOkYiLDvGyrcEmFLzcRfZUUC17JZvAcRUb+S36Nf2vZNHBfpA3agQ9rQFV
yjc2gObnjcDv4RSHMZ+PDxdSgDq1S8R/3srQvLF6BU/aHNI7RvLEM8zw6BVWD9Of0YI67t2U35WT
s9u1XS6++L5+cDEi3lsG0HgFJRxY9FSW+DjtQftTCj941SrTkX8OivTZT6adrFMCdyD3cRKYA5Pt
lcwbY6BYLIE9KK3SO57M18mph9toybWA611JxGC7+/pJxwsKROEbiriDtEaX0dNwz3pmKo7g0j54
MruARIw7fGDc+VdnczDIl9Q2kAfFZgE1oOGdTV7P25WH2a7PByPS+VvyQVLtPB9o476aP1gaptlq
pZeYBGOOfjn2u/zcUvkIs/lCArNF8iV5+w1X8X/NjTDxxLbpo9BU85Q5H9SlimfxZR/Ozg7n5NR+
T4+OMcnnSxmNCIGv1IlLB8DRzACZS2jaIJ01Kk49INt6NpmqWKsZ46SLuC8yvWnpXRHJJp7LMmqo
c+ZSs4+OFWY3ZJHx9Nu+mdIQhhxU0X3mvAO22SJXEhR/k+u+LxK+N9zPtNnqiqwSmL6ykII9wzjt
YnSV7zSIXtdzQc5T6fN1/ATE8JB5JHQjGvDjjh8xFEer0JMTwS2lafYVcFVsqpWQTrP/aRSQJdhh
TPob1OPkAlokDuJwIxk7LwsbC8eKpQTip5R9UIqRXPIEluW73DZNeMCl4m5Wc9cyDDT44Udmb3Gc
PNObddd0nuISwLYnxZObpDLuWgT9jJoz3VY4JSYXrI1t9lDCXbFnPnVSttanVs1Xh5/34D+bEfcq
ZXeBbyisM9F6gLTfH7Jsl3lVfLug7EsyYdKLy/ptHzKvXvs4joQJ9oARrhJuomZpUttjaSqDMpdS
cWWlPhy7SjXD+w3nsPLCyIHLDVZ1gDYPW486ie3TE0Ye0X1BiSTlXRCsqmOud49SHQnXYfwTvgSZ
vzjKH+Ou8KzqCIoirbKcfPi7EpRuLZYdstnLggTNXsQgJEYt61yVr1RBPy2KrkSM8ub2Vvx+L+CZ
h6wbt/VmEuuM8k4Jsm6C27S36Pu3IGBt3aR2H7piXLDifdqEyBhd0+nZQACVfeeXngs3cOVgZFpA
G5N5pCiyDwHKfhKh5LVE8SZLI/7HEz1d/uwu52Sf67aCL4fsT6YNE9mV7vykNvstPm4kUlSRPt/2
KVD0i6PU8O1c6J9T9X8aEGmxUyTCL5Ti+SXMJQsVyAeqCVFWDmFKB+9nxqUaDUyDuxADy/ksYblS
6oAEhga+wtaVetl7FCen7MbnFc8dRd7wnVeCfQq67u7kPs6nYAoM2T2/kkYsYXrAhBMKvThuaJpc
rQYq2IbXmOUXnWrvtasgR2Iwlq5KmcmI3NFHydXv4xsUSFnMrMZ9jdrDHeESwVh0cIyRSeUQ1Qah
1/B0LYr0FpXLoPGIRpG1TW0vYh4WpsvayaLsDHEk9X6DueeGsOnyhxq2krvjSHdz+3rDQxTjRQfW
axpOzttsfYsKWooEOjZbnRW35HrEyrpw1VhXX13H70TQthN1fvqPptaa+59ZsRh4RUKCQmns+m/X
b5hQXo+lGH5aIsZVj6xLYzSnkjdeYDKMZAUUdXndIKZF87J/mCXvXI/8lJpiSjE+twcmQaQqMTiO
Pc8MYgdg0MXzZ/KWSJDsJaq3tOZcvoG1FhW/8JxdJcjWaN0eB7PKoXQ9ggx9R3YV5t1wneR7iAFJ
VyOgl7WwtsUb3t+zfTO84IKqja9g/aD5+9bT6sEgkQasOAMA4hLccA2rCKsyqD8LRSifUP83gOoG
xlmwenszSgjWeZ+or6dTbB9BWpdkqYJjivNoOKnHU1VlnUgGItEbbx3BNBl160SCwMZ1OfGsbIZE
+0jR3j3t1+Q0Z96r2Md5/93jdES45em4WtRcMI2T6EhVp+gLG2EVdEca3WdIQnNogS2zNTo22uiy
dPxX45eTrA/2n8kCcszr4DXbu8mH/LRDIbl/Dw9/jXXlywxiI/tznEkS2kdMxYhLnOYRfNg/5Y9f
qsMBqyp6G/K9+umcw8GUJjalLwiqX3JgyRyKqyfCurWEaqNtFMtQlPZM2ZZPcnUDocwAykz/qG8O
1ujULFfKCkzKLZaLVRhzCtCn0FpQahTS5jUySljQnHOYWbLROiDuFgHTHxVsBuTfHNXFWTAKEvq3
S9/o5jGjeaxlb3OZelPbzbWVDZse2c8pCQgVEWwrCoL24wNSadHH5E+l4gmJ4PSLWuFSsglQfxd+
OBQRkukxuDRXD/3k9E3Kqr+0i1T23VAQbsAUTRD1QCb5GcUkMEdaK08kSOrb/6aM4zGMFlI7yhv/
M+mxUP8DDYFj48zdc4gsa14NH4GDN/iYcMVgoq6Lgd3KvZEKMRNZL+o+zeAmcUsAxZ/mf5sqiA4P
qoaMZ0NPfEpDy4TXBL2ax2o0OSxWCSSFNsvVz7IhlVB0RQhk76ZtoRu9pMCaragb2tc1jbg02lgu
2DFRm8V1h2GeQmpfuKBUmefpfTt5xXNFkZXIMr5XvK/wake9krgbZpaM7nterkj1M44SRdvacukk
lphUiIy7F2YEmfJT6ni87TPqcCeOofBj83a5bpio7zt5fRtvpqc2ThX1RX/aFqoCPK87XBGmtRqk
vqWOa+ZB3KTsoCa8ZtgSNgqvW5IRYEukvQ1e/JCfNzaw6tmmXEdLfg2uavCSbcF/HpGFgKSHq01S
UTEBjKKp7yoaGt7jMwY7StdTq0DGy64ejOApx5GUGt9PWIaQe+NJFeMMH/WDSejbu5mFvhAZ6TGI
nGZvjmFNuVjtKQWfJnvU/bnibDE2RrzGMpja+eaaPliDHTBmR+H+sRYVseado7TWq5+dI2J+zG/Y
71NTZfqnA95SlGV6/ob2fvPZo9EHQ32t5q1C/aHj0QJ0fcAcWErp55WvNikOdJMVGyjN1bcv0xj2
mSqj8Bv3bIvgOVhnK4/IXG+TkDWXvHDaqtRmHiPv9mSxmwGwihIbrB7Bf7yWRn14MuveiedPM9E4
xOzRK3c9+56Lyw/0Zx4RfYEZVuoNCOKBoMbcn4FSiaYCz1n+cTmTwJXPgKfd/acS9XpyFAw4MEsj
R5jx1HFYg0qvMiEqc5mu0YiNK1yfzA3NL2xfbMHdGRw/Y/YOcGJtI+pAb1ZIsCJgftxJIUbLg/Tw
cwHWaUWjZ9r2MB6ordBa2tq8+u0YpKoE6TXAWE7a1xB/KHpNPDCmlbP/m6SOIFCjY+kyPPlBtbIX
yv6r7QTBXbFDRypNr991/455PameaRphm8FFmmKHZFTOFz7z/RxZtqQi0LMoBf/gS/mf43sS6Ti3
lwS7N9RdsMnAJcFBrO1obODQ7HYrrsCO28z8JqSNCcerP2GUzMdtNqBH424p+Pawd/gUuVVymic2
YUYpP7Shz8MrmucHlstZb1fyEM4A/bwEb3SwTN4BQk7DLO8ojHNShCIxTxVOBXw75IX7nJ3A83bR
//tW92IxHdpptmJEZy22lf6gXQl8beTrxzjWqAXetYqOVgqyXy2K85gjwRuU+kY7bT2b1lAG/Zs0
T/iHqpMWlpu6LL8D50FwWdXENVir+KKLSHbSEXjyVbj6x4TQGZfB9DBYo4+kOsMFWfQrWzC9o+qj
O40Iyom0xsXwzHpKj3VUWs4yQhVW9FxRKCwxwL3GQzq/ZWwq931ydrrG3s6R9K9QVL07TRvvhXTm
/8xbRtW84iu+J3et2bPG1hQa8UwoNLiynspgIimOukeA/pnUyu39eMSavuEImMYhZQMde8WdURuT
yp7DegnaXaQbOnbbjakluqsC9R/1kkaI6ss7kJcFcFwy/XZZ17fcP/iVgpm+wP6xprgVu/TDpc/N
jxpjFspA11VwtjiFD1jpRarM5hRLQzsUEKRK31LT7Ug8BMna/jelC0PPcH6wpbiLofmczCSxbqqV
KkGyL+9pha9Y7P5Wxc2lB9sISQ6JdHgWjdmo+uLet7aRsIzUr0sZGS3v7L45IEcBLIBd4/+GNwrE
ZTkd8dsjhWAV3i91gypfvmZFJwF0FyzuHNSYm0EJ9rgM2wJWo6my3uDTCkiCa47eRdDi5fEhCLA+
TQECiUeZE3czI9o+D9PTHOipS5XTHPsU6mgQtVs8QeProJ48mZZhmH+IWqQ4v9eabWLEnPDCQZka
4oTFdzEBIGTO4NRcL5GT+pcJIUXIGUcyE1mM4vnz7OSSDFgRnv61rfK9BvVh+9I9scNcOBIUpANr
VAb2gRHYW46lTQxbmacOzkSjuJJS6kHyDqhvTPkAtdURmTd9edTfrGOKI+k4juzZbBVVjCIrqt8d
9VjrhOwi8Za2Qu3XxTiGUZ9TbQdFXJlMOULTMcoIbYkfgLQaiL2ejH2CbZDAqhdT6Y1AekOxUera
YseoOSYXmjOJeD+aj/0tCmwM0vTJmWrPSSLsP7Tgbv7rCl3DF6H2buutVAVZvLICh4pGy0vnSh1R
cd2FAejHoHoRYpffsNGNG/QWY8KlniXwdWAj9eQTJm4Wp9SCJdnmbITw8Cgyu/zpg+cXy99Fl464
3F/SERswkZzMSyoIAsNKnesSY8pO4ZEVLAbAsYC+eDp75jEUFA4ymMke+irpMZcl5bag6gWXKizz
sEykQfYx8nsRKDsqFTyFlBkXg0ORKj5n2SUuQWs70b9qGMnWrIe25gjbDZ8jh/TwoSi41w6cTLxc
LAEArunSMpLPLfGh7fUoa3/2Hs3St4oGK59RiIFAb8ZvfNxy97Yqp9vixmCODNeULP57AENjpuYc
J0oxogTxJr2INL2a9nq37wHkMa3hpiOpOmQJ3tD/rnx0tTIi+6n+rwlJk6X4lUF+2vs07+44uasb
IMchknLnMWfXlK+NWotJmW7i/slKd4xtTXCuXrUh6jZNS4YicZOvMHID92kun4DMHJ8BKEmFmtDQ
ypCpvhrlqlI8Y+vSl0QLY2svHr7krXfTlAF6cptdJtFBsYQa6MEZGK0mvaCFe9kqjjv4VXrQ/JSn
ovMxCRmYdHyKo6Z/31eYwpVU2Db72fZHzBMEGE5y+dnGZkrXU+3W0UJ6LyDnxD32PIJSVul4RIs6
vGKTJXJDBpilGryghI6Rcf2W3aItiqEr3FKlXI6P/xTE7XXbd8eofa7AY2nMDoVDos436Kjhyru0
ssWZe/t43zvewiCM0XWszhTqJ5NFMReW1isIC5pIHq0NRn1PXzPR/vnpQSfgYuS4N9FFe3Ihypc0
TxImXXTkuvyb7zu96sG2BoqfczK/JF2eDOmpwXLJ9Y3COdyU7FafkDr8ae8DwiJZfT3j5Cv31L+2
ZXZSjJMPDN4/rji/W4bTtSkGibfJ2AoS/xm140MYqsjhWaCT5d6dCv/RLrgmhAh4s5ugbAaHBvse
+zODhBIUgkGRnCgFylJutwc3nPKFfUNb/hXH1QWaYzAJQzOMuHHVakV9kN+thVwYdCp8Omtp1UYl
axFa8ug/g8Mnh0QqgjNxzoV+lrSwk7/b+IOjyYM/0MX5CJr5u3bgF3f76ffuG5rzsfXKWGJXhxpu
ioWeeh2Z4nHNFuS1AcvPYC0uFYQKnnq1DvTElMVwXXcZa6hPmhC264yEEhjN93j1wArZmWmalvif
zC4irGyc1B6SLmwrgciMpciEcYJKukwDPxidIK7mgRtl9knuMK+Ldii/UN977FvIppe/2ho748kg
fX15fTmMMRpbzR7wSTA7iQaH7gabm/rdgOQ2aOvJQvP+1m6haurxrdYWz6jazRWrJKUoA6adIj88
XQ+NQ/GDygWzXId/UgtywTDusuy0cqZTsrQUOsE6t9YMR6+jGx6g//DMMqewQjKvXxwHxwJX7hZt
snB0KvEIeff3ja951/aoKgacM21e+LTbE8Oar0Vft54p5tsJWJCuD+fhWSOHx/cyoVWWXdShFSU3
wjg7gY9kSjcKhZy4r6JUJc42GdNG2xE7UVMkJVz0SiQrv1r9p6Nzm7IdHf4lt+tdOJsXzFP1HNes
xzJDntW1FbdWMpBpvYyh+X/n2dy3Vy6o8FiKuLnugBiQFOMdZ6GcS26Zr6UVVcXY301ns3Iyplq5
zNhNGXd8n4DHi0So5Jsc/cgrfpOaNrtk1pTeUuUWvTJo1H3pjd142cJA+ACc7ziQMoBuGjhmEN1a
ZmfjkfRBirkgmw/okfZDaJW/yRsy42dBkrdf6CUZuuhPKpTQkIOA0VzDccUqwAZfM14XBdullwqp
w0gbS/otb2cV73Cp9/C6Q9O3GeMT76JGGfyLzZDGWqSAee2kvkJ5nTBng5X7pY/eKVTu+my44J2x
/JoxrakKd3XC/ZhsRuBxO/VPuhIxEprMx7laZu72SRLY39fw8bPTep84xL0ndyeStdZXLSkjzzSJ
KjrLWO7XKwy1jNqmz1S3Prl5cZa0zwvnXpHWLRyavn/hdh2jQJMJ6l3i0G/112KWSVN4793070xd
YRxd3ulFnPLqHYu6h/t453bzgaby8Qhj4+2shRGfUiPODP0JOzFqPOmtpk27U7qrKZHIF2vH8A5F
bZHt81tFV8/8Dy2nxYbNabbgYYHVVa12ez6L+hg71xni1L06m2KagXaFNQrHSmPPC+7Jrym/bDXE
24SuNvg+l1sRtxGoh6ohbcjoMEQ2S1InZ0yd2EvnyKm+/meszyb4UR3m0I9tvSjskjYs73aVYH2R
Z5o98NzefynNIdm1DYRJ761TpxqdCy+x02zERyoYV4h0a3Z8vtJA8dS6o6TGUtblBYVC9jKDLUQo
WTOkQK89poeTV08/MYfEi9o8x43A02h3nE90k/KfKeLeA9I5BKCQD+Xn8i7nwSspMgQka+Je9DhW
0GiPhfI7PLUweY+77wV9jCemD8ns9mk3vC3JPEu1vOlIhZyjHjqS73yN8JBY1NCvph58ZLd8iJcN
S7hpYkyXSxGbvq51IO0/FVXwOBLok5qLZzzMbBd8IsROvnSVmrdkUTW+1ekT69D1Slz7cHEAY8vp
eBKTVkFsGpm2V5wZ/HQYhJ9vp+QbUMirY4GGfDLhhFTK4Xz5Q+AwHNVavEZb1AlkJ5Cec5ZQcFlT
x9vVrFEeLjGwuHNLg2wkV/Zuz7HvsdNA0DHKnqZiVvDvwMBK2ZX8kI6v7ouTm9y9JpRs0ZlZ/oJY
yqVM29R28wY2jETb3KR1Xtt3C8RqAl9bmxqVbmk+Bf8s0qNBQWeoiCkpRlLEFMsmduXVkbXlsUQ9
0tQLMPb2gKINGD1ikhKAg2t0nTEuy3C+B8qlFObeQi8u1QgN/BIPPpArK1qFAG196ahpV9qGn2gl
Yonoj0qX6yXGPp0GyjyVOu+8+oNmvZ5vILEXpb4kqjToJhCz3TpOBlFaJHSwLY6f+hY9BRFgFtG8
RxH4B6nAWotsjakn799lyxCtSX4qjF88y1SWjYUflXEfo3MGr9J4e6gyxX3fT50ycOL/4js5iMfi
x/Z6MbnSDjDPx0TAD5UiyirZZZESEs5bYDw83rg/Sk1THSRMgSdsLsambN8ZRWEdFjcQc4UyMbgr
pS85f0+TjRqPI1VvFjzSsXqzvyg/u20AYr3ppLmcUZhHHVz2Rva6jOihyAeuZtoD3WPUDcywitkR
RjR05AaSYFfQ73HTRZ26dY2iL7gT4Nm3EoFe3k/Tsj08EcvRduF3zu4dvfGXXWw+XDQGEw/mGd85
gazAbSSNTi5ZKiVj6N0jQnO8mMG7fFyoxsrYvXKrN8MdQ8O8JwuPjcOaZBotfx4EITy1yivqwizq
Tr4MbduvEtKnmcr908LifQ0d2yBYoZKQJPqtOB3674dgwfS79KEG51JhoXW5eVMP0OGU2kdSEdYC
r66L3nECM0uZEFVxiYgghFEwDc7cFGmdLR5OvvcvjzOt6IMue9VzilERu7/UlGUAWEipY9k0thZ4
gqHctVhKIPKIHeJcEo5AXoQW+gQIlphw/d3S1z1HSUtA9JV1Zd1zaVwHSjyoeVLKASH08UHYliWd
cR4stT3nnt5so+jYlyFhR3MP1wZB1k0bvm1LYEJ3h1UXkNsGPxqYZ/BUP6Kf1iQUzGYk/353jY3M
vHqdNCpD2cpwlLUaxyB/CEI4Az/neWWzLG1+rLo1acEUOU59L/0qKe77B/cvpcwSrR7tyvTwUF6A
icI4dZGJj0gJqemToa8vcnvgg8H1CgGxVTrFHM20GmuBbApIf3BfVWgPOqR7Ao6YmSRga0U5tWiJ
qYbFP/jB8fyroFnWWEEfk5u0wtdEgBauanBWxnyuSjA1Pnb0flh9cSBj8ElVLdLDkeoSBMsMizu9
FGcYPgBmEMB+TILs5CzxuGN/HtoOQZsTwS5glMwMGbXAfECkE0UmP0fIVRL0dboDa1Yk9werxrC7
QEGzZSANbZNkiXOg/giBrIPpCPdKxslICBna+5R2Ph0yezUxn6y5ZHeUkWYNusXKeCHoBFi68ixR
psGgAiMpyI2/mgM5Zj6Qb+WRScwvx9JYGZNV1m7OY/u6z59vzeMhBDH5eDHnpCggv1T7V6C39BGL
dvykYICpNcgWcK4OG2YoDGQWB6qVzVlK39eSmHU/cOG1Go9sEzPm5MUITBegIWEesCBaVPDfvSM0
5RtuztsUGPJTJZRB48yvLQjq3cM8W+GYqWj8Nbax0Wwz2o47VR3d135xnVTwyt5QMvgGS5YW1FB6
TwpRs3tG/YA08ihkaYRnGBLBRyIft3KcnPTFGkl6LOEZvITSL6Q4qHrGo0dKGLZJgDdhq7spLUGz
Dl/tLU+Q/P6maVOcJBKhvgR5il8N3z+rOkgvRQ7C7JntxQOvqT7fJ2v5vfz8SRCX0jmJ9T57L1jN
Zi6oBtncYW8aCk/g+V4+tFrMi5jxud84y+wdRFb8Fm0t6vTq+uwXubuekwQrmPwnQ5uaAUn7ch5x
Q0aVLFxfBbeEEV1bo/CNO+COTl50GcZWgP+QWfP5R+8gpLGSv+GymbtvU2Q5dA6o5TEwbVCHfdrV
S92oXhsA/m4Gvvq9klXSqlvrjqVq5gnxehTnhKDcii+LLMWpgItBur3JwAguiaCPyvYhJqwdHRwu
suoj/efTPDLlJ6Qtw8ts1LpizkxrbxDzaPSjfjiN5rSbR0TFBK6cCQ71Gbvi/GOpPpTS5gFy6ktx
Mcu/vBf/EJpIR08uozuECQOE2iyUbQ4mC2V1XoFhLoevKFeQ4zpu9KJl8SWgmVDbuJd57mVbfthQ
+GcGdymA7Zp3S0+LHr224O64f979p4+ZncPmhQhi2LZqVyr7ToEdaaEL7dyWgjqpVl/SsjEM96rj
0qlQwWVlhcIkSKN5qB3bLVpOQD7685wmtGSA890xmmzlfkkTMh/3HT86S/abAe2EnL8XdeUiaU5i
IBcjOVabFDi5Idp7E6iO4NVPd68uV4UtwXMhIItwC5nODh5WMFvKmboaJRKImaQOoEecSve0Z/yk
CERb/cVUzpBMZma4h0eaMa8Yb/fNHQz1XKslLF3xMr0pMQDdn4bx8Q9VmWbfiZdYqoIZDUY8Z1u3
QkwWhPqQ7cf7U2a6PIt54m6WOfKEtYrJuUbXufek/cAoiZdhrY9SGjqRsg8HMhFB5WjPCbycf4EP
vcFLAy++mUFz+OejrNphg8Jkw/KrZKPnoPM0FwE3tqESRsMqeR4diT3eNimE548FcKGnJFa/mbgt
EtOUzqZiE9uFdqV5o8nPvXRJL3ilWZ5NlXRrDg9TMhqTp0GERhAnvh0QPbZ9a1bJkL1Pd/je6fXH
tdZqTkFaGCG5o9wFTqnpvEVBi2096Zmf6hVodp9HCEAB2wL35/uM1JZaAaKU5A3eyu5OPU4LZTWL
+NF8RaKl2CXtV522/MAFKGxg26qHVzEp+WU5AidcsW7C0+1GN/4tsv1Z19pfooPJSYggL/bQt55v
bqOvdsglYmq2mQX99bY0tYeLD5LnLIrVzVuUGXaOOo3ZoONZfTyy7xXAXEDXR0+5VzIQv8KTz1O2
IuDlEn7x2XKEU3zK0XaBMrNCmH68TPjJZbZGrx7WB6aeC2edMZqY8e0J9NZQsU9xgocyhQbPMKEk
KrcHDSeXMfEq7qdeiwZBwl4VQqDWOOSLbStVAUCgkEh0zulbLDPEBOeCHvwe6pMO9cvV3ruGp8te
KUGU181+1n5MezNV+sLWLtPDvGfbyPgnOskUdbelzjsLfahoqz0NS8wKbnyR9QAr5FpiPP4mAnHb
RNY2gl+ziiBWmU6LJoAq/yYelDI5T1ewvWqEipj2dswDr0Js3CL72SLjISimnNISqWWT9l0DNBOD
lF6cCRJJ0/lM2SbQEYSVikA5YX/C7qXT4KW0Tfx7YvwOSi+6nxHrmNGwWZ6zEin5CKKzIjFy5dHG
8JKqx/+BFr9NFQYdW+O2xocPNOl6QMEEqs7ywH1+apTKHvNhGKmFBPvvWtEtcfjJ3mDF2vxlap3Z
tXyPGOoJca32/NWXFZpBzMCT9Z+7YJIgJXSjeBip26z2QGKfCAH3M0BFpVJXSsuUEoIvSBtRQOsj
xHCS1kPFYC7KCgYdpWeFrLI1BO+tQVVqXtq9q5KOtd0GFWlO5NLagXm/jGLJ+h4GB/qVdsyORpZ3
Go9W1Xo7L9KrXdCtYNpvy9pyl1srv6sebGHHUgtBmED+zhqHQLDDSWVRM2o5Rt3MJda63QD4E0rl
ECyj9bRPtqejmde02fx9Dbx5TsjTVUMxKycYGuQwNoBT7BqdBJR95VpR+zN2seOG/Eeu/22KmDAK
J7mrErdtz3FsAuue5dldse+7AUeYEiN0IqkYdNOCN68XezJVBQHAzW4nOEZ0TgUcOfAInDVYdbmz
36XnczGGT2hZ6ZB/zAuTfMWxArqB4iTcra+mE82MAknhTcPjRM0xPomujct5wQepSPybh54ErsWe
TLYkOKXu9UNLfrMSYt9tWiHd/HC5Ny5k4BGF4cSbm4uZ65jpk+j1HkVIQcMGEYZWLggDT6HSAw7K
OPOjKUzpYUVpzhpI/594Id20X+/rZ6gKY6ehgVUYDgemLosGU+QgOHRZsrR6dzBu7lgTA/vNuhNh
Eg20c1opjJpVjLra4UmIuP3GRNPrBmo4gSpIHGpAtB9XeRTyLI5+6qUV2MZWqaVRj3mjtYdm1P9i
K7EgpBhBoL6fBKDbSV5ISFkmuJvcyRARrNAgD80sf7LEIiy9evmec1ZEzINtVozDb+S1afbnEpBw
INO4y5hIENUvbmf8rA4Eb+6O1BRao94J0nRqsK7KlTDTkFF0pwXzLjIb94dT3Wr/i7cfUHrp98i8
XHHUpMT7WjJHqXeIIFeFidb42hIoIRir+JGOvyfJnoLEygZBL3S6LznMJl0gM1kG3oxgMqCtLoIo
tI6OY5OxQdW3XiLKcm8677W7oDs1LAr5SmjnYdRKw01x1s5LvBNOJZJAzmNEhmW4qdalt4zIhGuG
G+3EhemFZTnlAAbWfsHXy49EYmkBITxVfjyhlK97Kp2974u+NHeRDqibzl8J0E7y92ZWtYgbGpnZ
OAQ/sT7PEdYIQrTy3GlgTbR5D/FUxCECkWf8ehihq/F2dlKRwHchzeRcWGkagDXIasKJLuH64uJS
NyI6957sdj8l3y47QLqFnKzYV/pbdpIvQMveoNO3BaRUb3/XMs9gSd9qIJz8M9sX0PrmgW7muvpl
NpH0KNuOF1mXEcLaZiE3kIBp+8YbArQIwD4uPXho80SLgnVGp/xctZmKB8SLzjR3XtWGvkGIrAuF
cP1RitOl5G9c39ih8Il7RpG05xU29vWw+BffbHXeMHhF1Bwu7/HLNZFVVNq4wJsVu4ZYi76rOgD5
KwFjJnYYPenSx6mTv+E6V+1sqPKWnrpxEm/92m+YzHjPKUI/t3x/p6uMqe+wdNUyVt4GISAYAjY5
tEGYykkZVQfOuGTOLs6wE96ORv2DW0jeTS8dwHuCdaOLuLGtmgmsfqKBPKKCWLZoQ2slovW5bQ+b
1LfM6eQXhITfuNRDWJXvOq8zEf+bZLUzYg8PXHggGiy9Y1JpRvBH1sK1/1nuT9xaEXh7+W/khxaP
m6IeJqUe14dNpD1oxLWcQheuNUNyLr8MUnMzSrF+es2uSnLrdOI7WgCU9Tu5mj8CGsc9RlnV6bCb
WxCaXumU3+1jZ0pvQ36L4AvQsxXiTdecKx4uQeDMWT7Tf7AkXin9iNTnBZgaFbjUjEpEBJu2/+Rl
ST/iuBW50IphNH5PceySwuwUxmMr9Nq/IhBX5JCsVtuF6/HJyN01ediets7QHsqIVmcsi3h8sI8H
WE7rIcPLlQhpL/RCnSWpPqaN51jyDiHUkMlTKBY97T/jD2v7Ure7aHEf7O0jLlWNS7DFFOdH0CDT
0w+VNpPuWlnFwYtHgf7hmKVNoz+UCHM7M/hh0EMxega9Vvd/7msFf/J5S2GF/Q2B7eu1mN+mmp+a
lU7EtpITN46t5Fya7Ms5iRroS750Jw4S/1F0E6OkH8oyJT9C9aAzMDmjsspbdRIv8ZVzZtBkYXgM
LZRCvdg8LtCKD2CF6c+uaqKfRnoxnPFPtfsl4D+9IJl6rEvuXFrE/i3/UC4IL4hERJlWeqK6psI9
YbCNpkKEewh3cz1wgFgw5Kz6W3NE8zWRfA/g+dPp/F0PmbTTLXBXosx0m+rJWRoDyvCt/nIppDC8
GHcJeuqh+3oBgbGGZkvjXr63TN3ACce8W+CFM15piVtANP+dHuW05d+mydN9WniQMQao2wmMGc1q
Nl1beMilnPLzotMpsexxB46r+CWj4R8XVe8xmtN+Azcbnb1gg7sHnmpB7uxXtkiXDR/JoFekguYX
Ars0TtWlHW5wE/tecZ0B83sI4BbCYm204/vnVCZEr2vlD37FlNCbasU57jdB7R0G0lHd+oxNfHI9
9FqYd6ZsFMDiHc3LUfd+a8zELaX6GTMTWW6jBRJQwzKl3eZGwJQ9SrweXXM88GjfDjtmFBamLqWh
4jvFSluWneDvaHoOt1VkfLyIcvp+tofWUpTFr3phFtFB/7ZG4ZYFfzvGSjMTXm1SJp04ROlEn0io
KrD5TgVGCRj5OvpfRjuwNzcYuq1EzMD8AwoGxX6YIwbrBglUTCJwQ+xj5MWeb3DMkn0Hc0rEfHiS
rIOjMywfAhed+tkX38zihypZTLo7VIKr2WhCvOX2jkszjx4jo5YimnNMh8it5wUEdJYWxWhv6DWu
I3QBafyV0mbeHPZNyWahm/9h7UnjxRROtiXTVjiANYnpMc/k5XNmyMpiP4dJHsp+ZBaJf/zGUjDt
vTYijH/516gXN13snGYkCOuKr2MfE5DOl4SXAXG4OhFnbblS65gWXo3A171OOqmpyKbEmQ/lrY+Y
ljTPzjGI7iF22kWILY1Y5a2Bl79kKZkfdueMQ0UeoKSaZjkyfoMtu3ldmRhIgxFweohA1/i/Mnqj
/NTgyH8+r8nTQGts1lqVwU4Tiiq0U5lEbznzZyYwMC+/4bumu1JULAiJKSnzmNIhqwWeA/+YQxoA
CfebypliFfWbMSB5+I39ta/N2KEANuot5pUOIg6eTqP7X/KlgD3B+EDy5mUVbcJEshKgxBn7VLiO
B4JGMFZ8ixWcLSQBCPWwDk20QErZG1It30h59OjKPP44mwTibYxUmu5ATSg5fa035LzS/q7dztUD
NbzI6XmjfBfrd0napj7V6qRzKAMzGDOGIpqyNKLwSLiY/ojou0PA/RNMZoTL31T+H/tb3zqjt3WS
CEFtx/r0Rge5R3LHjbPjCdcMSvw2Y/w/x23wfHhS8Xs8vsvcgRfe4uAPjFAlCYZGbT7xVtZhdCKc
1P30z2cioCClf2yt/hSJKyrgw5JT4pvXzzP0ysDP++6igc/OKmfrIg1itBqygubWsQhU194Nkb4U
8NZBzPE51n6k0hRcoZYRLkXuJReLgHQzQdGEBN84kpAF3edmVegF7SV7LHC0goBgsRl9TSRjajET
oZjoHx1lkSNsCwi04MSSQwQX3iPLSTPd1s9E4/yt47srf2A+oVXyaPPlca3yICdV6/62a9KBexen
2Q4t3A5e5qj5hBarV+EbA21IANK+J47WBLg6lUCrkRw4oBSCL65xxME5tYZ2T0Xx3D7R3f0Qe44F
C/NSBxVzNzeyikZx6izBokkva7ynHqYpihC8fXSwVoC4Hy2bf2S7tYBY5yxzLEs5kzyDXlIWceWH
Z1m4T/NA6jw+9zdm8gNiPiprWr6QNO+r+5yIIgI95GkvSRdlCpmDEKLHQnxjiWbYqbNBP2gYn+1B
FTxK5lNdKdyBsPZAFvvt/mbA7xaIcRLvOpgmWZm1ndOXsMnjXLg60oVHeswH6U8+L/MRK9M97Euq
Tz9LFqOghaBtl59j7HjZfcB5qDPsEy0oCDIdFN2qsM/p3vPZHvOL1DZiydiw55CjxinxsapQcvnq
2iXWAfsOo7K9xntcrCQwH4LmdDXMl93MVHcYkvoODkcqN570crYr2Pst0cPx7Z9pYMELY4UzAal6
XQGYoOSbUzlSeW6YmkFcDpcsmFOSjBZWnUFPjxf74B0Q8FUR4EUIMFGSxJQXRnB/i95jsXTAqN+0
9hM67c3qVPCmBwBxcMDplk1dA/2cKAlmc/sNYWUMkzLU1R5pxYYM9riwkgtTJcjQeWqsXSKF3RCO
XqyqVgl6ORqyISlOn2cwMsI1IWkG2SzpvVNzSBLctgsGmzwR//DBm+ga8zup2Uzr6yu5jYvbuNTS
3Q9SlNTzjLdhXUUs/OzZy959nfsxZ95HPkwULESlOn3gBaCVAry8ODuhxGtco+z9covribnlb+xH
/YIgoBidjonnKaGNXQ94syoAfFFAlD6MpoO+r4pQ9twWG1PiYCyz1/yOvnjHStlLHN3FM3vz3Egj
LK3OG+HgayI+fkaqu2EPc+hEL/lQEAqdrTHd7i0+hTmVqjigmjleTSh5bHX//26lx73S+nIFItop
6e4VbWr31y6/22T6r14DKCDEg66mT8XigNwswxVHq7GXqx+hHHazg2+wP/koyhojgGKGUNLbQEiH
HzsIrAfUCA1/zOC4goTKqwBlOcwuKk9PzgkL0ghQzRNvm3c9NEGZ6DQ/IvcwGP+605j1MGjXyhjF
E2yq4i6+wT0MygDHiEGwRq4E6C6kFjDopunBf+5r/QRcQEACg/0tGwlLdaSG6mwZQyPnv9c/b37U
TyXa3dbvGLuVknId+23c4xercuowqBnBaCs7MOcLYMKDv22KDvjmsxyrLREwrtapVFt9706+Iokc
+bbRAMxwg4YPHC0qBfx9adT4iC1eAGP73FuhmEC8petI6F5LxaV+vHwpFqKY5zHQnejsN/2ppGeO
t3txIUKz9jSWvuVA3w0IkFkO1wOVJCkvEXK2pjPN5RO+3qt+55Uxl2KurfIJPTT9i5s8bZ6Y21PH
SCifx9RNu1ky38XMZCs9KutVXKg8QUMwFB/25gTszI8fkpDAoAm+tw1wGUqJV5xOKQ4k48m04lPk
1kdCvDq2NeWbSBPYrbP7+ecrGv9UZfUR+/Q2Vjzzox2bkwDUcyrlgD4riQRd4bqBBCQzThKSyyhE
VqUIw27W5UhRmc0ZXXeAxn2+MVF5oM981T340TnC+R0yecasANsof6EZPyP+1EoIr1oqvNk21b2a
jwUQYSBpyDbPxfIfHiXSVu+N2oECkaLbbPmca1mRzK8Q0X/YNaHx8vyYuPAm3+/3yohdGg+AyTR6
8/7gVy8+6sx7yriXfm7aYhx27+VfnAvVBxFWs8mnMcIHFcz7u/Qm3cTs1pMqZZ1fxxE4QoxZ64n1
xzBfwUwzCVqCbIfiIWepkA5eoaAXoX+ZEgjigTsBQrAj2k6TpK5c8ZcG48wW1A0Xsxq2rZOdGE/S
ziXaheEKeA4TXt7mDiDJ/v4W+CLBcjmeEQF5oGpZ2CuZ5/BN8Sen16FH8gzrOtBXMfgbSnTeVK0l
XDBZqRiij4bir+EqrIls+8gucsaXRj5vzKNo34Tiq09sukcj1qv0wLAKPk+FSvLpafO0+IZKBOVz
kHZF7ArLu1rZZ92dsh5m4dbJXGUJ68u9oCyLWlhvQgnz75yCOq33PATD4fzdiJS8GAVGZICyV7gN
OjfzD03OitM7R9ViYMabhalyLMJdiiViG3J++EhaThubAukNc9EIsNwIWwF1vxXA515p9w+HFlDX
dxDw+smXACibFINEgxumKTXyBndfMA3xwgvr1v/wyiqjxcGOV0mHRGaU+crLA8zZg8AzCh+4pcHj
AX8B8bNH87+EzXWHdPNb+QvTmbEU+V/HZ+0b7RY6/c7wipZhk1z/CrFX0et1KvzKpMEAxS13ngJL
sgtES2zg65KpKwPFM9XZjikH449FLRTRv7cVdIClTxlQ6M5V8s+SgguSCcbuyurQDCqWyo1mWFN+
PrClNw7YR/MsXGpcCeAqI76Cok+rUEr5x4mhIJLIN1Z+KGMr4MkOe0HS8HU5kVWbG0UkziNsl+b0
r6IzQZZy4pSZKEEUMq5aLqCZnlUt1DaLFx2MGEikPygkA4qGbwg9IXAtnxfvDBj0mVU5nLc+q6Ga
53KbBYnv1+bRnyGNnm323usr+XHn+dQW2mWVzITwPsAaw+U14qU7O/zAMAePWcpPOCaDFHOu0EI0
MWnnVS3BFYdEKSYxXD6X+yuz+wcNfzUcOOHxUgQU1WIqg0dRFLnd0kMhmI3L9cHhMgaI6/m0MkDi
v5gLnPMBKVIGJ34c8+KR/64w6swxH0X+hfsCxiW5Y/IIbRN2yV5ftJyBcR9pj04vQv1fdLhiTIaP
g2U+/A88Q83bN4scvbwCJRt9+jKb9j3e1VqvxQOqYdoGupg1bFV6MD0Jjmix2natihAukrli7U/v
JYURohsxhMR8Dw8jA68fr72ab9YPYNgtES9irlwzzI9b4o+S7aIj0QmZUBgwTTr8JtbEkSI/kvyS
UCvtnsB/lDBKotQIDQSyhS8HLF3enXZalxXPmQN+uTDT/4QqXVSsJmsnKmw5/5I2hfutZZiJauXb
Hmsu6oiZR2YavmApGseky9r/GJDUw55F2eoZW/Vceg4xqne4y4m84qJo5/rOtSgpKlVuhEkl0lgq
Q7Cd0GSS9o6mFR+5Lh0z+CswYGdQeQUzq0xgm1Oh4jbM7BUjzrMi0MbupRu51iIOo50zeL5aot17
XUfh9+k68LtwLDQVziaigrdoS1u66RXZNdD6OFRqoM2CDis+t9OazgGGIvxwiBY0M7PRQLHFTG8Q
4YPH1RCBImsKKVUf21gzg7RTAFki6TQ/2/8+l0rt96fp6wegRCT0NCw4uOIbThXOIXbhmNEroEhj
/O+as2YksWYMOhiK4R+rVavxiEJdXs0HFH9wJZpu9q5kTde1zW+3gSNnMIIHSWOkCO694GAzg1Zf
fAYe5jhKXIhN156Tn6wnrwUOmP6ClKgt/qwlJiFZMacjt3Km4DKyUFFUNh/+y1/Cl4Ed8rN7gwEK
HdWvrVxSX98Pa4gaUJoCyDAdFpHlRlxKd6Jyw/crU3cgMKX8DGeR75NbdPAZpPCcuL8NAnrYTJKL
DHGyP3uJYouUI6RIMCaIBRlK4wTyCuqtg/tPJY4X+v0Dmx/VQx8B/WrJNcgbQ+1YqwUTcblcXa72
LPqvkJ7qfsQlCTdqqUCBKHUnZOs5dyXxVPL2H75nhftA6iMGBpfpJurkxEwdSursPepZ8Qn7OvSr
E0wQ/p4+xR8OouaK+Av/xq4LeiOI/XZBLeN1RwCZQ3URmgyZmGVlcjWbaucEKTDgACyDq+RTh0rv
V1jXAZh5kFaIcwu3WSIJ8mnJRC7g+7PAa2Sfh1D2Lk9+Esk6xIcOCBoRQr843Ns+FEnh37I5Be8g
/tiBBMDzo7pVsdj9CvZVNKR2y1Kd2hzrTuiRUlD0VMlzSsLVmx9mx+PpLNZe4C6WXZr7EM+KeTEj
sA5z1iwf4LfZu7v744VW3eVRlnB565WQHh6N4sUaBeRMjAGuJ1NwHVgx6ZfY1DZfVwm3m52l+2Pe
9FAuHVWrHOno8IJgJMinDktrlZLXfDz4+esyWFB2ZjHd07NhPeXg4aWgO2PJiauuQIURF30I9+p5
bazZTafZDsh3ixwruVHK173Bp9qeC/fIkV9J+PWfY/a/ePNF2jWpf2XC8SCkoAtk1B8xAp9p5Q/4
Xue7/KxhhXbeCZD7/E2wulSDNtvXRXyTtaMSueo+p06BDtkTjsWc1+bT0lWLenMEQqbtWJgd6KG4
SSr+dhKUZ3Vdl9kkLaks6PHnMLQ6RISzVTLz1yXY5AU+R8fJtXKolAMNXyzDbcLAJ57MRJMER5iv
GY56ZDyuBrTI37evoWSubmd7IVFrJmUq/hhaiEnQ4v4tfkopYfYr/+FMyOyGX5bgL154y8MOQmd+
LeyeVMaoun3vB5mP2uBTmiWUCTswaDMDKz/4Bx4SZD5UphvUPlENeN1aWKLdNB/dDjw2U6zaK2XC
WYw8TkBrTzryZQklgZzI5T/ikCU1U94r9BQwdGTt+TfYkqiH0CMvKXQRQk5Ua4Kek6+q8Zsod4lT
joKZI8bAJ7UVtRMuk9x4wQAcIk2afCgvAFq2HqpRspSpgg5rnLxuUBhkCssLQr8uNRUNXe2euxcp
5w+aYg5ZUDcHPEhx5+yJKaRnKIQ4x7GcM704snS5MxaIKjSOZ2Z/WNnIAQaLkmMWBr9nO1UBbiqv
SZXRUxWRi4At9yJ4Tjtci3cGHtwUu5UaK3aWotWMY3yE2mHX7DJ4+WgwLRVbrTzxG3iJBmaPDsgA
ogJs5a5aw5l+HCROiY6cZpfYOpK7W3kGuPwMprgezwE1s5eBxvvYv/14AZwTAFHdgkox78G8vcf6
FoVukWUwUsoG2ibqqebivCd0bAjLaSKlPI1Nb6qqAaAOduzzzqcfKYN0tL+e1KONHEqB7qgX48Nl
xvxLrLGV3NGpFFNsaHTmHLd80jypnSTogROJeqO/VU3mFcJdDf3Y16wSfhjjHqmZNqIZ7CKQ7hug
SrasGAm+qVPqBg6ZbnJs11cucyOuCD+mneVabwMnYX9HRno7mLkU2GesPkG3Mr3BdwpYIwNLsMmg
an8BJQYBZwPZ1ZYXBYjNoYs3oMzJKdQFSfo9H4C7xJ4XVcvxZ7+oD02v4jZMghk+JW1WKkQZUkAM
tROgZvLgaF49rkfMQOPY8RgL5Qp3VNW5FeH6wX8Vo/Y9XbNbCgV5PwMvZyXvacjEAvdKGj/OHxLc
pRtBH/C16DqE4fYWAlUwvYLJlEdFySZ8RxbuSQ0IpWsx2cV/P2xyrGUGCM7daO5Dm5JKoGh1kgRG
onloC/oeLR83zX+/7keXMkXwLB/O4Iks73vaWxar6/f6gxL2sXbQS4okzYtsEzEpj0ccWnTvmqI0
G7v0t6atsVCap7DijFJeztZA0+EbY2xFklhBsFb9Y5JaCEt7k3PIUx/hqqA3OJjsX3oJF3J6jYL0
ioSzRF9oId7NqIqtCKtue+SLC8orfVc1NeeTdYLzIB15DvMUJUGM0Fm0uc8zt1vzWYkRoYvU6id9
c9E9RmstTHsPDZrDOFq2ACDe7HAM8+SlvbGJsZdCy9v21BAwWjpz5QoYCBCvqAfMmPWBvAY3iUwd
YxgdgMhXkURmaUEesjUq59Ri4CU7uSzxjp033Yg3fWHMm6qMvWTMy9bSzY8cFwTnY5vAwo0Ovc0g
z8ROalPZncnBVNX2S1d3gYpMkLQQaBEQ7wjw826luJizPaiSy6MxzHeSUmxuEXGqvTW8Temn53bn
2siiL7vjpRrLcaw+sVnZuQxamIQVngWqO/b8caYDA0duNylBx98HsPss3h0zO/nAQ80UYWwD70TE
yitS3zfe2yFT9fT+CU/ed7yFvHFPtqAf8D90iLDQ07QVRi3rQjBPgNtsKn1uShN65+xfMt/HS+MS
m4jl2WFbjFHWR7co9szcrakjy+3kW/XiHkafqHiA2iQmEaREn+SpLbU+ay6XjH50gcJ8D9WYUCYU
1c4UVopfgoryCSx+qvex3WwzXz7aGwWFQTPSxM/eA1ZjlA1ZvBEj8Z70tYXJFF9TCkdRI/XccWHN
TSubD5tQ1frSynwLFrK2lvdxcPa1YQjjXN/ZJ1c3trHb1SFACRVF9GW3AR8QPCzbaVOw5X1RMtOL
i4HlxXPJwEdjtKY2XB4EuKGO5w2qUxorC9pjTvwG4tYod55hx/S9vjRVa8hvdLe5Vl1mBJX8iH3v
j7QsaKcz+PqYTg+H8G0x62ZLYR+mdDmjzh1+/Cc1GKEMUdzwjgmyWTOZaAvK2sEGemF8b+sKsq/n
ogVffpBiGNa/ZoWlnRflQQF9lh/T6qX0HHQoWewUYg/tPswoVvrTilujpXuMa6BEgMMEUUNzva+S
g4aaLQzBtj/1LcuacA9WlK+7VMsa3csy/yXtCtrEhQlXqBjwxEqAIddssaecLfaosqXZaFPwtVqz
HbkUQ6/zPugznqM4u/OsaN7hQ/Ld+PmH8H/q1KShVb8Q2QxFhvZlSQPzma8PshxRp9cDOn5vSB/k
bl938tjW/zHffD6FebrhaK9NXKK9hn5j1tr/MbfcuxDWPniODuwYjG8iRurLaTWBZUZ0RSU8pQ85
aWwLd+2fmnuHLG+xmONOKkrOCesdpLbQnXuJmYG9iynqGTYLa8o19OSWVs+WlPIn4iNIo5J8cD4W
3A60oSumaDxqWu0ZM4kDzniGa+aTPtoHNR6aOKRbMKq6K1y3zrA9+YtkVhauwE9WnnXgU7j9h4Ft
KeEuYsA8itos4UhoPcf/edhxRaZhqTWkrzayOo+RN+XYQwAzZvBbv1mett5lZCsqZJYwVTldukAR
OH2kG4kCS2JuaJ8X90Iju7hwiStJFlFDQshevcm/aSmv6JlhJHRBm49/xnMzUn3fPAxZ8do8eDce
Jrbx2XxPQtivP2WAmPw5NcHh7sHBFLx3ZFW4JsEZgbuxyhj44O9qb/kYVL0phRFT+s1eRL9vVN88
3dcuuNjNyS1klV+hmo0x49eFRnr1oqitYLYd8fGSuRpEZ/Ca2fa4rf41lFezeZEdyYdSIzNyAvcn
F2AdQmdvgpjcMq5ziHAiNetcWwGdlxxgNGsUCvuTrh9IAjb04xgqdBNDyoiEYan1xwa0m9XPZ/wo
PRtRNCM8PI7mtIY5R5RahVwhzW7+8MnSyTqmlLSOD2FM3xuBvYtEGxRI0u5LlgmXuLWfb/G6Oci3
h3bD0Bkhi/uha1OSWEtytw9LUaiXBlQSPYoKA+FKtCAl/uX6Dx9b6BQ74xTKiBY8aUCkXwwWPoXj
2Gg1VchTegnodXEElp6kGiw4WtdlQUn1CdE2wfcyeaqrtUcJH8Ba5O7+gRu/pSPX+lC20weNvkub
5HZgZysUJTe4Sg9Ga2FJuA6We9EPcUsZvpyhOa5a4MKOh/+l6CloJ2fviIoFQBNEO+L0yPjbPSYU
l3tLxh5tlT6QWwYnGAOJwKxCzoSIZtiSYgRZZa5HkzOg2IZkzS/0qAUncz01fbAU6Tpxv4X25ytm
ItnJ8EfAX2dT/4e2zQdN40DY5iP3V0l7jYq101LPden/EOKiz3+QafMnTlfqAzKBGde8lcye5uTu
jNhAGNUaBoBK7CSg//bXAfsW+rrmNiNO1Vuv83ME+S6pKh/zCvfX2/FlU/vimJNE6Rr4CkZxX5K1
P6RY1d9hQNw79QcFJKPjPe6yuAu9hZp5wa73i9B3cVYnz2ZwgvKhDlSV4uyy4iHa9urcgNAb5kUh
FDe/UjtgoheESTNzJRSS7qpa/AEh2PFsWoBSGGHH7ub2UzSnzwNTj8YO06AYWujbniAqLEFfQSOr
NJ/vxJkhQBZbUnA7WuJH8wQU3OfW98IVhXTRAm2txt09GX8WY+d5fHeQ8TyWJ74CNCAgvHxepxXm
K+jl1Qk8wOFU7fjnylrd3nStx5Pmn9dvvDTNANKeY9Tw+YZWlI8+hov6KHkouVlluDz03EUgqLuR
w9rmY9935Kv8YiWZfhWDWe9H3ELPVwOeIZMNzsyWB+4QLKl+3PWaOlm5FZpvbhsIHMbVJKeyiuGV
SO2zElsoOSe0hjmUosTtDb9Qxm/Rl0t9ms4N74UG19w6J6EIoF4A/IIIgGaPOpBUAzM7Nw0P3W8O
QiuYyi+kNFIODzhqYRk2ztx2zLkrtATRZo9bqk1PrlTWYJDqznPx3kf6I75SEES2vJ3WHcJV4BdF
WKqn8KVvmvXEihQp4NXyCmYNEN3CW+geg8F1ko9ZDk5neDVHYIiCO69Qd+Su8OeYIP91I7djKyTX
yzBhmTovInuO+f0hvYOORxccmBFIUSpSp02NtXrdiAsbYvNgODc/cYxVSGSxGGrbGrQE1mG/VwVo
KEHpCwKZLaMxWr9duVhhFw2AHwOpsvlCd7+AVK5gtWzQzbdRZ+22KhkytPFUmyMe7E8Mrltq6oIL
PTzo8KJF4InQuAMqSjaHIDatNaJJ4jI1SjJDbkOSh9R3PT5jalhabUTJkuuloxkG19sZLcVVKqEz
6VqJ3M4ITxpTye6Ckx85JLuePqMskjgPUex9Y6bbQ6Id6YVNK/djjAUjl9u4oFT/GOqDAg2b8Pxk
9XnraOm1o2rWjRejL6xc+dclIZGEiP4NUpv8+XpQ6wBWKdjEgP/kFXoBxqRHqBEGuJXx6cDkcPjU
scyPu2LHuO2q+/OkQjbYsf6+CuC4zYqd75PpVTpi1TN/p5J6yDeKbm+SohTMhyk/ANq7PQQCCkmj
48fljFjCaO1GLJH5gMtZkC4OibA+9BcnC4P0c2OjVnix7HXt+ojcCvAofvK8I+/r/PUSU51D1F6a
pnNs4ZTOdk9G6mUqJGJxSWJI0R/MWXluIpUnbgOsArQsF3WHey9CiVtTLUA1ElMQHnIh9eSPBQet
Pz1fKbmrj3cQE64Yb0w2pv9ZiLv96iAuj/Vgg/lU2xT3bGyQwAExwE9uh2AOzkMNjJk9yafuwA1c
cbg0FOZuRF/yUXVNpoC9hlP3EfAkJXT1eFzNuHW9trDfB1BU/9oly6vhsJfQM3Subl92TA7ahkJf
4OfvFF58YAXTVN4y2L8riKFQeQlNzbMRgTPjzIWXtXtkqo9L/2v/6ETvdP2TsSZ7kOta3kNyqoGr
uF1E/GNDZBRRyhefUT0AxPo+p0Gk0/Tgs1sESdnLNnvmAlMWYDXpCtenQ0SR4PpZUmbljdGpv2bH
ZJ0UkYCssFJIy+72V8MPLVM46M5MPCZ4bihJ9N4ZwW3Y7zFsOo80HDF2CZYR/enBtTB5dSMKjEJC
k6+H1g/I3Yudl9DrG/gpgzSHBxXp0s7hXEgfqCo/CEvBzNQhANpFAvZzNaHLdxgN+uQrZyOsMXxq
SuYvYqpzJAVEu0NRi4lm55W2QsNEUvurtPtlVf2Y1XKytzoA6D5g6heRGAF8HjGfZQQjpKbuVhni
qLcgh15YbPsWICzCTBhN0SJn5q+k7qG7IWeAOvTxaKCk1OQz+2+SE+RS1SOuEFPYkElgoGXCyMAI
MI0SuOvDNW8Nyf6VTKg6j3Il/9vthqDjRuk1axShCaa9yf+Ml2q6vZLdojP2mvnQAb7B9A68C+Mi
OaTgKqZNIukhcHHcAuGP7VMicRK2QfJjqsRuM+YIboD+sL72GvMlBpLGVsmNKxA27/xVzfbdrH7V
9zWH++hELkqUlElGyuEvXcoYeGFTQB692wb5qaMoUbJljLLLCZipaa3fM+wfRGHRnrlug+NQb0ia
WS/kQ3VLsxQNdBnut/YOfk63kdrgvvT1LydzFNLhLEGDp996pxVPq4hrC5IFCcDjc/aR8CiMyGo3
27he2CQqxNn6ld9R42S7Z6SaAvlMBu1RcX0a9DdHLANN5XiT5pUzRPh2YdrSCMv/PY23vXaapaYm
veOq/nuAgbaT33GSIcJhFq1nXoRP2PFUwhA9EemiL5FgwiNvzQLnbB/uyfZ7jrTeG/NRKvWFa9m5
dO3pyYOA74Bsv+1kwNBQLvuOM4TulVOHnnR1e1DE68I34TlXVVQuhqhf+L/vr5YiSEN5PRtfi335
LRBxvrdVs9RlQoDEKT3LSbnCqodsml55LUHsSJZwGfkQlk9NV+ya/HLShJ+F8LpeQBHmBlsIjJSf
exCYi1sFU93sj90dQYcFvp/mu/K9Qicmx+Oqd56gv/tj6OMAEu+85uhHnm9TuZKtkKm03OvE2Vf/
g2W1z2XAH98P7QIFgyiGAY1QbvIBO5bPtVUi/GAu84etakW0ZxoMxjo/RxzcXfZK1yhb17bNF74t
1OhkPOBDQS6rRms1np9N5ukmzmAAeg691nm7FDnJ9KSqcNT73F/Jn8SC2Ew1/6w3lVs7SpHUk1nw
2ss+3p8u+6N1OHwcP7CLpgJy2awYdkcsT1phDzYww+NPh7Qbb5zjaJzf7SSI4ijjxiCJ+C67f31J
4MvE3O3hHL+5OWuRwwxJSzzfnR3eJQiEgqnhpLtWwLpFLbs6zUNLyBjuJeWAPSJvtlZ37NQqkNzl
oubOCV7QNnWH44rJM9StSWF42lGGdXPoNrNk0+25g9irQ9ybJv0dQXlYiH/Q9uVrMddnUvLUxORx
8dsqfZ8g0NRQ7nGBEws2rkM7Wlk6M0FOmkclgOUHIDHPkTskRmiczOrGnYs70/ynbCZHAPlmv6cT
6Z7iEU8NwAclocMS69FmUodSdKe3An79RI6Bsv4pKVIzAzDgJcKYQEKPHoPAamypHWh5bTNT1Yr1
8W6MA+EWbefBGeke0zenLDdCv+RIRAvuz/63Yt2lXx1phWVkUpRh6rL6Jj+7Aqvo1FinnkECRQIN
SzQTk0SYtC6ktQaJ+3/SvxrJBtdJY3Loo73BQWpta+TDaNX3svd5z3tHmZuofwK/PIMJa7vhjTM2
2k7iASqc1JY8eByoM4iN74xl7Ir2SJdyBcKOiNT2/QNNcfvG/xPKrOud6V9QW6XrFravU7LorA6Z
JLad1PAlQexaR3xK5N8ik6/BqoooIXBzjhdaik2UcAkmGXfwbUInhOBzZe40mUPxyqOLO1v97TGL
sK5BrUlLd/NaezNdGs1QSmBhmuLC9ItvXot1cClZvN33y8IIJCO0m8L7J9y+iD3J1+6Og1CYjgK+
ToCWIyjpetNrHPOLpYcZ2+wuZw6EIy2lD1yBime54YVgOv1YF+ucvYGMkUzVhdkGGO7oi+OwpqrD
luC9bwUCy6tLdBL9quQOF5Cr6uS0fNeCtLhn3Gz0C/LykF8U67yOpIIr1+xe+sCSLx2kD+nuQztQ
N30Cb2qABg7P8lt/smInnW8/tkCKjbGJT/2ymtHENVGf3t7KsJPsPkUNRmaAvPE1Ld9SXDRCA4xv
JKoPyrjMVtV3ITj23vmwhM7dKCuW7J5OBcq1RZM455gx3NQv7S7IWSU7P380b1rvP5ctZnaKKA1M
TgBJBrCojWuJYWl7zA6Q640PTGhvHMOpWMFKUsAQcLzjwO2j9MGCKQbnYvB6g0ytIw+FCLPy3pns
sZV0yqwQ76sbaZ5WOrSzJazXYRrFJuht3bt5NrblbvOv4OZXMc1VtYSsp/DRxNfA4B1TXjnumSpD
tgj2c+S2NUdlrLT1svK5LJXbSeSZMis6iTJ2pp/GaS1F5tedW2GjfFt8SOz1Z/uE/OxLeEabA7W9
SZQFzFgasZDq0yE2nPVu1RGEp2P5AEIX7wgdUhg310MTrlJZshJpakqJLsQ/elUSlKf3all89Va7
jRS8JLwX0881f0eKGQK1WiIuqJ5nxhzEjtfQqPNz5V4/O5fuHRctOQt/pEWzCgRI7W7vbZjNj77g
QlvYzg6xryYmhvLEgLlfVN+YreEjr2xylNZHYB5n/6uoXBRbjbZB/WoQdDbjs44XFZnQdwueNFsv
jdHG7oipNCGg9GYeXYRr2kDmFd3ILYeniEFfZBjqo0YM0wbvqG4GGnjxWowp1FYm9wPaYYpIjsyf
24D/nRfQgHZ7DRHKdMTzdTYaGXyhycaEwWXXZkzcgC7YaoKacd8TrZ6om0yDywPgl51K0Ux00pjp
DQin16K/jIHVRFTdpgM2A0FFIebjLDG7smc4pK8D1qakvFWXjm8uElRcVBJcfcAnJoI2ky3CHsoq
A2ZjigW+OGMj34AsyGDDj+GECcecekCzwAozTVYtbc4ZgFRH6jkRxaxLBoprlzqTBf94cQVSMAyQ
ZDGr7O6l95Lai2PHnmhWAe+zsX6cA1jI5avjcp2LlXj19zdimZ/B7Rk31+/2FlCue1bkWHGndsv/
3V1HnZSmoGpSLGJiA3Kq/OEKxVeEeOSaolTe4oB+p59Cf7yHtfczemnKbGYIEgT0lXW2CEeMbLv1
CDJdshU7b39bL5EcPLuaG3/p8dA8Db/4dnOPMQaJCHttPmBByk5JHONNJQpiTi/FjRlm7B6StIdu
Yng3RAgRXAMGeVp83QRZkAzcefEZg9A2oAEBcEuVkTBCRCZVV/kkNbaB73jR/cNX8Q4SMyxxfPRv
ZxyekqE3Qqv0qYqh8ab1uLdODenoHzXrS4qbSdFw3L+OMJ16U4N6OHLHjV2j1Ky3/5mTfBZ8o86P
AVQt9toe/d8A6jr37FuqOsQR6e4RYeAcYGr05a/1de3jPv9bO9+RgR6tXWXaGd9C+mTYqBMjOHQR
/3nVAjJRv54RrUGo7lxByNNLLwDI3Z/D4KBEQQdrpl2exRW6Occ6P9LerO8biZsIeDy3Xlg/yIGd
+lQ3Tdik342tOgdh0T1KaajUOxB4WRZUgj7bzGO36ZZMtPiVeHKupapIvLnDKf+FGJc/Ek+TCbys
VOb8CDSgp4gG5oWYuMuQAndzNDRFSsa58dwBw7+IpL3yFmX/zzLIF4sp1tX9yfnCIq28LQaqsIPd
XxL+RH4w5fBVIVIi/KJWbqKXnjvHqojWNN/yN614tLChI1dbelcWTYFhO6UW5SrZ4SVXYuZT1koA
VfY4ylSmhF7LeWm602KZm1OsPeYiQPgfe94mwybCmFYpK0XvWKI1/SJmcUN8r9e80oDyFhfV/jBg
JPh3yqF3Bn8FUr/Vhitf8GgymamoSK93FRx/bVUYFTb5g9hoCGAMiHYmpdcfw5VFsuJBiyot1b8k
t+SKX4ekZeauyUpOWQf5sThM8eGSMUiV7R+xTtxE5i1NDrVO8oGdqJfHeB1ETTK1P0gJwRS2EuwR
xUnYGUI4v+ftfGSggvoZ2yx94OIHaipPVeUaKA9IoWlc8Qc9na48t46lJPNn1jr2L0n6ilU0ZR3M
3j7voCLAE4u1hBQSGsL36YYbv8UJSgLsAhU4dknJgt91zI8So36fXVCEeNU7UIiMb3BQYDsapgjG
yvIP0k0QBuCihkFhbjpwVWYW2i/uwQMn19drpvptVeL3tK3MAGhVpWBS4LHHZey1/dalOHIu+ubA
GULhVYKyDO3CM3stxsm7i44BppkEqnplLJE13ybJkQA6oy7OJVAkRw9wVlRDVXkvsZe1IKbFN5Sb
8l+JKOKhlKqatpP0zpVbbNjiGZq3xI1FhDqrHN/SCEAFv7KNnjNdHwhEQ4ke9B/QlRxFMWB+FSLq
VdN7cMZ+ZRyNNWWare+q+g+LDTSmsu6bZxr6iAysrJTZY4IlibnQDr1zBvHuSzlvPzPaN+PVC1VF
mBiP18TvT+yYGyM8Zk8Uo9wVsofqaluTp2uheA0ZHqLnKMja24USlr9b9wVy9Veg+GlymN6qlOJU
lCmIFFmpwIVVPM2Z4/u3eZD9DKopjNQNJOhWQupMearWtsQSNgFEVhFBnTkeHo9D7O9ew9q257sk
+m2zJqIsmm8awsIcDuSnFaof/NrPz0J6jB/o0h8E+USRQS/eKTxRNZXaGErCuZZE8WzN2tFguIf6
JIEDI3QXf7XUPgcT4dNhAN/aPAB2XHLdfHlUV1U7Ykz5ObKZOJu+cSQYZe3za7mQ3ObayJifRi7g
7q+Ed5L5vi7TcwAT1NpiF9expOm0Bd+qS2a60xKITOL9qIoNNzZVuFsbeqA5vhwomG8E3FrAVn4y
HcqijX5+QUveIYcvd+xbTgv6fWCQ7eS9xwmN+yn//1rNyH5VK/lEwrhB1souAv0qeiP1eze/GrF+
wDkjYXH7eai2eg7RsH/U5hjLdeG22jE2tJlxPaOzydfVVQVLRsCMQHtkN8mk40DzHBMvsKkEyP7w
8FtKS/G8ghKy57m31MSmoR0OgCYGRoNKDzxD43tLBnL2l3BFPYI9YzfpYTP1GYQa9sAsvBsyfryk
94mF9cTWwfzPcnBH7pb8ah6DdSJF5QFXOeio+mbebrA4vMrBp384R/StSwgiXEKFR+VFZxS3HFfn
7RPRQq37291ruOnXwyW6JwOezfu6KgZUn2LkLabbPI5RpLxnUD+cK9U1d3BApzwVCHjonu/zCDU+
sWj9BojV2fVW1aa4sQYaTvtROzrv1hZmJ7iJ8JugVadtrQ0yJKtNd0hqPXZWzoHBSffASWPHXWQL
s0YbUDPOTnf8bdvHWwUfwfn8UjiWZnY7EHUPe7/cEPe5PTgOwlzW7Uxx+6cz1q5lmms2VbIF9gmm
pXoLkA/s8EzYG2y81uRv2ZR2DSNlEwalUhD/Iqi2txGRbnerlYhPbtauVlfA9cntTUJQ0CugXDbA
BlAcoHhkuHFnYTlc9yRnT02FpJYXB4wf7xlMbO8cThjwtZzlktAGCepZMbwINuGsk0GVOcHI9vvq
Hk8TbRCnj9UThqv040NeUK90wymbTiMsUpr86IQsP4yvArZpo/zQSA/29qvmGQMAMHNTduqr+HEx
JNiK8WJeY9if1/RLW6MfiBqbX/HO+y7nmXYa+ERFVJeAz3RXTnUnLlio5fxT49y6ZX6imjPsXjLc
1xoxGmgNtMLd7QAO1W4E/lxpyHtQoiBmQtGzxxlJt5zsi5n7nf4/Gnsge28RmGsonFclUR/xhEtt
bkvnuX5YNIdHAmAsWmnojdPQZ/NH8OTNRy0F9QBTpCOK6v+t6Miqbpyo+pFTW7OILYjSGjSe7lyc
lzlUZrzEu9O4YqZ3BKpX4nyxESOS6zIjrE7xchnoq4h03w69/1D5ds5YblFGfk6N9ZY/XQLU/MgW
RScctF4v3bFYT/B0eGvMYO/CdxNaqfFFSrkaKH8Ix3fYmCZ3xx6OxXanlg4qh6NledSgpPN+Z3Ou
KA2qu1B5xP02qLsL5BBaoL6GQ2psJKxNNS7ZLF5iFYfUhhOFffWDiuI6U4HoEszZ3KLwqQCaEvmK
SKsR26KEMMUfQdIM6DhJa7P6DoJjEYPdVGXd707JM+crF6YW4ANm3oSa2PzQnCn/BGyzidQHWsl2
zP1nxsyEs2349VwTvVyAS31vLksG2AudQd2zQz/H2+U3QW4MNDmtLkB7ixFEMjHnW6Ej5SkeVNdI
/Hq40BKqgDtwWhq6GX05Tnwk77WG3e1KZaWTKGNfMSsmolt3NILSO3UGob/buqxD91FxcTfBJQ3Z
85H6UqT3V36vNsf6xZVRvkurd2NBy8mCaUl3TJE2UAJHeGMeBxoQAJZiRF775pFx1qMid1rxUc+L
Usa71xO+pGOitpUw33n4X7vFzY3gYRT4ghq3tee46aGezcv2qvv273oCBw9ZGW+VLKddaBb3E9Bl
feBAJ+hBdKXroHQlgyoJCPCWsKlczw0tJwyWj02rv0VxkVHdx2XXZ1unBia5A/gybwr9sJLggejC
e7B5LI/a5i5lXeZiRcv7V9Cd1HDzpDaStjxo09ssRyp91ictw/udZhbYmWYa/v3YiVUhJ2wNxbGh
GTMg7DsFjgeaudVbYF166CO5YN8wWw5+12nXIYqhhUjfCmfNlsEY88O+JFXaGPWV4I54WvQdyJxi
2l1D3E8JxddCq6T7XdAzuW5w/mL5k6SlpWfPqRy8xnIVey6CaETmC77QG/rdOXDpyCAOxH+67wZS
XVZVTU/0HuebcTjNJn4Jm7wANY0lX3vhg0nX2O+pGE1slo7V4d/FMj+1KVwDInY73agqylEDzaCj
1/IrLyDqtGLA2ujQE11KL2iAcZbMYKhli1cV3drEfR4xg+LAxhpG+oQdtG6hK9BGe/6AwJYP+B/S
lkdSdf10zNmtY94EmUYJu9r3kXFmkP7zKw2iyrmjGxaq0QjEZbLRqdwo5AT5pAtNB1Uc+0tTgQjj
qR+qEwLTYyFkGIz0hvBrxO/4I5w0r8HwP71nyDIFvZDAikOwLa1vRgyCtiwQmGxpsf2igq3wlu1H
RV1N4HCzLiZTjyDdInCl7uxy6L45IWmJIgS6zwhh7PknJ4fe54U8FAIdJO+D9tyVjJGOCgzWno2r
cnHZlVq+DtTMAJOy8GO+H38nkrGXegldW5/JFjpz0R2kd/bShNlo5BrBcbyczPZ7lMBrckLM8WUF
wB+VXw/ma22zFmMDbmpsESRIBjBWxfYtgFwH0C5JZ2Yg6xGwUXGynqstI3WgwTF7xO+m+R5zxUTp
igNFsa/Ig5xxLhw2ZSiADTS2FjQVtDuMQ1m/EvEKqZi5AAKC7tBgUdYcmZETmgc7Bs/qehe9qrgt
VSg/CUREBrg7/IxJfewhazjE4uQsc+ACBnnmmT2pq88SDWKMJE8X9K6mhtGQ2QUzm906tnfmIkjy
1nKYJafBLVh0G9tNHJF6i5LWIWUnIu2yrBZsqcis1eiwmaCKPFK6zkO0j8RLTAzK5LT1ugEg26kT
I+7pEaD/OYudCBuDwlrY6NAGGaQ7txURCSGyAmtGnsv+rgd749E6KznqTThkVw8IzS3koZqDo5sr
OYyTKDcr1dk5y9X6zIaGCjOkn8H8ufq7hvw6uy7lLIli29g2WiPr4PKb5TrP+a+xJeUjdcACzz0k
4qz8gLRnKtdVyT2irncr7iA8AmPAFGYJWqciGeQ9XA0Q56+fPYFfU+sM2xVCbmoJaM2Duywqb4hB
qBfrFZ3HFc641KSTB6Jh0iDYVHBaluyvraxEmnT8btSTVo4Ewut3/BKLK1wHjP1DH4sPsAn1qSIn
CVJ8ziSohg384rlxPtuo1KeVIPr0/avxxw0CTPmp8XiwDdQEJZyXSklO4WT3Yvg7tLp2JQ0mHNlX
XY1aISk5D2+4UewFYjHvU0o8Sqf3L+TVZiz9sEHN1tB0jz23WD9xLzwt/2sGDhIPiZpROJjwSeTA
dqPpZNg9dgzZzkRhSWlWl7IQyJ+byN9Dca4PS68ij1cGrNxEpg3ftrexNsF15NElX+Jxpj9VbC3E
fxG4qaTo2pJKXv3enRD2Cwk6PG7MY7py3ijmLoCrIHuF4bhZIznn8Gf9IGOGpc3LFuvNV9jrkQ8x
L/Mv96Hqqk2hDBy4vBzg+JOf4cQ1nKfK6cLK4FmOPzP68JFc28CA5xqgPEC8MZqdFNisdBj0Pwuq
8FZegszWR9CxT/OjMjuXSGMzhyYfcpAnZpze5+BljW0jFW3gnIkx/AXGNyhzGNUt9ZPy4w/tdyJQ
/O4lVkVBx0OBTKEBFFtle4YTOMSX2Z0C8GcCE7ktoCJWB4zXFTh7n9GDy5pKD4rRfwPl4INnrzci
RkRIcK0gQd/NEOwhq/VUVH4CUyjh8ycGquHeJ2pBnUBzkfaVfq22g1XUJ+TKRwsA2KdrthZtL5xS
8nlLtJZIFvWaKMW02xfAJ6dT0t+d/WrtHYgkRF6VxL5i+SnTVEW/hu5HDKW7XXyiL9gBOI7LDtD2
jTqSZxOm2c2sniA4aLiCR0BrlGQpv+LrOlVEDUHKtf96MA6/oiY/gRbnzFWV1BwbQMvn5u5gWzgJ
KY3ORhkfAjQC1aJ39zO+8ZWU+oSaohtcASQWVBVUUpMVqL6NGc/SypxEwCCyN8EWDGgRFuqioKvT
fFGFzzPH3itM7JSJqmu/Xfc2slUdTeJJ3nJLCwXAkSf2TU53SqYtFCI5yUilEanWl+KsGKgXoG6f
sTomfoYYTCZrXyZTqT2FJ20icYrikQAXvIq5OALcAKWY4lqrig28GI/jeURhsOz8JZAMF+goQrNR
PL5/hj/C5CeRg0/nZzIVmtBcsRtbiL70ZeptwIU2L+o9Ge49ANspsE4dWXmhX7uFHlpuqWMxtlaQ
BsOcNHOa5CSIrRRrKQ+t802Kr3FRyu6RcLbniqfY+t0flRxBJCH3ENjF/FGh5c+GH4i4oAPdh7Bv
eiGCJQVjyKNRlTOE0A86x5DXrEadFxZaV9H1fnub8Fe0hFDVlbwTFv41A61NnxN9FttBHsZ4p+pg
eXuUEKYYGl3P+BwutabmryuDnETGiovlv0f51uPNoA4yU3M4kj4aKFHUfN92MrHBhmZPzl0Q76z/
GEDdrnrZwlEozcmyJA84qKA3E/JmgXgy34Ky4ox5EWV7ZNib9ZJFe5U6ozulV+cm0k5USkJ8wkMt
sFkHQwowL5R9HHTubtVzRzfK7PAW4AWtDP3Aip+3DuN4wTGA6z7pbPMUO23zaDUhsvvRUpeyTYWh
VKX64it5VPpkLX/3N8yPjcKcAuuV2X6yVrsrXOd4j8lRR1QY+hINEpagNXilFfdTN6oyTWtxaEPT
60qJ2+vRvPZZzwG2NrOQFUBr3Y3NvCLbHU6rQjrwvkKdg55+ok9o9o/xv1qgxsnjADit7RO9BW0R
5LDkTebjMblumPXh9/5xt5Azdty6dlUQzyqz6njn/ubN+C7q7gb8nv4fjh+1TYqQHdfzOpnXLR93
j3bJDp9Vv1RnSD6/JA2DyBRnYQanKwQGFsSpWHdw1OaH0wKetrLkFbf8ifUwd0aWHV8324dNyKmC
YeEqfr1SPozdSnuvCDo9rok3r2t9XzFSHJU7lrlS2JcDV71Gao6zIAVBuiCFpaoqTfeC6N/HXRTt
gTvlKZ7zPs/QEWVOVNXn186BfDB2V4lW5kqsaTyx94d+atj7siVLqhcB3iZvmZnK8GiH+zFt5sfq
waoF4p6Ixkmzl9mc6m/sMjoea1Fi6reV9kY1t1IIYgKQtOV6dI6EKy1gWK4tcFOLS4S2VYe4fpga
ZC8J57XiBa6pOpobu5sPf/BNPK3Heh8KqSoffzNdnNfYYd3WJEvOGXcPrabklUJLAhR3Zb/iBPk0
jkpNfzUnGs0XmeT2oZviJfPkgbZWpQ4RNzd4zNxj6/4Y/3NC8f/IBSIhfwW2T9UhbZn53fpNbP/g
ryAdY0XZB47mV7tXMJ4vzMxlWvlo6gI0T3bqIUI4k/4cuI6BCF9QMj+I8CxCFiB7CK3NNBQS0eHw
2zZRnsgC/QVdAL0BqAgEsXK2lPwz0JiLOU36pF1ROfPhdVJqwoS1WOQQSrWC18nJySxHmRxYIWDM
/IWta0VCxv+GbUQaTrOocNQnOqhF065ZKIuDn322977mwfcgQwfO8QrtVyYPWJeT+UuInlQa5bUn
LbNFnPdQMGrp47DQ6P3nqJAXsX44ryZ2oTxUnP8rfPKXznC9BSCsYWakkSLRi1vmb340APBAtwZl
ZKFL1d111ziXMh3e8veomRJFu89ZqQAelYx+q1rZotRSpBJaXZXq0l6h55iQ6MQDdt5dl2QBYQty
7YEjb5rSSwOoMw1uUEth+1cCQ/nvSofxyhOc/u91tV+ik120EKpMuFNiSH3pGBo7EK2TL1p9EK/L
bflvWra43zcw1mHaL05MKVAxG3IYzM4mX8JUjRdWrc749nJdOHDIJO9HRFnHqURvobuygSFfNu/P
xnWtvODtaAUDRTIdsAhekumaDHa8bYh/s6DWuMRW2hI2e0UHQJKAKdAbIxM4oxbW+6a/Hyjdo8Cd
UGc58snNVk/wwgJhjYuSuAyyiMxguhWOQGEbwrXi0GALO0cTX9v2F16Mzarg66MqBzfG/McmWy3S
Pd38F0BKu/tYzVxcqAYPMIVF/oPDu7bMztZhZZbAYGDNe3Yhp8RCiWXPjf/swjcmpGAlK1zlVh+N
f7CxgpCOtTMMCq4WKDzUA5W0na4j9B+efwhxz67ZZqPH3AAepgypCAyEVmUmvJ+m73J3y6yM5KQb
RdfkHg9GukWD8Pcy/fTyrAVYsfTWdba3xeSvUT0VlWnPg5J4t86Xu2kjx9wDTzp+T2qgBSZBY1kc
9kV37/6sA6A2D0PrgerpJfhDdo2m7v1v9y47GM+jsMl9rbCUfzo1axk0kmTrSgnWEhxRv2/+5zT1
1GK7C12hURI30RtAo3C+NTa8P45X1PiDAmc+Gb7n6A1val2+LkQAgf/sJMhoGHi2BJojydG2aIp3
Pg9mb8JK9f4KPUzccb+OglEX9QUu+B+0b//+j5rYF56zNdv8nHoJJtuGtSM8vB/NQk50k8EndnPm
/5G8Uswg77XbCtbxX/u1Vxnt3go5grnsiKWaSqbIjgNZZeOymtE2f4ZabHg5tJ3yUN52EWtp+5KT
Z6JiGp8Xx+H2HXJwb0cL7TafLSyC/w7l+Ku6/eoZWgqteRcXLDjoqIi/xHIjZ6SEuknMdSqB9lF8
dvcnjtVaZTOZEv1mrFh3K5MRovPF/SaxKqw/H5m+bp6OWoz+dBHgyr3Ch8o9AT/+ljuFJacEn8oY
WZ44+Vu1VT7K7ZRwLYkUAjlPb9+Xrlxk9ThQeSUqqoJ2dNR7lk5Q6rxtcJNzn3OiPSqqNncuxA+z
jFpFxUioyeseXHBobX+aYeiJXyOU61gFbViNGRsSnAi7RPT07jQ6xZxiMobiPxsiVEV84R/EovYW
HGcAh2CChPo6V6zvt1WsgbJXb9ek/+SAIzvsM5dxHcMPrkGeOrbPtSdFbBta9PqqlK4QvW2janry
y7timx6eoODmgKcBZIfkgAVcLXi8NJYwMaRNMqtD453KOsRRkzF0he6khrTmJnBuM79wme4nl0cH
pOdrgDLbEp7KHNKRPD4NQ/2/7uyELHsRUIiikSofYSCHf18t5Amn4/p+5F4hOegcXSPIhYDY/fJx
QPXaYRMiAjedDn6PZ6SSoVeEjvf9ginNZUMa01m6vKvNXHhN5CBmldEDgh2ZsNd1XJdKbPTASGPe
YX/1SqRIk+gIlvKWCvVD0Drn2QZyT1S/3TipXuTzwetb2MrF2V4R3KbJvB1HifzfBM8evl5vaMxq
1n2GqUVianQnWMNNLmCKBPdpTRBjsN4yL3xnMPuewCj3PiZEnIO4t4iJTnuHoK42G0Naeigeq543
8cYdQFz2x49H9Fb2v02N/wndXQE6tZ1HzPLgS8jJDu8LDDWjHnDg9nf17+9vaSQmEDGyt6EYAfrw
epOfUSPMtsmoxoHwZCgnl/ewD/Dxnvfo4ScS37egNxLrsHQnMU3ZkNiA6lakHFJMLuPt8RqxaFO/
BapFR4gB760cqx5nUCfeqorJWCsyTcLxNTECbyf9JOUBvMEu0z21nh4MxIVqOempeT1LqvPJfjRg
h592q6WUac3wDmMTKlajmIO/Q7ZbSLIrkd3sUyWYseIgNrBTngdYOCLWtey3IxIGZFhYHlU+DHQw
yZTjznkq85KCiZt0U3A64RsRDz4pFXa8OGPwNkPMDgPA9exIOCzUmQ6OT/nGVJ6kvlZB604NegrM
PTgDdxtp0mEKIefO7aJnhq1EF22G86Acx9uIOMxnTj68XGa50I7X5A6MIEib6MSB7zHA7cT8kNXt
Rha9OToIKn4bwNvk8F7cNVA4G3h+gQ5kCse4VT2im0BzPlM+2AKa8xtVG5dXNzAPjlwFkFGjn6Iy
lrGN8JVS1TShE34QWFO1kQ9oznQBHAemkhwfi0eoiR6AqWeQyVbJFVb3NVwQC5K7/a/KZ/HXmFsx
kN/MBoZ32PEh8Q0NmTKIhwTa9IxdQwS1lHdqCAb2dVGJyxFdQZ0H9cnTpWWKzP0ntyHX8/0uuCjT
0Jd8IIwZgx4iJJX8vemmkrPfD8mDS3t/LT5ow40xv7u36guZiLKMHswQPSqyjy71IRGa22mQIuHE
qOOS5r4QsKIwGF3NiXBMsEJRWAL0a/EQf4m9na9Af1Tb2UYIishIOOeOLXzkDasDzzPXoDZ15Cgp
eOXSuAkKMnqcPx2pvedShCHTJC/1bod7lIci7s2AHZmHmv8tCrn5HITTtg7ZXLrtXMMmxwgvTO5r
BA5qzV1EpJ3iIx9kSwIzgxxKHF40NbIFSQ1Fk4ngOeZzFlk3nLmrj+EddxS85voggLRa9NX33/4E
nijg9EUpMAtITGTB03Y0pS0LK4z6zoZ7bi+3HlTYSNbZ0ozw8llxAx/mhHNqd3Rih7s4myqK3N8i
1Cvn9XkmfT6ZTSXkFZgr/v4uBayx65Wjr9PELbPUPufmwX3+p2aCjBTNHVL3nzxYfqx4C73xJWhb
4eEuv4xP3cgQSj7JR/6GY4XCVGUnabIZA8m3a/a4n6Lz5IaAgSV8EM7HbF0VMNa13/h5loJ0KQ8a
CT9KPGhYCyiQ7ChXjYRyxuJiSr9BFcutUuWbNr70rx7GhjFSEPmuh55ZfA+ekn44jluhXq86mIXN
3Xz+w8ceyRpZZQlh17aOMEFlTV4n1i9sYwrEVdKaS1OH9LUgL2w8zePD6ODGoZYx2XJKHTEQgKoC
3WWSv1uyA2ypgDGHSiAsg1xxaZSXPoXWEvChdMZ0ZVzc6B/Fh9NNFLvm0YjTEfVBU2FkUBA86HWu
vUoTfP1ldtFMXVDwhlO/we2mhLtKEj1KaPm2F/wP1+0DKr+IA6NyHUPjsr0/WBEYGcSH/yN8GS8v
xFvUXww/VXbUsJw6ACjpkFWcUOqcgLWTfCofro9qQDwfC5AxBdsQaEi7eV3odPhFqQeG9XYfSTuG
qR2xNLWyZgUhHxW8KsEJ/ONdxXADyjtgh8Uxi3oikVWaGkXGdCXu4ke2JryjKZ8O/cFDi5PIah+C
VRDCU25lIjWtRjJfCy4Sz91ehXavdyPZCVajWsRpUz6H21b243WCMf8Y4U1wX/yAMLSECk0k4n8Y
X6HE7o1xcrTw0t7H/HZ+/47f0vbxRE/ZDpPRqxXPDj0TZLzuiLiNFAvlUBEcEK/sSbAhA8feFeO2
EF5ROrzWTl0uJth2K7bVE85r3b/rDwiWGaRTP2o++XfVWlo04Xrcd48xWUXz0AIrI/pjP+/7qdft
4KOjunHzC6TaU8EnPAksmOH6gKbdGNJSYTtZbNM9kDTYztb0NnAeRnD+jNfmIoWT85IVFbZC8Og/
85Gdl5GCXdo3gLAKrfprdUQg0aBP7hnoCBC5/FGaEQe/dLS8pJKmIfS5j2q1ioVVuW+RwbYy6u8x
Num+/yx7AMGGLOmy8SD005bBlDbYdJPqgIgmvLTNTUFHacwqoMYT8zumQjS0CDG9UG1M1An1YAWg
rGSJEEV0Fodaewb3VP32MSEnrBSUe6Vq3OLHvQbfux/wOoyvGc53DN/OO2MgugeBytq0aCjLCTYY
g7sXrvWKpmP8pLPQ+DlxG2/mJXkaQ3WisIGHTRDtDMMeQpy8JS1ea4UMQvl+PJN6WztawOsif4ov
NF+0d6ZKlOreCbczwpjBv03+vf4p/Sz199Hl0naYRcR7SnTM8pFuu1QHXVI/SDW5lwblY3y9r3+u
kbsQdG2Xbkm42mJS9cbf13OjCTyATS12QMdNfebKrmFwWt1dsxiiNLRj1eWW4UL7BOhdr+ENyY0I
dBBO5Enr0w2l+IpMwcMUr+tnW3B8qFCWFurA99LIkVSd+EnmXHe1Hh7xbGbRCHDybRO3U7XWGQQd
TMZPg3g9BqRBrCytVQpa+gMjp6p2qi+Me+YoNOPFu1RR3P8KyWp2Hr10A56hQOjWdStwrqn2HGFO
q7iEWAaoFbXAmSO4/HIWyxriWqhCoc7LGU60o6WDJwBuQ+rXXwEY2RlgddE25EWOZECd7f9KZA4O
l4nyyJiQlaC/4ZB8Asr+zVuAnmc2AhNes/Ox4oTpWYK0Rdi4OhItT7Mb+7xJUWot8glP1eFpi1s+
K0vc9kcuydnpnqUc9wihJNHfgEM4WlCwRZ5GI2P2A1sPoyB4hJND2Pj4B9EENIwUr33h2cMZyPEo
vvK8JnVT58NPPusVtIw3tILMeFvn0oXl1cGYZaIzBzL8hTReAsMzB84LBC2GOF4fkn8M1+fH6eY2
eNAgcij2AlXiBZMPvRuXfjPxusp76gjQ2tMP5V0a53kcuycngdTmxfnzmAeS14PKvq05l278FUCe
WHjohniS9I1jQMkWy78O2UgGM7STNghNIWT3Q2jI73yj8gbDEQZSbXUFjEJ67jj7cCVqiFrllRDD
1GS03FR9JgqvO/1gJm5YVXGlRLaMYuG2IKUgRPSnV4hD/T1SRJlgpI4QzX+IzsgvVQqw7jK63j3k
O2pZ/sdcKCStj8YSOu+wmRaafnto6UoNQnYmdJpmSRTYqB8hFbkbd2UmXNcR9dfCZ9uzfchAXx47
6/scy0RuCxTjJe/8hLkb6f0uktQjHrke18SUj4471bfNVq1mgzJSvbNySDIeGfezP7I7FEOCA8ye
KJLZca49ECNmoOrNzPlh6UvP078h5H1pyk82OW8TTBdpf5w69sY/CAG+cYRAFlGH/Uh3P0NKggAz
fmAE1PpyNNqsTrxN2cDtSOuF2nSTlhW3snlXNF3dlEMg+4O5YeHodnlc/FWq3o4/kSElzn6E5XkU
OH80D/fCfe1+dPbx4M3sgfGEgR1189a3AlqRveAsjvTgG5vyKzkl/ZBR7Qqv+2mfzHcs4zES+bny
r2T+s8jpAVhu2zbd8q0ImTMCQRxB1QpiMhWtqtAHHwUQGqXoNx/yc62Q7Ha40kzcVb74In9+AQ0T
5HWyZ1pHBurIudPwN1fM/3orjlApvNAHPgvLItkS4Xl7QmsHD4N1zRWU4QoXnnHmgydRvKbpy+tv
8plKcgaFcNK9NmC4VfW6CvXg9zZNm1+FjVa+21NLbHlL46U0H5zBDzm5x0Yh19emohwrV6Ugf0yQ
Nb2It045Pww27z892b282fvcMwxDCIxpupmtLlQ0yMB69CErk0hiXvSLev5pLLfce0/iMvZ83TAB
+Wbyad7avQPAnFDJySIfqM6KwXwZX0SqaHsWFBhrdub8dKDHB4ddYBrn7hdJhjPSBqOOydKYOVNo
jwVLD6Nt0x5UFszY2ZUVSkWrJilz/8F6tRIEv1caqm3Q74buRMyfkPEef2Tp5PkhfVOnzm7iVJ+w
Mwt6KXFbkf8yXrkDcg7mdRiJmoDIVvjqZOBTUzNcswc/6A1pqQQbzb0XMi0+U+cx6qm9kR88LS4X
zf7VY8pdOQreCQTG9xcK1cf03fxIqncN2bWubIoIraNcShFlG9+m1at59pxJ0U/VpATvDP3jsHDy
7FlNQaciJC5pR4KfH1/+klmhrMYb3GDZZt4MVKUMwDtnHHaPkQFu2MhmTvbIHGAiVymm0B+rDshG
1+FhsjrW24dqMfywwFInAXOATCIxH0oa8nu6O0rSNB943z7bjneYRUFaKM1ha2SjfwWCzg0AcRMk
zBi/LTljYqtpEmQ7FBYwp10ZhGzfYEkye0Cg1XJh/H8DnjyF4zH3dQnWXgQmO3VuBj4lu0jYN5Dz
HrGJJOGJC4Itt0IrH+/xbImy4x4EvRwuQA9AtPAvJzC3hDrwMXngSZIPk5vwFREUqDKC6k509hp+
e2Wvb8ayTTW1kOTDNaD0YBS77PP5SdpDfH9upmqu07iH0Cq2FDPZ197VMqiUOgTkalZGJPIIDyLL
3e1l/r1LD/upkEozvfiemQEVfgjuelIlgCcXGVjx1XlEKkV87xR0lf2Ajegi21gxi15VlLxVdrgX
Chfuj0fFaL/Sr5/HzUZuCVI6EqdVQiLAPiG0VRCYFrjX+eO3jelB4Dy/zAflncBk2YaJ2HT+Eni9
XTmFqVS642+cH0LMsuP3DbvEO6YiLQ/2exU89yobRPvEDlHohNcNTREmTS6+N/kJXeJvHksar/s2
lIR8U6SIhpU1NDycZETokAnqkMFrSTs79Ww3BemK+0I9+FTzWsJRLwRZiytFFDgQmH8a68vmpSeX
/Rwhi/0l09tP0n3RYaqHo/1flf6KTdDnK4+yjZ4jZW306ImN8adeZo8PigPIBR7VCE/zoNEVMZiL
DVBh2qj9UVToOnaO4UxN1VGNxs7EKHMm3aHxFPXZBgDmCQC1zXJ4YBhLM6/DxPQIgQVueSCtGR7S
lzdJ/yttbI5JdM2XOXqGY2hxysoyWi2d4yYQjNyF4YGnSgfj8uh9RnB0iUSn+kGdbmUnlDRcTRjl
RzV7FFSP7cSUL2GRA11r3m59wajB2RWkw++GALLmDrusonRLfuRJty1v60HROc3iH0E1pGR3E3f5
Xbl5GP6KJVgJmHenf/17l5TUeVUmp1acW7IjgaP4mS3yFUjpFSkJLqiAuHHVSkA3DfMUtXcg0Oiw
GjEgNyBH7d2ioaJOpFWfFoGCTOEbI8tCMRQfOX/XAy+zNAL43wKMiOuyhkKDT4afC1zvOtPseh11
F4p6r763bD1Bspikk1P4Q0so3VguvdYtc/IF8FyMC8eZMEJtLu9SttIZT6bfnF3F76hl+sFCqa8b
bt6/BPpRbxEwKIh+5n0xjIeUYB9TRQvxOBRyWMZJ4x9OKbgbnuA4oTqtGIKumQisCeZG37U3zAxL
DGSW38kO9hhuvZ6wW+o29I7Rl+aPW1UR2g1dbjCpjJioHig6BdXrDjNqyD7TjAw2kLRoVSvtDofV
whv9DSRtU0KUXws6jOAOueN5VvcAz53MrSr3UyehJuEz900nnv+Zgkb+fAUFU3weZLVLvgqe6uXX
GvDlnJKCYfWdfJ34Mc0G8p+TYmtYEC+Cc9LkrqKboQw9YlQMsM4k+EJfJFPr6rYyciRKxUOMrT35
fD2MiQn2QKTeq04nVcb15P9Nm9neACG2FaDu+Ks5Hbuy8gHiMnJGXwkfcwtx6BHPu3OcQ5mXzfZA
/uF1KK+NYh1zdi5igNKmLDF91oPUzP1f6zczLYd4Yz64OgAztWjv/oNNxE1LnHNc4x/TxR2R1iaX
/wSxBpSTH3rDZB3PKOjsgd44m+UmldVx8nQecJijzRa1NdLMOqLywKjEa0lC2VQnMx85aIcT+DPT
CIVL5+QdsCx4r/+0lcVDBQIVKATeTLqO/EV2SloQO4a2AZrOlFugIO5wu0BCUV1RSZeC5r7pougZ
QGmPY5yY6kM6vjo479HzSS7a6LkfvM7EJtvw1OJ+KP1r/69LOaxE/RMKmDIJj8GiNHXpfDLURhQ8
aPbQtrSOtXeP5JmtvWARHlL/CbDcxrI0ErH+fp2j4QXNTP/cRJxz+S/ycfkBc9HcAFeM3cWM65Rw
CK99wIsVad1PM6bQpG2DmUK32QwyAOfaArQGmnAC/Emf0AVL8YKWZ2f/Prz3AMqrW4c/9fVtTlqU
TuHpa+sSV3Et1hb3A3oEldESSxEV3TNa6XJcb0kXJASkv2IhMh3/LbwkkV2lGjYKXKemBo4MW/2y
3QkAb7UlhDrXNuJ5G6Gy9iFSNJl463JhAp9rRq9YA8a93kFsM47aTzlCzBhqPgR59l3awbKNr2ws
ebqtczNvcd5g2P5EOkIs9O2Aup77e59lmXIFPFfe2fJv6vvqPUvxxUCkHf7VrTluWCSdLe5yPqco
lH8o4cCaP3k1gWbeC4F5R+9UZXyxA3Wbm2WqiXeuSPBynysymTrHZrQUONED0zdA3KF8OpsY0m1g
HiUQBEV/whNURrZrbGXFrohD8k98bG2i913VqMMv9bRxmNA/vnr1jrVo+ovuLZP2PDC3CMNJ4xi5
kTmLpH2SdOyDV2PGe3kUHOiN60CISEMQaWPNKKAoscPfa5EClKNeXeQskXq5iP2RrXY1HqrfsHrN
P25jztByWag3pk5tsPRUBEJcEJNSJ4PtJv29SLvig43pG/bABjpx3SyaSPOEaU+TkAX1nY4xeitI
1gkIgkwjqPz4S1nWZIhroSXFJTKdRiY1BZNGaWcCAkROrzb1coyCLpFIPPJFQKkqcuL1Zgx6eyxB
X3j2U0xBg73BJyq4skDfNmVThe6CsLm/Q0aaXNW6UOvRRK6zYhRoaotG6FUrKQiOIVJMZ5PgvFoc
w2BUId5p+4up6U3fPy78aqj6paXaV6x7ENFMoT7dVsTWNWCoGOJODxqbUR8qE0OENrw8pj/0fuPa
XIOMzYLrPvmrRhi5icE+zn4g0EynN1bHSfVQUWImdgXmj4VRi5feEyaznQpgBcAlUH1NxF770Y1f
HCjeQqgrQ04DMBoNI6C+tFcvLA7KX66bMRc6ZOAiKlEctHQQQjk8bH8i3xkCt22sOtEXxDHUWfJx
DrPsa5M3+8OEW3km9YQny+Q+ew4r0RrCs6gZGsKauNOFSyNv6gJSBDg7epo2zDqECcRfQZJYaxaf
K0v3O3HS+kiiWOCN0Rri4xlNQaVvmnCMNtV24ex4CRMAiaPBre/eoJjbT/k0UbYDC/xL/oaksw8K
yuYx+j2JdB6eO39BeFj5KtQcnVPM4NBuHJatKP6SQeLuD/Bg4zIUPryiOHcgih4OkBZvEsKA+2za
6YzYmw04b2yQuU0bHf0kTDdJm1L7VuWLBRF+/Pbcfn5sX6caNN60/v6SNJDgdVLwjROg+iCm9JE8
SpGKAoxI08+TmoGjdhfk+xka6XpZVUWFszuhH7OHSmzzh/w/8ggn4GFliCLXCqIVd/gQVYwBY+D0
f0Qt8Z51dorTKTuzsksURsPLv+PaQphcl50wUyy+IRB4OezxTLAsIbkrJklWua1aoZCvNkVYH3EI
HJ0uWcCd4H88SkU9D1jHJpToM0mfaEXOUWyZtac1/5GVZXFJPdEkBTF8cuf+pCWYvTS++is2kHGa
gDMJZE/0k8YFr1nIUaUSgixVo8QAgbsQ6/cospx9KSzQ3MlZA7CzIdJw3WsF9aoqq+n4u+EMP3kw
i8dBOIZaNMFwQBA4JlnKMXOyr+Qv3Q5+tLVS+cz4Rg4LHJ3ELJYznhXGjD74HuPS0qqyJK1d+WyO
6i4XmH8PKGV9ZksEtjS6/SqMzTzqMzzNlOJn4KuAYkWd+kaiZS8e5qLAlYLdqUdDbbi4iRhviePP
He692pcE4czm1TO2F8g5b7ijl29Pl8+nk8zzMNy68GOjjNuN8PBY9+skzCnlu7nRdp0efRNLCf1f
YqwZK2C0jMvWbdABQAiPCM3KvBjGNWYuDlK6SB/GuO8+qOgWst8J5BhdiKrF52wkC7jMSp170JqC
OT86pqtARaguVr++uGI0OjCkOoc1z4tgKH9o1oBizYp29f4NSCTcv1CRC12ZN4x/Bo24nqF+g0MM
6vEMk4WHsHRRF2MOlboM0TFIluaiZokbQOQNA995N5qowVtO18ecLiM14ZLclTsij2vA9ZYwLJiF
OqJV98sDVutITkUB5/SWOMHf8NHU/5jyAVB4GfmP1xL5x+UQue4MlMeghQUxMyUUYishkEx29Q8g
wZfz+SXMs2xCri8HWNZB/RPrpiZaFyXv+M3KColl7ULyr2JukqPl+WSzQOCGYtoCfTG73F8zDauX
KnSslHtfIJE61yJgYMVwFL1kIovcIh0PGwx4qXcRULomDrEWgBLIjpi72QO69NDiEi1aD3w3igwm
PdRVG1xOtNRBBYM/4c+GFFLN2RJVKSsGmD1rotg413QpUkop5qhqMzbHrRVha+z4SWQfxDT0ZGzH
o6YxGWc6/G3M/kpg+d6vcEKTQCvMaZQJRRpaczxsvHp+yvSSOadXwssj5r2EmjCEdtaT9673Sf7D
P+8XhqRC6O9XetcB+uqOs2B930hi/J35r+AdFCPraAVL2eKCzvKb+SIpiboCmfZCxUgBQA3Yi4Rn
wJdyaf+Dnvm2QHe8qNw0amWQdGNQBBvp5nMY7cxvREWKlCaivx78PUqW/o1I2CXen8KorVcdB6hZ
sdMiyVsqD7mBPEG/0b9Hkki27ZUwGAL2AHAen6lRTOzVshJnF0OYnpTni0XdoUPPPScdbla4u6yv
t5zWB/p/MMVsxvajgOjXY0aJIVG/XP0ngd7eeknorm9KXF1LLvJ7eKOitMWByqTJ/0ARgQ6K4JvH
ttvesFT9EFsNG9EiF2xbQqCjRCTjecSA8WDNIvBas6aJRXGSf8Rr0RWJ+DwWbaJcc5DYLMpCqY7F
rbIq9PM3EEtwx1f2N9YFFf8fUIfa1of2w6QuHhHib0dx1TeRRrH2E2pVpg1uN0uOVcgwIjbuUF0w
PfgZ8w/NHtJUHJkBerqpXXDzXtFsoP57BrBarGl7toaxz68Y47JTzzaNWLlgDIgn7GvgwcNsb8Y7
qjbXP8LkRLGB0pf7t7kuSRgra12und5tMV0UpdAvCXsOM5Bdq4MhqM4Nx1hXKh8G1xMZrQb+gEt5
hlfzyQQyId6mr8IU/nWSTCG1V2pe0z2INmic3fRil4zK5eOI+3j965w71cLODHdVaRUmOmfA3MMT
QGEsKHN3V4NyBsDb/VEPlfTbaKK8cL7Gmi5uLzhVjtLYzFiSoBqWAQ7/OCVO3k5QPzfWCkRBXGN0
9baafljlfm4nj1MPEiMBDS8wH24OoNTQCCDAtnNaOmUj6iI4V0051odH4iO/yu7Calzad/mhR0wb
PlL8v6IHSRTf6rR+18O4/BY3y7TfjhWex1e4CKw6F4mQMvAcemhy2Msn8UwLnnMwXGq4vF2swM7K
y0uomkEpryMTQ0NpqKkIU+5omZlAK2GDDP9BuGJEM4ieumgBHzfW+dRM5ru7RrhsSFMrc56d3orp
jM38HB+D76gTH2iiSDsijA3yEgAltPZM0v7LtMfASJYkGi+kYTpk9h5ZGLSFHlvooF5Ako7pXBtj
S29NudQi7Wfw3o1VPPmzMQq2mNtHuk244BYnWFxzqMKIf/7nqkft2KzElY6u8ZFFNrqYYhQzKNi0
tVeokuLv/NUXyG/kzvU+fj21AV8faFLGuVzqHJraOHwxyMfcrAfrfhRp+VrH3G3N6Bd8H1Bo/9Zi
rkpUkhqsHuUZLwuvBZx+x2MiriLkx40AnRpyXjzrKU6md1aLymtQvCKGRnMF3vShECJhVO2KF7Ne
Yj+n1JCJ0BW6tF2Wqz/ZqK2BCBR442cW1wxd+zw4WGGCYYGQW4+3d0bwK+XZDrhumJm4h4rxDmg2
P09P33rOgZdW3Ca13p/N9f8OMshItabfsaolF46Ygi1W5xdvDLnmuZqTgOqPcv4x7R5UjGkuT6O8
vmiFfm56cCMgbbjOvqe/6E/78gcbx+31anEFyl6ERcZe1EvgENPOwM/MMKGWCHcxE+dYX8p+4Va4
x8iWiX/XFnO2RCQ+SkTuiV9Pltn9cM1KBVHGlvaBKyONTXUn21MdlgP3RssxbRgpsgiXWQzk+l1g
3FwEqf+RtOKGBkbk0StGrCb7j2IK6VhG+mR4wZpU4Kpu7qWJUB+Hyz0mWk0Huro4j985bfHmVIOX
AKVKrCQR2f974RFJEkwI2q/MPh0PN5AOJM3MpIL51q8/9xjgI6iqIfaReHAh0KynzvfGuDWn4w1p
ACv8swTLQRuTiMQhjZw0bOb6bxlxYjQxU85lxIttK0P+T+Ts8E62B+LLkqENBeOx7uYlB35ktfZ3
B6GBJSj1NabTZ8CYGuHKB8vstNXEjqGhuFWl4YOUCaAbKXT56nfyREFgPFFU0rypM6mxZU28T30S
o/0Xppzw3BsE+wA4CXIOAx4z2Rt6Qv3SiusdiLUbC1f3ryucYtHWh+qQ4qnP/iW5XhxpnYhbou+i
MIccVeGDkknSCjc/Srg+LUCbr0AyMsja77rBwFU5A+mfVImUB6sMKh0t7mC/jDbOX6+9Dr6PD7cF
FBov3J+Qr9aXBoj4pKmtQtuEqYJZDdFM+xtitjl7PixLfhCHUXb1BHsWVtBqHGkPEUQlGsnl9WD7
MU++aLTZYJSniLRNfIq5R6W1veCvK4IbtpOWBhapEozeS0QPl3/xaAncOa1lKMncqGBh4vuPzG9D
QniS48+8M0btvTQd1rIp8UEoAUEG2r1G0CbA6jTJxs5KO448GoaiVUeIhxz4udhnnBbDER4+WdcP
uvbhHR6WsWjE23QGXPl9snKjESf8+DTuNSnWtCmV15P4qXRNLfJaqN50p3kQxJOzs0Ifvb69gjzc
byV1DWQ4PmO18a3UWlGTteYNEi1w3tYYn34/O0mEotum4Ms6Qe22p0B6EnOzhV/DeMFyrQ2WAMT3
cMsczeFsGlUxTrvfE1wu7V/c82vj3vGk+F6tAsM3Kq6SU6rBApEIKc6gdjhElpwi/7atObHvgQYM
PgT32VLB9bQtXW/hCf9zHVDkW/3BGdsOXphEObzPpLyrKZiK4/h/OVBqQwdc5obnugeFhkj8Hiov
X8weCxW7yEyW4bmimikSccLB7BcE8wfJNdceY1fthUNGUJTI5zWSIj2/burLo/GxG3Lc468/tHx2
HSkvDbzfEHRI5r0jSC81sengzdCvYPR8oLt+cMw2sZpVTzw91atzGde9GB1WdBFAK2TR3UCChRfK
HJ/o2rNWe3ww72NrSEoUnw2hM3SJO66gtKucNeaPnhgyL0Zo32gg+LTpf3V7ObShYTTwMNW7Q/qA
IDZxSvEsD0TSuTZddB1GYmy/JdDxTppy4MWXDXBNu2qcdQ43FKsbyDNU87j+kwAqCZxFGiChR3sg
XYIXQRCbLn2G2hVScTkyqHLPaE6TvxnmrlPGQqI2TUvGT7p2Ye1EQT82ln8ewDxe7Ufx5n5fchAA
r8kMY+hzlVvA91Wr3aIpRJZvifFsG5Hgk1/LmHBwOcDk2aFMaKzzKrca44mLzUz7rUmv5pDU+KIl
B5OtVQzrXakS/1d+F7YLhtCmDU7UaoqCgbJ5cDP2AX5NHJnWMO2WEt2DHgMGdcpQMkUsbJyWW6pT
4POO1wjX/QDz7lG+WET/Y3gFjfxgT5Q/5CeiCsBmqQ/ATRj9WitViXUyt4oAhmuumlDi0cFMlTso
10vN2c9C/oKH1B4apvo4JhDB6y66kpKryj9QBh/ej6bcnKgGOErJeshHU0dcQWj0nwWwqEkAys7Q
5Xo1KorflS0IUJ42FWeO4zOqLM4bPt/EgUVOzcBZUV9R3pPv0q5Kbz0rLSYore5d2IKQBQTLyI0y
+r/uw714+QCc+5Y1rH5FQ2R/RPVLu4PUbcIPAFEYfObWJRSu6/3Tn4klm+zJbF95QFrNBeI46ikb
XkBkl2pkI4hgn4lD0GnM5AuyBzvr3y6IQrIJzfFVc7KIHoVq1l506HvVRwGL8HpIZqkG04Vm59+T
tG2WKWlnR8KFNZCNBJzlyMxqhg2oFwE+HkuN0rMeD2SPhWQqx3CGZwzUXXz8zhmGPKlZmL1XRC+D
5V9/QE5JN7h4N2vjm0/t4DFYq1hdFwllbJhtYCtLboOD8o1+H1Hp3GRfekaaWkaQrl9AqvjgX+0+
g8Hz4aKa6dMyAfWsYuKOphUKdE04i+5Q7DYXqOLbvnHIBCNwlSFg2sEst11jfRf9Yz3g7Iy5FAJH
NxnIEWAGoc4+9f/4qRjfuvvz8P/7GmTlEtpd2crz5U+otpnOM0SI+qvzynRjPqorJ/VLrDt7WHQh
YqAOBlNXHgYzn/7lbruUnT4yYzGujSugwLl1hIjxek1OdB0kM/R5O6vFTZG0Fh1R00Azlr1kM6QT
gcCuzzecIs5Q/vO4Ivcms+0IxqK5OQ6/zcHZWCT+P6uOvd40Dk0Jf2dK69FDg3BaBCWPMzyunQTr
uRIlO2AsjOtkcQmsQ1sC+DD+eWAR8Lr0rPXW1g2iCPYEKnKa3vikPHjWIadD8t6X2u9F0qJzi3Cd
61FpJ3KtqTuN8L+/dwJK0RAEfqSTfJ6Z4kQjLRkH3vjUOBsR4RHJk8dcKN6gLP0BRojnrPMcn13R
UQkq96k9MWyAw0f11tKPc7as13lOJcZJVNZOlFbV/wncTUNh10KU47clGRgXCEdXP/UhaoIf4I53
etB27/am6OSt4BKcPOsOEtBAN9DbIvl3vwei4g/ylK3K1jNpR1RsycBLqs+qMFeS67oWiHF6qgoF
F4lQvfZHNofBHmYU1PNu82QyWgF78/GuWkAj3d09dN8waO3Sz6DF5mJFMq1s5LycidzzVadO+1Y0
rsf7iDhbfC9ohTlGzRBe9Su9JYI/bgHO+DOIuY3ESEGo/1zDJghnDZW86/yRIU2bE9m5jauKqDF3
q0GJ3psipoLSI4LhjDQzSFIsSqBDHTwL1817MDHBDS9+sYMP/NciVzoSjMGN5UFh3rA2ZUeaVgHk
PNjwge5ytcDaUHaOtjpO5LZ9Wba3sL2aQOk2sNjVm7nPuEYorRmqiB/7cKW2eSZxz4ljbcPtJzTg
/9mFILM9ebeaDMzHhsAxKNHHqkkrBi3j83kxpY9xno8NlsoNDZ1q5vPB6X7JFOoVGMJKhWEiI/1t
nO+4nC2TDNTPwFImezeKn9+KuSjtSRm0lXqhqbn9oRHvkdlm/AGmoRsH7+nEooaisY27zaex9/9q
JZ0Nywo/rPId03U5USkalLlLeAC7ql5zWtk8w9CYubczp3KOH6M7UNPyRsbQebEH19CyP9RTq4Fa
6JlQ2sF+NTgIwSt9WCpWPHQYGVHW6YZ7oZCCYJWdP/rNhe/8xhRtgiVa/7RV7n8g8fzr20c9w7DY
ZS6AN/Gwl/ux0V1IPNCufheqO8JS3Cj46tUb2cQGFwqtckjuETMtnRCcxx2xe14fP4JSKm8uhncX
Fd+ldjg94KqQrkwiwmLeLDwgdGfgBPTQT0yt+j/U1YHxU1cTT/x1NjdkgRA4C4bwMAK2+Go9YOOO
hzYrCVDHjIAKIErLml8uFskbLp2ENGPwXmlFLxQY5WlYM7ejkg6S8o3NjxA2gpYw024rbNvKJiU5
f/Mk7aKc+d/LNRwyk2HhgDcKm9ejknUM7xc8HfgXR0hzyqhU8hs5ZwZ9k0c2u9IZW4Gtf+3oV03y
A7uk9fy/WSl1b6BBv/zhPZ6n1kBO3/sGmnMyYbeoeLui1FG1LRziyLGHy8nTVIt92Lk4iwjTNm2l
Ky+tunBPDG6BtQ9XcjQR2++cQrG3PFtYI+fwDYe0XTV+cCF+n2PzRQfyyjJFZ7MhzeoK7ihRSSo6
MTRa0hcJKkBDqS3uSyEgcuN4FN6yvTLtfiOGuGKCiX9Nb7FCfxRWgzJyKXoy+xfm6aCF820OPZxQ
sAe2jY/VzsJE/2GsTAEfxbiBSTSkd0lj7CIHNWz+fqw8/uxQUoFe3e3TrOhevIY1gPh071LeCpJ+
3VOZZwzu2sqttcpWxdrL0sPqSm0pUFSiC36xlSbUNi2TtGrkJZU8RoRKk/Xclwa/U4hAuIFAZWNG
dTOZ0VbghnhTB0Ppk2p4aE4Uo9adgmMEHg2fuANm9HuUEEKvC3RZFU+/y4CVwFB7AZCJLnP9MTKL
LiNB49tk/BwyPAe8xxQqPZyuCZWYnA/HkFD/IbqD0+KE6326cCGWshh42wNnQCi9aY4Y46dLGYFs
lVmS2MFEGjt8TUsKImf6F1IcnDxscSRfjwe7WKoszwV9APF3jnyyFoVjWy5pBY5nRWBLpjITIHRJ
1waQYF1TGdcZWW6MRjaqp2axzrhlzQrs3f0q1BZY/CG4TppR1ABk6hshp0LlksC2jFr6ZUuL/mGH
eCTpkTX7hw892EmuKT4mdYY8Gg/YAir5aboEOU4l1VxYiMLp4NfmasLT1Wy2hrkIlPGTw6HOnFOm
eobUjgt9+Jwzyo2ihycflGuTICUhpv4BThNTSnSDa2PGJZcvs5JuBalaK1T507u27bPQglH/baOr
B+zjPkTXSGizEv53BPN+gaWOE5vj86lHDOAOR36Cei5R8SIBK0g5pauZ61FUhvvIwNVhlz0JI6zW
Lm+fmYxKajgRj8fdOy1hXcFIKtnKUIq5nDCtI1+c1ZlZoAR1TnE7rmY0FvH7H6wj89XihrigKYqQ
s3XcBG87rwcKDxZvO+lB/GSTp5tdm0ye3iqNDikkU9/nbRYRymL1N2PPyzv/kE8jzQvJjzuYURCX
ipX/lL5WmJ2kkGBHQjhyUaCDtxcWscs98Gz1pR538czpJhtpXFzHA+NGH7PzH6fMR8vUDIlR7eDz
uwb6PECUgSdnzLGwHO8Za9S5oYzIUMVNAvJty8vhTrf6/CjxshuoCuOR3yhPbV8GerqvkdKI7Xmn
FamUdwFkkAf765+KLI65ICV4fvuHmdIw1sa91lZR3Myo6HZA5KoVq3y6EPU65h3VQa+05K/EXRju
GTnbudsmvnhNTnmREkjcH4aERESVfnOn49oisrAVIzrkJZBdo6xpwIpdjmI4iWvidbapprInN4WO
hQQMvyS2+4veEYytdBmNovDeChWfxUJlRxkiqrPWU6GLkowpeYIpeYq/ag0h6t9EQ7bnV9M5CJGt
ImQIxyqsRiv07Q15nN/z4gxUMzBnLdGGiyRNpfsJnjK4fRbVUQOCv4pphexTdNbD1hgax5ETXPct
HLx8g4ec0noU+JTU+6lxp+LL+++2MAT/s6lInZyHgA3XqM88R/yXpwA0998Owsp0+mcK5dQze+Ug
ze5XgreNWwREm64QsyVKukhCtee7aIv4b27OT2p32Al4iG6XGrNxSGJmIolRSM8EgxNH+T0YZJY1
GCdHFv7l7hxDcWWk5VWTIngvH+XEEDkbayLO2JUfMt1x+1HZeRYmUNXattnOosgBrvWkzmMMLWaJ
uCC+7Lebh7k8JnPN1c3LXGHSoaASra9N4mIXbD09TF97Phtvr09oPvDxbrajiTjnfOJ0S3j8zMtN
f2l9bYlTIYNiLKbqn4ZP0J7KtDTN67gchF2Kke6441M5XMDohtwjZYd43ntfJ6YdMoH1je4QDGyA
RiOJXszjj8gIngNL4mQgJmEiXZzd3XgNHu6xeA2vQAIkRU278ihze0IMfIu/vPkmjLaunTEyWAXw
iH5pI2CZRBy/S1AY3S97Adg+10xlnlswirXtol0nKogv+EkBgyhESlHyW0WeNetIf4j2Xyi6LoSn
7VtxTFB5Q1LA/i73FWXG2JK9Axe/cbmi6myE7eO4l4rcLt5Ix+if0w38INJpXWgxq/bO3p4yIraT
9U3ubSE1YtABFjJyAWq/Rdx8FsVOVuZP9xxZ6eXCtqrW2olGpmtZYMM60P6atRQOwjfLbFt+Bo8G
IonKq4OVigNh7jmTt6a/eKJ8ekTk7cROLTEiSl/2Vyd2MdDTplYL/z+faM2K6mB0w3Xm5LHSMqJi
8QVhF0QA+wG8yU8mOi3mcb+im9+JXH3dODIUDeOrTpmpQyDgD4tNPgEm6d7cIfyl47S5ow0Ste8f
9qEjEqbWeQx9wi5z5iPj6454+du5XHmLzFZMfIcvJgs1UQYAAz2gaQ25C4HfP3fugd49+PQBd1u1
lYFSE9LKBSt8xo7QdPJrKYh6SCY7T2J9K5RKQEu2miuiAImfqbLmTPaZWHx87KSq421iP8PPO2aF
OxIrTO44CSXbBLQKPUV6nwTO49AWXOw6C4UZV7exYAZbmcH8ExNvxBZG0LVEJ2FIrOhcIBbjCo1Y
S+ZsOo/2bdHP7NjeFZOa57xL1Z7sZUgmWogKCzAM3HJF6ErB5aVqmk9huTFAu1KlG5XY6Yn7Qe1C
Y5fFBcC/ji1448Ons0T8v6l8FcG86l3RhB4naeDY7gHa32NYkIjImhGsSUK0dGH40XqhQ4YIy7Rg
H2Z3QanR1YI17FEwVORXKvCGv5ObSv0ppN9eyfQVQubpdDxpSlQWJPh8yiA7t64S0efxUup1vig3
dfyqJlQ60wxR1sJsFc5/F+cRXNfNBEVt2r1MCGNh7raeR78vjYKclWPJ/xB4HAQ+ZZ3Di/yDaI66
Zq75bJr6/eAlJ4F72NLyGbbYD7URCk8trm9bBDeYyqb/DYRsrIfOIoDiqrmUA8nXrvV+1At0+v7c
XFZuBHilbd9B7hTeSsxECCShdiQ2Gza6H9sRv35bnZjBZieSusVXB910XDsA54v5HDysPGlNfWIO
XarkfsNw+nqVu3psexqW0Gitv2bffsnxQu+OccDnOUhPx2BH7XuU3drxDZiX+yyu6jktv5Iuj3z/
KrBvnReQ8Lp2/uf82+Y8wa4+aRzi+7EsAjlylsmK64bYFVA1MC3aBzEOkVvgOL4OrGSWfP+yTCNz
q0eZuDnDZ5CzdkyBr5zdeiGMysROYxnrZAeWT1ApqdXuTkjl+HWnuVXhgZEexULn8dwUQvuczKj6
AystiC14RuXGyF3k5CO/6yZG4ujYMWgNm/OFL8UehzMetCTexBVZSdCk66HBfO46wDo4+7p81NKP
jSC3ALxrJXtf4F21eV5oeZgpOekvTwqXmMHyF09nIYnzPMZeyt6lYchcjHnyNMXzLQZgbuaHr7s9
GJ2/u5msbVIeZsCOQ75ze+okmXQgp+/o8r8U8X2LqSCNt4fI6s/6z0cqjn0oxov5LSseQiq2nXtb
5MuVDae5cfiYBWH6dapVxNeSbP682QYosSjQ2Ev0lsgnT6Pc0xYsoqLdd7xtWgkSkxjanEGB8VHZ
0pIXL7bnrZS2D7V6mkYACHN66GEhJDOF1R0Yyv50GS5SkZinQvlbP+83C3Vl0YDW+kVFf6BAdfko
2VLYHEW9X4W/7A2mZMGO5cmaX9XQu3lImZz4RgFeOa+STXvcVTaA7fOSHJQandvcDib24C4v1yfd
7vSDw9PyDVyzNDX+1V02YPZWpgO6bkUQq5DhJjb29wKC9HGAVcxoJLA7B8iPQE/M2YJSlffxOW9H
91N1uaMl50SGby1Jwi9qBRp+AG4aHeiN8jnqPYCwEUY86xv3FvYvTWzIMzdm0vB6aqrDDImeFpM6
vzUnoWVBWtNIc45Ux5y4yXHdcWkxsxZpVsLEjN+SnN6bhBLnAPHQ1RtHdRlOuU6JaDXrahHVAtdb
hky0ZlAH+DtaWxOSrmx7BGWYCya1uINPl2c7QgLQOPAg2/A1e3wzIw5pv3GJCVdj4+BUekhzU1fk
wHYQVhV31cJ6it7ouqjZbAfzNOZs0yT1zwRYdpEHzEinHRoQwnUO8LfukpHeul8jMtZ++utsUZjX
Vha3qnQJkFZeCTvNzN/XxCzZhsa9BvjQWHTZRyxBA2+gWjXfk5nP35wUIZntjH5/4G7s1C6VIdc/
zF9nxZwd1g889LlxMSnXkzrq7ZzQXqbNIofoFklb2yiQzUDSSxIwNQyvHCuAstQUISlrEqeFErpN
dl+yI82SNokmKHvjs5L6nBULJPkjzi6pCW0hpkOj+T8myT4yyxCa6bHqng1oV3wl6+BrXMKLNxHk
df9M4g9FecUR88UVEJ+3RsTghj2mVvP4ILniXeZTYCYZza2LoEd0V2pQ0XJIYPDXCDbpebvW+pim
swzJynnFXMG59owc/4Mwb6LtCPVkGu5l0qg3Lo26kjMqN9Zt0n5YivK4tDucSnga11EK+ObIR+YE
VWieVB2MygukCawo3R9MWPZjil7CnSHu7smeM1l+azfRUM5op5z5KeT/qQ18FCKsQhiNYk5SIHGg
Vs+U56nKtc8iRnsI1El0uBvTCENc1tYitiL7xokIMrVCg1osk6bKZgp87IWS2xBmATXd25/OWP6P
oV9h4h/wb38i2ch1oDtrCri/KdrFA//fxKeGWnO5s2P5XJ91QiGDmDVgRjPOWK/BWDXx6l1og4ig
d1bYhJEmiG+3T8+XYIeNCaXT3Byl8YrjPuF6e3SkH31hc6g3eiiIP8cgxWAZLIRhahwGjRoBsO1N
MiQmZf+HzLNA0SlMpfFMwJTkPaIq67q8gw4qOedYyqKLVsFeGCMosEqlnoQUPkRLOJ2ch+sxkeT9
pih2wRoAmtC5azLuxZAnQNuZefzxgTjE11sapgrkYCWlTUbgs4n4s0HFUtCYguRwKfdmcxCMo3qX
ciUbLYkIbcJYxHOAnY57MdDQKLHBCuJA73ZsLIjn+iaiGYzCxT+e36Y6AmrdfBjNxZoOQgyquS6J
3xS0TRMxAOqaMPugBydZbDl9I2OzqzX0RaXt7AdOic5PqD1ubWofcD/wEtt3M6YQWdU4vG6ItKJL
+KHTuB/iAWyzlo/MTKZ7/4eV/BlhMqtVjO0Pq+FgnHCLkm4Jbtztk3cStAVVRzym8cwq5cUrcmcW
W5Ttq0kRexJf0tFMr67EE+qbFVh0z6Jo50CaElDDGWCdKUvQFJo0riYfcKGn7GIwdZpATFSaSd9E
/IEsGOXRFOcEUPfSPbC/7OjR2Y7ROi1xkBvIE45+3ymIAxJqdj2u3AIigw0ChHitoa48k4WOUDm/
aBxTsbt0vVuyYIosccIHQW6uJpv4KzSx3TwaM1XwWshjnABErofAcrTOk07J2/P7vzVHPRdqwHrL
EDNA3bYb84+QUDXQTjo1ipM7itne4Qwt5Ma1BOnc05QNnwZf8dUR7EVYURhOnZVSNz53RN88jwKD
vI2/D8Ff4fPBvf55YOsEDgQUUTTGqeR29coeSXMgouXh3sKVOuBCN4EjUM6TPezs0EYKfUA6DQv6
OAGKvtd7VLVeEeZJod5lc+9dryGWzxDIzw8KRlT/Y6HyYTe09xJTJu09ahMLHSJ2l4va+ocJhQZM
GMoKKijqXcuiiwTAGK+N5K/aPXKwrnttV38HwDVs7GuirTZO+mBzLepmXstjVNhi1RFt9EU3ZCIk
BMagBsSBT723lgx+FOMr4p27kMAGE3+3vODrK7JA3+EP9H6fmS7BS61DBvBQBpyR+bJYXlQPMjS6
kezqNwOFsEPaofHfxv0KzuYfp4Vb2Me1O+Qw/+ZZc4hgfFz1X4g0sxEnCk+4Wp0eksa7ikL6IShU
GJpTkuiU92j8jpF9+eaKGL85gMR/uXjHbtYH9a27HrT6yuvLp5aHQXPifIUXwFtSy258GSxWnDZv
OglAM7D+ixI7yq4eS8oTKYsW1J8iQuqrj3e3CBpHZWMwIUiaVejqdr8GQw5p8mtHCTLrxMVtLcNo
yr7t0pluL4vsC7yeumbjqTay55SWGdEyI3K+v4wx2TOlz7273vp1VCRP2mtPryRSxb+hn95aZziM
mZjTysBsE3FTCB28Wc7pfEHFDA8agxEJs6Tt33wxLAcC6VFclcH90Y3tSWqhJ+pDcr/zTOVj/1h9
mRViulKXP4yjMJ/i5Ev/4WWcf5A8qzrO5NTZ51JpgJnZohnVXWbGWoGv6kIaV3vxPJBwsUaHPlsH
LFW7ZDyPLxVay8DRfVJm39Kn6oBOxfT3GFJXTp8hCbdis2F5nWoYL1EIqLd7r62aAKrjIj3OvbKJ
TouZSvW4zwgt19IQI/ccMK0XBhbY2avqbqzNrb/HyPKH8mmP7CN98h8F9uIEmlk6iNuxaifE/Jsm
1CBIp/aJSIbzCumaRgepQon0RCRN1Tf8YBc7ioPJdPgQMihfzPwBuY86MXOQseK4Q+xwt7g38dpe
nHBwiDG2laaMA928FNYd97RbMnqR6gmEvw4rrF8sLB2cTzITSvfBgrAkQmlrCbE3ahbPnPu+gh/q
Z9Dw4q01JDE943FZdTKLlmAgioMp8+jmQMPAg7Re0wvCVIjjSguhXZXn5TPt5oMvHE5ul5Q4dt39
dmffZnoCAO9zbKdMbaDukEEWPM7MixmaxDJ8ZBCLxy0GLwRNvWaqhtOb/hpJomU7IGH7Gt1Jw2jC
MFKLUCurNhZz9srQu7zTMte4DAmDOua+ZlFjyyN98oS9OYv1E/iiyitWuSJj4bBDWHVDdSFE55w1
zJt81nd64Az3ZHbgGGXg0xbGXFgEUH56iwIlZwj5Wxe+GJ/VsaADCPlCegA45I75INfPe+REp81l
2AW5MGpAuQHX67ivn4N7OsgM3CuFdrgsnI7xqkRr2eM9+JOf+EsWskyJcl/X4eszHWg+lWeN3RfZ
yiIt1H9DHlYen6p+VVWXwKJE9U52mP43997FmUNFgS9iHoRVxL+q9q9W7HTwv7p0Odc6OniGxVo6
TZd8+m+AZv7+67bPsSCh0wGkFj2kFr/RoFQxB+PXhPMjV5jYaxgpO6T7BbJG0kWQOAPgstZQ45A3
Hxkbrkh6N4iJXg0FfIBtk6a1mxVOAxxrkKvn3n2fvxfitZe0TjUrWKOWwrqnb9a4uDzXBlsGAYwH
7wpSR1lbyw1Ofz6tLUj9qrdSXx9D7GVs0pnXiBUEqZwI/jdhZdeCuAy/SZJazCjC4qZ6HnkDKvxX
qptfslSX85WqDxNJHiDSik8jttqhFkZwjdmoNngJvjRl3sFIlkIAl33IZXsU/RmiCiYUuzQlgBuU
+qmBy8pucy6ZLOjQ0fVKtmX48IZPRH2W6RfeuZACDrrTXLHpn/oSehIkq7u8993CQo0yBQvJfWUl
ppyOx8aFK7WkybIptobdLhyfp3xZK4pnMuyj3JyYSyuzDNyqBuXstohNaCtsEvq51zO2vhOy+5E+
QhxGlnlHqVVQ1mqSsuqTuz2teWZNs5L5VekWK/h6HntpYd8dHZP02MgZrfOPOqZDLJjvfFzJ2WU/
F4BlOr+VxwGZHFe+na55hkVlElkDSLaELuP/Dob0N8sRpIaZSblPpo7FhmPuUYM6fdutL3sJekdO
zwlYftFohZkzp6NB/4vO1bHAmFOxwI8tixXWw47DTB9O6jM/Y8lfeRFYwVMe2KrPN47SbyXQczoq
kEneq5XMpSuk45JNuajY0G+qN7ARVydRGvW5peY8DBU8m9WeJLilIJrLzi/UccBouk5pPCmYizSl
jcLf+OS9GUqqfheyKElOAD5j+hpr+4PQNGj1jIVnJzES42Y9AH2xH6HnAXtMhJbkOhQPm+3OIiJ3
hEIKEmTC9Ejs9OP8i9Q1YiFO+/Vvbd0TR+p7EZ1lPo3b2RBev/qORkubkJR6RfDmIIYBbg3LSXWM
Clwp3nOwLPG4rona5LlbTvW+3vZSickg808sYKvFCxRy/R0uG7RlJAne0kM0A1g4fE3xyGmSK7s8
R2J4Ouvr+gJYER8fP0cAVQMumOBHL3zXJBUx9YDmAqNXEANZkuOrDj97udH4NxhiYFek7RfkMzfG
KmH0GfI3LzqdPg3MTjQTz0+HhquDHXdt/xSmKZosQNBwwLETtdhBXnOXhTsSqIq97A2e9FYLSg60
xj5xXXOhb6mprSt2btDcZyp9sxkrYbeeyW5LKbaML91FGHYEmiQ16sKEKpJs0W85E+rz0N7D9nT/
K0B7vkxFyXQJaz5AGZkNjZTFo+OqUwFlCkzYEnxrHuMSWp9YozpX75UyOIkMfiRwqkns1m+z/KWb
QeRWdRXXftKKDDLUpny45swj3qmX6dqgejHHC3rHqwvKbFfZ6FyfcIkHszrIDKDyyTo0/rCbA8jV
UJSN4LMU5AUYdrrTTSm2PxuOEg2GExh0GqDhHlLlflSDPRfieISPsy1A7pkE1KPwXlvQVB0sgQpb
fQl4Difw2Nu4OFdyoG9cipxDObYDzheSdIO7Y2od6zh/hpsaRvkV7oL9tn9xnDQrg1k9S6V/EUvj
/aFdEUnGgedAIJNXndtjgmH78Tz3tZ/T+semXoY6y8jfgh17DLCEqKWdIG7P6fbPlKON9Eg5A+4v
+jqDI2km9nTvG9yeNFrOy1jNQ8iBPyVlakZKSBR8vH/Hh2jdivbiWvTnkwKFuNd4kh9xOda/KGGc
wPMQqiLGY8TBn4LYN6vxoIqD6UHE+g1/vzPa7d8rVKyTXHnDU/PcUO37KxYVR1U2jWyxZGobdhCj
xCgqK2NXyaz8zsHQ6d2o/cK9ky1FyGBAPW/2WRGq0+UJ7uF2494Y7tKtJM56Lx+EzNe8hTiha31A
+7Ckepd1iO/d4kvt0wJd+EQVAxKSBYUzuyp9PWmLEFg51w8/jUe/vYazIT7lNhUKun4cb/Hu/P3J
bE2c3MvxXXEskGDoaxWegvp/OIJ9QfPm4weK5eJDwWIw8cCFrOGqgrXlr9WRPsVoduwZXKZB7iF1
3ExnSKQcB+LLchcUHFhf4Ds9j+BEuHwIvuqCDVPiEywP8W5Yg+/U3ycdz0GeeYfeifD6hSen0MkJ
ZlT1F/7zTNUZjQ2Tfwas2kI67mxbomfBGffs5nST+uQcGheLeS6fk2zzWM/76z6tXNP0xBTohIhn
/hZuSfhOynMUDIeRoMAt4Er7BWbPl77Sm1Su3KJ+pggSZcNZgm3OUprvIoQmDYdQjdfNcdiewi5k
3grXe/6TGqkCZgi9wNd1cJC7qFWkP4JTvVeweS5fBCPyH9lr04Czdjb6Ogh97V87r3+iYVwt/8Y3
eiBcc+Dxs6WoACaKz9O+YEywBmm4I8jC5qN3NAwvgXVM5elG80vX88tLjww4oiNBbT9WrtFPi2Qv
1Asnd9BO8nFyvzSKy8XF1+ugW4dbmSVff40QIcJkQz1oJtfjJ6QwmfAv2vKlLlsA+y7LpH9o9zA7
bGJ0DYrDGZKYvesJkix9qqNIZSv/STZFS+ecA/dbwDux1VWlAYcytaAhxLDUH8TqrblfBI0il/uh
AmimvT/z7iAD2mQcEd0z4ecZG9SUMxVpGvCLn0QHIv2+hl3KGoCSHnq6hAxRKR7AfxOyt/lhn9zl
o7zWfDpDDOH04dKQvHdGy1yVhkjSXX0jcEohoGeSgy+rPbIyhnCQe9yaRMmIzxuIQqz6ePQg0rNw
9Q3SC/uPEXP/E7VaNilMISZvOtecw7ZiO8LdJoSTzEtZEqkjX5HIiHZQyk8EaPXbhVk+M2lAVhJy
ONohr7t3+FKYUxWFiioRp3IqRuSm1T//yTJ9LrEXduZdom/+J/gAaSokEz04f2Ial+46Zu+AhMCh
JyWIOzOj5HXes4+6CldhOFOCUVceUFbQwbM/1sml+h9SFwXzK6AbbojcmpQg0fYeeUd0YHkrruoS
qH7FyhZOcz4kr612HOs1n1hPhiupp0QgbO34UPdChWAvH9xkznrUqp5hpM9/WweN4BarmSiv3ctc
LG8H4AuYpjR/NyRRuJgLO49h4lTOZIoTAfhPjtncyMfITsjNHOwy2awgKqm7lMwtLeT0uPENqYA8
P0a0jUqi2v3gUCE2A59Urh6biaLe+c9XJpVMJkTXUHELml6C7UQzrXVkehfhfFy44xnY/vtdvuTb
n8/NV6V0EB24R1acSbZUGmXZN/rnvhz5IYo6OKcOPheH8lRoHOj1wvrOsV0x7hh81n1alRmMLRys
HXwCScByoiT4OGpiUU7sJSqvKMcxkzqx7cjXTp6pwl864+ZzVCqS+haSWCtNigcKwkdm/oJKx7eb
gzQKpkY6g+OuMH50HRD/9rm52Wmxygbw+8fguD0abe7B+PJNBcWcdddRvmynnM5ms2p0AAwTGW0U
K3YTYp/pmiygTwV5QKvTGSzHx59F4nQNY+AKE75GDiyeEwKj1t7vzarBDK1HGStgrP/9rC1Gi2Oe
Jl6Gi3+Zr/S/6ENFxUAqhoDyx40/+47YCcIb+bMurPA8zp5Zc1l2J5rqkGKFznpZw3W1RTkjXQeC
iUQn7bJuwEc/pevIN2UibbmYO9/NBmlSso2iV59HZiyJE/Gu0ayWKNIEiaSgiYfgacuyR8lsSfy6
phOj1yAqwDbFhQXpZEZXv/glVvleaNRz2ok4cldh/F5UvfY/bLpZs0sCVAweOsnXpIFyO7nZU1IX
xdVlWMYjCVeaTZJmjGYAFwNTHi8gtn6tKn02GsZN9V4F/8VIOYS7aFKTTqnEH95bh1/kCbr+0pgs
LFk8qPzl+hKrgD93YPhTu8u5hWYpurTklwFE77wNXtpwr9FvCGRI5iVS/1Gto0Zo1e3JjLcO9sBA
4+J/WLiDC8vAiyvL0ic4MGGEnps0xmkC9VazW2D632qbmLG2ST87HS54m5xak65Un3rvg8DBSjnp
9QyZbpekXz6CWY4qNne0UjCgUwAY7m9U/DwuWSFiYR1nxavR8n9K3Gs9NXa1ZXgkywVIeGpiQmeq
rd7crfPcvOa4ehs5fb7gM/cMsdyW4JjDjQxeFZS7aOpt79i8nMy7Mr57JD63QSlNuDkwmldhNyYc
w3KURi++uDVJpMbu9rMEk+EfNbcqj6zlfs3mQ0a8Qrl+YwwgjEqDLRt5qUmNQz3LkG/ofCDNxajF
PI5dJ1x5XITb5Xje31OnOm6XU5U+x3eojIoBLus+GFH/BhxWzsNXEEzpUEOnxi41NfA1J9uHeAMq
qweVHhLRl+LkM0mmB3h2Kbhhp9uNpHGk/gZaHtZQyxmiRjQZZ2Zq08DO8/BX8X4PVVaF0WmBfcGK
yuMHBwW7mG27HFDOi65LC+RR4EIJxReUr48ReDuQ40WKOrqE0azVcrjGdU8fiq9sxzbML1zv+52e
3/7x+oIqR8zp/dhfGej04MltlDbCeMKceY27lOP6me6mSAcXM5Z8iVuYygq77tjVg54spFL8Tz6A
dTMWGHO5TJCDfH5bu2bRjZcIk4j8CvoaaaFVGHBBBizysj3SeywD0eAKHNV9BCpk/pSZUZoRbRT4
+Z4SrGrhBgN8udXQTxw4RAOhDblEfcBQsW0C8Uo5bb1AJv86fzBQo3NGB0LKH4X0SsuayDn02d2F
yJ3Y2oKM/YnEFd9gvgVnyvvJ3l0CCzpAVdMIMnBbe29EH+m5wT1gF+cd8KEwuGI8MrwgQxWsb7o7
OvzL03vHnaL0+N2uFEe+6Y3rWznmPYpVqevVqRqh/cKAX6GpMw+i8knHF2k7//SjhtyKYyFe+f21
kHV8IIPcp7QtwNJRBwMKa9l9oF9B9aJVKr/vV3Mbn5nZg8wPnqyTWMw6fadvN5LST+4aE7WLD7Ve
RzGh6CitfJSmV0YwXSylGH3/Muj3ujF+54MUIxxrP9USB+tW6zMvduja7wmHprZkjs55Uw8z5cGx
MGzZCA4Bwsm4/P92kNqXqTbpqml8g7ZJCCHwH3WfNgJ61lpPxgVnRg8yvz7UqOX220UK7Ufh3Bkw
CI9xY7asibC6m0WOrYnf9RohT7iDaNCSAJD6OsJx5pwvEdARDTjec5fR5d5Fc4pVkFgq6Xj9STlO
96RLjQoxHwHtDd4hkARCCY9y3Y528wqXpjSrazi/rOS8KX5H+utYzz/Lp1sXZyA0Xd2+8COt/Goq
s4uw+hbwtvw+t2cTRMBFVP8rMHPa2K3c6cLyE/sEsU1vqRaXq9RPBes1zCSxTwG6pMrcCurJ463s
N3K0elIPe3a1YM60zE4NqQPKPRTQfCjKwwfc8GOFfa40tUC8QnSVoRK2mcqTYw9o3esCDAGGV1kV
HZWkgrIGwt3XEyC4tggPWffpaU7ND+CRkHOclSdkxol4omPtA/WJ7/4t3GzVLmNt6kt9rF3QkvYI
hHJvRgrbkn95P7b584+uaoOny3nIPlbNXKU4KpOPIkjA78tZCKjaL+0hqivQGwW3onao+sPBRHkR
PJGW9pS1Vd8QGDN4FQzIguT0H2wiZFKjhFDgGY71JrdOYZIkuChFbjoBmi7nZ2vzYVR5GRUoNBBZ
tBKNxS7lrLPGZmuurflda1zhmIJE3FxAzqCkISpd83i387ums0O5QjJ2DTwUuBzrP38dKWTiMfo3
HXFXdT5iO8HMT2eb3DrRW6r5b6ZkYFlWGuNgCzV18kk9rsjX0gBJlt86zT6WGfHbnqcSp4QvcuZ+
97ik2BRl4z/Orj+ycHO2V9LdNkbloQE3PZRsoohxil4m8kzeWW2cG8SGUTdiJFIdJBuq/NOMWVbl
urv0kSmWPnwyaDRwoz7nR12ukGBdvd5WX0hy4Y1ejNoZWb6pKkZ1j1B0c/cXpN5TzF5vM0zrI9hQ
nmDHvatHiPCkHak2TuddK5uP0mVRBVtC6Ar+i6SpEKCyGXUyZB2GV3Kcmy06OIn8HiaImoxyOks6
1JWGijQp/omYOpSQ0UchZXlhXCcOSFqdNrrprr2cYEOxiXCtsu570xMK0o8UnvG6/X9izlADgKEG
uBqC7baus9aw3FrXLZUS5YpY+3HO648xB3RN7MW0MfSgAPoZTbAJIGwojgg8sheZS7LgHpmkDYGK
mkTCue3hpK3PMpY/J/YRofHuxQcZulNwTr9/+Gkhsa1oT7QmBB0vO+ZIn5zD0MXW6irL3DjDF1Qu
4k4c0eMQBTrGYaze0mrIYQoxsk20CXtRA0hAkiyDJW/b8ozIt0LkGTRnTkm3e+shYzAKGo62+3BC
sGg333XnQFeInbVySDm/8gUiunuYQQ8WOxv8ddEsVZrHjE5d0i4WKpajUeFjySNc6fEu93EksXfG
I8k1HU0G/CW9w54pJ0uM34gthQUeJ4umzRecZrhlOH3n3+SqQw8U3wWcjSibVRHJyv7eZzKWWOM+
eGTmz3MiAaO9I0VHSKZg5SRoLYkQSgsQDQwIaAmPB8TgdLFuwioyj7r8mo+OFRSSLJT/ewtZDCBD
w2hvktD1KOk6RWypFjmPslZE1cjEVibYAglj0jorhXYTnJVkUTGVC+hXgC/mv2TBjO/33aRAYTvz
dGkRplfN6+DlU4P6q1ixL5q0wzrFuU7lYfVfE4d4rKhak4la6eQgVGz/CPk/uSv8dSn+rFW64165
f7Pkv5goawhG4Brl15+VQwuG8EfLHI9DnJjWcvEDC7zXBPrFiJUmYVOsfbEZyihE2/Tc2JQDn4AA
oTwxVYxrTCNTDTn93oNDZAIpd7TnT4VEr48h7CY1JzETLW4uT1n5I7gNoeqfhMe2kLB7AR6Jc9kd
XP50DgO4BZwwdQXpXQwosHbzwuJG2JH8B4EWMcz/UOqvSg5zVOMVgFNpAjyC7t0vt0NiHtrUh4Yb
9NxaERREH9ceK/AicwQ/OzlzvsWFPf8PXnC5b2tYVwOhIg2B8hwIyMPkg8430stvwoyRNzqxm7On
U7vCdy8iqeKErxO0yj8ZI1UJogCH/LIPl4xul3nWaVObbivcNzmS7iRGHm4VSpTzqIwOJ8sApn2r
ULLwjnJUpOrrOr/jWOjTcaNAGqKOPXH1VhPzFv3+kINkZPRYrc0VfVwrQQZSzCrovWpXZ33yDzdC
X/iuMHDYFzdavO/g5Rg9k3xJGSTECl/YwR+2GOeavPb3MEubnMs90aXz32EwYe5M2FIu58ulmtNn
s75QZC7cwf7Y42kMYztiYRqg9pFdKBnbu3p5bydtUPl4sOuCVsX983zekZGXvZHTMHTewlJZ3Wym
4IrTv+wz7ZmELWARGKMhfEKZgEpoiBqpgSG7f2kh2/xaXvSjo63qMKci2PWc0Zo8l63+DSi3gf6O
/iv3V1lKXNNcDv60g7kbZ2hdSMaPsDMoee9CjKW6UK6miIMXQccn0Jv5NcT2CULo/bFKHJ2Jo92q
imxtX40sy3K4AjxYKE5i1C35LaaWGhbm1w6rG47wip0W+xkKlWivVFnveXbYJu8SE98UyV35twXm
7fjel5Cay6vleBWGC0IQbmeH4+nBQFOX3vkl2hecOmloH9/A/G25rIvZcxgQy8w0S9SMqQGA4+J0
lkKdoa9axW9x2H1fBjYcI3DrkgSasteaZxVIqlaL4BKTBbSsq15ojQY+5CJpKxnZYilm0JDoVmUu
MQUB2cPY+8s58hg+dwrSRc9gsb9BF5dS84/pMIp3rRTgSlNiz1/Z3WjNI8ph5VzG5BlbXGT1CYaA
8jkEXJPiV9+4Q8DMKix5qQjJmO+ihpl4dlAXgZpGdaJ1dpajjF4ywoeJLI/q6nz9eJATOexeBtGQ
HHAqp0nB9Y9vfTT3tnAJNnFwZPKlcm9h+qcOwX+aC5GoVbzI70o/QVP5gPAEOdVess3hsB07zJHc
xFqOq4UrpA9IOMqVu+8REb/27H1AON36pm6mOnKGDT7l0ta6swVqfwuPebIG4q/ip9H0z4KjrL+A
sKeIQke5P/FP8V3veKbZCmqJ72mL1VmobhIeYJ7GrhfaLHsAvTA3u1UGY7ZDAfgne5HYr9p3aZVR
TvZvzvI/kPFUi22rDvhd+TjPNozq598uCqmbftHiDpHzLKk+nJ1JdqENFkduKasF/W23AIIG05jh
Xgk6jGqo1qZlKabM6DMylrVZMIzTdRil1PExON8ilUuEixQrL28LCF8DdU8A+XYxJNnn/GJPUr/2
rlctU3z/xCgzgjT6fye3VSDKBl71B+Sx3oKbVhwAT4Ze3yu5mQF9pi51mfa2Hd1uQP3RmFspyrwM
t1VEjDJqfU1TDke+jivlA+cSqVnKlBdCHUAEoJRaCiBO1TvurIy5xrSjQaDLVsJXDG66e5ZRYQIb
Z+n+GgtzObEkxxZnfuqq6apfby29k7VLaJOHsPMU1AojzTxEJSfJUb+vMZxYI9l7UovjVvSV4bHB
APu2ubbkipQqhGbRCYcuX5PmOK8DSaLVMtcxXplOz09phsR15t/a5Me7R1tINdjoi0/rR7wif+vp
mT5rQ5Zunet9+wCvYyeejNwey+05cibS09+Fk5tYVbL88Mmb+OYyPcfLAQN4Qf0lsTZV6K39cQNb
BZE8mioJklEvwgAczRFLMLPo/OBsb+m8bZbNXu/O24SlS6jMAhj8klUe7AAF3Rj195X6RcIDCwvj
JLk4FFWSas8+mIK2yOjEd50Ydh7tJu53isOSswo3zNEtqu6Vdp4wZAXFOO0iqtU7jeGRs+0c00UD
8Yy4lSQX61ijlUqd85EYRtezX1lbZh7VaWucZXRLDj8sYZtIvSdqBXYdsu2w1kAoS79QidU4mIlo
Lyhqpqs0x+mOb1wm8hUA4WfOWkd+fBBTpjoIxrFE38NYpgjxgJ08vEZidEafEG3ovv7U0pWccVnm
0ARb1bgeFkr+8exCTRJtRbdfzv0aMUuMirKou5E3yoFJsy3kgB01e64sWTooNppoZ0JNNRVtsHuZ
dlodwONR6bnzElJjdwmCsnIUDseNSDpbp7Y8HJZ88jiKf0OuADnjilOE7uJzgZ98Ujszg2N7KQxK
YzZ4ymoNJuHBDLnVzXb8BOASWxkoGQPJTz9Jl6v2FXs9fvZNUW7yjWKD5JYUbhXdkTvXAbTP9/96
mnvWuFS1GOvzc9rawUThjNazqtYcLvtVVN6Q+g04eQ2rVU1uVi84I6JS23TzL7Y/eIz8muM+8VZ6
09rOfyWMDSeBIIMqwas5i/0R6mjuo12shSUeykTcB5ptjOheFdxBl3/gcztEWRmMKlJg9E8L007d
/m62N9SemISEJDENvv/RBhh8IOMJgitnX5vWNLWOJlHx6Cd7fvs0IgMMzPPh489AS4fOb+x/xC9z
fxm/uf39nTEF61igg17pgqx0NIIcwFk2XTNfotjVY09O3ainHAzLRQV9X8WQGVEJD2Cw3w+jFqnR
VRfQScCXZsSgdWdpIVbtW6geiJR5wlhRgqlPPgvQUxe//qKcFqIt69VgaZSqf/6txIMZZ8p2O0H2
wnyTtSml//JuSiDbAtCu3NfOlEqF6Otyty0LMi0rFVUfYC4iK/ldiOJNN7Hnnf9Gi6uVdUuTvgBW
+p1tJ9EK09o5KXv9j/py6HhLFYfjTO8GpOXi8WtkSoPqaPIxisUbcgh5U3nRuhmOQ0ngKJWFyJRn
9WfaXUoYEHPRm+YrHke1mj2KIAD8IFvAL77NWT/G4nTmDbRiZPlvAQbPHF1tpxcHZ9Qv3zGQ5+1M
80L2tKn4Z9ir0qEfJpAdxi1tL6tU5T0Pk4ggJokhPn1sYgIaVn44NV+BNNwH6NeSnf2eoa3HZVTg
iFMyYxiXKG3RpYlUtxZcHkuxov8AsIkDi//4Sk/jST2nA3MHNKfd5pZIbcbkTvIi977brnSoqbFR
0WHZZT2nO8sjNxqcqxqIYiYkvXOduZ25L6gtkDOIfmu4Q4nxpPnS3FSTMGu2yKRrA99ibZ+F3zQN
Wf1rlu8Y0Rvm6tzFAVIxtkYGVXWTaE1fA4Mu0lDRiFiJ10p9yv5WeXB6U3Azmfx8x1eBy1zavOLz
TCP9UWRrITYbMtOeS2Ij8mG1qhu/6VTFDhXJ3ro8uqfu84W9ROVSwLEoY1PCmDk0M5VWu7t/1mVY
47vp9rzQK61yqrtd4vQE8gDFA6A0XqqK90cqcnpQ6lzAbcXIxO+Wz0p2PIXnJ7uud3b0G6QbzTlR
p81rWy/jg4513qwRSDtu8Dk24nsG1821VQ+cvpeBsIW/ElifFij3N9+xZ0vu0bGUsSfvDA5XnDVS
5/SgKZEFFYE0wNk7Vr8u34NaYNtTbjkBXFRe6tDkyoXUC1npuvgCLOzshoKOGIlRJw4zHZTqJFEM
hm9SmCcnsTJOx/8P5Q3ihit3cEHbHxf6mn/1YrwrcIB4pIDuRP77K0m0aMvedqzqcPT+PXcgt0e2
kCY5NsbfkQSIELJO+vYBX3w5zJY4ipyKbS93B9N7oypTYFY6iu4uewMHNHBdfoDjqLw0QGyy+m67
JKaL0RrxIi3TQxzqptUD8iBDSpFHfcdEJjKqCqxb8xFPE4Z7RNzmYCk12YiVi/8FLUdSaOe/U8IC
2Fy22OQseVh2WJ5xX9tiA7hfWrEg4xYiLFBXUbChc14zCgB6smzvdUctk6L+vbgZYVEqK0pnFlT5
nLfYBzTeDSYOReYBbbgFWdrvoBPhEYwsGhb0aTvnGZqBA1KcXRt1OK7H+6dfpp5p6m8vY/kHC9Bn
t8UMfUq21mD5Fp4rrmXPCGMbD7VwpBl1gDxmpeDtMkmFldC6dfU1hlur8N5YAd9Ql2NPmmmC7SLb
NArP6jkT7w2UIQWGWFUqGMP91uEcdwcgd/lPs1RYEnbIfKKFxI6CrmWLC0xcv06083QTWLdR5Hnr
I3vjHUAcmV+8XwuifG2obrT0MYncpNqmlnit7trkKEM8HuJFtBA+zp1CIeaOwolKuNkrbMhuGezy
iXMFgCwAuKF97iWaLNXOhzwP7fvZE3cQS88wm80wPh10oCdL/fDq+dwgCN6zAfvEaRb/L/QZLzFG
WtvIT2A01uyi2M9IFUzGEpbaax2qwbIy1EBc7nbPGjRvY9dwVL8jcj5JqQzhEAXoBcyDwXfC9aZC
8ZgpMEJyUNvK8yu/TDzCwyH5UdV0v0LedvgA16CUCinbhQzkMbTqly8Q49iqipDD8B/ocMt8mSGz
j+vlwRefntKDLx+RUVeUmYn1smOKb1bpgeL6ExZhu74E5rxTI0ChWyBr8oDaC9cO3cowV9U6kSy5
7HrOX0nt2ss6+Sxn2qonZ8e2VNR/tefbgZyodBBWA4Gz5HSpRziA6jyLPRBWHuHkWExPCZC1G2oV
EA5NlLcA4YKcmRL0lEA7wQAeVPhpop0YMR9asOkjySp7uXfGyKpddxx2MQhYGkAsD9oZfDJVBvTk
qMISK+gzHjhNDneNhg1IXjGUItRQ2lMVzaJ1W/2QI7MgaAPHOJxwyhznblb1O4PpgCVzCnptxGq9
PdN+EMuZ1QDfhZZgt9H/dUUZWP7ekVCv3ska5ccN8ma/oD2XsxuAjkb3V4MSbTyfkJbiTYd+xEw1
DB88/258zPaRllksVL7BhHBLZ0BUimHzKlpjMBKes6es/LaUK0T+wLc14VaFhsD4ra0am/Ta1twK
ns2AigBydlydgdMhKpOrrAW6fa+EQWyzVIAe9PKGOlBJtaIYgCAHXPJ96PCWyU2a/AgXUcTfAfCO
XO+egsvznHg9eNoO/3jEhCo/Q/f5ipReQ2ckYvNl2PKjKm1Zad0g6CHq/Sr5cmm3J2qHPAmLjO3V
0y0yfeoDZqMB0aUJ7blMHSMvicSuey/Upp4ekql1w3v8XS5cJvApMrrap5Ah22j/rg6DqYqnXkKR
QlmflaCQNca5pflQKAUoifH761v+qhqo8oBBUaSXLYF/cgFIN8X2cSFx2Zxk3nHzMLPb7PBlqp8p
MyqzPm9Uh156dYuZTOEttkNtoIXjknTl108WkvJeEPOhcnX8sCMvr8g1BoOqQyf78i3vIgWEXlIg
3ftDYxjBcQIQxV3CwtBXppjNlmBCVKy3y3pRVp0WuhubRcezvKv6j21fnoIu9f9jnc9ydIkKddLD
+LbLwy9lUW+QlAAPCdYYnQ8QXmXfBoZEjePOoWNzh8YLKe/LKZT1zz0ktYv24/yOeNcDa5JhcJhz
UDHPt8HVCY32vU+VCMsmNkKYbvbyY6OkNifnAwUBE2IaWSnWe8g65c20rc4e90LzS0FWqGzSOy3l
J27Qmq5hFya2jgWa2WoDow08/tnoDddRo7s1D7P2ryx8+vsHHIHvBLWrm0+5Z55SO9iSVitOg+6b
V7UT4j9IN/eaVONz+Tv5/ht67JECRlgQBOukqEtWIyO1326d2aoPyVpmkKkTQK0UVe7lC9h5NAw9
3tJe8Ve6m9/oZwe0bzc/UgRIFisTwSNshDiH0mNa003gVD09jzdlZmIZOsB0Vtcb+xxq41tiXp5X
GrNDMKD61uC1cP5vLIG+vkcM1ma+8CeztnA8ArauKICRQp2GZOj34XoKheD5W0rQSGye3tK2Vthh
b3P8xDjJFahw9noei0bbF1zgy9wYNKZnh57dgCxH0Kwes9TYY3LJxenENkFg/R6b6qsAH4eaCD3O
u0rh2XKDKoIramDsu/VHTq+q1uAYdhYdmWSSpBbm7QJ35JVD9nFSnBjgaX0BG8Mho+2791iphW9t
scOZ40yZHpKOkBdDrm81tQjlxQ2h/RPDwSYI86Vgy+08WDxQw1mQ9cL4mj/bIZOisrMlTRIk+mic
HE2iIj0esukAJ4HRmUW0uw6PwAOL7+TW4x6TXYyx9T5Nqd0f0LnDu300GVTZXD7ZDrm5Z19vqoM/
Qf03C8TpUn8yt4lPY2gyegDEQISJYpykQgQvyk731c+zjLE8gEiuvIkSuT2luIQZ/XgQEmAz2m7n
U9Ozc7O+mVdR45YUbHexm+O4ID0e8HcX6djB1h6mQPo2Cdhr/1dCYwvgbi4MNZH1wl/EFABw7mTl
HGYqzj9R08Ht5nSQ+07GAu3KoyyGnPcYAJoFSFOzjdjiJ00qeDf041k8DJlLKY9kLsINTp6Ii5Ro
+rcv9msXAyzaGY+oUrT35B81heXtVtPdRs6C2pj3Mivy7Ev7ve2YsqNbvq6EHM6PAsTekoYWDRer
KQ/riA81AquqdAdNKOzVRNROuPoygkNItAKrS/Y2LlLGGy1jFJJ6t9YHOso6aX1RY5QiwmR7OYij
o3pylvd9vI0u/eezmVrgSH+bluzUs8SV12B1OnPJaDlTTN4R3Vwlaz+KCjWAwt/6sPWkf7rbDdZw
zArPQbBG0fSQE23bOST0bjqqClzt9q6SEqBb8/ROjdTXy1t4MmlrrGgCXmE+Pzh6u+SjiTUf6eKW
P9ERywFdjwAHzt5naS6DTdLODNO3R6eryZAzFAksVkW6KK6qqzklhMUjoc+6r/39h4kU8wPqJnDW
fJ45MoS3l6LDzX1WdKaYIWC26yMBN92h9cwab3/XMvsYvMR2EmLWksB0GbVytBUwduyrw/TWQF25
exHFnb4s4VIzLzTF622j/cOWtcceYx8+XJjXqfNo/lvcLy0yRC0MfdqLPMtLL0nddJl8oK4x0a+L
jhEk4qeRte9qvoTZH4xiVhJgFs4hUhuCbWh694B6O6wbBkHWXO2ntjzIyzM22v/dlG2oW5VhaLwW
+t+KMjLo3z6rw5wSD9BpmZ5/otBA2zxOfp96seMcQ+ROKJHqKZd6/jzRpx/MnFkqDVwINCnvPf9x
qcA55ayF75X6TSABeQvPWrbjwhxPdJhrgFgLb9tM/LUdbF2i3wpHY+47CVXqB7wRvpv3FNNW5b4n
91m3YNZvnwFonYUfWyi9+cdt8DyYAeRKIe8A24jD3ln1fVAu7SyzqJoEPhSPpjfZK/Y8n3JJGkgx
eG4ujJDyUz7YpfvzRV4sqORMWwgbtuU+wpk1nLnH6R8cuOp869yUuV9q4zFhs7B/OAC7CPq3BStQ
YBCQi7AxRQ8yEqGt+73TAp6xeSNKQrIJYRG7i+HYbNHIPJI/Jh8QFKhOzanWb3q1Cn0dw3EBWwmn
pulZgQBEzNdbmIMlSu9TqaD0AOhmW2vaSXmvrTopFI30dVJavldC5K1IqxvvaD7VYCbFgvt01g6A
8O/FqJn+Sb1XRjPSCBiNddsQOt5NOtGH1Eaj2hV1NlKBBcZQ+75wE14XKMWuEhcZsDezHKNfui+/
mXXa2PBKsQBQqM4mUyG2qwU5cnZmXkJEds00863CZaJLVvtRzxPDzUywHpTDq8asp7PYNT1PiK6m
WySarz6yEWYMYXm5cf+fxKhSW3UPsheu11lSQNz2/46ItSdsiUWx5zjBFQQGar0nkkbbqVpVvgA/
RtSGSFHDt8P37lVPtIvvJPpKCx8ic8sNyeXVpYVjYlftT8ACrDZtTzroDdTTtCpiReAortDhhlpT
dJetO6lkC4TVeVGCvMwO+kJkA4XmwpBN4B9nWIPF5wrwnf6YQB1hKLaxvBDObILwSO2s+Jis9sIg
5HToGZ7Uik8F8c61TAnbncjxsq3BVP5liGGIQtjPJAN2KldRZwaoK/Yu/X6MX1ghS3e53oQnf9kY
IgYixWvlz0Sk8n4OUcqybG/Lm8TisCATP6iyfTtIAhoAUTeFbhOBH7lMOirWJv2vPMvUikt8RdT9
tHBYS4DbOzu3qRWPJW03y6n3i20/MYYEF/oaxF+Z4xN0ntHU7bMtOp1LfTOlipQ2AwqC16m3VVmD
c4lHQNdUyGK57rYezkBA5X32nHZyq7bytByNCgaXXJkKaDSu9mx6+aetCVbHA3YunKZLWhMBnoQ7
ptGjIvK0U9m4t4FyIDe/5ynZnYnTiWzr5hshs9xHHFHaQyUc83N0h0zy+uC7pd7bOYZX8ZDvQSKe
4UDjzJ5nxsDjgSiDEMZW2vscPXCKJqnW3092CJWfI794H3K69YCpewf1Rn973iJgLGx0I8BFDJmZ
fj/EjD8suP5YfdeEaTECEiWy/OHXC3wxvp7lytHDEU2v2/6A7sgoCl5L/QoydtBly4sSbGfefHW3
f9DDb0vyRfyBJ2i0+NxuQe5631LIC4pq3Z0LZTRGSwE9mCIRme/SNy4Y806n7U7RMis4bZzstZUe
4+xhTaTVX0rk0bSx6B47JfIjt466N9w2RFU6FfwuJbdT33PDXERT721FBuBajLc4GwOXRPxeQu83
2kANHkMfl0X1njz8cG0WDzPPiuy5ve4Dkxma0d+LW/ecWaBBjaSzmMUony0YzkKuI7tqYss9o/RV
6wVyRJaY8Eud0mrfKTDt+n//08ph7UTqpgLuxAidWbirElguqHsrKYkHRPwfHJXDDaDvh/1CY6WI
xG3Eoi7sPNU9VSD5un2DwrxIOfNwwLL469w0hJTiu+J+LJkQlgUHzs4SqI3/sUDYUha1TK53+b0L
5aBVkFcRO6n5+6yIdLaf59Y5sDE+iA8Fs5kw4XmCc3Lz0E/933vJ+tFVXsEyZj+HtEg6ErXKYxHG
yFMBi+IeLfpTiX1aZ1mHHYi+F1kpegQQBVTjAf3eLsmUfBzmrZokybGMhUe8/HnMt7QvuMjeWYPH
37RBVbU8ShfhIC+tmMkE3a7XOAu/pWBWjTS52lelc6bAp4DccssWK10pis3nwg/uu1OnvhHrwVTY
vroXfgxwEHlV+gA3YC6pWRDmXVK+deA5XVdwhE13kxPDTQxEXJfLf56yZW8nSkqbE2udWcH3+jCM
YDL3n2HfM+9a/fmsspoweDK86EBRnVjag4txq4hIauvlkqqtWQw65mUm8b32TJAPGgotac24ogYe
aCRQ80p5JlC7aucgMYhlB2z8GIq3i3cbdoYQo6h4Qi97pdFaGCvTfNO5GeMq8+ZbddnsLieF7LwH
x2i2FvuTpzDzHy80kuYSU3FE878wLdvLZ8IjgH+GDynZm+xcHp5AbmXXbGmJVuGvAxymIuFyJoCG
XixbsCvCgJzlPHktoUv9QadLGcW2As0mSUEIRAUgS3iPASjbP7imWPFEwirARSqfIJvE/GytWBpG
e/OhQbNt0ogmJQ+1rknz2l/Gu+6Vv/DQtcYmQHF8p8SqWSbDtT6p0zp6qBACjIrM6mriGcG5Vzvc
UV+kDBwmru4q2zXLzDFvYkfwfr57Rqf2um+3U5diSLJwPHrQxmY7NI5/pYrc2qRtb1RF6YmlRUmV
V7Bu2Nr+hiEpiKspkMgJHJ+EpZVFYTVuFpTjT8WcHZPGrbOJezPiKsOOORk8YgtmNkTlmZTLOvdp
RNlvb2fXpuzMZ7E24c7G0prhJUl125iyKcjdD2IKVR0X/iLEJ2su4h9jsO+xkbmmF1Ll4y0fafcn
je8y+UFBDEut1ep/Ih6sab0LbLtXsYb8wgREznYa8ZCn+Sa9Wyi4IfNJzg2CC99Lgnb4QM3oXPwa
lkL+Qv2CzmN8jbiqJhP9BT+P6z4Uz5LBscVkjMCW+ejLqcgkb6P9WAeIDZrm/FKawJIO5na947jt
/2B8LrHGkRmLH3DekT8scE+F3nVkmyPgI/UVR6HO71nUsMIe7g32jt5OSoQU5dtNi3+JkKPHLhmX
bTA2J6VwXO8Z1DQZOUNGAMvqFr1dyDsYHuU58DgFK3L3aCA/5a7I6cJLxbiEIFoG/jLqYvTZAsm5
xoYnUOYuC9T/4Dottpoar5JWPjdSUUuLFFy+YtD8FXxdLYLc4yxcaqV00edfH2Yk0vnfJapE8SYc
UtqMrR5ngmnMoixaCanxIx8x7mxeoDBzBlgazDwA5kaGCpBNJLOhE7zoXNDP8QqQF1pnuwDVJTfp
T+Qn+CTP9imMUBdbjmKY29vB7BYZ5iQntp+BDkgYDAyqyCWRWJU6QjLGHis61MBUfYjrmUqpjEhN
Rad+V9BY9+J05TNYOJdcyDOeNnhfa6oLXCc8g/E73uV9glBJPv53bobNuTFBtPzj1UDSNAEbQiD6
/yYclLqsnan56uhLUeErvKSvo/WwGkMvXRbn5PlAhXzoAR86f7hr8MEVvvaaAMCJhMyIXFkrDRNV
kiBYUDpG5YjnF/ur93bwhfz5FiOfTLVNMW6ljMhNaPeW55yeqvFRzP9tthLcGzIMfZbg/dPohUbL
e2L8K6PpQd5G4PPLNl3UGdNIpVH7RIeKdL6XbmXEOlHvb35ceAgCKUN2MT4lYE4Y3MTkA38WuHge
+xUbfrZawYyxzpJBQUqDUX6qlAaZdb+tY/r7A4e0eiuTzScv42XLWNfbz0dqG3BgyfdbwdDrZnMd
yzEgWLK03goMiHp2mI6oZ+8BCuHP/879pYzDucInEk7KVBPCPX4Ref+dE1rDlN/+4oXtruhcD4RN
Q6eS3FHlehyRqvOSF4QXO1/SYr4ZyJu4fFekGlQsZEqMS9sijh893HR6WnRvNPXNXce6RdPdxBKJ
dAJowuFNeJSPeZzM1gQg4uopbGFHGSyCmJqvyTv6cz0U9E/R1iEfnBilagjG1faPbxgSd6XwQwPl
W4CjCzx2F1+BugjBckDjJKl+Pkuiqj/JLm6yI+fZNXTb2QP6qxM3k54ID7cdTW/otA+5lrZWPau9
kgY0id/vll28B+lTNq9EY70EG7UKV5ljxbl9qrKD4uyyyf/66fR3ZoW1bnDyanO4vzl4pIo82vjU
9n3JoFOp3xmuhi96dxrHYiP/1nN5LdLYX+Bn4xxK1YbUqUYxvluI8Yz5auuJc82/ioJkt1DMC/KR
sooxHVT62XjNgklgNHIasErFxLOOHQQDffswLSgolvWmTl/k2MaGYimUl6yh8v3NHF+eI8y/rmF3
XTqLO89/LCMEF8p0kC7/+FHaNSNwwCJSzKsArd3Y+pEklP9ZiDwNYmM22heyvkkhwQoJsDwb2eES
emo36Mdpfibw62uNYmWHymcbrKTKCSK+i7NimcbGAQrdkLfHlJKDOIZQDF7QfPYo2po4A8qsTump
1rfTiiRkT3xIdg2/EEWxR9XHfIICT1oiydzsx8TIQZjgf/rO47mRNBwGDRjujsn8hD4P+v0LOWfI
I+3NlkwQ29xY2k0U635Gz7mH66yDQQzsdgPYY2WJ8BIHs6j80DfDqYKd8c93yhWbSGoPujg4bsWk
ScXAQsxnomfCiTAUw4s2m0a+HgA+BMSv2RGQiJhATl8ZN5SrouC6PSfJj4Qqt3FdVnQCApNGhQEB
MWMXnH02pv3lugEBOjZVc2mqXnBpxvcg6y1zYugfYv/qOnxlPv/NRHYJebfJnMjH5dk7jQTbtw8e
XXfIUEZRn9ClUQuPC4vw9sLkTKLLZ3V4SQnCVcIhowqMV1P/ANbysQdZR9OYLNVHWKv/x53FfUZK
w6ZE7SB4uhzBonrWvEZvU5UPAZ05c5HQJqLLWQC+pR4rKpgJezsmImbIVxaFD1bBFwRybyxhIdxZ
c/+BThvjHynJGUrq/k1BG9U2KVdXyBv2qX304AC9Qs3cPlrsG58n6r7ZDK7GanHz4+VZDKyogn2o
OKSODqfdA6KZcDm6QvJ0s4e7Oi7xmmUCGl8bGG79JEoJE8S2wTd0Y+UFj+c0AX+3sC+ZodTIbzwF
L46HRQ4/0LC5QyMPnHjYyfb9bxKBwF/ma7pMFiNMXRyu0AYiMN5wdN9XpH9Pa3rxe8MPMfo6noXg
rx52DYV3Pq48fQEc6SMu5BDZFdJV1W5/SoKCG/S3dI8Sk4sW+AlpA8P9n6ZL0RVaO3lcjxWExM69
m3inYjKKRB/G1qU9t5qdiTfxtQIziEc1WwoeRGGs0kM3yFKj/E5h2x79OXI+jikrpMJSg8Z/r6Jr
7yDbI84JZp5sYrJwOTUiktIknenoo3m3dPhs4p9NeNJFwcIHsr4udLcx4QNsB4bxw7e7M5Z6/wn6
7JcSYqDZkHwfkPpt/HJN8uzW/0seM9QdP7MQiVEJNQCW1aWAi1ug5huzXE1CaluPPw2jU0oYdoAM
SNYN+XJe/BMuyL+QoeFJ8NpJlEydZNFj7jxGOSsgthyBb5+tLtTkd/G+3KPqb+EgakOCLMlIX1os
rGLItOtbKDYDtDrbtlvN/KIflCeFJpEzNJP7RXxyvNMzmrIEQPRyos7cYriIbLd+CmXv0qt3tPg2
D2RFccQIEVx+zQRBSIsAy0bYkMAaft4oeXQZxmaYand0EG9Ky9LLhinCMuHDFcUiJ5b3LQQo3Hj3
dHUMI7SO0b/kh8B0AZ/IFnPq6eHXFYjeUKQI+hWzr0aG144ktvrvXQ4QJMB+3AI2Nce8RGHRwjrD
wLTL70gIqOwnG3ADG5VXj69WQXujLY/gFx/GI/wA4IYVA5rmhJRWWnR27hphXXmFrWU/brCT+bVu
V6hzsV2hwqYgv+CRqaUAu056obyeDZ6BheShN1GHhtQ86aX3IVAhClr1kFpyLLd1EvtMThKkCda8
7tISG304hqgovsjckMO2ZKpgNTcd/SI6Kkj+rscITfrng+RkRhdUkvItu8iwNVIlfrtaLjm8KgVT
QeyKAm1SMfAI6AKKuGR6lSIOd7fMrfefxTS4q4inMRHa/CjFBvTLgfN5jh32G5xH3Gq4xQFvvp2B
FJ0sjbaDaNrTWZbG8rLsAWZdDP0/n2Hqs1zlH63vmIRh03dZsqZqDGW3tqJ0XThir4iDMKiZRB3G
KnU2jDDX+O3Vxo6DEfsB+9GBYHfQC9gHO0wntSgRQzZr68QzmU8Rtjph6cOz2HrBJdokxzIa3a68
lwVb6uxuGXSr5moOoQrP6tan406ZwB3x/ARAQl0ncnVDLUwfpUbHM4FjlPUCLLmIQxfrxZLQ3D+1
h2CUR2uHLggOKlIvxeqLDNu5LOT0OVR+gyxhV03XonvvoigaULqkLfGdwtD0D+pAjG3Dsa9LiQnY
E0ARXpDKwdFo3q1CKUuJlY/of9aWq40I11jilZB35MlHYLn/KUS3pGJ7Zig5FGI7hRp72rtiGuDU
f/IvJgh48/oclzt/Zwy/SPP0lc6RtO8CauilUVdPh7Zbh0Fka2N5A63bRk/z2UO7Jw6LKRA3cxIE
WrO+8Cuieo3qL4ZzmVJV7j+rMSOKTG2mVh79WWZorir8qfeR/SQmTrd4ZfePckbkYsh03uFfLp5V
3vFPjR3bARmkdQBzRmQDvHDk1eC08QS0V8NZF4dCLO1fyCVCRjSiqz62lwIZVhUXZmvNC/NbQ9wT
w+ToFu6hUyZTC4/P0C4cxUPYzPRZze+3cHWrgnrkDo4aC5G7TvfQdM3WlS3o+rs4y14bhP9oPwg/
uZrC2mo2bm48gl95KoL/g/5sERBoBKyfiOgCI4do7vVgHQT05Totwdsju3qruDaOSD/xCypGXeXO
Sokzgu9b3qTubEEgBa2e/qgfn5NB2a4OdOSEqytQZl/JA0gW51DXuM9E6gASNZtem/BAaOqP/OWJ
JJWgMABQ6zA0Yg+XfuUgOzImpv/T5MxVJ8tGI0bGmMK7/zdDtKlXmDHV7HE5HhSbrb2CbDCFieR8
DZuzvY5MguVhU54OMersfNlQwv12xsgPKc1n13BKtH2XX5y48r/0VTkYbCc65QP2O71souh60Rmz
JP3nPtG9sW060m4nGwTZIx9Jwn4fmutAXzMFKmtMymT5DS9/fu2Sj47btQfmNLELIkG9nx5dJyIW
0kSSI9VIsEAOVS3FBYhNcmokoI9DNGHyVTS7GRUEiaPqCV2Eob0wehuLfcKLXulSdgtbKOGOl6NM
Z6SBoYi+xYSJCn9Ai7I/hf7yEC6r/Oj8ed4+fLwvRiu7JRd/IRXR1RR7w1Oy3RjjSfFTkEQ+4o4a
Vb6FcFf2NflGkPGjJRH+B7BNsS2PGGy6te59dR5Ez6jC234gqlZTwqlWEjgB1WHeFfgG2qCFDRNU
79IoolWbSmh3gVR7Au5syTt5iIOvbZZ+vcfW8i8EeHdHNINiSorkR/4cJTlF7XC50cMySYpctVYx
OEBPyxSA0rtAqrsufxi/+551bfz3GSmFYtx4tzxVkEBDiQsudrbRuGXXeib9Q4VhxIZs5CRR1aLI
Q3j4sAQZIijZVktUkulR/ynGLiVQUKpgMYp8IovAH2K7ClnDG/sdY6bSaRGkqfCmJjoq/gMYXO0K
KkZSuSwH9TmaIKXPpmN9rfN32ky9YDNc8ptvGnGpJGPZ+hiCJWRIEDvdLOQmSrSLnbn0Vy5U2uP9
FCUhVmOm8rPz5x9y9nGEz7D6i6VpllN4X4FLdCyoW9ywDeGRiNCa96LDKEsteO4gb2REVy05aRU6
6OLcH9sOrj81T1OjkLvAJk0O9Vwdu5XRk8SlLkb7PuIPnJxQTtXa9MUdCf6nJFuyGbypyEhLLNia
BaZ9WnJQZqF/zvqH5rlKTjhisM8lkM/pJoukphonS8ESe3+ms/bWZ+KGKvUQodTp5sSnJv0vAkfZ
M0PRprf6vwrDOq3T8AzVNsWAnGNI6l+5Q9SeYoSZVagSq028mgDoM7nt8T5tuLyWfpP8u7i1xDLQ
DPVdsgaCqmFGfSNKfD7o0kV9n50BqwZSNfyMs6ME8LY+Fa8CVw0K/nxs40L65W5nh6tPi71p3GUr
cdvo0WtcGjJBlufoWAumXGu1OAAWt15Lq7nWyR0joPDmO8WW6dqsbAzuygX3Hj5HyxtN2979FHp3
zYBu0tPgsmdfdFoUKW9PHqPgdDb4cRxhuwButl1CEG4bo5U+ew/UHljLZvdAl53T2VzF7g6+ttIX
XT1nM939KanvrtNU0J7JQBZPmU5wR0w4UrYVbOuc2UG4FYPbTfr6u4zdQwe0gZHSrpPbbo0l8HpZ
V1R2GOhxIWaiNtwsNc0+JemWO5mAVSQDTno3du8p0Ep+PVFQ9pXPpwQkcRQ1n+RtMzdHGTyQCYgs
nWAUEZ/ohSjFRaXP0FgLMjJ/fo8P5vhNvfl7aRykMxOoigqxGO4ul3gdOoWKagB+Rx7pX7WN0zbD
xDlL7nxnCqeNN157G1rc6QbOT6gLq32vfRGYV5/MdtJX0d3zNlDFVmPJHG8YfJK51IytfalE/xmx
RlKoxEYc/L7nJekcMZx7KJBRmpL4uTbsOCcs1EMWoky5kvQE5f6pSefMYY4JKu5Ec5rGB+ADdBgV
duwqhEhrzGUyWfSBLkqkCYlDVT3UY3MGtfQ6mZxQbv53sjqwW6fSu7BI4Lc1A3ejUhpwFF8Zc63g
WNo9oZpjOpK/5TelRKclvePtwxtNexU/n3uXM6I7b4ABeOS0B9ChEso42DfPq4RNepdJfickeJXU
c/Uc0ZjNWgpuYQ15ev8tyv7axGOOkmdatGTd5iGNBWC0S2YB84kTL8NT6nqI8xQ83XctttyKLRFh
cbsGFYP7dDPZtLvYeNptqE/7JenUO8LyifvSaZuLRYO99aagacyeuFAAWS6SaqLVRe8sg8wXaryG
zoD6sUPlW7+BFZMMzn0PnVoSW9e2Hf8rdkVQqcuJao8jpkr1O26JHzVvrr5Eqe72/Q9ubizizZi2
QxmwSZ3hItXhIsxfhmiuDHDdMPK2weNwKwNx8oy9l9PzGm/moY1V95Ou4e1OT+RKd+k1ysimLlb0
ktV2jn34HBHf2Jgyg92rc1bWXugbfekPVYPfD/geudLa4Q6oa81ex0hutXuNleQJWVeH7pe2smG1
qaw0vEavaR5DPbLql1h+du9JwvZQ+Nos3we61JaM+J/d3hEnLG5ySZMpXjBwr4cv1cLmjpahjHKp
FqIPrAFp8P5XEuKQduX5Isq2xV/brFEsQDGGXTtD54GDpDKqMAldzqI8NkEUQHi0ZGPhluBoikyH
lSLeF4yfhl5bjrOW66dEFDQ6pSOeLrPdc/rmNJ7458S5QuCve/1NtxL8oVFnPv/2Wg1oS44Yx7kl
egqWUbg27UwrcYeKZj+eBUqBC8R0EbMiliuO0uzDkWdkP6S7+ouZKa44cN61YavbPotUB//tMdl7
HsK50YYK+R9a9GwiqyRZIAle9WolbXlXeTEjpErHiJo0HNSPQ4JZppXmrUjUPaoaD0IuIcMdquo4
XkEu8ro5NZyMD4FWRU+CtjLVHGBU20tWBSqpc5LHqbvlk+AA3q0OrKWQsVuw9VoGmq5HDcpMxoFE
4UHOm1c+hpyVPkWXAeR8Yerp2h9YizjDErU1WFZ2RhYSZ4kDy+dYZHOd8Xw0KEvqAv2qmcDufGgd
BiEV2OQEBdUXQqszT7YCAOSiH1A+9vdkP7B6E7NHR5XEQyopKpsNFcrp72Jgvfctu8iG9Rsll1zv
PMvP7qiXgi7oVFr+yaSvltz2+FvK5ExL2YSVyu5OQHmsyNIaZCpLI28z1KmTo44erj/KlosWTrAv
fI2XR2lkF9uq8djLcvUz8Lm8o7+lVQsROVwjb8o3EOzRwsCwv16HzL70qlRydJ2im1jLXYiAFVNt
Oy7MzrcVmntzSBCJRHpXuDFEe0CuD2V1J7rz06qZjkmukOzlvWEvGNV58u9WaTPLP93dBWSuY/te
IbUqmDyT6MrRkN8CABjtMkZnNrVEXzk1dQYdUHF13swTWMa9A9iN78mMmCn0XZRIIsgTOeeIKM6q
CEYLwbSxUoAbWAxXW5kLUSkxe8KKIowAVLovh4wr9aOeRE6pxJRPFLcQ/wSVDyUSijRtGPSJ/Jkz
mPaMTbjIsuvcRshCyLzpXSL/BDjzBqJGZoccC8JZ6aZ79f25/PRVL//qOeiKQdNpB7SFnuaDiERo
dLnayex9uqIOwllYeIBayzOI4mBt75wS3lWnETrnVhwW8JEvvOeWPtopklHdZqMWycN01v1FJx+R
Qs2jxcRStDcbZs3vgnfePGEM8g36btbSAaO0zapV66yxDhfbEtHi028PBz1lYkZroSxd31mbwe81
R7X9JNnXkSpJni9xcIc9Q4FG5d33/Gt7GsBm1ca8ZF6W6SsB9Qy/bNLrwlAOcWfXnkcEEZIZujHI
4sOdLqRz3KfPhPeV5HDNXex13e+lpPm1QFybryBkLxLG3w4HMubO7obSt3RPAwZIXkG0chhI9RdN
t34galaQKixxX22kYjhrOaSPvOeov7Hr7yC3uGThipJJb68qLCbH3jm6KqnrSUoQqVTzkaE8VqKa
2YFEnR54MICGlcHdyp4J7UxtYtItjsZfNq9ul7yqJLoDq48gjhkz4oK0ZeKRg+1S6herTuv9Hup9
qw9OAdcoEYaeb/U1yHX4dkkF7qGfE0naFcb2JO8GlCZmhK8mGfQWIXqjIPwakKfMCOmcmF3Sel+y
pJwZVMcmolUifCRyZr0QpE8f4+sPqNbpneLox0aet2Qk9pM8nxi3O2QzYkm9bAfTJdWc/ix4gNbm
QpN6Ge08hibC3pLpKBMXjBY4/b6El0w62Zsn74vUMDjsxUUJrX4l+PwbRkBmhN44+qDc45oALuhv
RImKYuQYZ8uC2+tueAjcqMzlf38nHgqQ9DcYsI/PC3BgFODBw71qEbpQIEsJzYNL/6qZbbjqYPtQ
H53vIy46nSsBrL/uw3YTXebVs0lPyY2fxULTD3lDMJHSx5Ap/qfK2PYDMZBY5biAMlfZ3QGgyMJb
WUt71G5UFSKbhEptvlSuy/yVKS/53QT4khixLP1Ek8+pYeIZWW/5JQRFjMvBpHsVDl14FtJUQKJB
lRbnfUHPa7R2tI8ci1GoiDPDrCacZIfhIiIC8r5Vni/a7YjCO5ma2PRTug/VjA1+NyFV7tCWCWpQ
MC6NhixIaAvYW9O0Pzo2ZY2kSqr4he0igeeC3I7uKjLcQ63mRgHXmckzlmPU1nLPQmkVIeKscj3c
Xlns07FG5XwzT9KJpiW0/kMu3wkwvYx2KkS6XeK5ndhJbYwrdXIlNxgWJIB1MOGC+l3ZoCCxoS9c
XSCkrIfOYhoMItbjQ5Th085bw3RbMKU4Vzeng8IB7suo9corYnUy+Q+6LATAFnknDoHdjh8v5EkY
zrUV+LZ/depLbxHvZLPk9tOeYhwdCtCHIcMtF+kBReqnJpbbVCseov3peGeC07g3cVEd1e/y2Lbo
Gn8TGFiew5HPuS9SKYjUCopwhU+6idM0ksNiSOAaskUVosSOmjid8VA2iFJ4XeyL7hev8pwRkIEU
gbezZm0/py3yH7LZ+RNYJg5hpU9ks6NzlY/leFrPpGrSXTAtR0YrMoD5GBwV1Tpu5YBt/3QK3+Ia
Zd/gd8IXI5p/sCGllOqDTL9xVGPZ38x4MIPoiXv5nJUcIbtLhn1xSQfgA/yqV6hgg52L32l5cYdf
V9PQlNEKFf7tuggRxGnZJCNIkvi7zE++bNDMt4epPdqvbKQTGSOTOFv1pmq3QfgbvzIohXAp/Q5A
qb6iDP+zXeZmbifco+ClPc/tlvksfdXWkBnR3wG4eMU5X8u2zPumDPcKGcks1YQhK5AzVDmmEOlt
gfUbqSK5zgghQbR8pDa0N1EjZLDkuT/kF1z8DOiOIT13kyr2gvu5wt2ZROVBVlu2tMzL38EqD40k
gY2x9HSsH0RDSZkGUUAU5BbRCEE0xYBLlWedkon5KnNrqNWx1YWX4+cyBluvwfBpD3kNJ6tXF45B
ma7eQNNMan/wuMfMK9JbUPIKcsZBXofEwAwS/t1EF7vtCZZiDykcXv7LkzbbJNjfUOE/7PzxyIEH
8pVibrPSTMH7N77z74TSsUHczZvsbFS19doPfZl8LaPELL8JCSbpwX4GWv5M3+AZl3+Q/ykcYnlK
N3ovAvGLOigH6z3fM6MzHMcxm93m0IP1ZH86E1nfG05RE+jo6S+T6QWhQpoEaXVlhlS2UMgB3Cd+
10kmpWekeBtMuIiag5Yx/0EZeSihBJSvc/haNzPw1DB690YtXrRunYRtoA0F+ZEpusnSY46EeJNG
OJpPTP9AyRQkf+Eyi4r9NovxUg0PmmFgF9Z8/lnIKVvWfFeicBaa7Z+V23Rk03zzA6pUOOXrdNv6
10CtYI53x7soLVrT75CtBSnNtAhdEP79/tcSJZl/FU41KRgh+G1BDadupYmCJKN33JUtvYdjFzBi
Z7s/ydUw4RUy/0Os3uoVnBKMDENWgiegc77YxCmgQqT9zJ8AJqtFYskYHWGlTyZYmGOHrFa8JWFP
+jU0+0i2gRURUgllKp89SA+r4hsWVkH6edAlhwBGNQUJe92+236+nhrgLMAqjeWy8fa03UyKYk4g
R4FSlJwjpQITJeWizPAmseGC+xiTusUgCxKDsam/KLfIAAqV3TG5YggvC3nUgofu9cL8PVVpc4+z
OAMlNxhQILHuwzTrOK+yVgNDH/rBqd2X72pDOTLTxUlsdnjSHPR/YK2dwsjBNsW5G9c5n5aVhsz6
KIJtgLvW6W+MiimSFLuCf1U3N0IDLHUEYOgb0YnForKmMvw9KCTI38X5xvJUkHIcwKLGWgykPmDJ
jOQaGMHvHhNEzTRf8aQAtzb6h9b4h10AAP+GAM6UfFu+8rwwUMDxJsoKpiTUE9t482RyjtmigJ8z
aYCcUbah0X/fK8jEiCK0I2n/JyHLExfr+vdmb02dYguGtrF21N6C9FIKjZaZK1/6N88dqw46LKMG
EUdf9qfo79onTa7VFcK2lvh44QU1dDGMnJe61QLTaUlUAgS5Ie6XVEu+vktTKDiOp9nOhP0gP8Rc
Zd0NrxRyZfbrGEDM2e1tB6zeNsdRx5BwaCzncAdLYqSEUs8/BSHbTS9hPzGlzQr3Cuj+BnKMgM0R
KvDGwO6o8fhAw07674fh5eHttfRgcztgq7CBBnIwjd8PGSKMym3fUt14JPteKGCJa0zP36ooFKrT
GoPPB3y2c+0UrDcunc33mTTpJymJqHi9p1k7cYgmfd5tXo5nRHRHh/87FVRqfA0OZHUJMqfsIGgV
BOav5mke7uRn10W8lzcGxZIyqxw7ZZoimJe0Xg5NwtMLHxYEXSN3D5Kn0wyQ8i25P2GvYAQG3zrd
SDLjJ8X/4WAQubVHURZHloEorD/q5wCPiIYREhpQ7bEXiJPcoNLXLBEt14OxOAG88uMcqLrDQNZv
1zDNmehHCN/xaHiocr7hF1hgZ1HSteaVu7xHQMoP7P3MPqcadOCf80/9m5jzskQbC8jMfKagSMqO
ndYJIhbJGLqKJUMo6LQCbUl+Poz5xsVGELGzZ4ah7uWVT5/kYL03ep2dQBy2MsKUvnDhCFqUcPl4
qXP7rIcP6FFkwNuXEn2LYHcnz5g4rP52Buy+DokeqaTP0RHVGm1Xzim3sgHgvtuJfeRoGhqK5YOU
iXMP23qPdadtXlK+eMoA3vluYunDF+eQdUHotkBaw9jYfwgZp1KPBUc1fe3ePApe+YZhpLqLsK81
gX276nafHqjsZ5rLoUNOu0OdG6aMRJFA3H5ZZYk7B8MTtXSDZ8KHnwUdmCI+iH6JznTtYV3auAtz
t6AnVQCLFCazQCpLeJytHs4bcFbWrk4jX6Cuy59X4mMFeh4okxPCmJbE/BSmjuwxShItNd15eyAg
YmTqMDSS0KLBPMcVNkMPrSKbtuj1qJDNxCvgwqGKceZ6ZpE8VFj590sh3mCzgKMNr2K/SkV+sLQm
xb2LYxlqQMANg5pY7pRiXmLBvLaCpBOmIzlkk46Al+l9gxyDjeN8DbRM/eyVkzByDQYlnVXCRuUZ
IDOYSzH5GZuCis2lOmKYT3vv2xZ0Yp1Iha1zyZH3l8EeG6TuPkT3pm7UpmUR5eVeHIfvzY6N5IXW
YdRICxY7fWMWvAv9gA+vSUfkTYaTW8dvyH7qTcjKSKEzPHoGH9C+3kjWMtVZGG5qytJH2zZsP1pq
67xqNkFzWGUB9UwH5XhqCExuN/I3WqvGfW28mkYTYyOos8WFjN/LWMpUAx+GJIm0F+QUfYQNFeTA
+Or/f3w3L4C6IEo+5An8Wzlzwsc1ka34ffzQ1qQ4coa/XphaEJYhvNYtzrDhAfFJ9B+DHHf+bVXo
qJpdv8aOKFKA+H5JzHB1xiWOfBjL8zNSJ5p7UM3nIuUmwe6nvOB6q+zYpRLl3FFpYQuVeqEZz2LE
MvHKQYTWRT1o6t52mwpJci3BgL7Dky2Lht32gPc5NcM+qFe9TIz82aMF4RkyhgiDQul67Wk9o+Ar
AIfe6agueAOlo3XgotaEIOxbbQHqTj+4gFrrcUKMNLLFMy9DsOFlZouB/qhLfDYzYfuxqwHSy6JW
/Uwm3brL1cRCqrdPFuMgLC6i618HbR6d1IKYiwc0STv9fD4K7WAV3ZV8DS5voqRqFgCn63p8/RyC
CqpQj1b4x5DLxOaaZ/X+Z29c627Lw3GgBLzJwUmVbFB95ZMgenZpMmq/rVSNxsJ/eINwuBnKVDV4
ZKP9jVGXmqlF+lQyZnyRxEAoGU3GnUxcL8AnMoO49bE0+lWa7s+jp45rekMo5s7b95Ihp5J4qN4P
K6SpdO2HjyUwF3cYxL2Hgoo+m9RCDp7kzbjeAVywuoG10IUwNI93EA0XOviBZRSmDlMehJcx8TSX
uc+u+bS471zQ0+3PaRGn3uKdA8WYpXnLNMLE2AyBXWjSWRbPixm0STn1fmvXEaCsMkxQMMKYxfMh
mVEjvZrZWNrxlmEyGW+gke0qfgDJdFzo7WyTpZeBRfDBED0gkx9tT4Hb/gJGjBHedFi4n/AnYkXX
kfscHGD0CaWGNOWuYM6kEDD2VkMeQBK+04epLCy44JHZfabfZ1TrEAlEeOSwsfh86KIwBdNliETG
2IelxzNGKFwsXpeqWyCv6HdeljEzZ0Qtx2+lfEH5GseeFk22++2NL0A4m+wqBLwwVYKnVq2cVOD0
qxuZDCVQ3C7qHbGmGmnYKq0Gvdb9YKeZ6+tGE4sdUrKfnxMiXIB4ISERUsXzbnM/klRLDDgL/g03
I3Apm/dIXY1fKx8+VuZtGZfvMwbTcHBlzgxxdxZUqrKnsuCl6kGIMSDLbo0BLG65mfhYXEcnEvEU
johiAl8RnTbvH+53mZgTTNc5njUOGA+32aw+kasbeUu9YoaRA/2Qk/vrkHZBrlpnD8SkZetqDEGx
eqO/3o90KZiIM8tuqGluSJ4EX3fmmwD/2l6Q8GT27EVm30a3lvb7DsduNie10wrbuflI4GHbYSuu
8f44EZHpUwH2+g1w81TIdOzuZkIJvqf/FtKH51b74ouuw4mvY340Lj1Y4l97tMvnmizGqAfJQmfN
lTN/imbqB8PLoQVP5kXJ3SCbFjarbUMLos8b1NbJkXWItOudUj4BVYJ8g6Nhc1GCvQOOwmQp3ujL
QPZgSJJSI2LCAW4wypeDOpZgEzss0MptwMjy1beOISy47yUN8tNvuvFS1oSaFba6EaeiNFhs2amf
8sirGeePauD+DkzYkDXWkf3NhDaSa9T+BbYHGP4kReI1vxti2YG6OhLFeFP3RG5JovlkXLombcBW
yyQG7B/5aDo0LWGwwg35562rCyM4XvzdqdU6elgeAuvHoi2say9DvRbRkswIlQg76m0QxWIljz3m
2PikuR3whhbk8ck0K1+20WWFO3YzMskwwT1CPgLQO1TmPmGw4PoEuvofW8dhhrRiEgJRx54IoSAP
0fYmEpbtzcL6TjtCVYOlgN/ikaoyxd/0Ohv70UM/IJx9FXlPXoX4JGQsQgTK7AeUW779rm5noYiB
zUr7HCKMlO3I51Dx0OTHJAWfFWcdHRwwIKVYFsg5jTt5G0pvZn0kYRLBLyjz9iCLXRvHgPOv7yr5
5dMeC7k6L5z7758TQSHaZlr1z6AdgUdW7M+Xo7ezYInkSpeq61ubvZ7F30MamgD2kFYmq9WHzP51
3nemAxyGaEmn1pxdKSb8Bb1tY88jQTsxqNikYLO710ph6jCWHuEXIsqUIqyrMrKfVDJRu/Q/pmqS
Hr2Ngcwbrx5Dvj2D9ZokiXcV8tBvAQn3k9Gppukz3eaRNVrCYP0QqO6kRklUWuFhIKIhFY1B+MG7
O5QbuTKHTvevznUzrM3UINvajlJHnZONMwcQx9ei7XV3SaBCGXHTaE/I7THeoc/YygDTGNnE1MT2
ojsiD0S7VwH08x1EM4q5kcmoRb2dX7suE5M5Yei/253EZRkrZpLbyouzc6Ko+wbnutZ85v+hK/gg
UMK4SWbEQBgXTOlyN2CoA1hD8SQIa2g4G8GsDOVTQLxz0Raji31z4fy9U2JXxLqn5E6FjFytkBYl
VFYmUue+vi66/I9d9DdCuZEyH5TOrKRPXwmuLXTuFuuF0jm2UoECzaW42I/zCO10/Y7k1CCA3ARr
eDEkZFKW1dRJvuhyjL7IM6DpXmbINpgEBPG6ISCq+LN6aCws4zztD5WJ5v2YQTGERkyubw9yiQ9r
mvpNhlNix1dZ7Kg/dYXeBIYk26yO8iiDbhMZKhp7PxD1YimSfsDXm3Tpj2fiJzc6I8mpg/hn0U4T
X5P0dYeBu2gsVO4W2NBFp4Yux5QosBkAEvvj2DOcGVbi3lrSLkx/49fW7wsHR1PE0LjbxeMPygCz
0MP8a6ydDPgmaEyZBO0wN7U8pKR5CXECzjJPUrdExTKz/UpSQDChAUbzDRXAV2UcWP9qd/VCN80a
YwYG3QQ20DS06Pv/GkxktF0RtuYHxPPWckVVoCByrKMpW7/uj3pp47o4tUDmnPYnAWjW1dDyqA+K
zFpRzBhZU2siiC4qjUD8yvkVfAjiNrXNTeCK2chlWi5Qre5cjtxk5kHC5i2Mkt/k5ZxCQLBSjkLD
/N/eFwKWV3VY6wNclI60J17M/ZuvasT7NYwKBGsJVnbmcphU9Ct8ITlEtXGHVlnsyrX/BL+qmUG6
BZa80F5b8XCQFZR5Q69W+u2RGJWfRQ4ODchLEp8YNI1zh4OJ3dwSSkbtav8zRire56Niqvclz+v5
w37p0PHm5PgIdcNjEzVmB12jqpmRr6DAUeBG610UCzPY105rVMEL5t23NWr8J/TMmzDWtc9miL0p
BJVEI6AcZqT2AD8r4YSp/Gft2LayK0118Y77c/1aEDk7bPSySbijt+HxKVkWW5RinfSacC8W2JG5
F8y7ag5WSF15tnQTysKJE3lhdGOMgKiMWjfpHj2p3nQW1Sd2rhN1HfMCaaIeqMIvK2cHZU+jaCPM
hGVPKgW845cEcHBx36VeQmKIAJzJgIpNE994FIBppCPamU7owfGVe5V/UxoVOR20YlaLW23jlGba
WpmXG2DA+6OP7+xD7AzbOOQXo/B3o3pIcVIASVCpw8ZFkjv1oeEM0zmuM/Rfka3TKroRY1E7HBdQ
lfJVL8R29TmgmAf7xCGwipfKoaCKtay4wTSm5kP5qUatbCklOIi2VNtAlyJwwZWh0esZA6Lcxynl
8Mc3jsoukUxdhZFaAdDus0vAwa7/Iz2rFUs3b8myJkaFXWHOfgH9twVaw95rMFJNJ4zz9TDoXAGX
Nuek5tx1MoGGvtsuAtNnAmH0T8vMD3OGam/ckspOQoySX4KtAUFKJLSHX+BhD/gODeqhaDciyKrH
RAJ1q1fe9o7ly9i61D6jlvk0z9D3HlWNX4qge34W6I5QdwlVgS3sT5IUyh70MD20VgBKJg245Fr2
+igJpheaKtvMyt6jJzo+FfPFUE42mFlIuggN71vU6OWcpYBA43ZDKWkfHOpcWsvA2nLEW/YULS8x
vrwqiCKHa+U2H7iU7YoE7U8O54YEGIXjH9PBwNIYcJSRhZv/WQ+YtfM+IkLaP3iJwnReA5mWM7Md
pFffpB2xWibZ7GJbeV75Mzjly+lQhhBeqo5ty+QuyWMM25sDx6eEc31MXrDZTw++6bg5p39QdA0A
loPFFJVi7rZpdhTss6a8afziENu6wabIw33ff1LRvK28ONrqtv2xyXy8q6AWL525N7NsvrNs6xFH
JC5Re+t6NliI1xJ9thT+mIytNueAS6RGMZ4O18uZF8Quk0JjW5cDa5Djhdve/IqsxJkIv8vRLxqB
eaVvZU/SXEIXREWAjohlk3ZXY6ReRLPUu1ZdDxm9HgEN5w1g0fMJt96ctfbnT8GU3KfMVGfwF7zp
3CaNcXIKLwPZnJ6d6qESqWDllbkelMvZ6HJ+D1a+WSsWMviVbC8cisUNJ21jw8njUBYmHbraNaZU
2mC8wo4sBpPXedOj//9qCYLWNCKEXps1swW2sCXv0NWpVodrZBGtZo7JeHV1OflUUhccB4GazMje
QI/6VnkQmERVBaPHTYqQ1PsBGmj2g9qCrDmb1jrbqCUZkkxLH21VI26YOhVK7/KtReOejStvrhom
b8ptd0jv442KGH32DLTnzd4UN9+GSgT4zhwDKPRLH+Lgm1mAi2B2b6Qs44nVleRkO4Tdr91rlIEM
eZumh7DVYh4fmkAZNv6iFJ9gvi1RqBDu4cFBvqFckjyu7lfDUhdWSTbHS10rsVyfBICc1RSY422h
MwVw9WHX15LWkXLEp15IzWfqVuFMhSYsoGV51enUJ3F0CwEyeuvUD0Q3qg8ZwVA8AzyWcLzvFzZF
z0l+6Xnu+R8rIFdcyEuDHriLaTvndRGuSFRNNY4P8PHlxUwISEvA4gCVQCwMaAT01QYkyguUUoiT
Xcmtfz8L7DSCJ0xLrs7sIAoOzedrobgu39Yrr+dv1URtngdn2McT79oC2ehiHXOCHh/43//VvH7i
OgKeKyshud9or5WmHwqbdogE3Vv+IUL7bXSWB+lVO8Dbi+l41jYIYEJakaCBunrfmcb8TLgJdQHd
ztD+E13dhcoBLljrGE9AKdOjj8lxtywV8mf22SJEMUYYZ52B6C51vdjomWizTrpi0HtVe3KJ3u5R
7jbMJjBWpIVNH75leY+GQHjgySE61JZStDCc0abrLIf+B1UCZCq7HE5jvXodsIJh+OrT9bRjxS5H
8ZGLJ5/78qCMxr3sYdH5XqJ/H+7JHr1jPpwNbu7FWVkzsDGxnlxss8KEsVfVn2JXiBhEwzdFjWkL
FVGRg70haNFVjXfUyCt4nbnfnuameT2jwARSRmmnnnsRszu7NMeZeyladLBN++ej0FQTYwFq5s6m
QUYcqGly2dIQIDA8puuu7mseL5sw0UybDyrUeQcPYPZ79kWVK1dMSvURsvoXq0qYaoNJroc44T6h
X+1RMuJWwaG0v6M9xcJW+H3VoJhU1LvrCRKkGJXs12P+EFVoy2n+eNrdUGuc13z5Sm1LsQ+Jz0LG
TG7mAhtxCChn46xAJ8LMOhVc9K4Q/U8WePVfUw3s+ID6SWf2eTPCx/l6Hl34bd7RKTtCMG9HOBGo
IVWSGmzX/+3TL+Nu1lx1XI7KM4v/Wxpes8IcDjOpzvGWONUoPnCfwVJmiMrJFOJp8x6F9tzdkTav
uH/WeJxp0flLJjlPTnfwcPVMpmGcZQkxUX6RJfDuoQf+ivc1pd7cW3kZBxBj1opYvFCeCCdmuqsq
T7cKIAIu1Z4VPHMY4yRxZdpX/WNQzy+PsP5vj/jjP7aAWud8lJTNWaUC+gAnsMYUjC7vBpELv/GC
pQeQ0byj5UeUxMQWhayZMnAzbv4hfuthcqQO6d3aNuuZNOluC0BoGtVrU0/yj0Odke3lSV6y+hqT
4j2aQ6xtzd93tHOIU55GRbKYIULhJmRCvGpIolsBkpZ93PaKfHQk0jQSDgj44+6t7+kDkEYJO20Z
qq/E945jhEfNPXgwMRznLD+INehOSexDgJeF4pqsgChvJuMLQAG8OAUNMJElw5I01Z6cpxr+4ZEu
eWI46zgO9yegki4Do8h57lKugc70N1Bj7h+IlotR6syEmRzdsWrGi5tLdURIy+zISUb6pf3KRVwL
fWpRKSVrE8GMYGDp69YUA/YS6FecAI1T6bGGYGUQN0jzd4iSlcGiS0eL6ispjXnAHNLHwlq7gonq
UWyh0eZYkqaC5nOeaZaUOLTGpusMtB2upUSMQqyeS3m8QOB3MHq3amSG/2SVT18+UnjKIj+k3D73
UgJgAsWjy6w6zr0GJPkyBTvmv5LVXKtfzvi+g8XKIUhSSnOdEcJrqMhm1RLpyLW9Tg7zTveVB61w
k88Fn+uoSM/uPsxLRkQyScAi8dEn9vmzuCdDUdzJY/3C0hrVaXwB4cp593VwA0AgksjhD7C6EeTO
6lyheBhIIsK+DGx/v0zR34NIl0uP7Z0qxPbNnmwz5SgpTjU0bQipQX0v+8FIHyTLSTYnOMTqzP1H
d3+SefWzLpCFtFRJVgkVnmB8OjgGtM2apwndaeyvxAqOEOg6V8OzMPYhJoMAm2A4aWbZg7AEUUQx
H0dYQEn6uDH5aTmtFZeonateyoR43CF8xyOMfvn5+SXrRYhKaGZfjnztUpC7F96l1Ap0zopVDeQM
KxuaZL11C6XQgZNsvfZKYkY6Gux845p5CefnZqTc1EcXiXiCP6bLxeWqgGwrWld7Vg4Iixc/Ab3t
bpzP4qXDoIBd2A9lntu2/rHTxq/gjtAygjcFY+jCgRqM5moP5n0bnY2kMGORTQ5OIZPjB1Dvfo96
UdhaJpqTTcviIx+/iicRVfqIvc6dxX08pflUxRT43hVtqRlNKRFs9Wb7NSSLM7YSEenqSVjODIcm
xKoBtAnmsl2z4xtah5sbttUN7DHngek1mwGvPU5tYXyLcM9JvyqvRWhNl2fVQAWWDg3K6puvaSrd
cvGW6O4OspevR9ctnfNFpz01z/MQGnSBTNmsoI2fwxt+ci6BM2BmxkzGM1MPVFO6qUyuzziOgUae
okefmwn4D+pVjK1UtmsqQfB8sTOvMIioCzqzYBC0ZNCOw/txb4BqdLao66XRJvvW2y2vXVaPlA0o
Z84p2h4inpmFcGDASjUK2op9vfzl09KdY6PoJdfXAI0mrhxjDJC/JZB+ETb37JwVl0unuI9byGAJ
ySmC42EkE8eCvXULHP3k8y38qX4hZ4d8zIZyif2MHJ2V7+sQlHsK85i3N9uicEfDW1F28v9qddR1
CSN/hiF5khEtrcjOIw8em0gLmwE4HeiXjnq1/OdN/mWfi7Eb29WzN0fn3nqNL9Ak497ryA75xG8B
z2ZMT3MZy//3ksWZNLsEVHPs8hmfSO1dUWjtUu6pai1rGEP4eGM4IY7LUE+/K03eKY3PW6S71wtY
s0DJNHoFlIXwPwyZgmVfokhYNxI+htWzezvl/lFuqB9p4jojGAptaPAVysexkz9jQ2VmKSORl/qd
hgOLDP2fhJLXmwKp+zaYTQz52Jp2B9ZKtwbRTxI9VbA60jbvPZxwBbGABoEHvh+RKcaXRvv8Sbzo
Ajg+QW6096n8Yhfx48+qc+IkW38/YwCDN2YE15w1sQUsiHhgxgTXtexHOPTpZTb3eEwFMDVqit1s
hEte+MlSf7H3jFIqOdxsS3LOyZ9qTWB7hrPwH3RXegrnL+rpVmjneJZ71u0mC2YwRK/DqBH0Q7TT
L1FoX5iv8gorMXRbyl0W1MweVAWaiMia+vVucCzQRuA3Fult6KbLb2ZubT5LQYW0D7Q1ClL1F0GV
lov3Tc53jvxRYCPiEdoyvPnVuiQ8II3MAW9yj2narXi0a3f5dgmPSOKrpR7y3u8nYL6261hzEhgJ
pr7Xp9g6OSVASxMal7wKeABPiNFnfbcojDnh8/JXXXHXOMufwPhicTh2fHiDra0ve9Fdrj004yYb
iIYjheCUd5SSVfG7W3zFe9gqc1V9mcCdYfvKTYd4ahCnY9MtggAVkkphFMQbUI1xn3mR9snpJZOF
NkkCXLzp4AR9Bf9GY34gZ/hRqqUZy5aCggSv+mXQzcZSlEv5Ya65KBdzBckt+E6u72W2uN8ieo/V
lsqPn4DATl9z01rsImzo+qMfTK2Gb2bUA+skwEt5F7gkRVKfNWznbwRuoHKoJjKGR5Zrp+KkQNdr
OYBdS/HoztxulWJIwhomHOObla0hOntdSyuXBqeu/6yDJg9tg3efZNoRbD5n60TsKNv1cVSzqlRw
yo3M6IiaxqjWITAi56x8Cjbr3H4NJ3Gk09Zjb8V3aMSTlBGNTwEw4vM0n/rQKbYPZaQ2GHfD1ePe
oGJoFpzO8BJMpjsroaXu7A+X8pGunPsbadANe30IjQyu15iwJjE14pKWF8OfpJI42i5An1FSDKbs
gQayQmQkmcSmrOyxmnlz4z2OlOJKXmbVd1pMDttxuiKxyLaIhCkdQ6SVbndB4f/+IAX8emnGBkYW
uItybVel2K4GQUfD3BOEozOrf5WbhI1v9ZNKbVhCKFstf2QAWCDp8NtPMQPtHqV8jLU0UsubXofd
Qp3NyKpYB271uCN84v9QGip12K1oFnuNx7X5pIWSrLpbJXIdikihdoduadPBgHjOyIYTA/Bn1J2d
qVI04ejzdBHp/kfw+mCeC5Xqmzl9cf9Wq5ugwB5hZWqZcEcJXmVScvejwQUvz2/YcIC8D92wNQ6W
2SEQmRbFzCqk3S2BsQkyBRe4rMlSuATcXL4EaBSK6Ts8GbNGPPE2rFMzyKpeOxIvQ2typA0z0rPQ
t54w4L9A7yu2ZNgXOTPzUvfnYWDBGEkX6M0dhUO8g+lB0jfT2fOLkc0IelKL+cVljvTEKHsV08yP
pliXL2zP/4l0WsPRqNlmOABcCr4uNwJVirQW7hp46fYQJ5DmPXIcXFDhcscf/JUrJ/eCOdN4Gkak
2tpyfTLAhaOULnf8PfPa6YAaRpQFzIvOcgGly7mDtxjpL0+mpkVhhVGTB6gj/EyggFz6EDQfxPNE
csE0nt8xt1FYQuNGS2uydBC0e7O4AVENp/UB1UEWvKkdGDH8xX24IyC35m2vjJpYxC5JoPrhYaxc
hqIJWjYRdUiLuouo8gK/M7V4qdK/XyRTvPgBCNX8+mVNHDbZlpKHHrXmdNU+G5FbdsMW++TejjN9
b0fGkSGHNrMJUJxiPFS3N4NwUmadLsMpBja39JrUM+pjR/47w8GvvU7s9cHyRGrAKtqprbLflVGq
GwzUV10IbKqv06a1K650AE6zNFecW3xbpzHYr/etAI7E17+7aR5ax6c/5bvXvhMS/FGbX+lbm4ka
1pxk/oJ+BBXa92F67SdwYzFIZSaZCAbqAkWSrEh/Qm4pHEv61GNJ4pg5hdKv6dGBUkeZGoQK+/9l
MjPMrcfh3SVAhsH31NagadXcUxcYXopmyBXNnw04RQ0+STKqafQDEDO6uh8pinVNgyNtluAbpySC
rMT+DoO5x9dKBd28V/Y/AuNsI/FFwVZoIhI2h3H+knS2tN5clyTQRxb5a849dTNxGm+Fcq6KDMA9
OR6s0xiyQfETENywYW+ZieB+ig6cBNAYyoMG0m0xBtt1SdDOXo2W2ASMQnXAYVE5xP4wdrETkJZ+
oL7oNt8oAXlpJtuRxUvIlIETC/s49JN9NEstQbJtntOXy/IKTH7lxMyljP8nv90We9epmCbedYJr
17YTz3UwNurGD2y7nXiULuFft3BysjROij1lAKDmkBG3R7IruJ5lNEbwW3XGKgPBLYRrhqPGmNv3
6eDo9rSkKn7SdJEqJZq08sEdgPIZ4oDmn9HiRUPHx0lOVeF+S9NhE0suuBeVnWUe/4bBdRyJh5YH
bHIePYumFzG7TUruoOClUwYAO0macOYSfwUg+BiAGI6AyznbqJBpsclJtoUS9KHTcFOZEOKELnE1
2d0d2E5zAb/6200rHM50ZQYS7MbThaU5UP6LQQpEUApAsKy+A7TCvLrFxfv3y03OcOY3oy8j5igv
ZE5GQLBGCyM9sl8yW5QZgfUGsBSH8JQgO+L75yzZEtbdbIw7Q0886N9Qw4Mpx9CAOJeGCp6D+Ruo
u2HEUuPFEzQMAE08ptj3HLbnfQ6ocOYx4pXIsD4lrdYrwSRK1ULz5kidR85v9Qr5k0YAq4s+L+Mh
9bysaP+HrW6UGDGXlbnyUjv+GkhrZZ93Eb2HsBDqdNwm3ov9uZD0LmVVIbgjX1PIrea3JjxXwW/c
glgABL0ZYm++Q1n/vfpazaoNb0/+LKQiyoc7hnWE6xI3Af5jmke3VCmTi72M5bSAxglPP/VYRxAP
ckR9ptGmc5mCNy0Ze16dwaqL+MWcSXsnX2gQTa4KFAFsGXVOPUxoBCQcZpK3p81gILb5aAh/5Tc1
+oz2clMov92kHWXc1NNbxBWeGymBa5PvG4sulzMYv1eqDyNCf5xGzCvL8/p71pBhcjrZIdOsNbOu
ZfBdegiIYtSoAp1ieffvRaG4PndgcNsSvRmL+jjwyoQoKbw9BCep8jqs+aelggnpxhumUSSN5RrK
g0sK11NesAB/OYPwxik1r/+CIh89yVwNJjBmlnEW6iFk9W9tBNYoy568hSpXhAuTr/5FSX3im91z
TtnlfFW4nX2Wm/FplV2NwyHqfAkLFX7rmyY/Td3cVgmAEhrIMv+hRvmwNPHgSc5+qiuyLk6u3/Cu
PJ2o7jqy75y3Of8l0angfuu1579r93F3/h/FDN7mgDpYWN029OU/h/DiKtrKxs3kRfmBke6lOecT
8ZZp1xFi7N5pf83i5YtNBxg+wiSIac+R+fOCjLjcYS7qfNdK8dTLWDG5d2ber/M/d1Shy9fRGqy2
WJWwl1WcBiRVsnSh2sfPSmKj5n2gAhJVZ5X3k8NmPHJi/ZhI/LL5S5f4wqneBUbrLX7yS+iILi6x
u3VVTToWR441Kmkz9rinNkcQWYUeFMrjjDk/byJdA82+W6iLnJWPfEAS1d1obyICYiwF7hwruKzg
CmuWIlHmICD12nFWX/ezQ0gaWcAMKCwAFDDJ5iwukBMG3ILQqdtlirJbXqgcVI6bJchYHcs+4uXV
umbBDMSw1T7PMFaKJN6OXEf8uYy/+CYsZW18flxTHE72++8ix7YLIBI/vF3gKFq9k66tu58bdzyW
ziHLTfMHZNkNR/UR6iuEzFpkGajMPz23W/A0YlKwx3Io4wGb7RedvOCssoKKu/5bKm7rvYtPLaBO
z2Td7WKj/lmUknnGM0lhwpPQA8PhXCpFdOow7+qroBPW9TKcZaL0jiNOAVtuUVmqYxWIUgLUXJuf
P2Y1Y7T+CT0GzY/fkWcEXv5vLvwnrPEvmjhDhDSoaZ+oDOAIZy4OiWR6hUPyNC2wyV5g3bYQDGUU
ODSuFsA6Hr1OAVD772UsW7hVwMf9iGDmTnRm6QY5KXbDa6EU/Pqu2qdccv92As+F+rLjP5nLG11h
kwe+bgdgKYYpRP6zQxsj0OGDCi7aIitNzmw+KbaIWepTQKJ2hKP3ZimS/nYUaSx0gb62dM1UvIf9
pURPe/6TGDfNAwGz+MiGQYdpta91jfpByjFmdFK6qDcgvJ/Zy1I3I8By47Gln2LMrtHtqAN//Mya
FYmAZSKuSJEzoqnSXSbuzz94lDx1oV19iiG7GJehGf5k/2dPYsSaVl0FCzBVv6jBZ+anxwBKi7WZ
39VEeE1+Eid9uv50Q0iD7+2xqC5r1N6lOMbUOLOVg5OxwfrUou7ggtnMHPszzBHASOGKVAZOBXWp
ghoRcscLfJJJC+Ogh8r9Kl48Bz/6drl+4ZHmeOK35GSue7jDWzFcFbQaHji+uWgEOa8XO7mxbv7r
iZU1YFz3ceoaCznMdYAxdjrKF5t7/JTJ2NOoH7TT9BxPpr5YsyZgIf6+hKuwxQa1TFW+O2oVlQj9
o4N1sk6MSEtoI0fmZ7RA5p5e3g6g2jw8T5zGHDEdGRbPj6Vf3nijqz2wEYGNEeeZ2FWUPA4erWRx
zrj1aMwc1FoO6N6gKrXDnB8kcUycpzsfMkE2dA0RYxRP3K3oBo37inwB7HXo5OZHqvM94p2p/0HT
0vCmUFJPRkWPos7Yns8RT+M5JW5XYO3c6xuc4hUcHGrF2YcY3GAokMm2peA60r7ELM7rLKjQn2jG
4khjs7x06R9dD+J6cI9ywL+d7hpOdEYdICfnazpx1QyQb4pAg15Qz9Z9Y31B/KuNlgpb0xnsN1jr
9iX+sjkY4yZA0dE8bODXyJC88ZWx2M8LF1JOFm4YlAqEjjh0B5+ykXWBNhKPWsUcHTHzmb8E8fr9
74lA1qTMhpBq+4jXB0vfy8fk6h+ak3toy9sXmiGutUy9KebHkLCRC2UR2tKDsyn4464kn1ZnLm9Y
p84zkUzBdi04zufcT5nOq6mXj7DNeWNX0pEQiYRDIEX74GED3u3Et9+QeGDCYyTLBTCAXR4ctn/m
GK3quZe5MVxria0FuT17J7Gz2jMyAnQVxPCcutVWHGJ/HFhdslliMTt4gDv2arWyGXyS2kvJyl0j
9InZss1qCpOawa4vYnDFHu/E7RAKmNnqXrgfgfRXSrxiO18Benw0NuCgOWRyuD9pohblE0UIrVPR
buxzPEbwXJX6C4JPGdr5wNhHRwfDszlTUOpBpPAHeErd3rNe5ZIMQaao0gfiIpLU1va8iwiFM4V5
mPCScTT9CC/eeivQz2YPEvPhnZev+e/n1MNLYb8PL8EMCiqb5uuNgv3l3+psSVA3FtimpWyiD8V+
bCFajWPsL3mG/seZLkEZ8lur1fjZL6wH4tmFnPDMP0/CGy4Ooy0vE0LmrkkT1g7JXwGkgQS9WzjA
9RnlWUCRV14e87GBDEmgfLUBmYoZ0zg1XXcyHM00lbYZFrTualI6xiK6cdrkt2XL2VDSkx8snD8o
AtIcgU2j1qHuoOG108ijt9DI/KEHs1hIZu+dOEZGPiEXmRIwaEMir4LhZeBbtpmTGI/aQK5Q2dJu
X+6LPqA/ewEqIjt2eFgRpAvl+GlcNl5JWoAtnLTktG6HrlhOiUHbPOAj+sK0/oxBhTRo1gLeOqnr
I0+oKt/OVhwTQof81VqmV9ORIiBySwrt3gl+vDLdwG+bOamzoAO/8IyeEpNC/QTqnxBmEMMlHKWm
eB8uyf7wCE5NxEFCh+uqcEPwM1sZzHbK7+DD5wCqeBTRwEOjR3xpB9yNuNIlvtjstSptpnUhF1ro
R5vqA7UywnF3Hz86vXHAZGP9FJ3hHM2JqL+mei652YLBCMN4IqhNgDYfmz9lo7eFaDtJk+Dh4a7k
g+RDjg1uO4y7sjNBdOz+GsIo6qued46xtzTeFecUBbpMGA4uuZb29fQ/4dsKd5rWfYq3Z5Ma/Wgn
z5KQWbMLLIj3P3MOnOxDh7eiHN27te2NizwtPSyhFNN/bdDT+UB0RvNdx0OwEEmZ9lwlDR5DdVr8
Y9QXNEC65tJIOXfOu0Z2YRmtSQgd/rYUjADQZ53dQgAkGJTkgRMS59cLlTjIPdMvnUlbfGt3Ke73
0Ub29M8MK9JhZOq7LLXd8Zo4MZIBrVHaj3DrjoZZjWZwahMLfC9xtlVqx+fUid90F6XiWCdf54fZ
twJQCoNWZIX2EMnMlNBxUJfxgMq5sQrSPxWhM31mwXrHt1zPTi8gzYfaYDEasLRM9PU0bpwbESoO
lgC7HvUFbnJU6++96AKbg/hwAeWVtbhkz6/jAK1z1pQI10JNcFiJvyVdwhD5EofukinmUlUVwrgB
pIdULT4bKaAenE5mBBdfdhMeQyn9W4BZ1piDG+pHI9Jqdw/BkUnoW/NfEjKRj5LWs2xMqHhZP3nU
JfiJr0uo+R32qShHIaFPhKw5E8zTOrkuCFJdv7p/a9cUrsD6lke3g8EIw27w8Je7svlZX7MSTobW
lN/UkuDA0a1BmZq2fjS0YZ/RQVgPI0cv+s2JB+JGnqVT9eGMiHvAjsRCjT0w0iQKDYSZ8u/6GYcL
a/WiIaH9+C3lB8WA6sh7180j3XswIT4Z72m5TTGTu75kdHhedMMk4xgZPLpJuENMBIZAqQjW8rxN
CB7J7iU+V9LHz40h37x4baiB/JjZyIsYLOgLFVmjtrg7hA7LGb+uXsrh8n0dqBI5waCpK45cSVGv
g+jOvAHEPeSiO6JSdWGx65tZcsWY2JI1MTdp/1nemo91TFpEvEgzaP4d+krLJerWWWJSpoOh+/Oq
WAH97d4J6/gIPhomRh3qXoYaWGzYPOF0p8BjoqLqMW0qAZNhBUu1g7TrWMoHcsbyi9vl9OZJ2uPu
8a3gXEWpMjZe7H/8Cj5G2u3xDJwiHLf1GVKSrQwu3v2skXmmKZ2HZ60IxV8u3r30BD+kHcOdh83/
++9z1C+Lv7fQ721Hx4qQyMm1yNPEdPOL/v2pJt8I1T1GtQbslRx+oDpDPghOSUkbWDmCKyQxAqfx
6mjY9kWoMtCXHFQwolbbzER3SqO0u1RlVRRxCT+qLnGre7K3YSfwc0f4m6cK7AV2j9PZzkHQRG+W
2KhaoS1nbQJJb/CT3DANo1AD+j3pkgqqU105WINGmXDXboE2gofEtYDSMMQ4WP07Z2UejrsnbuDo
GBYpGAOOctvnfm2S+5bAROuPFBn5g2fkA3AaDj6sVogqXyl2PXdRvPqQOfwrOrtt6e/C6YsSf4uJ
b2kZPhaSUVSO9AK9PX+QRiYPBvBJfP58W093EUJokoCOUDzP5ISPxrJj3uQXqxe1lkyE62pGkuZf
uY/Qtj7CByjBk7LRGBQs30eQdqf+3rdFYsMCl11prhXaoXBI3olBZbOkw+8HPQBBwsqZmPsRzddn
2aq+JfDo1mwKNUEhrJ941V0kA680gNcHjt/fq9F60Um73vhXuJYgq/g9fu0aFHqdE/7NtExlvGnF
qL5Poexa7DPxeVkuS7OyoMS3tEbeADJxxoaBULuQytFayIbqaCKDYs4OrXocDSayfUzdp/Mx5a0P
5htMpJMwEJuXRF2pa5FmoD7E0aNI9eC705hJIaZbq1h4PTDjoNcuw7D5IVaxUU3qGI6WyHOY/Fr7
a1J3PkKL6aIT7xD2os4lxQBjX3GwYtYK98RhEe9X/yqKp0sFyQ4ENm4pHfczK0VFf+Iek81rA97Z
mk4SN/AxfOIiU9Faxo5sZL4fYwSN9tH/efQKFxOV+tSv8S95lROjTXYwDmQbBd3o7Iv1AE2R6VNF
ebWGErJj/ENdpVUSZe4x4O41hFGTTg58x0vEDNsjKCv3Y9GGYPGmnyrXoeCnP1e1Jbvyk4uTqvjB
95TxCT/SqNDTgF3bHjOX7SseoR1aflqgVauWYyYR2UiUaOMGrPFzCRb2XqvXHr3pya7emW6aj9Gc
4gVOp9r8nk+P0gj839TCNwfZMIMDi36PNLgZXUJkK2RiifNvkAC02537iy9qQ1mSW7F2AmvTdjBD
zsAIb5cYsJPGWxmLD5J/OprqGwtj81738DdHv5eu3/dLQGYtP3c53EvNDbKdKaUvdD313SVgZl6k
CA9r0Ek3QYZyDSVYKX3hoahkfEqbB/ITLVSlXLCcWogkKxEzF5Y8YQl22AE0HjbJTMAflvRcnq89
qNTzkDEolbQs76bEEBbyTs/2OrsSfgflo3oFnGilcEulRF53ijoCPs4vHmIgj062n+s6fCV8SPdu
sbcoSioUQsKt7XZEdLdp8DKaAoZivz4w1A30KufmQepH8AmlmLZ58kOB1Xg2hGLO3izWgWcTyFq3
xa2RljiJgW9DcMuZiPsNrZIhhAkzK4wB7PhUHNiEQ5CfjnknXeF0ifg9flU0K8h6k5oaz6ItHfbG
FyjhhIO+2Jc8n5iJyZGKX8raOnYIvRt+XUWJRuMsmSadXE7P4KH5z31WHa6F5Bad4XMyFJo+IjbE
WNxZ1+NNKvWFd/xo9inWRDSO6DedGitlxXvxu8Ob2wCLeaEVsylmnms/lCiIgcDW16UGlNERoKEy
xcYmK81NVeCxsm5ALg04PoMAZTqPTpYRbhtm+wcQpLmAvErNHW2jzx8XxzkoGuHl0InfHCLtidGf
F/rd1DLMFQpoUi50t7perkH7cpRDVXDruKkPz6aq1lMwA2NbKxvNLvCKlBGJDUMc8belVLHhVah6
0ubrNtilrf3+PM1kGVBpszJMNfDzfzM9jnI08/8/KAejKhFxz1aXE0EuaTxlx091MzYZkUcniH+3
nllQl/SEuXPy0LUPC6fVhgi8h1qFPUettp1uccNzl+XTCGO2aQHC0iBraZIEGuLtzDVizg7XZopw
+NjkRQzK9AOUCPThAtA8zX4QIKvp6dwwDIqVnWqraQQib3XW6sFetA0OzYKKxgEn0KuLtGbniKKo
q9z75oYtBnlQXOVlCJ7muwqXhQjavqmLkSjD9hY6cUfmCzFnZPTWAl3QWTuZ5WsseqLxJ9+7rvWv
4XHywD9NuEfW1RL57NDHDkPTtcT4DEMsv3scXx2BRPmkoTnphI9pJs9pDOHRKbJtO2YO/DGEvthc
CKXFOQeS2/HgX5AhLXBWY25IDTAB4nBfYANmoAmfkTwiybkrAz0zH4p/OVLWvMeqkleIpI9fqRdn
YgWj+AzHvJ1S8es8Tf17Od9UcjqXXJW7aCzFKZY8lejqjsw2iyWv0ItFbg2TAsMsB2cVP69aAhpC
xPxK57JAMqmlAWDgWolkZehZ8Fzc05IQ64OFbdKduo2XvM/5AN0JS2Ry7qvZnCN1UHSUSIN98+Ra
K4FPbrFuqNyUDXPQ5NZllu9Hbwu9k6WS8IHN7j3QwFCx8T2GEMcOrZ6eANWFfwrZDJhsci1Ye3oB
dNqATb4dStXfARUtVrwQVSFofOf3SJeKr6VfGe9LCU9t8tCV8R9waJTtLpAgh2KP8/3iZ/4onaBn
NW1YfDsmcvGJQjVSFmLN7i/DnfxmwydHFyFOO+GQQSL9W4AUwDDEoLoOpF9BxqyaQoqurPLuTmx4
/R0xWOQ6koGLwyYhiegUQlMmFqLDM1izc7XTPou3kb/W9GgSYwNsLvAtv+V6ZngAMhfemfJGHmJZ
Oz74T0BsADrkh2/Yn70N87vGZU0i5LcP8y0O3h06ffXVAHToXgQFvuXWwevlI/y8aITTKFCxf+bA
RqZxeIdMFb1wktDbKvExR1Tvz/PgrpyfUlPhS6XQVX2iNTQROwq/f3a9raVlNrGjRoFigxBQv4QL
jSlIzKaZ0Vluj706DcVWdL4LxEbjcQpGOe1aTwui0tUCYRUWYur8pvRR6kXVd3U7BLtxBDsKhb8w
ByF0yrtrdlDvWMhmKCWBWFdtvopmeE+SJVLubwncqdtPxgUNvVw6gn4scoIrlj1ZwiWxu+me3BOF
Ohn1NTg1gdvf3t9bulduZ9ukf3XfJWARlOQ0mNnwyGcVGKhdSouG2QyFgkWvzynuYHuBOwxBM733
JE0RLkzqLU4RgIZO8lKFVbthsqVEU15cuh8Al2iEBaOua5K6XMPVrLUgx9iM/6B55ZE6ajQeCcis
f4G6W+AWAxk069ZL8sb6p6HMT/uM80jlm1Ax+RKETEdI/YakhJjarpfGEls8KkPvfpsdpnAbES0Y
283jS2k8cHwhWqqQ4NDDwQ3P2BC/zjE4pfhTvtj/ZbYhGtNqcTno6wGCACJO3R3bMgKB2vFDfix4
7A2aOg6xYwPHGLTRsnGFT4drDhNeOfrnSTS09dwqkp8NTiVoOI4GJa4S00cqhLrce17UwIJNA3sp
8dmjAoCDIL1VN4NxQK4vgsvGxck/Oqn8RMv7mrwbfDAkH2m2TOsX9HZ/ZY5bJJ3NyHcK5UqcMka2
u4VS1CO3iHs+L0ouil1kPahkNjoYG70QS8f/fdoYUJwA5v5RTXdR/4y5Eln6jtRpU4VafF1X3ShS
I3aWuastVE2ftGOxAv3nM0ev3aOMeb3KjVi93eu3BOcAvEaWt9IVh2WTegwhkkEbQFJMTFRWGmXZ
GR6qDhxm3zGr0HVDJQtz83aL4Tjg1wjSefWEEArheGIO0ePGh2GFhs39a7XJbAj/asOXNJhe1fQd
FT1eKk/dG99un/hpN1T8jSbkt8IIAod8le4nrzUuC+83Y58jJTi/YiZyd1lxBehKYETbuaRKpDxJ
A1dAELh3B0Jj1t4eo8dSJjeFeLm+oWEe+ApaeRJwLA42sATmU49yXvQ/YNPlMoUvZP3AbdGneMeq
9vs3IICuqb92B85pJanFhKc9GMV6snbBaCjbbLsErk5vNREQTDErzveR5C1zaCQ540A9SX1ajd7B
KxG1zOVdL7lk29Z8FxspDfqhsGEVBM+IkK5nKvQ1PZSjWjPHCVh0IAVm2kKD3zsef5o8Kim++DbU
gNQcf8BeZrIPRUCebdxFltamPxspT79BAcKhaKxZEycacEJQCwuA//5dbcUtdFlmlAKAFUM7VCWk
jNVWpBKw3ylKZ+0WyqTvej7lhHVWKp7l5GYopMRH+mJfiULm15RvTuA9+tF9RUD8yIDiK9VmqZx7
oUi5lLP5wYXQr+I0Z8lJG3+gqN7gAbcIQsZ6VVCKI1iqMtqx+j9iELRnDUMWuBmiSRJnyUkpfO7p
J+CT9IwHPFhY72lmpESQ3l7Gm+rlILwUgO/NTUYvTuMmiMmIiD5TZj9V632DEn2TTeRGBycxyDb/
p++UlCl9rQwf+1UtPd0YxoGfLkwxcjX0xCTZIhBBCV+eu9b8zE6LcMSjWqDExi9Tzj2hqTJt4hNG
AcA0OWeREGK0FMfQ5A8/dNEqQ8FXpm7UqkDCgszQQLUHxbfOVt4KwonMZ8g3S4e4u3zIAuafHGxA
evS++DfCnwYs6smViV8TT6Spsm1E0yh2lS0P2zunsKzNWtAQ91T1V9Aul+kkel5Y6O8tidLXHsxS
I7yt3UJVTTq6e37gkl+M5nlIU8Ey2/AU6fm5oDdci32aXKOdkJY87mOTfYmTgrCLf2ml9LRVpJf+
4RrckE/tjCmrKUIUHydwmoVEmF1UIDA0LXH5W4nQORztGnKIfDAtw0KZWX1QXMPlMJ1Nc6HPYQaS
dsV+EG0D07/Ms6roPgxUp7u6Jpd+UPM0L0x+fPOBFH3mtuoeW6caU55bx6fr1sPO5vFYKM2qB8NW
mRVPOEKspBrNV1DNYVOqGAX9l6B/TYxOERbpowBW/PjLm7rhey3aqR/XZYHivmahgkTKa8t9KPFi
mVjKoKKI/91jANvT2SHKgxpzwQaZdP8f8yvA0N/9yM8LF4FGo1a8MLx/YwGT7DM4BvQf3lWrQETv
WoSS/P1+CMA5Xhm50JE35hPC9zePicr/2pKosENABTGd9aJgYM3AyST0OqwkUoQkEmiFgYL+Sx5l
qkq9OfyGW1qN2linzR82Sb7BNl6HTA3YepXZMh0SkCXxbjktlbZ2Sky57PdFNpehJ2rSBPH1HSIe
QY4PPAX5TdShoXBec0FlHNmTpJXl90e5moiG7C9yZAwvB7ALkEAnXeqNjopzqYFTvbOx+HQ6KnN5
Gwx6CNLNfac5m0hhWJnADYP31OE1DU+QavzFZHa21iF69+Co0hwMFwqErAgfbiaiVJ+7A1UCjjnN
4a5M3WMT8BdVoKNBOxZ8YSR0wjDgvoKhTLfjLLQRTcx/H+Y1bH+HKHE3R8iatiM5srM+/ou3k3MK
SWS+QuHvfdC+ZCpGUMSe+brqtE+4XNxtfqCyQQ1sXbHBIx5bm1OpW2iic6VICLh7NqDXGuXfO+Ep
l0EnSo9IR0IR54u0fpHNFA+GjO3DLt50MGZA/6ZY5oM2Y8xR0fnpPAosOto275cUxC2FWbfyLOBd
kOf/bkAsA5pwLM6SrZ88KsmXygE9mdAP/sU3sthETtdQhMYKWL66m0ROLnfF0r8CiEo0HZlfgwRa
qwR396zYyVrPHV/u2QiZ2Qu/zR01BrzD4UFPtok/TTsZWQrXNXg8CozMMib9snrNMosrrqGAsfX1
9rhWdeueLzZjzoDgKVU6bKJb8gCI1mr3tFpAH+ebQrXDIARppGH7yZbLeiIDRE/8hHFfx5Ut/TmW
3nPH2kV9PYGL8tnGjTsU63Xb6luIZaX7PpaQIc1h/vvhODlHsuMvBNCd8L/plRpMXDBiktBGb6sn
3UqR4C+of9QBG8DxxX0X4NO4zMmgIwIeKDJHCdhZNCwHQQIzGP5d5cE+s86yJlXs4FG+ux14uaSq
TAIogdfv4j5xYzmkEThwlIl81v2Hke5z1UmpTP+5yRwbVw00xMQwobdJS7r1q93T8vYGgKJ0yenZ
eR1umv3y4zISyTZwk6OKOdpb2yJnehV+Dv2xML9psDQtFHp+27gzmNzvFZs7Xo2lLKibRcWR2OIa
S1tlIS+4XXB+hg1NIdY6+CgECj+aPDj1FH3JIz30RBk25XaiK4VyriNlUS6rjyULZ/h2i8wXerVm
rx2aPSBOTC9qD7DRno4utn36m3uNg7JDALhkjIgvaPPBu6HarxI7IWOhR+gYA1Uq92+KV1dFExI4
TzAvMDDQuSHJv5y1g+2mfsINf5h3d/fBpZu8YfdiecWDDJeYLB1YFR+rWH+J2YROF/d/uSeagj4K
GDpFdJXKugd0B3UtxWJFpRgOAr100LSHx4ugXCtUMtbq6WvuHd9FJ3eq1w43v9crkG1fF9mt3J6J
7+1HQ/8vhNG5GkbNqtQPkH2154unQazLi/KcVRKI4W2AlZrhv/ru5cRRxTZJ1yzt/JtI5pIA1XkO
sa/jewPGyVamDT0AkrSsuPf1+3z9nr2H3CJ0SA/UtnW5a1O53hKEYqL0W5V8nQRiqLpd9BlgHU8H
AM3z1MvfzhVyageMxPuaX8X31sE+hGmY1vBUKRvcmJyr182bEcgwYgENW0oNwtCH0d8DHLd2iR+m
m4QhRsy8qjQlUgY1Yi1LwGck0De8Qfkt9FdYR3T0PDdVYfKmEcbTfOoaC9qHeoP70nq6485bOyAI
LlzXqFm72UsK0cHZ4GhRfCPOe0Css0EeSM6XulXVrujJf4MT848cGZOYMfMkYoeXO2u54UNN3+nu
Bw+AMWXxyiq9QHqJR8GF2NVZRDUBRJUw2ZGWqmHTOrHdRYjoOhfdfh9eFtjqIukJXJ7wjuWdZlea
y9ZTUR3tRPE5Rok4EebmvcVCeLeQffP4pN+cgoH6tmkublWJ2Le1/ONX7OnxQaE6m28aS9tJ7D3f
T3rZb6vWIB0PJcbvwya7fLBSRYMmj10qJyabi5jy3BkHntm0I0KoTCvWd43swAZQbiiIVLXefJjc
qLyxBu77/ZS7X9rrBXPh3yWlVC/Yj2bDWqHag1ZV+JaUITL+J5ih37xFs5/cEpdLcV5d7+LxrvJa
9vKXNQIL5GsiFFWtSwyTlDzUhmvlTiqEK7sTaXQEe9BtT15XCpgpZd8N5RfazcPjuIJ5++3LbGEP
0AVIx6AoGulAHDKOZxumqtQE07xdLuCbZpKsGs9u0zg4fr2B/dAu65cwqosZS4zzFr9n79b/LDbo
VoJxd4iy+YcCJQeMtOALirntDd3DU2ecR+p9kInJ923M8ImVYPAqwQ7N0/tcWjuoAPCeTPyfoWet
ViQcvyakOuRgtd0MjktBxVH+CZcZFxU8egKc3yh0tQT8wHKU/WWPeXrqefVKnHbRgnzGya6Xr4El
Ub1eHycwxYF8fjKwH9vBMv1FJZN2YDpyY20m0rFCC/mVeUIyfjm6q0yrEQT1M2nHKnROG8zHK7KR
Exqm4BD8/cnLRr4vnmj17zAGw7uKiiyOQ631Y/yD47gGFbtUTXKZLw6OnwlBu3ktW7RpVsx7PiT4
ysetE2OcOavGOOYRJvYtRYflKhNgHYmTjao8ioDsCGS2tRy4glAqHd+fTdNyiHSYehjbh0WKpy4x
/aKuWJcvn/xb9xuSTfg696hrTIwnaamTtjMXbk5/9QYySt7mZTnimgfrH3UcISEJUBnZcsHZu/b4
mGm07Wacv5XEtfWYzwVD/FwR1AiYnA0CbYZ8V07mDQx+KWBMLsRi5xce0lJyr06fiSeLl3FbGDi8
uH+28TfsX/MvmZPEP1yEHwu+1MgKP4FyQfNLF4BXHbZQM0ow/jv2VqKS1L3MJsb+VcYuVXAqDnRO
RUmzAKF5Z2d8TokOcNVt6sXmg6oHnuoV/QZXBLH0tt8C31fAgmcplL6ciRxGOwJP6wDaRGa2eaDX
1sechTpO2FbDrHBvff9p/qGBKlk9Y50BNJSmMHfWer+ckp8otG+oQMdQ2QzSD8zF/pBth6getIUl
iGVO49dfrl9h93avPHyp3jlRVagiJlNFiqg0MEW7WnRHRIyLlkN74vOj9JdqHIhOpDgrcFFYM86Z
6ch/F7aj5LG2Jy+kCxWvRlQR3BB2TYKBJ8DfG5IUnAzBRs0adBjKaGhhXtv6GjQrPT1J14zU91XM
JsT6kKDXcR7yX7XHeQfGBjq8ZtCrFYUj0/jdfvqQwKnsM3Iju86mLEOUCCgHHXpUPs04V0kxeEjp
GrKqzg517RDSKmiQhNJFlR1mA+UKo14neuJbopkl/h231XszJPZ/qJgJf5m1H0gW7SidPMQCAhJD
UxYjGAnBoxeX537Wirn5rc9kyxDLAnjH07YRJkvPcbNfb6IE9YKrf+pZ7+UxtKVgljZ5PL0tE3s8
QvliqwcJBUHGG6fOryrGMNcUMR1Wd8ztNWJEziOrsCUEA9vyoBQdYdsTUnfOmDFmn3gppE9yjoLz
2YVUgPcoeiFvASNJE/n/sJtnj+N/YFyuBp86lLVojVXE3O6c1btAYMpMCk1lv6rU7zRxc3Qd1MGR
sxZpumAlE5Axa8uA1kQ7OTbpHGN8JUVZ5eS1o1y/lFZHcZn45cJdnxYGd8NXimqAr1PO7i38awQp
IqNziBCqJCf92ipsThY9O8G5Yo9GC2ieqi8vdGBzD7qYkyocFoF+DRID1vbrVDZNxvZTWfVnCzu/
Mu4ir8FQvwQPT8bSW1vFceE7MmPdaAEzdYvoCho0cJ2BeJtEieQUgTqiLeExyu404qx4Wrj48Ewt
N7weQXtrMAVoxrcDOb9uc+N559f8PRH7HeUlptNl35rZXk/Lg8Kc1w31x3RHwwYivpXOzXEV1xoj
/PvC3eeROTJtdkkBj6M2tbwjlsqOZhHjZ44vG+3UXo3yB2IwU9iU8d8Aui4OAMgimKyB01xBI7N9
LH6z1MdirqynvdfDETiiu5sgUr/85RmcZvekrhzPg2Pck+BlLeM2bu/G31ZeI38tRQDnX/TEK/ch
RsjBVa7akwmb1vSTSogi1gUhfqXyHqu1PGbBuz41ISM8G68HEgcklnPCsZ7AYYc/t6HTrJoQ0+fI
3rlmx6I9QhiIn/m7tF/IureIi6pHD+pbNF4KR2plUXrKO1L+UVwW/SSCxzqahtG9tMSv/wsXdaRq
eQ1PsM3hYF3FFybqE3NXGTin5+Wo3B3pHQJMmvpdyegxTMJPXHDinGtypRPT9lFTgojvpnowYJSL
adeKVFPxwVeVjPX+fNrt+ZEfwVXM39WbDGI13hm0e/NXQn1FzsSuG2lBWFby9wAE7a2hR87yARuu
YnvPt/FUMUaklSoN5BTOXgFc4mlWpnex/Q0zXBlIdfCDNbZhELXW9CuNSf9+Sck6H2Yxa2vzMf66
vLw1s6GT4opqybtRC0doInPWLfl6fZoFDFy4ov+HmFuRi3RyEUm2F2n0ddjtiGoJKVDCYcD90xuO
vNKPqbh74TRrdvP00WWcYNGVqmdcjqDSJi9/NkAOE25aF7UquCPzPgMkwv2/SVQMGlPwMmIsu09o
wvEBWX9kCETS+SWCRQZZvv3dJ5vyNZSFoUYuRj5FHYSlB3azxQv2fpeIQcegbzzaaTZc7KLTcm0t
7PWtuEs2jMudFRUeR2qOOdPI9rTb5QdWZ6yhZb89A+ez+akYeu/WEO4J0FhQ+heh1DTXVRZRSmxc
EGkKMOhQfMrCRMk5SdBzIFKW18lXp8jW8ENeyYmQpC0Y4hTD07LaWu7kXdGJIqiFZ7V68avyQljS
heX1l8iJCKDxy1ooavPtlm1RP8f3adVRxP2npBLBeJojyl/xTz6E8fJthBxJp+FuP6wKgL0XMX7H
PHxS9PKkjmVGeZ9HCP5kdKj4+UHjIvq68fsNtFCXkoN13tfbaBQwV7uEZd8wwyTL/BpkUP8dt7/8
MOGsQTZqoaj1iEmBxRTMpXZN+ThzaGHYwWXApcYDXh24vgnB2v3+kL2Zr9o7UwLqbV6rd5i6x4js
2IiNWA9jtW2XVlUYGjDb44QAojJ4Biiyg6h0+Rk66ywmL3Us5T3tkWnZ/9t6LRSb0SLvBoXLrBNo
kLz11nLk7UUU4bUKajeGBfPn6I2rawjCyjT+vSybFNIv/Ar/zUIrtAClOsHu4wzmXtwXeaCdur1E
QhGbR2q2pfoAigPiEpsxjZYViZWqYsCa31RPZIfb/HxnR8vaR+gF3RpXPxvn4H8dZDfuvAhM/K/m
35KXRtPQSukzkkxDZepgjiiN0MHO6meD/VIFozM4mM/i7TQpa4aAQ7kY0EKTRPEFamKlZib/lKcI
NmUJHA6fJS6nGUuerGYwsm9AvlmmBluWX8UyYoweqeDgR9xsMj9sZVUyL5E5E4QAzoqmHdI0p15h
2kOfT1A5c51HQa6TX7JM2xFuhAah5oQnyyJqPGpRxld+rmPYAhPeGNLrcwIITCPDw2TiO5JdZTUl
dqmwk4cb53Fv/rYHffLqNRGO2aQvuUy7OcBQ289GrroGHd7zwM1sBbspIqgFpiMmhTRUZ7ujX69d
jP6Y9RgY1WrjpMAhWzz5PBAdDUPGAdPrCRSXN3qYn9jFWk6Q+lFxNSJB3MoiQrs47/feLfGS7hHo
tmv+EZ1suqpNybTQlnqVNM5JkdqPgsKA9FVjbDW9twwI9/fx3d+OjKzzOLR4rliIQgYui1P1SzgU
4nu9GRnzcbCQESkJ0HsM2YUY6DAPH/fEhIulsnoMgv/ipG7ACNCXUjdHPlO8rBfPY/IhzXLJa6Yd
Fknm1qXIVeD3kiKJlhBUh4yWC8Brk+V3UdcVsK+i08sbXD3LniXWN7VWqone6HLmy2hoRgpcP1gk
1mEtn4f3e74b1Kz2+p8XHEaT0A8FGoUzqGd8nlWNDq6+UcLrt63YC7Rzx51HNCGJ8fZX1NMXvS+O
3MiEkZg0Hp7kZKtSZHiZAqFKrr9kp3+74JDVMcXzjPnd8IM58zT/Udr56uD/b3KzUJYNKqfmbVQp
wLpayerukOrjR/RMyEvTuTbjuPIv1P+Eqp3WxnPv07HUVu8tyMW1+WzMfck0LZ+QGDsWq9Ror5VV
d5B7NWfdYKIERTQlE2EjCuBwUeHuKoCIIwVEjSpVBsqn8TzgNZrvGh3JrTr2Fv5PHGwREjsagrOk
hH5N4zKqKWBS7pM9h3ZzQ8EQjkEsFV964Rwwd1hYFfIZHNlG5IAM8jqWHl8nBRZ9n/wBadFD3i+K
Wfsmk3iBx5pGHD+FlWwjMawS8QyAEldIkeduI2QRiRc3uQCpujnxi8R10+gZVsx9aeyE1BG48Cqx
2ZnWE5A61rvlSjmEzp6EgzbMAyBJttAr6eStV3vxzBB9bomlIoMq6XRZtVQ49PEKsXpplQT92tmO
s4L25TOCRXUuSFI91xbF+cLXDYCfmzkGeKvlhfn3O7IXyfUG0J7KljblV3Xm/wQN6GAdYQVvPDOC
LNNTzONsDC1ThFefPy/vrrgzsH5wG8hl3rsiLrjOjddEhwYzySZXrAqx0LhtbDrYteqp5jNRtsjo
fyAmk79ITRsGjCSlFgExmNGnKw2/BYrwShM5/5uaPzXbHeeyV+TAW4gFBG0Gvr9RCIlVyTC1YIxA
3rNEl2nvM3DzOBkzwIJaYu5tRQ2eF0KVxtv6VZpw3FWT4K29gQEyYeK26V7NFDMEdlls24lVrKol
U99h21zHlwHP3bMar2r9vTDIg8kTrjl+vVEvu+pUFtGBX1SC5zOQbJGsIcR55CaZQ3xSplAzWw/Q
2ZTh1oPX13CWqlXPTsh9a7VEIY4/bxgqDXaRdjy9NVbTeCdR6w9LpacEWOmlIn19mly9Cs76cWU9
NEJjgTD/IuBuxXRnG3bbhIA0B7ZjJG8j4Ue9JN8h25X7p8+tRB2IRDsksNUemex54B9fEWDSXG0F
uoQReOnyiu17w9IgtX1vCqvMrKVhdborT7UP+yFGGiq33LuCSD5c6k9SBcY7kN7brUPjDCJKzMQS
PFbKOH6vc5O6Q+5NOWV5kmzJxbgDb6JDkdxqOJB0PpDT+5pn8G7XYjyAukVW3mce8aHyEbt1hy3P
+/9rAdEoumR7H1LCPUDCMpg4xC2e9zsbnA4GpC8PsZSJoOlR+XpbE0uP1EYNKl5PQwZ6BzY+a5gD
DZH60PcLJH/DY4EyS3eF+Ig1/XrISvaWQfK+1RPU0KLSENuyNQ2gkIlSbOkgvx+5tqkpNCu5okBW
LomCtj50BUSO1iIG69liCbj3XqQZMKSGEgZqtoAuwQamdG7SNlTYHbCSbt2Tp7/hZKmU0dW7cWcy
2YjN0ETA7Mp29ldD1D0Su4CCimG1/X5WnbUiCXX2ruYCoarSW5aMoMkoTjSsTF5PtWR9ztdcBntT
gKYpMi5UIvcnSbA+iFssmrCtch0pfoouw9Ele7qAoMXRiKP9hV/wp8Fh3jCFzKxeE21kwR5rc+F7
HM5ZoS64PnvtP42uzVP/f2lKdZvSfTW5pZkavGhOq23jWLt2J+KbrpJTwnlvzfKJBCz8Q+E3Wobp
TSX+StM4t3RgFofinfgi1iAn3Hp3FWZNY+7ib9gnELBEKbu/p9XVkG6Bprjt2oQlTxgPYZNrhrCY
gNwywOV3Qb5KjZOUBZk3G9eno3XPUOIgI8ml14jLr/SbVVP/kCtU7UoFVzFFPJ9n6zXcKQdaoqpb
W4gmPQZMutFxE682ggx3Os7mm813nJvcy9msrYJNgfwMK3hZpO4oNWaafP5ZU7Azdv5dhaD5Z0bT
LJ51U1Clh3Pwh9DzvJOi5X5EhYvuPGT1d5RK7T8XJ0eGkDcpKr4GDF1LCikdIuNLKc9nZ+oI9CMq
hJiVaWngV8c8Bs/MHCWu9DLYbXoe7/3Tmcs+dHeatpQ7fOWrqYeCOQmJCdDskUYlz9V7siLjw5je
DecxsjAYBV7pJQKFwpQv74g+QBpgjdRAZrTIQNhUIKrVikTEG+HKZ3ZDXJKDm7uW5lF0yUd5Jz3Z
fJP3P4Ok4okK0ryfkp+X4dhQ663Njdb2b/sSiQ6HkVtuVVEPX9CH8FmM9NMI5CmHY9zsPWcMI+rw
5cDIuPaKVhEEGiSTDiufzipw3I2YluMnWlDOhV+29EdIssCCgnutPBCBMi2Bb371aGZHvF3lKgBI
gmAQdHjPPFhgwneSr5kGfqWf6jsgbByiC3eiSvuwyCLUDfUofJ5r5p7XUZC7dXxz2WI8w0Mirheh
nRB9SoWcwiVzyDORR8deklEKjGye0gAGYJ+ro6mKfdzCVR/Vn5GO5X3huZ5zFHWrP8SxvLy8ATcr
G6BZvGrZ13RQhH6AXtrie8jC8iqjf0Lsaurd0lx+g+sn4OYVuMs1g9KF0H5jmUGeZTXZ/Peut9UJ
g5JYymjd53Czn8rpjtleLEEoNGepHjyzHhlbOY59EYsr4QCwALg/UKsTQ/qf7uJfEw64FW7TT/rU
2OdjcS/WDgotg8y3MJggdZ/u1OzsR7O/UBlZcWwv9O4e6QE0BUPb6g6tJ3lodKx7MKZ08ql9/TlZ
MjHhhx5VW7gzcfLkNl0MAaEHEorL9BnhbtFEOcQVVRtn9gYIToIln2oQLv9eHrTJtgNAPgU62aOD
+jDuI5wi/Ij5gupobqsTO1CQbiQPov8RyeQM0ebvwCorn3gNf7soMZVhOtfAe1a/5i0AZ1+HQIUh
rNNSYnx+Ec2YMMJCyzUXRc6A69926edLj3QR2hL8EVn62Vu19jV6b/8cRU6h6HUXcbY/gU4cmY20
0WaLPQWurG4jAuYi+YD6joBkaBZOnPAd3X0n6lh3DxPyasUfO+pGA4RgMdDkkU/BqsnZg0jwurw4
eCaFmiBSVSB/ow4KoFRI1IKOyDkAqrgRb8fD8yAv2tRh096rsBPxPjxUoZxYapM4brXwaOSzJ4Kv
XrYitoYVD1hfmgjxvssgNfv9WfK9ZSpgI34M3h2q1mUrwUXiRe0Fh9bcalQ6qowD03wVfGQ+YsaK
dqWTVBxVZXYgEim3/KCtzgodgSiPDPlHbiEA6mleRXDX2ZkJ+gcMWHg0+y+63FJOVLFm5EKFE4QW
ibdSmp5PU54Y3zqvU8/cDkHKjjCY96IxWH1MxQY8Wj5Zik8YNcSAud9zWQcz1sGuosbaaiP7GmPL
9PEogmmIuL2SS+MWsd/303XUXw9xDrddx3/wpzY5sJ/7o3JoJzqLofgk7uoCXgpM709LyKRmRXCA
icUHG/uDgqAhPz2jiypqpKGdG8H5MpxovOyFAuXnexLk1WSkwWMMMI6aE1Q5OwS79sY2FpHX4iWs
0z39O1gRBX+8Z0FHXhb243iQQLaGuPpyDwC+CI67FsWWb8orQsFEmcHWPbEYihlbEv9T0Tf9k5hL
Ws+ZWOfxKXQSLJ8eiWv/4aqjW0rGYurDnPzjgHYoij4qWMA5YcwEecRr83cIh2oecyeHq0b8sK7n
WuQeflvyYZOVUbKoMvZDQp47WmVRzY5Bu91FQ4U+WvKCIiG+Pp43ep+fhATDqzmFShG5doLs0BXJ
ntfNav0B+gDHO2xC0KJcyzYSlc9ZRxp1VRBJr+EeUam1dswaYGNezUncF3DfpIBZYfFxpVViyRw4
lKKHf1WQLt35qas1fuAx2NcMIAB1A3QbWasCx5hzOiF6hrG0EI2Tn6PJMlAR6W89WIhCvwHyKead
hy8ZVzw8jIwrZppsJDNaZEqGi0YDkS/MjJAvvaXqJLsI9I3WrY1xmTRjgeKLIhykIt72A3/aWjns
UOoKlNB4GI9Emw7/2y67DqqtBohuEgAsCkQ0PcbXNKUNuf36aqgl/dwIpsbvda2b5W06jzqY23Qy
4KMkNdp6k+p/3tlaab1ZtisBlBkMvJ+H6X8g02gR9XKXa650PPUPMuoXjcB3OxDJ/tImfgRuUx/I
D/bL2KUeD5s9NLcqEpld2lBv1N8DB1/SjJqsEl//rH1hyZ7ooLgzd1sgKSH/E9yOVXE3OROB1Slo
26Lo+lOhDZydTHbY6KbGGEl/eFWtV+ZrEjXLf5UZebRaHWRsXEi3qCA/+Um98fub7hzWC2BW98/e
cJbHMDheyoLRHOnQj2GlzokMKMB/WQhtw0RvNAgbPJAFT9Brex3RLc4Iozaqh3lCl9cdtHCZojEn
p+Xt86+cGCyciUKgOWx771YDZKno36G/s2dpfLw+hXVe3sBVZHl2PSFcoyhY6+hvK1s8pmO/7jYh
zHo2jX+Jw3hmySp931CdgMRbvftrP2d8lDe8mOl7hnc1WUMly1eyMthgiea1NMvNZLrNo2efcoS1
uY1B5gdAITWKZQS8SsSn+Tb7OBUs5m0Kfj77GJ6E+05H2qhp06LeYRSWPcKGjcDB4S+X3XU0NelF
CoSNC5cTLRRkjM4Q7Q66mtqosVWb6SuXedGw6btMSnM/XcP/Df9aLqhtnlSYerRywPrpNaQEI9Ai
vQwhm6F4zllFbR5xQaMB83Ry7UC1ogsiXb1+2aZNrsUa8VB+BfnAv8xg8BaUkDo0CWigngwOQcO6
dvVDhxjMAdoqPRmb4qGRjM/7OhTJbL0+V3FTdu3lyUsAs6RDJ16V6IBaRUBL4tI+3ZBRsxKouGBc
nrGqSiSBmMQDgRyWLRqHw7FASHvm3353BiAUAYsyZk9++MVIkSU/DQlR+j8jN2+jzea/aW/yeIar
1mdaubwfSnGF/B/niQmWLB8o/LY0QHbqgBpQtGD+j85gJdQQNXcONMdvF1N10Hm5XlBEWXe2CUXB
5C3GeFa1vninKV6BvLOTrdefdDQvR81uGVk3C0dQt7mYeoJprUYlWPfjmAFzg5OqFyxPj1aWs17f
Yb+k5GsjrSG4BHabHstNTazQP67D4xJSnRvxGf0IH5wXgstjy/8qW/Ha9n4IQgvU/dJPjkKhGb/o
72SgSXG6OfhIY0s3MvDLM253sj9JO/53h3WfoDuKjLBAeY4sztwhJ2WAIMQhaFwITRdXWyU8Zhi8
3+3BezW50CVU6t5oUWwkJeEO1k0ww9Jn/8LcWTQWkQMj5Egbe76pn4g7b01z18+oK9F1VtEtz3JO
KkStDkYDwmeu5RwrRdMR5HN2ZzmL7AWu7GjCadUI1XFzZ2eYSxGXg+y7RVfVsrljlRunWbMhKXgg
+EtyvxbPp8XkfuzJfu0ybrudgIEIEcLJrTYk7qn4BjdZJXcugGRS92ALe7wG9K6kZTtIQyyOM5w7
njw+XWVm0NzO+Ehe2FJHj6kZ+8QvH5sPKh/jnggufY3P95WnsS5o+luKSCUIiBdE2QGTal2RrK0+
1HPsjQjGQT1C44I5M95fAxdxacRkMucK+42f+NsccsyA0/t6q96QS7Sen4hy5/4sdBwl94HNoOB+
T0JnEq0wL5OkwhMbjgb/g9kfokX8bUE/UCy1KT7znxFcHpckC075mKhtBZqpJe84yZpD9H3bdc82
7LktEpP8luiNScNr/w/IN/Ani6qz3vrTPoeOYttyEb7dKajqRHZRqm7+zUBOjI0o3IuIcg+AvI37
Lm2CHLr/+OA9r5m3nqyDadOavnNoWG9R2tdI/kUA95WKr/iVN964vN6Q7z09aO6suxvrclj5kpXm
WBag4hYS7TnhiVyW57BksXv160FkFLnmFVcA+9faVdZxUNzaxrxnT5WWIdgzSC+isnP6tdH4P7vD
hSF6XNuoZTqw/qObl9ZwtHJKBZaLJ8rS2wjsHJMu8AzOp7UKGIdk6PiFhhDPRfIWhWu7RNhnfWJn
zi2Cz/fVfq3P7rV9ihO1nBcCtWYVreoYgnXEhs4BJ5ZYjWKqKLzOm7l3qSdvCaYQaCkR4lcg2N2/
kDkNDwnZXfTQaXSaOEEIBEmjMn21LmT8PHEC4Vjwld3+6Pn2vcj8zgpf/vTogFk/jXryURD3e52H
TrG352nnzgaBKSqdveP+cV8J2jhuGxGwM95jTSiqY36TQyJqWxPOv3iIb6O9HxSl1Z7/XILgXTwa
e2mU3odiqc1fIPc5TTkU1/3zjmYlTgyVnAdM1z0SMJJQv8Jmr5BnBffN3s1lfnLpniYz62XuLsMP
NXRc1qiFr5Awq+67H3c2sxhaWKDdXkCfF9lvcZVtAWufG07WypgqZiwxY/5CepxIcg/1RfYuSQxb
uFKJjxdPt7tkUnaUX/tC+pxwT8xe5GEPIJnK5Q0KB9AxYce/sB0pIGaRmbr8Bb8V76NpXL1tsPk3
YqZ5chMrogV6D4pHk/84FhXKQoZFUBZbSbBui9L2JdLMNMSpodxJcvIFE2/igSVmimVGrYJssUuh
Pp6IZ21Aw6DkCUhltfSUfJ7ox5h0rtYxe/hGzlgkqbwoIX5uQHlrqc9U+iOnJbVOLpoAWlp7yih2
8pjU51NDh4F5RgX7VDed1bOftfgo4a0fCIOG1YKluL+eB1tAQwB+L0v+UuQbjtQoPo2pEzfZgFqg
rfpXwBZgGfJ+IbYdNlHdf16n7421s07MsAVVuPENj0BA0Xax7a8yOcOPOHYswoXe4IWTudnyj8yJ
GTCyGYYGXDO0A4vHpH7sapozU8vVO+51jcnXqQ4RUMjd6y59nBGcS6qqCI3H359OMNRlaMC4bZOE
n3gGe/JLhckxBOElNmew71dPfUXJ5OxQ+7csydoiFqS3zKjT/iMizIeLPPdKRqIt/5xbzRwNhNVG
RXBHTLEyZ0iKri7iAyQg9HPLehlTnPrpl7qJFhGE+z7UFKeSRQkfz0/ZpIsIHIFzXpP7Gajool9i
WFWfEakHw/UTnCz0dAtT9EYJzd9FaxgDR1rSmybGdBjvQ/jKUKlydEPKRyVC+1B2nOZiGunh+ibo
FHadSpp5bjd0VZrdtqUbYQRlYl5v1InnzAWzHg3oK+Deai3mO49pknzkdbZNFv6wgYUuFP22HHjs
x/jrzQwg4p4o1qbwJnKcpLSo5/wg4xsz0KZ7F/AVSEFGdi2vu2tCn+VXcPAP7lUoe3DPBhFz5b9b
YUsg+LTNnF+SZr0SHKeT/1ftlYtZ3XC+XPW0fPiH7vCirD2/tVcRKlKJvhCuAcd/uJGA1ATNVY23
eR+7rCuHWWormITiU9MYXVP2EfpV0MhnrJvthsQsHWGnSubkIT2y691gsj0UpOB0vjPGlFjEx1DH
7ERRv4NSybvzVhWnmWyyNeHAyARRzpuI3MDEqfxGz9boSL8Blq/6bg/fQBXTn3WuSDVkC0K/Ziuu
ZjD7rFqQDgubszTN2Xe84mib3GgziAhM52nb3xR/qjbp3Ac8qrezFnCUkk6aFR80S8JbLw1U3tKV
yp1qe4l0AgBzpcJsPow7vc3hkF9S6CXM3caRtNwrru+BeAiHfze+6G2utUwArsUkVsrU+OcnyAby
pvNS1Tu/KGzbOkHc9hTgQm1lgdgF1IEznSk1zuQCzKr8oOQuGz6EzzG/usMMbTztNx59HbwO8BlS
eOXKYbSHEnXrcyvila9Bw93q36qQPp0vdzYbkc9AaEd2TP8SUbKbIH4CRI6cfkYerPNUnjURxFDl
zaTAR/EZcJ6/D8b6HdeJe02sL6GeuLl0eiFCbBDHskuw5U8L7KP35rKbwK0zjp/D/LIuf/tXvdig
TZ8vVaha2FH3uz+T8zAGexl6ePkhcut61P9uiXXUDfd62KpwEI7RaYg7YRrhO79R3vujnq6R6Pxy
z85sC3jmfRaBUVwD6zghfkN/Q45fhpr10TRTgXAdQsBRs17jfwg6ecINcQANtJSplRw+DhQNANoT
d3K9RRRxcCez+jZRZw6B78Iy/5By/9a56OHhQzxPKwyHKh3ifq37ktipDg+rM79BaE0nLD/uf2A6
mVK8H0kgxgHAeOjZuOnNtlLPd4K6EWRuEYrSKwQov42eo4t4Oi1ZYX3fKMM9xnuFPj4U//esIsKq
yZ16hTko9kCKoAOXsk0SUDo2SYhLuxkFpIdhThaXy5zjeldF8g+JKADuTeClmJpT/rbGfx3cRIgO
/XdAiLFdWS5+d+YWCwX8jXkF0/3mKmujickKswvUlfha3n1QC3nVJ1s0sd574oS2LJoVOmooTHEw
pGoi8Hb6w/NeP/E4RJ7qW3JG8+gOi7InuKjwRbyVz+QsA8qDRrUK+t2OfOOWmwQXe3AjsGUxq9bN
OSiA6SbB8yyWt1QPR1TtYLvTQZxFjtW98mv1ZSW8eiYM+noozHBTcDX2OMVo1hpGMMPuoQ/elZ5H
r+J8kbncntG5O//kw9erdGGsbmX9RwNnPMj9EiWjKjcFAc8kwaj9wRyk0RBOKLIS6rVbf8KMPTaP
8aAZvpSLof650eHtcDmQC8r0rGs1aNa1+pn1VrclkcOh0dAA6u2Z2gJQ6uJMXq2J3h9t77J40rAe
4G1GFlsMPtTSJ34lpogm/VNm4pJNOQsGqyQ07TZom8nDSET+qsV6Vn9uZQ1NgwYYQKOU1IirXIJC
86V9fF+C+Mt+wtHKixq1lNI+HWPNAvQeR3OkLMIbCAnZNQvP6r2ISop7ea601nHNWcIxd+CRrP3+
93PML/YnOH0zh0vkFgVMN6OJ+2VxgACA5Fd9ZDebfBuKr9W+SFu3sl9+UIt8Nq2t5x0viALtvAE+
h6rXXtwoHr/j+nNPy5IOnA2VVk6pV9kyefQoiI+Z2oV/u8sPH8g6aNpxZB9ms4lntFW0iliNuzPW
r+HgsrI2uPNbwBGUC1NrgD8zsoXfA0Jmsfg5mSx5oFHCIv4C/kuJURRl0XEiuOzZDzV8Pb56ekb8
ifbUMGiByT7cGGx9o2eqyXlrc5S5hVOjCkd+jNciBKxG0Li8OgycSMj1QC6UqCpqYBEejOLTWbEi
EgNx0cHQNG0IyT45LgIFK5QRaZsmKdhUjhjpqfH/vbKr00F0fsiXxc8YYyFCBoT9uKvpAmU5mE6f
iLG52XdNxJ6Oq/wgVGPNYkw0wMV8ZWmR0cW2knSLC+LRVHB7xCUyz5OITNGy+C15jyEqNm/f/SIF
1zY3+kVT1ldFVkQJIV9z080m/+8+2xDJk1ArdEiA8oaiyf3VVAQAJlWPWKeOzgxzZDhRDBxcLC5z
vH0vaqJzGFIgQkjGPpHnfh7XAIWBOFbr+sbVAmELPRPvO9MhVtdGQAPw0YmndaoiA6MMcn5edSyf
VGnewaSSswGSpi7rtbXTdMi4IV5aK+wUOvGBzo/JkhiASuaswu6FV6N/yBUMfROrGqtCvXMmvfzM
WqsjXl1EP03IuyeDjv7H4IgRB0YcZUBXReCnOToUp7tHTDaYzjYOtOYolbQuGntbocWSwk3UcMdh
dhzjQQrsSfIv52vinrztpus3JmNVj3Qd5dTYyrzNzBpnysenP8Y9m92vrnRAGxKJ+Nj1fWkePI8p
BR3BkVNL0Q2lRYUGIVCR5rpYRXWpcj1yqvn2nwcHTScz/vuCIUv3asK1qZcMzN5271FdiaI9lSGC
G2nBSrar9Au2oGs4Wo1avsDPLtkctslcgfPmbQSs6IAE1ZBdmU1MOp02Q1KbDkaWPOVhZjFKS4x6
0DBnZ4mTSHHr8NIbhT3yowLhJxV+ZSiqp39uq0KpgmGnYCkEfYUmlBooiARSokZ3HQmfV6ZnRCzg
yhXscZrPivHGhYPr4HmQJAxQ8nZ8Ow0kCc8wEGQMYNzyuH2RjxwnDn5yHpOtGqUIn9a+sNtf7UD4
DNEFwUs128FJK2cibJ0NpE8PIrmsG8WJGvSTh5G5+50aiql+zpRwMPJ+K0kuqw+34g1NcvpLpay+
DqzPItRkEaRgRNLnoeSqM5u8qDVYQwhibNnNZ4mXXXxhHfaskMV8/ddhQT84z27NXEmlKjs/mMRi
97ArO7XhNFU2JRfJmJHbuByNR4JXsCNldIpfd6qkrceGILfCQF8+xKKxGYuBzG+gyJp3UTRLynaQ
96Mey5qlH7t5lq5dtT8vItce61jUvzGulZU+oyBC+XqsPAjuvLmWxoyn+boCVDgFipGwAg9kx/hp
8DWNKAuDsvYIDx1hztwqxGc1r2dRyD17yn3pYVZKRU4DJWodUkF1fKByYiOKe7ymFCHS4gEdIVpM
xoggEZCR+zAUqFtbLP3nqpLcaRLRTgwDLFw3xnRH/ozb80i+y0E5s9MEMI7/bL/5cj6HBTFsmIBA
nVc1gOMZydxTHdzZJmxRy/oh48cFEcY7jd/IsxDbEH6R16crt4uPcGWsbF8friK4UaMotGUUAQGn
dXkTE/fXKCbruIgqCVedcY4Qk2J/Eg/gFljWsq0RaewVreJs42rSHkczjpYv4dbWZsoDwcDHJ8ME
Y70L0Yy2qSAZ6aG+le7E79kzqKwQofsDHkXPm9H26wI/1I2vXyXrrNHCS64jMRqS2jB+2eXZgAuv
xXhAzOverz7o7uneI7RTS7Hm1PYoheasKKO6uSiUbQGto9teEB+Sf3djiKZ0zdOP8LhlATv1V04Q
oakWlrn5Oscx/UaDXYl7QPbzm+9sDLgYls00KFpMWuxEk+Ovam4kq7AGxwYRUTMHiUZ5SLPTxsEM
PtPuRnCYiCwlCq03JXkxGtRq3NdM2YGoyXh5kodv2nhXWfPTILkgDA8qzeAyW7z2zZg4ipQ/7xFF
PdF8226lptF7Mw0UY0D5Gk7ncXGhxL4Nrle/jVH1zyVJl6Nnim6jWRbMTIuaoxATnrAR1U8RpsVx
E9q0qovMHr1n3pl2Gd7WbuKNX+k13kjZ/SSRobKO+ZBjLk8Tq5q95lNPbqgIgQ9wOqUKkwhWCNFU
rSRfcLm9EQi1qoMGyL3aA+Cv0FTVq18w8s7bkEMeWBQV4buLvETGRMQM7a2nPWrVxLVpYzmrJaJU
tTCiJ4qo63/r6PAF868htVSjvVkJXMM7FXELZPKpRH286qrsKXjpOsiwD3bkG+QkSiNaERi8Suby
4YcnpC8A6URV3J64NS8/CfWsM7i/54ASujsOZxJviShWA1qJ0l9/ezQFBOc/BcezzETJY+/Fv+Ym
rG6iVMY/WDq4xK6S0TiMxPKm3QqwBfzfmaLojI7/XKauUGWku5+o8uxs9vDnEYXMgleVVmO5Md6O
+uPdA7DOKTNeLqgPqdMII+F/oPBqjj4EnMVJXriBnEbtUw3/GB5bmvokCrfSbgIFxznO6hRmAeC9
6wdPtL904VZ06YFfjZORfoTdO6cXsuAnhBzunQ9TjsElFIH5xp+EkXDfGqv824OrIscfnnn66tjO
pfV2ihHXVY3UUrJ7ljjJQKARfSWTjYOdU2sGwWLKWkzHGMmyfm5Wl7X/P1ICBf8BKs9X2JKuZaRE
fmQdmrsWnJWZqJo618Pbw06Ci6lalzIdMcLAo17flbKB69YswG4PRcn4Qnz7uke3Hkhh0F/cEQcF
kZblQR5PJThukNNpPvU0CnU2YnEDQMeYR5inRnKDfQytLNEHbBQyWyVxt43QJ2lfuHQq5apEzFjD
5aPdI8vQM9gC3/ZwOv0AMoJqhh5vyAPNYJ2e1zAq1A88/uCdyr1vVvNo1Na0+3MCWnuyMxQPLgBj
FYtQ3QPlUAzPjQGHdOgwbQREE0h9/0KQ9D1JeJyL63F2loC25psiHAhyfn1XN4WziEEzoK89xBsi
HOTOW8Rzx2TK4BgIHibofab2awjoO992ibY9dbQvq+1RXDEuUrBkt0eyLwOdgMznj3ant0dEAZf+
tyJKIJSaYsJ7pn3q4cqKp3XwqTt/aLlSTrqPsRbZLNCZDpNwRm51++6Rkl9/t7BhM4JIN+i6MA4e
VK/uC7U9Fd6DZB2BjpftF4kAsNiOrXuRTebsLilfgd8VUOx34k1AayAEOfCS3broUZcrrqUFMlSA
v+Y8+3AriSlZqkQlKBK6Ku6F7ALNAXGCP1I0zHtnl+BAEb+cLXIE9JpC5+FWp1GIiOCv4fkmfKe5
QhU0jTXD9luNTrL6bYDn51yce9mn6F8VhurBdAIv8ARqNUnbKjm+TGdqy9IkJCKsS4zCrW9L3Qni
EwI4iovHqgWPFUkDKnFn7n24fxXmFFdzovMMiVEa6vbvabCpK1gZI1mIicTqY6Bet+XVlsuu4TU+
7MYmYoZbKVrZTJRy8kzbg0EVX3j4+dnh6tRwqVQBiFsAjit5dOxInfBGNBzfG7izRQtCsv0t0UnS
kewZjP7QM9LocvDZ37t7YkfV1mX3AkiZ4W8WEEbMl4O6bRWDnFBau8/wm62iWiVld107mU765pDZ
Li94SfWgYjVGVu+g5T1Z96w/P0j4CTB1LAvCNirr5Bq9Rv1gJ4GFozlqPbABs0kAk2Q4J31ZzrWs
sV59lTZQJYawqeYcow48J2jNDm+PcxALa4KMvrtmfHh41EafqaP2dWp4+oOuM+V9oEw0I90b0eQh
sBpCyNJXJ+o82266pgGDk45UsZ0vKUBgyUo703+EM8zHeMXaNx1q14FixY6aABHwQ5JO1rvH2aLV
+BQEsHfG7UfdPD2zo/b7x0SX1qjzDi+zsv9J/nTEXv9V2f21ZPPEUVdlj+yg98ODhUXzMVskW+Dn
/2e27WnZGkxV2qhuNogGcLgKg8ga5p1VEHY8tQTBe5j0FS9ue46DUI2o0JI3SQcXM5ZF/T/LxBQ7
Jwy4j9hzCl6PPotmtSyr8K5qpVMLuiPGVdzo4RhJOWFj/8Cn30b5Hqemj1MhhVWuO7xXoDoixxpV
02Bns8eu/9mnFtcVFP/JUBTer/srrmBjXxd6WPMUk/0lrgMgZetx5lMOwXHbckWhqfA0rCfJTLSK
+/FC1Mn6dTwFnX4QduLKLaFjN+OGFIH7ZnRtJ2B6SpQwK4Sam6P5fQ2kfx3yX6ooGJRynwo0sUYq
GMdeFymtEUCRpSRfZw4xplebJJmc2FNRZ0f1vdhj1EZwdwHlQxLRV0XR8pbbzAJlv7Z0IzmYRRzt
J9inhctaQfXoVqxVDmi8kBvEodzulriCVZEY2d6lkqlZgJZO9WgcgrTlwRq4EQ8w0LjmYl+LRv5+
ZNK0icFT4UPaZpVSA+DV33RYeNZR3LuMovOiyMCQTThvfybVle+tOhQGE+ygxz2HdJvVgpMtDT5P
qFjaitYYzm0xleIPKkCJCWOX6FIbFncr/oEnZbJCXg6CucU7p1+PkFzsJNefg8ld4SJcuDjHBgtb
2sWabHWAiiSUDbQAafUlFQj6soCW6hTAXGDDT6kMXHui+4x2POY09g+ELc5jED5+Fj860cS/j9kd
AFGtNW2LTzwiLnelDgDcPxQOnaUd8VqjWbAeQHDMt76upDAS3SGIL+baFfoEtoR/xYgCUG4uZuIt
+3x8ItbOQyQUO9qQp6cjM4Zf7zUUxrKFPftLxer/L4ga5j7XG7cwpIn5uEOHRhRPoQZCqEackXiR
5nRNE6Uf4qpsZVhCwb6yfw478/xYr6qTbp+CVf6roRjbNmqRQBnHysgcuSno3rjD+UqHvvtJS3DE
3TGw3IRHjLOSB51QBwivzoAaKCJZ5ySuDKVJSczUpu+xlCxhVyZVvmrOm/elqxSGsX76Bs1M3TlT
f5kfziVB6zfaNK0xbIv61u5z081y4a39bg2hA7R2JAXs9XYrY8P4L7+bnNhTxwvG4ym7AgBr9ygL
p4byM88stWFN+B6JNKQg47CGxQNkdH6ch1yQySAeeHEkS47FYgS8Hy4dG36eQWmXEJO6HkH5pMTZ
2oa4nOsdIJtTicjzATLiZcB/v+tqaCI/KL98HmLz9lH6RqaPQsY2x62ZAKFi90+xlWSeIOLe0YGg
8liJsLJ+fPtexzdoscG7soe4+pH7EjhAl3N4q4ePAMfhFVDg6dc0icVipw8pZYIoQuKXypdlRR0K
2jmb0sQbabt95uxHK6rcV/Kbm7eWpwDE/ZZB12dV8GqoH21oI1agf609uJ8aTdYcyAZPo+6S8lWy
RiAuJqZUS6DD1CcEsFeWleFrRn4NMc8/AvGYbBC3OCS1/NxVAIFFTlN7uA48JiuZ+aSi9fnwN+sQ
aDseP6CC51n2DMB/vCdGFPAHB4TG+1rkRghlXTF1P8UtljIQfdzb1qPzZTDRBAAQCQ8ca30NfRLq
HU4jSdPpthzuxb+pSXvjX8C0gg/8/HzT4DCE9DFCIzZIsFOWj8/kzCgwgESMm1BUoVBGeJJsm96O
WisOghG+EtSzNRl3x5mhUzo/gzcjqOrsfe/muHyeia9h3DSg+KSTBQcUFzMvbjfJbgvBmc7nhDr5
vo68aUluXBEUABrPkgd6qw8kz1f/f2w8UgN9913+xxoyGARB3dhRNfKVrog5RrTzuwD4wxntJm4r
fWVu7zTk2p9WY22BK2qAxIaUzJitfT1G4ZVLKFuZ3W9THXML4uPUuoCZXFa90mutPqU0bAU9OONs
G85VNSmL7n9aL7cq0vHhkwXEhTrOP+L7LiXSLDxFze3ZYT5HFy/BeGZf/sgVccjXrUn+Zy5DE68t
d/pf0aKrXkJYE8A1a7sRwYVfED3VTbHn+kRlICsUUwlTgG1SOJnk3Ybe+Hlgqv7w6LPwG+B7yLTj
Br4YX50gRkLGuGQ15IRpv13V2Tyqb5DbOSIB+DAtlJDV51ux1fFxv2dBHs4Dg9uY8EfpPpQVDu16
Xe/xVhduBGsm/mnbgwwxugWiRqBLc3JFAVZQRvj23/8EqNHTH5lXaz4uI+MxtB1BlLAZtoe5Ug5o
bDLvo/ABo0q7FRBbnx8qY3se3hSjbMuhrsnkyAyFkLIz2a2iKLzlLSya2GI2kfp58UzGiQtXgjWH
Xv7CgXA7bDRVRpjDsXxYLPCt4WGdEoXvP8VvZBgyMGFio+h8a010h0vToC+pySTA707oiiyjF6/v
O+VxssrhMpu3iTbMHK72QH7EUd6P7MrOLFJsHv8irPnS/7HcQp90duE/1/3Dv/mBW/I9B3ikzKFY
vjew7itFu7xkfwBLcrGNbux7sSCvm7sksstRE9KmHPzkpO+vMqVhERxfGTOllsvGsOqfcTyg69pk
tUGzNjGZYyOxC7SsbLU4sgXzMnUzN/pXa08sZXRjd4z6DZ3cX+PkGWAF40QUTc2o6H7OglvANT2u
mjjX0rG0zcc3+YdHyXA1lQNcyup1E07BssZjcgLIQOB1tdUcgZ0GVQytpEN7bhG/lstZqJxmf8VV
xueM79INwvM2kite425G7/7lyk3TYDuDMV/3YOzN9MfhpVMOj32pTxJ5l1B/QsehGOWiT6mNjDxc
b+2ISOK0jknRh8kauCXDw5vPyyov3xUfQZsVcIIN4kQq70eiRgYzmVfhA+xWP5g3b6orGWnrfiev
4X5CdKTqz4s5qLZOfCGD5FQaatmlSSU60lpwR2f9bbcRpnwBlhdTyfzexkcTs1py7e39M8pb4yz8
IPnbwM9GFUxW0S2QgKkiKEWnL1ChS8eY9LEraignFBSNgCVSUJMMdL0/M4p/EQuNSxsvhN91jfMh
adSTP7IiGAtMOqAA49gBBqDnMlJepH5rewA945XCyksy1k+8nNLHKMzQdyDLLGo5cQOuPrI1hSy6
UPEJuhkhWG5J0wCxIDHxJw597vW4SplH79sOy70g1wnTIwE1XHJ8TJS1ukev6oCS4VWcmzL1bzcn
smO/VBdvaX+tfMQ+bOtOj9heXgm+DNzCtKb136MpjgcKXx0/4ExB3FhT1v+a9gJ9dYI00n8cWmog
H19vcKPpJ5+iCnjkUtAaWe5ehl7L1VE00j4LlyUCj+HpQnFrCYbtaha02rCR0TZEhTe9pWxrq9Lp
Z7LRiOZwbne6I0C3nsRp9gUqFoRJJ5jeHspIRlRT4kobOpB8UYZclvVMKO/WcRyxg7ArzIOuyLiX
/L7W9iA4iBwXIchuumSV40l+em1oibfxky1/Pxc2EkW89etlmB+MeYYvOfkrsNt/YTlRUblIYXRM
0TdS67UM0x+dtBkBa7r4MxcxVrZCYRvMzOgz0MCPBZ6jxjv4Gea3Nbf9xhjByxxgplkSzcXuiWpw
vREcigXZWFK9i6DaK3yvbXcTuTvO9k+l1i17a4FoiRQ1gLpIcZtqqXhyP7kBVuIf1Y6H6Ikximu+
w/UCvKToJuy/E9/cVGSEBOkFe7reYh5TXZcFsQLhUDsil3+nlPtVD1VgsaKqeKt54SA9cmGg2hBM
cJKzvcRxZE2GRrV8imIh4PUa5sIOuQM6JNVLLNdNZi6SU7l5npZeceufejAPfnqoAiVLsRhbvVXL
APrZvNmQlwFbn49gNCXqgZwF8J9SOKsSt3eaB7ODxhDGJZ6Ng8grNcs4GJiwXVQjbgOfxBLDYHnO
t+XIHf22PbB6+uYgWB/tQyKoFxa+zhqxBrq9Oswyx2bNeOBpjMz+WJ4Bd31heu1WBdat0smH6khl
rD0O5Z3lFUz4Zwlp4mwyIQTOiTPBxRbB8s0pCUAnhIDJdoIjWRU63SPtUkvj1YwLamDWJW2qSf9x
qFPehnK5cTjSF4Dw89mhPum4vyHjXhO+SWirTKzqScg+8WiAKCYMUILzF3bIOZbnFmbMh8QlKWBy
Je1oueSyIyhPh09wtY7hpeXx4xn7yphfD45sM2CBAK2ugB1nt/inkSat4Atb1/smpwf7Eox5a/aR
HSbYjLX8mVU0sqgJGRaisvOHb1NUAP6vN7sm8bHMmXapeaSdc0FKH88r/ohE5Jph0l6WQRwROTcY
tADnByBDFCwJtPW/C45hTkWMWshpiMDuDlSi0+5616i8VGJBu4uqpaYIH+Hcez6I8oOvbzIm/dEf
ADYv3YFlTvDkrV2ImFWwpRUpkFiPTNUFQoXuVGknQEOpgpMSa5nrfEbkFkswMQPUOwxa7GVuSXsF
CIgBiSTOdpjrj9Op50sFrE8Sywu8ofRLuOQWBxMImR5OG/B8sseWWkX6ZIdUUT0yl5AidPP+5Lu+
B+zH4gu5c3TSFMSD3LUHOaEC0tc6mtkSlmJlAjh61hcK3659b1I+wasmx3BxzseVOECW09xdyiPC
ggVVpHaeqtR0X9x+OF9NpPZIPgg8a0kXa79EzkOVC2aJONsFxGZxRfXkBFjgOSkIRetYZjjHXGXc
paEZvDhIn1LIph/CnjOhgLW5Qv/orr0y+hFjT8P0eO+EWKBIMoCB2N1Ng+5QBgMrcvNsWXDx42Vq
V7nuPesCEUxTozwMV1bkFwk38+Dw4PFNHZYS+2ikMrcKUnkqIZ2Aeos7PIQ1XrZ2Ga8XhV86KYdQ
p7A9fJOcl3KTPD+p72SFHL39IzAGZu/81N1t9BWqlN+RSb7PkVTjw2j28Ik8zZ5ARJOg1yYO3JNI
9eOh1F1L7qqkX2jxb35rjbAcGMnMG7451RprpT1oOi9wkF1al4/8QvV75VzjzaDs+gJznBdEYXVn
mol4mDcnBiPfrWtCyAg/qsOt6dTF4beEWa9NwHVZLjagODvEPcfQBOvLPsQG3s0YE0py5haMaFDn
4p9XnzomlyEKaCvtuXpDPP/jky1pZut2Oiyhpzsen2KsPsCpxo6W8GVaKxaAHXGwPQxlUhxD/8RH
Pa5nNI9qX/o+cbIcgT3NrPj2XqXMVzP+gEYfb67kOdfLzq3t1JoFs+i2d3IiHBRfb/stT4PyOvEn
dIRkkjFwI/BFhRho929zxL+F+NFZzmp/MXQOsgoycZPuGiDTOQNhC3aPPaxLjkOFDN3AwbQ2lkgK
OoxS0lPfLMohLXS8G6x1AsNXwsq4hY5N051DoRDm+ZYr91kOGXbC/MUajTyyLxWobNN0LIDVxH3s
EP7xbF7gUu6n2YhUDlO8jFX2a1avl5F0g/dhtL+u9FJ6EXKUYG1QTsunq7kGBJDioD5X65a8bAI+
yj/Zir/+CJBCRiUoq3q1Y6JplNdrKkv3YUMFeoAv15liXDT/4exeQBwe7+00rG19QDMBQURlsPq+
/gXWtDg8ewenpUwxjlh/WgmX465UioT1mBqgxDkDtoakuQBVukoYNvXJGthAaeTEzZcoVPhL7oiF
dqI1bjCARR392isAgj+H4W7dBNolA4JQK2E+j/TnjKB8Kj/8au+pDttVZSjYjkKoi3Z/NnYO5A3g
AbnTrhZr8s+wglh7I9mf2BkNkGEJ5GLFQloWZ2Na+2wQUThdtwfLiHJOwmR6WRe9FKhqE6eWc5CI
DZRbrykcl+HqGXGU1KCXMsvCRYpc0JlcqVllvdo4tHfpKp6hFQ/AAPS/6K6mg51Eas1oDZmj/4am
ksalDOUNAMA8bJR+43T3/3JtSN5BIlnW/ROSntUqwD2xaTgGbYvbM7GKOlEfJgEKZlHLIGQlUd/5
b7ugTjFllXkJl3cboqIFcTjPv3xmqXLu5espzcAhl3gqCtuiucflfxJxKUmYTVPwL+7S8/mMZbDC
hfJeNvC+JfKlv7v0vpaWAgUyhV2rpLgFOrsilV+Ir/o8LR6urE1KkcV2fRrY7X/OlivtsLqjDqRj
H+tFPrGJg2wO5qJl0GpNXIF6tVxe+dXvHDlKF94ZGfB8aMUEl90NrA0SAap7/arUGDwAs1yxXC1l
uStEMy5tu7KC3i5hiQramXKRB0e8Q0cn1HhDwpPr6rjIBcGTCoQB39rGQDGU2QZlTk/C4WVJqF4W
kd4aNdNNJ123lSFfvL793T/5SZiT9ZZ7LxpcQ+Ilqy/g8D6EoCviouRdxxUlEHJ60o+8nKZAdxBn
3MlFsPzLbHZ/B1wGp5v196tuhR2JiP3p+27/ckZftTQI1pmKpctiMd6xJSpW3HqG3q0lDJFmSKRQ
/0ev5ETSugxhIoG9Itf51pAln/PUYE2TOIbZxgLtUjSfjMZIS/Ycl5jE9o+1j+y1GqMHta03Bdws
G8s4glfei8BJQa+FrJLfIdIpSAzQe8XBSTlIhM7fuWFsA4bx7EGKVG6Tvu6DO+Pu2QaDF7ejCHET
ju6MoSSCJHqPOHa42iQg2+NgCLqxFmWSbWZNOVHypibSs+FbCS16vOoWUYmGrlmrLMP2na0FZKxR
fxnI+mr8l0oCsKeZBTRRqlHoAO3B5oBS57msoVorOmJoFP5Chd/GCoYQyH+UMabNzOwr8C8zvNWl
fMhSIGTEmfn7zbO+Oy62WNxrT9EYL2n1mbV02atopwvLBy0wKhF08sAy1u9s2jFY/g2u9dgj2SzK
K1Chg4IV0Bp9nXaAnSv+PfEMB7S1vclSzrEdOIM4IGGlxbBmRUgJBUxNBGlVhzs8bHEfDKPreneY
1GPOuWdPJCFjpMGQCXUN/SOFGoZSEz3ERRvh9S8+fv9yAR8w//tfnMRKbFeu///ZyIqDztjSQwHA
8R1xrll1V5VzugsRRMADLTXCC8DLI+E6y5uadRiRbKa+Ox/6J5s0ktCYe7wMNW5xs+5owN028GuO
3YWTtDJgcGi+55OxAgPVrmphCH0QjWoNhfpWO66TboI6NAUWbCgtofbE0/ZS7fTEQCg7+mbsJctI
cfTh8ckZNhsPO4m53zsR7CNMLARCG25+VawznhehFjhRJYGa6tyJMU1zhYZdpF72OJhZ6snyQ3dm
RwwAxecV6V1IT+fpEUWasCiYb2P037CghmnO+cL1TAgk5cQwr1VcJmFWLyqkHW9IvGnTtpz3kroS
+3zisQGf3QFjfz+6iNLkaPmDxCwfovs+XprcoWMvNAlgMx4xBVcwyPGwueY0aVfq10boaDeLtKX/
M99WoBAjdirO6AeGxmoXCASL5sNSu1Zv7Wkbv5YltesvtY9MosuZ0xflVLtuoA1YBJlJ9r+t7Q4T
qDxhS3VtrlJsCx4uCiy6pQnrrZ/ZMFX7Z39B5UiYj146NqsUUQyT7U7crKCAgBT2IVxoYV2P3zz6
fEJL+j59y399aKmiCrwXwQS23oTOTmg7RY/CecOHBt97oVvG8oWOnr8b+647NJQAspK8r2qLoFJm
nTSE9o2nRgUMfXmSP3tJNgJ0Gj4B6OLM6+HYTnMFOk0oehW3jYIpfWH4UuHXQXiJ7FZoI2fN6txp
JFX7MdOMpCozsVUtsJiMU/eT0pM+3CJjhup5CFbCXuaemxVptn3d7QRw+Jnzf/bdSRl7dPR/rJsg
BmNE0rMVOSeqyOqUyV4bJ429g8pW6Cs/xnDkpCqTgBYRZXxZOyQvoqLhhS8W2F8hfx+X9GQka2Ec
b268Zd7riCyG2OPG9ePMEimTHvjGM5WTPTTQSKXYxiGcwLEJSDFyjmPQckFKAZ1lOzzQi9DBSm2i
ohQTsCuOLw7NNGamSFXl/zSz1HRFSeh2zgfH3rLsfSPMLG6nmabRMFcdzW93Z20NWNzON+ganUf3
qEp+nsCr2TTviwiF7kq8g4oa2TZ2hGeOTmd4ifPt6UScIwcpHfB57uK61nPQtGqzLzdyY+JX9zQe
Tr7bZIeM1tJjr6EYX/kMftqQHhEph+uc9zSViGEJZOnfEkf1cpIxen83J1FiVnzA3eFqSF9JUawz
QDBp7MT7iIrEbYAzd6vKtibeH+HWICOKLwkRBBJS4GNfS0P09ox9kEU9KKbzkszwffgPgNDk294O
jKRncw6P/XwB9Hh5Zs4L6YkDk1hAAqmNoik9dIERFtg+umaPbdE1RnFleyTSqnkh8zhmAbPfXKkE
5BRmCghNv/qZEF6rh94oOibCjWjYFl8lATI41u9KUFNW6pmseEX1oUdnwN07prF6/nwA2otkFerB
oRE5/H22U/48OyLTFNYGr+JNdDD2QaS2r4hPPbFrPrbk/NJfMAqZPNQtbQLjBnk4KhP4QTyPEHRz
ejq+FeTwc1Y0Y132j3sIQ36pM50zSSWG9zJni882rYbTJY13imysZWptilPt9LEOuQcE8Ikr3tPe
kKkpgrXpUGOPeavp3mieypfUWe0R3/4U1IWWBkclqE1XgsmSesnZYEcIHpqgTI1WFCGTSXVFHgI1
FoG/PzeivSDvqJZ+g8pdjeCRW0MFDGXJPFHoLESScB/munwcur3KwTqDEMqVuNsqWXGbKvUwGfqW
NTHb+ujYVl/fR6hsjl5vJ4EDMiCbZJVmwWTf8Cwsc1fKaDMw6l4xrCxTebn8Z51nw4yCkbat6d/v
ZlK3tuw9hSE13ucoc6ViLMOPIv3bNsCyl4UpddIqK1F5xrZpgnIJm7oVoftCmm7KPOG2tpDUEG/o
UdR29WJZzTELgXU7goY9y5iPthbl4eyNmx1lToFw/Ha4p3XGuDWd+206HXyENfW9FHAb/z41aIPU
Uw8EcZXgAqUkwhjQrEBGKIf5FQHllnXfSc+uyF8ghlddtosHheQcJ3YlykRL14DvOm1TA1V6YQC3
tO6RhEJCu8no30vl1ZX4tLMkLTdkaU1Hv4gTjvZ6LRoZee0V951RL4oAPvQrhmpj9+sTFpeMmMba
7v29GYqPN2ahZxDKCRybsiYPNSSpxgyWSeU12vsvTzqAvGRKaSNjvzYJ7Wk3D4+TNuGKwn/p4mzc
YfYFnv+FZN9Btejivj/axa97pZBzjLytqRvkDzGxGh3sa5UCo/Ox39sZ1s/qNmtbD4aje62UISim
EmBM0KW/xRfrf8NSOSNV2720XhtVnrr3fRS0/ochvGrcwaUEpAx6hrXa7L+gg5GZ6e6LPUoMvKq6
AFajFA4fYrI1OqX+Q9op5LYTz3FX7FnxYyl9EKocq/SOmWOYZDKw4ANQEBSS4k5aKe/Sz0K4uIX4
ew7yy+MID7WsBXUN7dcHKNZ8Q9XrIZwSpo2oobFm5/tRMIernFyO5Z8dSS6fXKGYOpH1t4+qLO5s
8EIy6fB3F2qmbboXQhGl+rx3ypgUFXphkV+8wPEhuAYlpTWNhlXEaU0BQHh0Htmd+w7nZqxIqe1Y
lAnOh5pcbA47jzcaB+HfoehjZUL7+dnlHmmGyoLh2TuAlBFrx/Ii0AtEk092jh4AVIpJWbCoMKib
V0Qb95+F3VsTUgHd7+fKHoQSdkezrlfJH4Ze03ju36QenlZcuzJh/aC/1leN3BGykT6ZkE+12Rc9
aE2zqkYMwQOMCCeuiZSl9q+/j2azIXvn9zWfLLz6QhhBkay5TlAxFivz2Okaqq560+Loyj8bzGTS
9VM+whkvoDMwLX0/WD7+ot8p2U3wGg7j3Xiab6LPw/d2yVsn0SCB+SfJJ2YLBgNcGvnpBZzBWEIk
BAgxFiBlrbtATePW5fYB5ms5Y5R6mZOj7oXDEOX76SvInpOvnTFE/NLc5rV5X7oEXnE9ucMhlMdW
ndTzk0Gd244EM5n+RkcbvslRtGJETFL8FlPosq2wcckF1nBQufwDGGDM3kyL2KPLqx28W75EQYcz
vrswvXTt8OmhVFwmgJ7jt8X4jt0A2EA7Fs01pwP0dxc0R5ckGxrJsH1eDBKFR7aR+kLTNcJopSda
kxML1wlKEPK2GoS7ZqboNh6spHZAScPi1JY8g5xT7owj6c0F6cd0kuLSyR09hU6SQApddYT3sB3L
eezchwR8O8MXZ3bfTKd3u7df5sDXnm8aaFjxHHmtDrXFbr0cGDcfAXmQBtyIhoBRZHUNMt4mHDc9
Cm4N4siGS6kVU2ReESi1LMZEpLY9vHk2y8swaF9k3AOZZUn9h1XdEWFxooS1bg3u8fCCC2DYy2MY
QFF9YQyYUw54nYfIrUpEsin+XBw7hinnxTvQzmUWEiejWaXLCF61fGxJ3RJ5y1rzJndHSqcoGEBK
PYyKtVD2Xql153qDnI5dK9odZ8sivyJQBriGuNZyTxxVICChkazy4rgCmQGWWK018J2bdgrmtg22
n2wvXZllRsVr00sS58f3iyN5pfMwG+u6jRoGTEu30X1GN6wC0CM6RMMJVqen6gLNhrRP0DQlX/iK
YQQDeUDh14hw/8uBrSPqV8SqJ5ckmfDzYUEZD8iaFKS9pcRwCWVwJGhGkMOoJzJf0VFu/sYOn6z5
NIWuM6j3ndZD4qnFgvRQNQgp1+XtfeVc3+cN6j2Z+DmSV3J388UKAxUyJbhb6cLxnf3cS3X0xHjr
jDYzLw7YEI+crP+jFHly414C1bhY54P37/bpIVJBXLmS+lnQxGK3e0QYYeIZL152atPm4VaSPTKm
j/spq34XsMwROSn9rK63e6K88OgkVwITwoQY0e/ngGdDrMhzsjoK1DVUOQi584pOPwRqY/8mkBoK
Fm6ttZvalNz6hhsuNxb46Q59RcS0P0daps3YTTjb1UhD5j9bnShFJ2JFH/xOWXQwrh0NVDY8nd4J
x248oHotybvKnXzDNOkNLDcld5/2CwQNUWrYGD073XtLfbSBMytJhOR/kj6HYQfW3S8VG2/+eDtY
moXu2x9z60MZ2AV0dhoGvz7kFRp5pEw3liSt+WzLcGiiH2oeCo8V66Kgk2XyiDUkcMifTixeBTv2
hF1qSyeOV/cCrDYFakPTZc+bre+LPAgk2ECKD8vbM1SG42o0m0pLyTzLe+fiDBZJeU3IaQQfbrgk
N+WNRXR8ef4wrZaUPWk0FK/w/nnfNKs8gvdRuDjuL9AGRa3JEC3MtSqdBzmqPL3qtqxq+7FQVazc
VEXfXUJpymMmyVkT8bi0X2xMU42qeZYLmJbUF8dKPAdoC8/BIjsUQLVZDvYf92iUw0HF5vX9Dv2U
IUX3g+xGlNdAPJ8/hDBWmqLMdkAq2m2+aHpzBJGNUYriHoZIB14pyMUslJUMFP7dgoRF484i73Wm
boBs08ZDUBpxE37rsXG9rZCA9o4hyVWjPXt7E0kOzoK4dPiC4in8HtMes8oiv0TtuwiMeOLQGrI3
HMRG8Z8tFdxvE88iBhorXrKsXxUYZg+BWEAGiMEdbuPjoONAwEad27BPcI3pvkNxxicPst4Zcm+2
+vB2jHEGbkH8l/+U2RPIyEBuS9RYEMsJXTn8e9X7BuvkCPVgAd2oJTVMch9KJ1b3ydr/LDKoRkeC
dfKMX8gwrGRKGaeumZPn5KVHUcpJl9hfFbs6EYyOmpK45D7oOsz4RZP2Lqk8DM8Z9xarIlydkISv
epUzXfRwOR7n8PszI3xqW5tV/sFGcCknuB19z3nX/x3svEC0babt4CNKMWV5ZyfjVxu4lXM8oiuY
Vtct5wD7uNCCBta6dQFhqwBIgqV/zxH4B39vgd9DV18vCTh7jsJ88Pa//xy5VtvjAwCD4ofebVpR
9ebdfnhOXvLB/p82LeG71Yk7TsvRns3HrlpP0ZKvy+00F3KwU5kD5Mhbtg264JEXQT3atDD7DFVc
1WNXA+5gRvhNwW3dzRBWOgWDNHXp3J8GatQLgI8GpW/IMiGmsjRzrhbWME3V3y/8vB2O3fBzijH1
Vu6Cxq+0OWwK8XVEFNcZmLdIsNXa2W/M21IvZjKM1/aFIeK0S3/vR7h/laBgUaWmAUpLMR4czlqd
sO5NI5EIgA9q64f53DJe0zHg0mRi2yIkti8g+iy/eU+llrfKhuMYpjBufD9nxWCnRMFldQroMvJT
S9Zn25zzdaowbHSCJArWTRcfs8itml9rZb6EIZNCtyWD+6ti6M0A/WyIYZVTzfnlLYO1wSuidYH2
SaP/maSF7VseXhdVz/l1bv5wrG45BobMZEgps44Mbpf+586mwSNWoIt91/rjcO5AlkeELAsi0Q33
IM0qO9Wgb1rV985V0KtlAtTGwmapC8p+SdaO3yyV5rzAz+CHwvZlz/9ruP7ZN/lf3XJS4yUxEgcn
XdalxQVbsK1nSySGNzsTHL2Fc57LwoNOyo+fkfW7nxaEaO1K47hhRtUDo5TWlSASw9GnkWEtLQB+
SsjJj6bxdD2SnJJjK+4F506znv/n19Pu4Drma21WLolvDYBYgyCfKuZl/6NyheVeZHCYVeKqYcP/
Vi3HOMMif1UTWjaqMh4b9W4NUYvnOkjnldCiHnxDIfhH1hrSbv2udiR1Yez+WNtMxxxpZ8QuyZne
1Kh1FYheZAT4yXGMR7mdu/N4cJx1mw4/uZSJaMnPJ1pPyrw4gOtS4silkcGQIpVvVQdz+QK3EEnX
CIo/v0ZCPdvftCKgrSQ+1RAGoENWGMcFPY5+zrutXbakuRLPrfUKxLbm7HrICivkSCTWQmZ9SBnC
FzLNG1LDRntNDx7x0FgRJzpMg7zU8K+UuH7HVnpvN+g69UkQC+ST5CNURtoNHlw7l+PwpUm6gGDw
Sn1x2z6TxPK/RmENJGlDoGW+Ft/yF+Gz8rPahaobJWgmAjIl7ZuJW2KpJamqBunxtXsf3THVY+ei
kDE5bcsp5R+RVNi1muBwPlZ9+3fXcxNo+kyMsaB16aJC+JYTN2idKL50oTYgf4iin41GgOYHbJIR
D2BEguRULVtAQgByiItfBcPFWx+Qw0fBITdqkTowh7AMKxRzbmbocR7K2re+/JuSLSifCrZSjt50
UNZCnJg85RgSuGHZMK0OhSPBxCCvno8X29+fKweY3HzCG1Lf7/IjNIWferLx0P5gjSn3SS7MHllN
1IufJJvKIZpjNsJMaXe64uNxJmq9PL1ZRI0AfiDUfrYVr2MdqUuiJOvsfvCY7VPWw8MvpSaVl7ca
sPw8e1fqx0hel7t2jHJHC7rEWZqTYO3ZU1ThOrECY4niiCJHO4L7tugr0YeEZvB1c68fKew9RSNq
1Gd3Wn4k8IEVMZYr0qH9sxWlKIjZw8A2QPzvKgnc8R/f+nvjHLLorsVU4xCi9/YasDsw37axQLbD
tyWBCfgD8cCiOwQxMsJ1IrKub6T1r/pKtJNpzksZW54mqWo1TPRn13LhmjckE7ZXGsNAoT6vbxMR
odd0VVMbG5c0g5mAzzQIKnY8Ct5Tlc+SfbFlZtmq40udXkvB4i+zhEe7IIXZEs77NcokK+C7kQqh
QSs0ZsXTvih2EQVVOM6/BqhExFoAZR/N5MK4taHbjcqWdpHW317hfw7uvqOUVtQ2h/rbEFu4bm1m
e6ju0UjS3KOErYXCWWv9ZTG3wrB6hgNBLDXx7uqarDusgIXuMPOPjg+7ugXnZo7IRaYhBl0nz1xp
IX6DAdQaP4MZsE+557HyUuGrBkpgp+dXls/y26OGSdvh9hSi1OFJyuGgQ6d+eRx+r8JzlDQw5cW9
BOgXV5uuDDKJF6LSBekdW6oDMSTUaqlp7pXgv07MoptrNZr6d0A9fIYzwE+tlxw9eUUojsLUpqxx
tfPuTWjr8FCPYuZYXFxbP9IBaeuVujIEbsb+u7/+eVsQcWR1mnlXpu7US4HMMW07MSl42MonO+bR
MKsys64ibd9VcKiS036/Er4oYAyNk9pQCpOArbzs49gn31uR/Pt0sAgpwF+rzpZonT2eLFodBr68
+pNwVMg7XcWWhwUyFZ8YaiSFKpkB84rRyaZw3P4GE211VOmWvYkYDX6YvrekW/4X2HSPlcQCAXiN
MaYgiDNdkwOvG0W1L++16b7DCe0ML2uMrV0JoYmI1du3pqFGJy7o+/qXYiVm38jQWoj5gwo7/a1Y
K7vwqjXKUTw67Dp0ih2zlGOkf5t6g8SS2yzoeGzCF87w1Pf1sAGez3gdZGKtDJhlclLGQTnVqRkE
E3I49SDvgX50rCoAWYR5dgc6gXVQ74td9JHI+uaRFr3dq4GJXkpusHXFDHO4qerkNOTNxD0Jf7Xi
8Zs3nn0m3mvwGHAaSbkmSJSu6LYk+wp5pH0/6RbFiD1JEkG9GUUoxjuE47fitrdmWycgNEH7R+hb
Nd6ZFixlr//yk6QqGMmKeWZ25MNZ/kkx8WnZQ5rpfL8dIZTohWBSlzaHvPi3x4cQg5kIJ5mOPjez
oRW2iDuY42npgubJ3IQB2I76XXFK9/Oa35xJHRNEGTOhnSgUQ3oakiWSBi+qJyYwReQY9jPpqJJL
SvNw+Us3INKkqQLKFyizFmSACAV1DBLnlbXkfbjxLm7uvlphCYnN0YNL9mKvIN5ENj1Rn2SEO1sT
/oUGFHr5a+WkKjs+g/wPRG5f6s5BlIZBuK7ypu+7Zo2V0h95p3HCe6E1SE2B1rSq9UxyiEuRMcGa
jP7eteMikPVmXakqfNuKjSdJ6S1QBNsfhOIJ65bocWSbDKehKjkyBZPYBr2D7n0hm4PttR/+pr4f
9yOKi9rRvui2TY0Jy+r2mLaKdbBWHm2dVuSCy78z7NeJj8oiegDCFeq0G4ark9apzhGfzJfJH1ZG
msEcOiyzg/F6FtsIYQq22V5cxQxBZJSKsWeyE1Iom5SBWVjknymuxkLWuGRc3rdtm7+9UEjAWl0a
8bf3EKlWtab0WdH9RsljErpp+I7Gr5F/OHbPVdVHDoy5apEG0Q0Sw9BBOxkkJb2wqD4eI3zXN4Xw
xXqhvf4D1Kg9I6MRIMnXEDeEeh4V0fywOitW5uloMK2nk44Lmqw/fhBLgQLEiATwU1s7vejfJycq
lS9p21LB3YhYvryDJkBnEilgCWcY2rlg2X1mQvLPaYQiH3rdLXLEf4Ayzc0JvtI1HT3d8xRoEFiI
Pe6dMgxTaGr/eDwPG0eqN5yTMeCR9YcSYLwmS83JeXK3JPu5I82sCyMETCfxfO59XqSsYkUyEk2D
g19B565jQ/4t4OS2Q+BsyPTCw+TNeaMqTrxd9PbiayeXrzHvjgQJ6O1EZoV9E9lIFCr7GoXzkagv
umsVytTxpF2FxDPNKTfC+0tqZIV99nEUf4poqcCMCX5OZz7HvdrTww8lL0RWIQfI/ZcSgsJfnUvR
I02XvwJPyflwv7sjVMd8g0JTitFEZo2/oZJxtaSv2OfV5wmQo87nrQ8W3qKm3CJ9ZoEAebH0gkwt
XjneYkr61OBOjcRkIgEKfGG5vtR6WjJp5w3miL5SK42nDvNo++Bii5js7vB6m/TOmYbRWy4SSBxW
0d5Dtx3qV4CTL7ONjcMpkwNGJX9C26ma/NRN76TDCGAbFRpizryZCLJXl/eQM/w7J0t5hQd3XZtW
wk7ou2VyI5A/+Zph+kqc1pkerH0V6CkrhnBQnu1SDSvASQQZKIRVkY7R6UL28ohb2MDvREOt78Ph
uY8KVJAY0ry2VN5N4Hy4HSS4IvnZBKUhnp/oneEO79HqVKV8Tb07rOdyg1IQVl8e7H2qihBfBHff
09elIYRsOQWaF5JLSo0jvtbdj0ykaPVAxulvHaiQkoEB3VKae9CGowuOj53wMOCqjTR/YsBUcqse
46BNdAfIZj1sPMspm5CHuNoMFFvcotTXjP1lG5TKW8N33Eg62cFaW9C4HoDRpgT6NUGkhJDs2WwD
sQFHoDS/YAfW4JgFx3GsgXkQJVCsGoHu8e0AT8iU1cZNJXz2zbEoMZ3oZ/5pRW+TptI9HQfowMzc
zVe9G1DNjMe9kvv9MJDzRSbaU2BcVyKw+fQZGQN2UtBgPFzq/gyRgZ3X9jCZ2TTnBZNekkH8/2OC
78QSG4ikj25U/8ENl7CwpZ8iJbaOt8DYuLChQ4mpqsJ7yyOLHZG4vji8h/cCR/9AcXlLwwqm/Hqy
xHBJLSfCKTIs282ibE4UvXTwLCIhj10CTe8eyW1/4EopFslW68moZKlkkdQhoNREPIp0im0HWMh/
lmo8CRCqqfkVE7RHqr0ot7Le6DtxwXTncSgNwCwJZxj6s6YhLw4peLU0jtA7NLfaVwCy9C7xhMqW
IWysE6ivqa0+lVkDyY1KcgdF6ZQCSGo49701WEl9mC3w3WflmagUgZjXx972qjfr9O8LbPxhuQvA
F2oYnxBX6EQ96r/pkP+1xdiBivEkJcwLyZFwvl/ekglmfyNKU75Nfwwhd3zzV9YZ4Xp53qFErAKh
LXtMH0N+9oVIqx9VO3nqQ+zTUu7SQ2q13JKxVYavyIRqFd3mktv7jl5AHHKp6sM5f5iBpNpJgDZP
dxS2Ta6xO0p7OBrVNBuFK4SR8PB0xeNr1bSPTAn8HN4FE+MRRbNeYOFU0CMVF4T8rVYQP4fRpYhy
wi4RfYKCz8Eaoy28P3mi/FqQC//yh35OUo6f0ET/sYzxTXLR9cBTPBJgmq7voNSaucq9AmyCqlVp
qwgYs5gRzAFzhDgAIqObSilrZY/V8+NcdUDkpN+zASKpfDUXPFuC2bkf3WxFBiwi9b380VgzWGRM
M7gKpIIb0yoe6Llkl5FeQ4GMRXIiJbaksDKNaL94uxWJkhfEsmT/a3Ztd2xUgNggiYiQembLSH/q
/88gCsLWcU4zBU2RW9JJYDenIbq4TayTEtrE//UZqBq2rv0qoAkqH298MG5/04dxd19gynyCERSp
ExuE7E1lFQRU61Oogk12Z04n7Q8MeK3+5qs+62kHZ30WmuTLBK1sk0bGNxI+1S/nhZi4TEUeqvaH
mlSpHSzggXtGcWQJz74Kx9YuG0q+K10nM50lSvkcRyUhtYE0HCU05AVpGvY/ho6zr9szmf5tK6YZ
sP723+lyUOmN0Isw+W5Xxla3Nv3LM2wgo57XkzlHUEsmumi2+42pct+nqdso9x5vf7fyoMKiG3iq
gWGk/t1TmJeHZFTqKqWGXXNogPaSZqlLxItR455dveMeAnfaiQVYfNP5FARLFp8qRtjInupsON0B
FQsW1F3WRudeCfsfEwM+aM4faCatbqVrRLBhjFxReT6chOWOrjPhzEdEQxXuuSAI/99Ds+w2N+G+
ak9x0Xm0DRu7mhFilB/AAUuCCsz1XAQ3RGoLO38/AZKgzCOC8p2INc/yJ5H8rct0jjpjrNwHaBbK
H2ugnL5q9Nm/FRxHZOhWtqFaTqhO/z0LsbcJAklbkV+eKssxIWCqZt/xSCbIp+G3ZS2ooG9apzmd
4SVYJy6KV9q6eA63EK1V+mdJu110AxcuBl4RRExBuPiXhtLyR4pomKLgSTF/6CAkzFkVJ5i+W8MJ
P8H2NlptKUXHjtY8LeVbcEQfW21wWQHkndneDexxA9al4azfY87qlds2IVg4e5ONbvmLVDXAbYid
tavmQsr9ZIHogMYalyg44CRHaeXYnotCsDx+eGdNDygW53Vc7KsSm0Gz0noNDQ2NIzaM2HMIVa+N
H8a5d4F0atycrDP2DHJxPfdGNc/b2XO5mNm1ZiZXHzut8EvfC4wZEMLLzTjTL2OmyTcUMjwmzmjs
wgvqbJ/It7fnATKIfB5LaXGc+0uIFm2Cs/jT4B6pQrI7xhlWeNysyOuPfSfSHWJa58qr2wyLGaEt
flhTg25WG8C8ZOExPXQh4VBzXWwQKAIPEG5YgHbBQfdEt3+TBQfBg6qHeoPpyBnbDOmGHvEqzu4K
xL1zzZY4Na7avqt0+mO25P4vaxBvnwE3jnCV87BVRSNaprJ0U7pFwQ606Nwmxwzw5pMJ2f2YnKe+
jxviWGrSK6IPCVNWyc6rxEGKwtH3xhu1EW7aQJtk1wqF2EzcPEMiYMCkp5YR+XIamffY7Srp+w7O
8ojzxBFaUW1xwRWwqEbQTKz5Rse7v/Px+WRDj9E4Yojl4qonhtjnNDg87qK+hYH8YG2UoDPISyGW
KgwyD9F4+HVOabLdOodDUgpSKRqu4Hu2smsdrvLoniVZtIsjsRBFAc8nc598+2cHl1e+YJdpRccV
q6SJ7eaHhmxqm1OEB/vZbAvp++ZF7vp8/Wq2TUmgGvuiGVQoMAgSgje58WtE0/mdi02Hy4D9oADU
V4CqkJQv7yHj8atC/zv1QeEckGYuag4pTK3ZtPl0I8B5ZMD4Vo4rClBXy282FVfw1KFK8YuM5rje
xkGkUO2cg0jfFXHYcqlKoYpdg9Nf9B4XPq1XLgSN//cITxxlZaG2mSJGcckWjUuSncZ3kHh3Cisl
CRX+qvWEHvy0K5r0M90KsJBAlifxFRyGEik4qH6o13WwhQFHi6v9ZfGLt3//WqqoMrZ6rWNZQuik
TqrpUwsu0smMPgkCs2+7F2Z0AkKH1nuuYGScxaLcRQPhjv2ms7yVemGDlSkZ9WFSkJtAl8ZdcIHG
dcODd1ZrzStyCeAFopQ3nl9y3HGFH4YwiCntled3AKbbeMrTIbNWB7U6PtMVjC4H3JOARm4YKm6F
jYTXcDsu2V0+k5XQtYcfB5ypk2nTR5xlwC8X0ZMWE9uLl2tvncrQldhPIf6oUGGk4WiHMwLe/o5e
tJw9MdQZ6AS9Q1dejFjchx5sTt4LIT4DUHFHdVY+69IUDZxxVvzozkD4g+TliuWVSprYmJFkt3t3
u6T8bv7QJGxel9AMYw//jqE7w20fBWy2832dzOi7bXeDUygJq+A1sdBulVL3/nmpjXMo6oaoU5jM
qI6bbnvTQ8mjAtnK/DzwyLrCSzHwsESnXdu8BtjiqJxiahXGDxbZww+iIWln/3WlPaAFbhk26eC8
0INj5mmodFq7CHVdyCw9hPyuRbSe7DXuFM2UhwUAFYfYuTmB2TJ1K70xc9rPZT09WLVV8rV9g5pt
kvBU/HhGTKpWOpu4sHwDu0Efj2Metcg0cODsxHVH7SCZCiQBHpWPPsjLmiw9TSFhFzk9KUKbEfuv
Y/ELNHVo/owve0moGVNRyq0KQYN4QnbvK7yTks6qAC1jBjwjt6RmuhEVUpdd95ADAeUzWnd8XzPK
gejtj1pZvUHKBbp78yUC38PYuNB8krEkKQjdp5rlVTCzIf13+hRzF65RSnEQQXf5TTdl29y1Yuja
2V1FHsyn2BoUlhpKsq8i11yunSLxIQRYoAspmhdXrh+F/+5TD9m7NYdxicwVr1cB1GZzQOijjMVt
jz9BC5NXqDR0gFXo3RWmNz9YTquMzCMQzUhQxW91STIxko1FkCNuLjrBGeXqFgD2BdhdM1QRyLEm
IkNX7EoDO7EMHfFnMZbCiIJ31krZ0rSZ7N7Guw5K55ZFJniVfKS0XwBICsVFlm8OJlCBNnnr13o1
ongbbNEAYDWbdKvUEowtJbaaIdvB1FBm9S0Cxk7o0V0NFsu9XgzZJYaDW2WFZ/D7xX+k7Z2kTX+w
sVFKL3lJRl92qoygGIAAAFtgURMtrmKOgsQY4A1GC8Whrh+Yk70A9f5y6dsr8wEVVmSYwRk3P+Qs
XEyA9m92ivOZo34n7DU5CWWqYlvpYhv566+jZJfuHuEukrRhs9BfDvdW67dLRuWosHwfzOQOuW/5
HATcQ+1/IasqVgaeGuWGiM0Wo6AbRXelBQkC/4FA+Kr/rIQGuY6OeQ/qOLxMRulf4hzRJf6Qq0tc
NODnjmz4K25Jo0GUHcX4woKIkXYmRlltD3SfwGbzQ9LUNBLQQrsVsJd7GBYKUCv7vAPqPz1wJZHV
Sc3zlkW6XyfvZwFnRSD1GPmAqNty8MJWHKdNFCL8ESOZTzPSs/DYNT/BcBG4mReyiSh1tui1gl22
3pePSl8KxWyUb1riIkgPfN1sNtjnxL3rA1r5DQOQ4JdELpcZ4wBjdOuFSsUDJpBxlyrZunk8sNkq
qDdjxS63C5jq3GiJQv19hEtei4/3E5P4v9pITDief/Rws51tHl7U+JrFE3kpIJV/UKY42nfrUwO5
sq5DwYpezSI4TkzPV29RYLEzwyqyqoRZeDCEoWF1jxddIx93sgfxXEWSUKubYwUngVW0qoAm3Jqc
8IUzuhLwnR6HsEzBH2EVKqKZ1SyaJ4KdFLVpXrtJJ8wLfObzSDhRVqZi5Q5vJwW67ry+ddyiJPJF
2JVtplpyuaKuTphLVq+jgRrzodTdlxUaWUaYvxTk3qF7OJfC/8EdwFZtsae1mdWrnyZeeyenLoHs
L0qOcLyAXoP7gtu/3hiG+u6tdfHd+++YMKJgbB7btzt7gUrdK9js49OoNbIc5RmQ9lYE10uo4Caa
dl7Um4bzKW9kAvAlVluoN/6X2k7T1Z7s9L2jpAuAU48IsVeJquULs0aBGlyyPpdxoTFDnaypWyPp
GWrEWUZXaACpyL7T2LG/irWkZHMsMQdN1c7hWTtCgyqZGxZEcO0O2xOEShNbwGM5QEnppjtfmmPy
TuDhAuOMv8s9qJZD9HSN+0Le2pGhX/jsLJCYGjwMY013FlBMCWsRgzv1CFG0vIHG5LyL+XDTfXQL
6Do4QtsxrlU4Ji7HADY2I2V1O78tuMWXdXvF+pi7Sfb+/GKzyUeVdLRra5cDteA/T2nP2Aqiuf/V
7fYRrDtsPbXucDlACKo7Zcaiu/zk5EWyD1RclpZ2N6IwFYIAt9EIN8ExgSUOKOfGrMLWcXV+7f9l
1h7UMz8FC/DjQ6z2fzhND6/2Vl6gz7Yy4O1rdEs88Ns1KrBjV/8j7GpygD1Ax9sZG4uZfyYpo8R0
i1ngwHvycfIefZFlFxuRt2U2WmRylZyrAmmsXBX+sStErHfR/WgiWrQW4JRvNwmCZjblrzFDOVA3
WmpYrtnF/q41f/z93Ma5sC/xrirIbyZ6Y20sRjkhROeub96h0k5MnrdIr2uPU1UYEz9Pf+im6jQK
nMVzFgjJEGp7s/Wk4EVxx/xaBDZ4BfUVBokGbZ3Ij25oKFL/TXznClqpOeg35wPtIJH9OvrU6zoM
bmVpTxJ1K/eSZosLRVv4sAk8oPNnBdu1TNFod4ilUtT+5mkFwPhwGj25qIgkcBgUdoLQHM3+EQ28
nSJ/uGx2AdpJkERdO128mAAL0HwElMpHG6wUz54bDzDURujDeByiBrBLQwfr9BsA3a5VJ9DJjBYm
zvUVVKHfItBKt8JI011y8nfs13pJyIhquSE0h7Qd8WDu6P8RcrGdr4TlrfSeqRzhgjQrkaWaudVn
ZNuSKxliZLdqN+1nIcjKKeZoxXRu01K9XzmNQKecWNtG3ri6COxOLfv490nvVCrCJt6aK8eVOelg
eoyRfNd4LzywimAFzF4VLAkR8N5zV31mmM7AXbzTMlKkfs0s9Ao5TFw3VZvyOvJHVZB7cqVU9Ka3
Sj19fjBLCkDc3woQIM8SDtuTingjmUGY/d/PKMCK3tDcme72cI4/ZRIaBVI/zUU+ZKVHwVnbp/dV
WcqeVk3vycFvhfDbX3YQIn/y2CFyVh4B/WnLrA95ptYb1CctAlat+zXH28Z5T8xOGhbMW3N8NiUr
6FZyl63EYzzEpocngCx2YIqa5WXibCwPYwG9Xnt7U6bzPtLFpXMoCem6SPdlkZN1joCoT5r0S7ST
nICDdm06HfZrVTtyiG3BIa930Jxz/r0yrTRsejzk/SGQKh1UN5u3SBQm0yM2Gvz6cqWkjitmVNsT
wmdSFymozFq7MFCaaAgSfTWma0lHtnOSrprBwL26vz/mOOgDNEBDdecH40yXrIQ3xCxEgRWXPyYO
mfEYe3xFYrlk4UcSDthgJ1359wKrQ4sgeeHIVwr1T3dyKRN/8SFYe7x0M3PcL3j1wpy0H5y6VtMa
kD8uUjsvJJD9x8RVQFI5ytwrxDSqeu2SUh1BaXBBepobLxbN7uwlMD9S+XuUYVJG0ZyIRQuPKA/H
Gmvbg+LSnDkpOYMiHNTzA5SwFjrYUqUOCHcdbn15chZiaDjH9zAgHpbjtoMEM7jaEnreF2h33BV+
NP1Z7NPU0ZCSJTut7RVgNAFFmRor9UMUDjd0B7+RWUUso5Gy3x3Y9dUCN2PiwymVq5uEC96rQ44K
0ydZSsJeATr9AaZ6QAWmybWNGntxhAg5fgjjmBkfSa1N4MGewRgdHaltEdfu5sl8IwHZn1AAnPPX
tLLAdBRdGT+qCUuX0V8vKjI9IaH9nsCkiTt9SB4xZALWfqoU+SDv0nS0hKgkD+fpnskVbfYFKvkp
bxOYLc00SEcDwdy96YPcdkl6ZlXRjCmq3PUi8GudPvNzbONJBU+CBFFBRe1RayHX5PSJPl/UR96N
y5oaa1yy/xuvfzhybNV4meMMEfZ93ujQRKgrTgBE+LcPNAKgBW/4LAV/rtU8eZTcr0Ld+GAWvpig
u8I2Aikrp29MHg1d0/q3KRT+lqRwftTUiPxq46yYTxCE6cUp2X45NQLYi2P/THyxqU+GxcivHB+u
FNNuV8uKfDJE1CYUBLhxPWrTo8JTQMN5jsNQHpGlYWhTGhzUpm0BkhflibisAK1Ouwbw8YwCh40j
ifKav4lAqoDbRxNdi40FA9neyRXnJDLOZaxL1xRKc86V7wSaGj8IfSiI8Ci/l2gZIC1zYYqs54WU
miE970PeCH1dPsCDLW0J80e/u0aj7Tzz1wbMB1mOU2UkGiNs0hD4vYAFYeL75a0VQsTsLt2eajk3
D8p7oONsi/rIt0mmCpXTdm/9On4SMQvE2BytbDPJMe5dZ3xswmAq4sO8Vq4pILQE6gyNhImaawbY
xmmiKcqaaz67nI824QpEnOoRPbPeLgZVvJKkbtiGnuQGjAupfhW/qet1xoG3ESpodwbwCivfcbqF
dWUhkJcRoblHs1YlbFGdt0W05LHLiyyjI20YNsIN+y6tguGx/SKbe9yCcwji9HiUwpXX/7tss3x8
PyzyW+S8tHwzqft84zecWZg4IMmDqUGf3wIXs1T2wKN8OmHY5b3wdwFDijQlK4cubrBxVA3s1/1C
bVJxm8VQdK01/E9Wyd72+Dm/zLrm4SpukXR2OdF4obwtadZUAkPsVZF/qgkRR7YPRsTnpTl5z5Gc
i9kMuATSVYef4MaZN+PgUrsYmp02RkmUr6HwzS7ICojjOIpv0aUbsevehxEtS13UoKAa18dN/Vfo
p+SFzmb/61Z32+ObdLuHmk0NF+8vECgDFXqIhiZK1Vo3i5qP4vM7sg6RESftUfvhGf1ouKjJDRwu
N4Z2nNdHXOdK3goYb+T7vn6bhgBjnT8Ji1X0Sh5IAJJGv9zBNr0vg3uGTyx32PoeOZQlLmVkGFvJ
mmclldWqq9OSepMxR71S/1gPBzyxrS1lNNmf+5hJ0lDR8hiUeBcPd2wVfFF03jn6HOqSDFy5AkZb
icKS5ZrF/2hYatvRsRmM+3hPlckkhmpUX0hPxWQcnTf2R1HZwLUfNobaNtzHi3Pp4qKQm/48WpTb
I4BRuE/KfV0pHmBn9O0458L4QhRLYW/HbBYyyB1yFJyqqaWvPYlkpZb94zIM7jU9TZhsxpioiOvi
P/MVgLJpyVKaRTXy22SXpRG8VK/yuZBvE7MyaaElaBhtlZXTLqlfltNu9ZDx06ktrkks6hNOdKjp
/mrLu5qiixq9mphLuf4fySe0oypzQ5r1SYFSIWVg76O9wNMiC6c8flqqgJgKmhl5+p/O6BELeBT6
J2St7cCB2hCT0BaAP+ulVbTX7uIeUYnDoUAxLjEe+XrPpBiqWyfBWXvM5KlINWoM136ElPebAH6D
KL2oS5kw1Zt3jliTEGElusQn+Mu3wevYow9tout4iH+i63ckSReCRf01wKQi6e3l61hPzrxknI2S
LcTJCEa/Z+5w+jUAGZIX3SGFCYgMWbRXvCeXCZpI3pwTZMt/nTrSoZBbrzM752CSuuS1KrTx4DAk
RM+v7M/gORNpxFBBlz0IabfuylOJh35bJoj08aKYzKcgCJRDBhU3YuvZGi6A2V4brFnV1pDzuhzj
K7Qbb1kyMpXW+BwA/cqrCyxYdO8dJ4/yi6k0gbx4461aK1X1GYAP7/85Pm2+UOdZu0WWwtucDG11
ba/fnD7i8qFzffoJ1DMykr6Cq1iNA3NzApz8zfTTM9Hqg/QTW+L0J4uuJCN1tfHSQyZ5vqtqNgy5
+2jLloivqNsholESAROZD+lJ8TDMgJ0maSXIyqSmZKXXg4290Sry1SbBJZJXNM83fg3wbVzHrcef
azM2Sm7jWNA/rsQPVjCZhy3VxO6S2+WgxbN4Wx4We0zEKiXzCEQH8zeG/5U2CU+fhRqCQqzcWRxZ
rVrh7HVGpgE2MycF8yLbZAKw9sxjtqGlZhY/3FLveLdXkEYttEjqcIt8Lhw7ksy5hW3Ufzam2+v/
0oQnLU0dW4mA2lwaF8XBOpZsVnOXLLxhH8Yv2ZfZqm69dwEIXl9v1Q9eLfog1viVLslCP6HG0Psp
aCuJDzIf8eMSez05D/UZlURrpLL7FqPfhjKN5sP8TOgzifvNLMdiHamLpfIpGLxBc4+wD5T0P97d
iu7N0GV7OGHyd6R7T5UE1sggsn/u4xBAdltDdwmvdDyug0dC+YbpFVuTuKxn616HwEJh2+Ut7gPW
53TN0tzbpjEpOB7XHEfmUvFc4kgkiivvTMQx7H6vbmsC6Mo6iLav2eutjIstiirv9KmFjK1RynIz
zoFC+hFgGdtfJU2X7aqcxI4Xm1DfaYasDVhk4ZQKSttqLRrBvI+csZBzWxNC/7XFIoJEhtEhhlm5
/s4wAw+s8TTKGo4f8xxq/+3XE1CvFmEPeeMiOE+xX82Xen1/cxDn0Ao9P/LULkR1ITk9ItYRwNvQ
MQXyFNlC4VBm3PhD1a/zDtSAyY1C2S/FuGRO/d+Qsq/VVo+APHO1iWjYEws9yzhcxSpnrABlsa6u
oNCcuHxAR3PMJy38tQKjhkXSKWjsgW4+HlmBh1DZfxnjsrO0bdC0H5j+zND0pp27g0CG+g+qFP9w
zS4tJ75EaaXTcMSFz6PlSU6t6lZpb4frgk4NvZzVr67eDkrUF5D+gzMufjnOKgFOFzTZ/4XwcvVU
PVWHH6ov3G9urY7zNMZIrUXViiH6w2pNAQLKh3GkZ/5qpmjhZsERxVJKYCW9Aute5qv70uSToR3t
U+++lcwuJOQNBP+oopPqtPGJRSUK0eYmwvuMUyeBGLFayvOGWzELrXyAmmcW9YmMCpxZM6vHiS5U
Zr94ioMXz7kgpvcG85UppLZP6+GJZVg5f1X/UHrPtXhhddSNG2JHyh3E1U1GSS+auhyAbIduaGWE
nJqEQdlmrPjgIq2UktD+0+sqDLcbnEQEYJlA+OO59DvRMyy8rMV2ZnDjNSLQMYeLpFfwCxuPoTHw
mDIck0cxJKWccjTPPA9Xn1jACZK+nedugBCxhKC+lAi/0W0inMIOa+EwNFnMTVv5R2SVMwVLToR/
bqhryjszwqZLrWIykBdpWnolJUdvi65n1UZOWzJ3WWAnpEXgdFR5goqvgPgRd1ZpHMqSjzpQt6rw
d6sPpYlJMLKSfb2U49zCT7kna9i+K3JAFjjdqndXfUmAA84h+ihT1rOxtVyUJUvGBZtlRYadciFk
VezwW9aPvYUFsKaMrAAsaaz3hrAAyZD3oBWm6wKdKGYCsuD7Y1HXM8ykRIPAIJeSDiF+UAvGg3xx
Opet5bC2VVXGmWrZTig+SCF1eSIF1GCAn9c3Jru8Fp5dlBLQM9Q2Fjyqg/Svd96HCtl2sRojj0CR
AzHjdYblQp1NLMdKPVdUqG9cju+t/O0jYTS6KFcIr2F5AeRryRylIvHcp3PdZCdUiGSmUaxDW8oJ
eAF5m61jO/TNuhPJT5OHcDeTBtoktNhLgiOhatUDx1WwMfix3PFO3iSXb74e3rd25b+Tb7qj7fTw
EmEhbFyZOKjee+YqtJa+yadvKC2Db0Lpzonfdk1PEhg65tVxq3Ppx7j5OEz95fyeXA8gphbC1qOj
+SJR+q+Pl6y4YHPSfisZGJkiat9AXfJykl7WonrNVYcojsrR0ltzYTkrG/cjC5cPM7Buuie41Tjt
BG7xMqWDx1+SwoVDW2m1AAsykndkBHj0fK0mhNLZAwug1s9DUOkzrFqhcBQ1lonLIT5tX2wFlCY7
I8/SNwrTe+zT6yFbReD5Vx+WXjI5daVK78yQ4rPPRFDacfs9d8rOzT+H6NYe1l50vtPGFdopkdLD
Hd9F+/enIaN51PtWhk5lHQmMDo78a5kJdvrKfCBf+x3ltZBjXLSKRn6eVC1G7MnZT6smRU/+iOOG
Mgv4dVilE63gMNDwDUYWN7gKD29vgBYf2oL4+nwJh4GPL8INhkHoLlBqCaEaHQWGo5w523RfgpDe
U1ksyQTTGQRAT70DAd/ybgNUJunVer3rquszcBaQqG/qjvNUbeNZDxzmyujaHvz5TV7c1dNQYbPv
2GTJwW7RXGAKA/NB3fN8VY5Eg9J8IvT4GHOzk+OHcWZ9EfX8Wcdd8bByiLXTzlSRNaTisC3pBglB
RKOpmxb6r5EvJcTjG/VY1FdMwk70r8yUTq6la1222gmuZh3m0E+OBvNw+fg8RAYD3oSu/YdkZ+TX
bhSkRcr3oIleGPZm3BeIJE75okkQuIUz14UzWScpnhEzBMCaUtbjl/JLs9fRp28CTxPyPdgsft9r
EMgr6jUlg/4V8RBnJfcwnTpxY07R+H+QLdYkzhX0OacGoXY4r9u6OpCqLWWX8SgXwTwtsokbTQJB
s/8hXLIrhwRZj6KG6764rVnRxxF1LU22CPW2ePJ0fuI9dSbcGLTBidUhpptqqzMwFMnpHltJGlBD
NtJI24B+2MqCskqCdo5qebpcAbvb+2KYXTeZglIouASWTL0tID6EWe+8KikLHupT+b4UgCEKZ8Vf
Yx7KTlYOMXgHp8zz2/OHMqDY28sjRO7JFJsgNnqlUYc01Q9w4u4BZaHFBssVhKXUZm6FOvkwucFU
SbYjKIGhurw5QNc9ncYmSrn9NV0LR+JTXO9jPrTe63s3ynQM6vHeidlIkXcZrQXTBawDI1i72z/w
02qAi7PxpUUr0la8mSQLpwPUK+719+sVrnmgdaveSgZalUMcP5dRm6r5bb2RAeI9SrLBYFTUwqMh
KArZGmMPGKb7WHDYQ2IrWhaARaaAys36x7ZFTS01Rl0TbrY3OCA4SVcT7EfxaQAmuZFP8fMNZTYy
CMA3SpYhuJyX3gWfzYVoCuggJbYMXJs2l0MNZoKQUUeM9IsCIo0uTB8/2D2fWGN3yiAynNKigTVk
ICi+QWo4L6iBprnHRXswKGPTdKgENXSTOXpEgvX1WptbLooex/YGTpriIV6RPH25alHKv1+1qvuX
E18sGalXc0PwqLAXOtniOlEscQSeBD0UKS/FyoNyL3doVuilVj8zjEIg70Ad0F6FAvYMFLo8muvZ
olq32PRxSm6FVRo6mlw7gX3n/m3LWY8q/0rpk5Gi1qTzCOhwRHYrINjdsFw+kcQKDJkcKMBSUmW7
UWlmdwZnUBw53OuIxOp1UBoI3U8JlSZ2N2b9W7eCE/UJoUXvNbwCN/YIftpt6DSL3vs+M5hT2+hd
cbdBockH6aC38yzfCgGI5PUaO7yZHDSCi/jQNa4tZfFMU2roCQHp+KFcU7C6aQmjDMliuC4L8E8m
uMBDw2ZV4Gg7A1wp/g9RRMSiVcDS/+sgkXJSWpXGW9V4ByOu2vh341gOtmZFG4fmaDBuO7O2dQHL
49Ix6xVIrDiT9T5cPzxUsJZvOj6V5pUsSXih/jfXNNhvFW4nfPCroyX8czl/0JSByyLWyn9HRdp9
fBe0utc2K7KU+ZreUO+eS+GJSsRGYH3FCFxf7F/QMG8Av1QHl3m/u9oYZEKauiCLtPPRvOEeTvSL
XC6W3n4MAwFJu14YjzbHunj2SHrrGexcN2sO8ki2poYSlrLHx6c9bM1VT1Xi6SdoG/2+31qKcAOV
uYUdeIdYAtc+dfATQ1eXN6MpSg9nl6wZjoMKXONtsHT32aYlLqF0yTTZGYcEOsHeMPECmqkXhoDn
hO34IhbLb9NxigpSeJJAmArS49egHEsgNyPOHiEuEoKzhggmuwxgpATSIbyeX1Zqxj5kRel037bK
P8EOk45baOViKg7CjstADWwDIkKuB1WKr20itbAJhVziCOloFGEBLWDMmXGb1tAZIWFIqOzpPxio
s1tjvP5vcYRLo6RBn3PLKNGHHaD2AK6UJKOsZzUDHowHXer76NDKfBxJPUxDXpiXMjJTFedinLjr
HBSNZOr+9Ww3u72HzQ1CMLpPQoIDCecUBDMBlAmETsDNM3MVC6TNQ3ha/H10iOSVUpwWljOPr8fS
AVuum294X0qc2m0bZ0/8WMN9yfrjtlpRxcnEtRIT/bc9BGuSMANV0w/BCl3wMtyZOHKubTnaj32V
aEMlDRhGEvZWWSB7kxTZQnghbjOXk13YJ9B82zo8/AqCbYJDacqDKdcqbclUyqz3QuCabFuNJXIa
SiSvtcUt5HoDCbcDku8G/REtGucO0O3ZzpSAMCU90xAmE6q0BiV9S2nRYpCYpwgug04yNH+ByNeA
pxT9b3e6l8JUW4ZhL9AhhRbdDZRARN2U7XDDre0HR8lb/fxwnA3p8QgkJKJSKoNSpTQhG31l10Jd
SoM1C2euRp3+04cOSKYbyYNpY5zjBKsWNx7tPHKc6jD26XJZwWzT8f9osyu+nyGUltjhUSD2z3va
W+Cgr+n5K/dyi1xGnD0ywc1+e+VHrYm42lzMrHg0v8CgkxwWMNbKukd59IoSPUTR77kJ0uym06Dj
Vg7cz4sgFpZPDolYGooPP6trbYu9wItahWAxacx8wfr+O3/PlQ/NCiS9SWc7PrR3FStYprjiZ9QF
uxYbdPf7VsMBzHecacQ21CuwDbIE9fR+5lXjMbj+15+jBXrQPhZZ51WUcfP2dsPdmeaMGh4eMsui
9hQPhNQuIsSUM3MJCaev3OrqBeSjXsfXaE3akS/Gth0LVSfEFmetui8hmENG1v5g5VA70IzTYgPB
rd7NhB5Kj89GfaQgO81h8D/aH7LrXVFP2GoS12JKoySO56bDo50tJSLz9KD4G/DGL7owEAzMFEpn
HfWBv5lti3O+2Rxr2fdYJt7JpueSWWGmAeR7vVHCTOYJGbHQgvZEzwj5xKL1Qp78mlP2zeGUgy/f
YbHQY0mH5vvDU2kafuGziradJRVlEjxcYi/yRkOxOry0Pq1xhzTUNQMFwJFIWkWR+t6PWFlwP+RF
9xlLfp7XKYVKf+soKvy8MUspRvUrA5Rn+7ZaZjJWZbtxSxKfY2G97wWtdMNaSXLcRxi3nuotD9j9
NB0p90MniYvyf1hortJmo0IeOrWS/j4xmOzDjriENfUVGn2liMaHXCSnKxE65ZH45iDlfeI5YBcY
UCIrDe5o/0iLktMvx3LP1OAW1gkj9uUOtrucj/WeUlmuxTM6BzNzGQXYhyp5Jm62nhx7bOJsOL2t
i0XORqUxr/8cZa3GcO4QdokpLEKBAZFLEEUHVsWJsQHwJ/xx3Zyts7z9d5c2DaCjYjTqqYyGUxwf
k7HHDzJ8WimB7n8WCu/tlz21qXBAdpU69AuMZ6hAJn8kzfXk5X6JeglIaSVn1IaVif2R8w+rTrup
D8x9kvIKFxlRcw8C3BNp+BYZ11cMweP8b8NRY3dTcq0idXe9uYLtaMQLpGIPFsrPimViIU7UeY4Z
zidXkMPsLK9q08Y+QYnElqxJNNIFSQtDPgHh61TKqNQFqayxYu4yV4kttabYXvuvFYDuwaIxuqcU
7lkawUErYd46OK88t6CMFmk0xrkOCAoGggMnPcLAG3ziCrUXkMG11R+Ke7kBZLqQ3DAX68qCOqPH
dJ76hAgyDM/JRxIV2f71ImzwMxHydkmJot3Mbjq8r5PQYUNgP96UzgoU8Rlvx48M4yb42OeVFI/u
jIzVZOHdbcDRL4GMs7MP8/YfGlJVyAuNe76rjFbM0SOf/RvdWM4ggtS3PPe5BLlgI6NhB4Yaqjax
LFcTocthYvpmYsaabKvw85oBycA+BB7Zpq+0pAvumVfzeJrbqCNr1DHZvmv4XMDQS9GGKOL8xxug
ZNjdwxXQPDU1b/jo2l2CbRApmd5J6iBduCxvEpGU05LmsNc7VRkRuyxBk4szs8ihAvKxc6oul4rX
wRh1ACy5Fmo/STtUyiCj32K1BU65tuMDYnJXhZ5UOZNd2Ad3rb3KvnAuFafmYuzS9sXjGbH47U94
Muc0PR2ENhx4DjilG/WP6+cmknoxE10+5DDGq1/dfFOUqHilVtznsVncUTnYyr3d226AXLXVbfYj
AMUhlPkpmUMhoO61wx+h1al0FloVk8Zp0oLTs9qy3DiCytjiQxxC4TW3lfTBancu7xV0uLiAm9Ef
m+cLJ1OZJhwk3lvGsA+LV0pBKG6qUR5MC4YwnFpCcZx+gEuZIClGYYaiXrlJOFu2pwdGTC8JhX0i
w0WOvlUEFhcIjLTq8wnK0JIuQQFOa2sHqfjcv0K3BanEMXZt0G2yv4C7/iPj5NDV54Mkdfmr9gCe
82p8Kvp/AcdfBsCcd78fBwgdtEJzTadjj6eVs21n1FXiQ9gkT1kzDuD84/4uLFZHeTJ/TZ1jYp7V
SW7zPwfYRScjgPZK4pVTbob6boqfz0BhMRRoe46ocTPsZy3sdK3okBtkDtel7XBv4J+YV0lIB2xj
oacRPP8CLF7Bkp4EyHgH9w0p2OTojDRK6BjVKsrdjhlRP1kUfeajLZ77J1NXEg4XHCDgjipQsGkU
Q0zvCF7etHOMk+lqkCjL2EySr2YDuvnkqbHeZ+JIkYOQ7euqF1vXdfJYZfMDEmu0D8gZlFGvTDHF
FyPOuKFr12INdijLBuG1PxLVSgZ+c/d0CaWQgwOntIOHc1NJlYtW/bipcutbRpw7ETW7aapIiotM
dWXgxCd3n7DfgrHhMiwv8aRxioeMUcHcFfFFEs9FkzN5Ixyv1kwIDIGfb/uFILQothiXpuIgc+KC
R5H+4V2coq2eudATzKlo4ZXCBTOmm9+H4TWa1PgYSdFkf1PmMxEl9ZqcHeGDa7NKAPdJe8Va7p5L
8l+5PAj/lHaiJY6F0rrKwuXBvE/Zp7S9vlsO2InM8QKRmg4DpzoMDXwMwA4u9kdp3OY0h8Awze/D
q/6NcKIFkHyDLPQ6ex0FnL100ORky7tjYUJACT7uNuDKkWyZw6pZUhFrYI1mk3pE210BLGQ/GXKB
5W1EUTbvchFIdzYDcFZ4x7JDG0H9Q/jxCIIGUl7KjA5HluEcZeuJdgHDq2UKwNAfMLXQj9cup4sF
4uOiykMb/K+9FrnVNI94mqfC18Llf2l4r5ib1PoIICYzuyiO/fpCSAl5YBt0wOPeSCU3jVvRJfse
7OTZy1Q+K+1M8NwaWrJZbMXeHTfSE18umw74yRp+itPoIzngknZzCRLv3b5hLYUbZGRzGoMULZV+
LNnuh/uTGKYVfhGbV01iYs1cHDjUd65kgZmiDYXkNHnJ4kQDca2lIuhiwfkrxJ8y30Ehq0ZR0W8E
yDAD4ony6yaqpEcsvfBLSBJlRc4edQivfq1XmVHuDsG8Kd/wh64UrWiHp9WkLXnWfyoaZmKsb531
pTiqr22kW/W+AyspKU5swRBrJjBAqSkMji4OYyR7W8LcM3IE8oBS3kXSoEjC6UR3M6dz7XdDrC4i
NMZMYPA2eprFDz0brE6nlhbIS2gevNCRbuAwad45t0il84byrkIyX88dDPlBiF3z6sr9KOgyd+yn
6aXMbFmaKFPPsnEuwAmkqm6gArB4E5oc0MlczEc7jAzVUsp9sMiId9xDNYt6Lsuy34wOHBW5eji3
MakUSru6putj//KwRrrp+j8IcZ6pK4xVubVLv8yCUlXEtMmsRXFa0GibHHkkEvHw0Hw4fx7Ht/wq
Rep7zDm96xPF0qNEWC6mN4D27oQRJ4D+9yoNqctxuVij79nFLcYzHhzJ6Yf5IwzE/kFknw8+HWKw
diurd5mvCZd1o5QFTF+qwktaxCzA40vXlFVvLp59ABYD/dE/f/UzVKiWGnGM+WdldlEZmYHdFKkr
FNo2+IPnwGM3Ep/s7JAdjLpZJ5wt8hI7TgxX0U2jUB1l/xPbylFSuoN6TQYCrEUKLsVA2sOkw9XB
UFB5RwwSYDUCr2dC/G//mM3/ORZR42lF2FuMFBwuIjciWL0xZl7VdUTw/LRwakbq0qzfx8tfS6vV
FBNNHmMDumNTH/NpSASIjB1EcWPFk1nBWPaW1yl0Z4FVvfDJhUHp0gadWjrjfum3za814Ml0pL7u
KzWbiyKyUX6BbTWg3XAGNssOvXWDcmvT3YeN/L2czRL+rg+zvwun/u1pdoSkii88crgGoDlZcjLV
Y+u1XM14HN6I0qJ7VBdvUt6cKJ0kpgawV8AfR5BEHl8UACBU9OJHKu/n8hb7aT2tsuldRzaTR2SH
70ZBqXpibTfHXown95ky00R2XQXyYueMWDtMD7KA13SYcDp+lfv5K9vbVzmUgokC1FFbF46Xe5Ue
I27Ubih2W1midrS7Sy4G0BLZjeZ6yHLynO0bKdWcXQ+Rnrhzv01uE9aERKlUSGkDLle71FqTpDic
D2YXbtt/JmOYY3Tzwn/wVuG/tfPJOKV6K8PmtR5GOFerY4y+w3h9wsTXKmz2LZvPJc6pUNPX1YQt
qNVa5exN+WwT6yp8YW9aROCMXnv3jLt6XIcvwfGbYRYwBFefN0Lt0urDZL/PzAFA7WQiJ81pvquk
Mc87gbpXqL2EZyl8rAEDtbqoNdyPT8jcGvRvLI1UdE0DkhMC7EaBWDYflQwOLiv20imIt23x+olP
jZXfYzj6UXrjYIqzmchIw5H13DeL6MX5Scq5jRxeCMWaFElXiqzR05zkdObpA+0TpjYixGuj44+X
+opB7UGVsb346R5F+f+Klf4uQ7pI8VSwS9oATE05QP6HCAMm3XgkZpV84gxzZXjfhd4bDKhfZEah
K0wyB1QhzLKWlllkP14VM6KUdpvvOTprJU+92AF7zQ3NqBbJ6WyX2TR0QuY+CW+JC+UdTT6Z1Q7v
KX2AYdV+mYRzE0FeU/FxlrZkk2s9kO7TP0BDBFG0EvmeeAqsJT8kqyUbdPX6uqjNFVVCvgv3tHDP
x0bAHo2VLJ+Pb+xa4lcszsYoMq8g0Y953wpTWWKJKAJgLwo2Jm+F3WMJs26Aa54/r7kv7cVPS0Lb
QghNE6ATC2o1b7CfLd5s1UbRkMhnrPeIrqs5oXXrh7aiLhLVlNPkA37pP9mo2+UZfgWT93oTWTtA
dhpI/9wBfazUIMBifryFaj85Q5C4yjPviFoCYMwhq6bmAfqI0yvUuw7HLCZADVw2cPz+HweZpXsu
KoE14U/rSfAhQBQJbiGk/yeh4J1xTeMJiCbgJW1O35FWWAfVJtmuWyvISvM1XoexcqKm44Z0magG
BQMT10zOUqxUqmvoZ8XCEAJWVMidoMQF8HuAh2WzxsavYokSbdwusGKCfqxPV9WPW/o4edwx8BP6
NB2mKFWDrA7xMKlvy0fc7KiXm/S1ljzJE+Bn3hQXCsDpbLkc9wkkHjUPpcGSDo1eBNEFD8SnhZky
U1OBzyv10MMs0Vsc87qC8yFeLXb8LYqDFNsmtxnOcKvWYzV7yOun8VLXWvl+mUiQTHgQeCcKh9J4
ujVHF5t5om+MRtNV8FJ38YzEScZF5VsEZCGspdEzOl5H5DfxOXHuKlQQhTgIVQ4U70uGRxyhZBF9
itb1HxROspHau5WEgBYbC1tjsh4O7cBO/sYKn6pUIJwuG9f1ozES8cQJIXCIAAr6nq+sXHxlF0/i
OikO6Z8dMx8ZyyPfqAwdo0Tr/yTdPgWzGH50EjMsLyfe0jh5YIw+k5yYnOp1avhHxGzWE7h25CuF
F8K5Jz6AAxHBUFVljszR/Cp0QizRPQmfzRwGm3CXMEmZ1KJVKLHa9YwTuctS7Tygq2TmY2s/7yDf
lKXHHGDlxvAD2WUXZpGZ0mbdlDfZ55fz+nWhyG75ZzkBW/HA0S66/w4uf+AE2/+Xmn6+S7R+G4Qr
Nz1iVR4C0PZ6h+VqaKJbHCaZ17qwubCO80k99hWPWmKPh9o3J8Vr9TlpYOmInS01e3PV77FPp3Kv
G/AWmC7q/IPUTjY9xGY0HgXubGfwmrDThoS8kdG0znguZWFO8NQDUPhpWJpwKW0Qg9HCMoiip32c
s0XZL1SRjEqyzT0WFv5ERAk+n4Lv7QThJPa/qQV6mnw+xIXxUgtdL5YOX7ulvsr4FUurRWsjysMG
BxPEaUU2SE4RuvsTM6Ofn4qNL39hPK3LfxzTnuOInGwt5vY/uEbl5H9OhEgUtK/0PLlzpghVBY+m
z6hCYQ+7rC6N1+GrVcBaKByFa0DVQVrPrC/LYBboaS2omqKvT9UpnrSkFEfyVy4yLW6MNlNJQUYL
JAM5Y7RQ6VsuRbVmoCa1Lo2F5+qq2GzNkygCk9cABOCle6MJLfV85FLyh4tXTsn60fz/5IaU4RzL
IXzMYB31q6Wy7VqMvAGCkvpWFhPI6e7WuAmHh/UeA3xa5ZAujZCAihR7yvX0N7dyhOw5iQhfyjLY
K901hyysQJglC3sBufmyJuafKiimyWNgSNk6Pelu9mb5SieLtPuQ5wxCIfNBIy7MulBnGQ8GuRzV
1CubAxej5KR6uqNwlLIa9Hmv9n44hr4aoNvVn55T58PWE0HLa8JRiOszd9L8I9s6g7KOqDtxK/q3
dGUx+YDEADDZ+75pRZI9zdmyc60kZKpeqgeY6VVwXQzEmW8oAiW0zSnsMfZGmJ3FhrpzOohRAvHD
JggUJ8OWZD0n851848C8evABa0z1kps0D4hqfT5glOHZSzVigLjVbpbbnKNlDlFPafXWwSdE4Bai
1rnbseIHzeJGZ8XgnSvkt5yAUGdsfPM8QAXSu47PLhjiiw3+K6tM6b6DCpeNsOqipD+nNPKRtkI2
Qzc2Y+WxsW6zZSPy4ONAa9qFIgVtykr6DyKaUYV9IE3MNWjRZgHOluqbfWRKFP7TcbmDo/2HXfB4
Wl6WYrdMlfIr66CRVHNUH2rutVG716KiAXvjZz4TSOTD7mqi68dDyVVq5CZJaQDWVWUJkMmABAPf
xDnigC6TXdmRArPtY7CWuBvmzFBJH++tvhqfuZMnCbLYmaIgegvBosYz7wujtgSKoH1PU1WqSlY5
LAVCMeguEkZRrRRq3b0adup/7kwTb3LhMt8gmr0m+K4qQ0csUnhNLmBEnAQcJhmy/GWJkYkjcFEh
jPkThM1utQYUpExFrFJpTAfsBa9JSQGJT2XiXt+vJ582xqD2mQjUpIBe/oMTYfMhbb2kSON8enAe
uPYsKWPmDhow4f9Dx+pYlLSvSEWdibyYHQwPY9L5lxQWJtHPmNSS0n9qlzrFSZuadzDaluq5PjXv
5Civjw6M4lPobpKmd/U8sa10AKUrjOB5y7PUNXIeJqPZumbnKRKWtqYHKS7EBgRGMRl1+ewf/1Kx
oo+XlEJRGAWygW4KJ5TLcNx54ezo/SlHjcekfV8mPhb4w3BkoPSA97nE9Sm+MdlXgy4VFcOsJYSm
wlltaIvzSoNS7NGHw0cDFwNRE/TzhRfmiats3cLtSma5N8PjzvEv3d19aLdfOuvS7DrRzuFQN1rc
1oCxZ96oOPmbegANqbebzG9AzoiTlZziRziLglI1nGx0/vtSGy2wZ2XlqLNJlKNrmv0Mt9AMQaw9
yfcVv8o07YiGSu6kHcbjhixCPgF0g4QHFiNNKyBxQ6h9K4/wpd3SJGz9AQqoDSfNV6hXYZJV3s9d
r0PlnTaJC+4sgp+4QSt50YS1oyTalDr19SPYEpLewQJgWTBCyhpCTBKvcjyMmGrDLWKC9xUZd7Qo
NYmQekQNwxDFmcF0zKvbJkxfzm0L0RKd9ZrUoKLrWWkqz6AJAEEhVvhAE05jYwzO45RV3CSSX/bu
Extn/GvhIUfEIspNSgPRpsh2gsgdeUgDyQha55GwdZxHNNE7bD1K9OXkL9Kb4+c096SMWJkA+kCc
/OIy0PfzMQIOAmoDwPTt4GYe/f5FYOXwWBcHk9MnUHRV3miAV8J3wUrKmmfGUcN8UmgOVFvbD4Ej
O9CdwKgUrnWgsJmXTp9cmWBekVfzob/fOZETw68fhFv5SrGqXhqgdyrAXP22HQ102Q+i2YqY5Ngg
lpJKvvgn0OeUHBTp6yokCQsjVGWBflhmts4VlmbyvKDx1XLTJUa2DRbaLNoW6UwbzQp7QmFVXduy
8oGRlxUGIHFjIJwgvC97UH9YUtmpeJTu+CAJR7vm1P/k5gtXGlntpnQ84Ei4CVmdeHKP96RScv/L
el5u+Uroz7JwCAi+OkkV33BPvjq1f6mtn6IFVgkcppixrN2K6FuSPYsfZJ8i4c27xB7TBspp6Goj
l1H63f3qUrnPhjYgdys1d+yvLAmJx9px8FNAHY0zfvqky6L+LQlYFwqpAYyOnPJW2QS7E5Y9uIuj
51o/4vihv0btZ1EYxjvmyrl8Ofs3+429TrmBwxhXGwCXK0CQ+5+p4GpaXciUW36eR6Dr8GPpK9Jv
ExksX8EyiamHhjRRx/QalNRUC2ReEPJxPtNZM/w2YXeSqvI14z1qNxeIbltEBDt6TV3u9W6aT9TO
tVSeniYdbHJAVCbEP5JTIV2wzFczr5sPCurO//VChOfGoJ79G44eZBDaJxXUJ2NKM45deWGbz1Io
sffjHydstUnHzzyjJRPEpjeiJwq5cG+30+UwJ+X3gCxS2tAGlT5H2TARH//fLSB+yEhoCRq0DLdE
xrglv6DHBK68LvChDC2XJGe/45l0nIbgcFWmDAoBtr/VJaveb6y65t1YsUPAqwxh/PS/6EtZJWpD
niFaLsJRiDGdl94LP+c/ZpFaymBQSHol+DnsUieu5o6jbdRiw7a3EHL+T9UuU1dsdIykuwgstEz8
42fPynAy5vi4XPtZDUKAx3y8Ykh9B2BfRy2Axm4kgfgEWry8Iav+nmDK93zx4EhmhkMwJdk+ATi1
U3QN5102YvcWXXQnB2HmbGIuDPymrJye4bnhI+HP7sjqV80abmtTkwP+mIrmKlm1FBJLz6nsAe2+
czMefaLeYWEhTnWgYCm55fTx/b405QIKaLaxDWL6C/VmMCkoGPLYGWb3vkT+04zYxKL/SQ0kj9ws
OoZlf3MSNM1JflxPELMowM6St58bigM6gptu9yBlHCJB125EeTNWLt/oJRdmqrgSfv+cK/3BXeDV
sYfBozxSdcJNMKo+e7Rhc/iT7eWmj7GIUHo5VZIpRfYS6DZilegpekw7aO4QLpP0vjxefeLVfuy0
kQLfnCMXAfyMuqkmYlJPTcjSeljsqlTItgQfVxbCpdWELNNdZiNd2VrMgcqj6b4WEq/er5qaTgh4
BiawCd4PDqtSxeLnTkBJgQ1l1yeRMt3DFiH0yIN3Tzg5v9Qfk9p2xzMtF7m09pEORP5LAvKktcBY
5+KAE4RcmMOxD0eR7ifBfHYE9jzs2baO2pkbAhrZ3YNNwBkY1aycrpdDtHbt3mffmu8QbbCmPC+b
QNz8z9lznWv5WdDKUjjpZ2C8eXu7ZM8neJhXYR9LPpihCeX8XH2HiiWsonOnsQ0S53zhuK0BfqEM
AEpUK9zxR+M+7bR1C7zCjhkEuDRwMLDF+d3fTVmwPHF3RPbN0hoe50P1YgzgFPZpLUpfLpkSbPIx
OsbJ55KaZwmp7UcEujUvoCf8OGrZ96KIhfv5JyWjeKE/f77O2t+SMvqVPuLoFiI94VUTXF66R4Ny
3D5PZ98IPK8Tb+u/6rjWRXaQSZYaZ0qoiIoZk5pMfPBwTxi2ubAERrscSI9CQ/THmpOUqZ8YxI5J
FPy8PG/qDxbFi0Ds+LN92PBlOHtT22LjQRU67W36l+lFFAcdPdkvHZKr+bvH6hCa+dIR5BZjPs49
1FVlKHuxlg36Dh1LI4MYsz0gQ8poiLNltTE1OEj+7pFe1omECXyJnK8hoxltLH7P0r1a6sGJ7kog
PhxNDm4MzxmtMdCdE4dUP11worH92Yi/dRkB1MI609f5sKaTwW9EQ5a8IfZxuI9WArMx1iDDRafC
le9LkXS9mugppDAovVO3JCm7uv9K+UzxUjAnCYI4zt8onyGFx112XB/WC9+sdOL7QzUaVKUJ5ZIv
kIITM4Ex5SiBOKtyyR1Xq7PoWv1Q6s2H5UByWpbVmkTtJMlqwKFYiIV05DwXUoZpDz0jNoX3Jwjc
266HNbr0R2yR+QaGkkgxzMMp9Rbmfytxki1Q/PrIPsFK6PkQ7FUBsgoiTjmJ6VMVIBlAXPv6+pIu
ubEcE6gRmHvjaxtqRO2HlIiCIMqxN+l2MFhIa1ChoG/MHKVayNuPpY9iOu3ntq5F77Chv6R8yCbm
hBWFjK/izzUdtQWpYFig3RTapSHoD7v0ZIIqUu5nGURjxqKKxdZCBwHzx3fQucrjrXKoh8d63wo/
dtdf7Fb2t8CF4AOMNNXVzod8/ofI2yyuesnxDbubB8CPAq6jPrXwh2SOevlpRQjR/8p8gB3VdnG7
DbSUfPQgFlUUY86GFGUvofmPR4o6FZM/c9yDzCdNSin1a4usH4IHG0D6hCPzWurEwj9PuUdxdOLF
MIPGsJmfU5+X50PieCOcbiCPaQlO+ta5JJY0foQ9C8qpigUYx7Y9AGfjaQubCfCgFLhZEgCSLttK
GioYQaiBQqKshj6CHvAojCTlwArgliQrd4TBs9vLFJgo7tV2tnWOY0tEgTqxkq1ZMev3vuWyrIvw
JHcVKLIEDQ8OjN3HZOb96FLGi2TVjpkFQ7be8d1aeC3gtV5W6eeoC+5LNW+W7VJFP75Z5r8vuo9m
W3cxjryEC4VTnc2VWwavA2Vz1z3P9pStM8vW19yBi6OKgz4fHMVVomDxNHWn61aZfbqS3TnjkA09
+jgHaLNBVSCCLr9r/+v+OAYpG+4wQSqgy0WnAWRJ3k9UMkJljdwVVRAl3EUBSm3xY1HBbyCZ9Xvt
OuKtg8cRnEHTzRi0E5F8i3nh42WhAEDAI0pLN6kqOuoCZRc/ZsQKph1jZTBsCxcIs7kzNlbu6aHQ
eCkA/QPNsa3xWtWeXVIlLJMaOhjbPFpMijc5txV7uBvIuyluSsPA6pE7M7r7+6+Tr3yTd4NDgmGI
ZebfqvhwuJTzy0QlHCwwi6UQ0m2xERZ7jaHqIsXyi2Qj1/akb4K2apPViBV0R6XtDGx6UylrbIgI
PSB6qUvWKdLJO9RRAh3SnTRHLluxImwREBpoIFnnl2MNvL3fIgp1E/Qsn3z/Npa4XvR5KJrjh1dL
H3VVMH2mwf/C1NidEAsb9ez3L7ChgHJcRhBTIkDww+94K22TkG05dzZsZSW+xD6rgwTR2ty4J6zD
2bQXl+GPpWsDSLL+vSappnXvAu4rrUGUQFwCPAxQgLcL4XOEIVFD6++MHR6WqzmuGQlIbeRQ4GBR
Spw5UOmm0O4txBdRMr+yeWhRYA9xOS+QQUOVVwrFIHDlHXx6S4nRxQShaJnZVhmnhb23tv/ekxcF
jgWzFe0uC53O0kLUvv6/7gPT4OCl5woa8z0YFu9BSCIopYMvMgQEiLngsN/CgAKm6BPEjaQZH+C1
Fs3UALD6G6fxCs8FmqEgYc2e8xQau9ikohFJWlj8tcUpPZ82dzahgZQHAm0w21+PX5eqyl9Q9U3P
xTqDL1fYr0HRBlYGYp67YCAjBtHp7E4UgSj+D/HGv3I49PNkIjNaKi5HrqOdDxSndnKosyI6d1lO
ZiX+2EQOBKn20oqCmlfBP3LEX50u5rQFK5BvtBKYRFLM/fdnvxKnvRkQS/NwXJarav/XKYgi1V/V
ApqeY9ed+r1RxJkf96DpMi3Lch+UbWsSOpamlU4K6uMHoqB0wNB0STK0wMohOuANPfHghAOoCJFG
iilRNyrs9o4hCIBNJwwE2UxxRanNFkx7XVED8hE5AspD8f1NOVCMfSg9Ye019USZoe3JAS3CAi4T
8uT3jGWWDy9gRL5MW2L8OEsQu0AoVIIblfDvyYvwnkNu4hIxDJmdA2XWPTCL74stbEwpWQsyUWqv
qaAhQPXd8baIM2MJsX5OQGdmwXqFK3UpePcCH50xhIuaJ7ehZBuYIXUCH7KJPppkAurFM1SXQC3u
RKgQ8Q3o5B+eFIfysghmr5du7Gpg00MFUCM5nyVw3uvm3uKWDqriqfKSBmKqgaoHEQEFP7z1PIdj
fX2+iC5do1UVNCI4FfBuYhwQN2kzUYkXsnAwG/uuOk8lqDWQXHjkinEyyGdVJ2tUfcI/NF8Kf8lK
PZI7NNw211SY+F2ILhcYwpfEsRoR20S/ZpavBBeA534Zeoaw3KJzn07p60aM6MY6suty3hg9KTVJ
R4yyLteFn/045Sxv8psgYNdLFPvW64S5gRuuuUNy6tvBtHOy3RotRVYQMKwdWkVy58laZ/+arERD
q1ZuGSiKxICsawBx/nLZYBWS+m6tDtD9SJXbOskouh4EzQg0SbNebWiSgCWCr9VxtlVdVFVloEdn
CiEEOxyQEmsaWCj99Y1YNgGc1UKGjGRLn07PU0LEpZZ08gILU83L//OSNCYNuR0R0EgaypqwLOoz
vTwXHIabQHtZBBU3AMAcDoJxac/3xGjgUZfuGIdNEQk2oG0pC39z2JqMiorfzZjfZadtkHRZ5zzX
gj7A1HHaUVGxqgpZfw+SSOewxuNR+FyiweUvKH3PgV4arg5GR0vaY9XXL3rMTWcXEdg4VlxwnRG0
BzWSjpaZ67GL2i/zR9a5nxTxVn18hMUTuy+FNRETVKsaI9nEf+jclk4IeiLTq2WmrpbbsgqapKhI
6OgkDGYuTMvhdcg0JAlHCAQOi/j87GbF0D5B8uopeGVipHoOzNhsHH3csETzgEzvnlZvdqSb5a1Z
IGGQNIAaSzqZ8tm3ndDOCOjoF+Kya8If/Ze8oZolmAB8Fv2SdRy/IMK89MfljiCpXundCr8nsDMr
FZxG/3p4Q0h7Do7A4L7czjHQ3yxh57UwBM/6yCQukh3aG6F7znqJymhhFa7ywhTtx/k61mRVUGAK
yzrIf5ExowGTL5M+JSjsDUDR2f3nygui2TuXaKtMhV3kOuHp1dhEFWaKFDwLcWxkVb6ZsW5J3Kpv
wdsg+d+oQWkbSBybHeaJqkNuoVFcmyctnvtKp7ChANn7PeEdoHiAIhdXtZgxMty6ZtUmpeY0ifSH
cZqtA8f16CtK/qz/Io63CCRb6SZTFAD+eDLOHFJHoZnlC9uioG3D8cfSzp1ia6Bxs01SjOpkMQrF
zMS/YOgi3iJ3Gc5E2EQ+7PGjx/0OpgQj5ks77XLffvrY1RQff+AX26CVoISMUmlu4B3FMf+YEk5g
ezJGp+nStpxAD2a0IhHLai5idbIQ7x0EvQFtPTyGMIitHh+SEb7ggjMcFTOzO8Fr1x/PZIw5TxXI
9Y9Z7ETQKLpetGEutAXphlPn3jrKwTHWD4FyenkqVnEdcQyCYpL2RI8+mYELqPrRO6nhBLJW29ZI
UrFUVu7ddc3xc1Jx0NNQ4CYr9zJQdff6CnQaEooTx+GgzYt5Kh8kytkLmam2yvtjhTGh6xw5Zy86
xhxSil/lggzFziQyEDtWO2HoYfa8fSme803c2ovC1U4Ba9mGE7XXGZb1tXcNqjcweE3UvA7L0PQU
qK2Fth2wAW33QkXE3tpyVRnkobtO97CdflGnR91O7z/vjZfLms++tNEbVzOGe3PYmlc8n51m9GG5
97DjOmY1KhYWVCznFDdWEWVfwgWaGXjOFekSOvK5Mb1HB2xXFMkcFRtBAGuM73TYtpTNg/tsmCXh
su4wqQIJXGP9a+Eodr6uX44RxE4hOXkquj+nhA6xB+OttUDb7dPuXVPr9WEHxws9sHzJsORD0sro
g2vytNrJNuGOuwnCSLaGrGU3tI5rcoVNDnuts+H7+PRuS/ZtjESuhPdZ6T/nNeJVA2gvJ19ymG+I
mJyYgAc1omlB2hRsT5bpb8T81kBntfpInsRMwSKOofUyGZbCSPaYiCWOzXzfrWYqp1Y8SagiJeLJ
QgEVUt7+G7LJDenq9XnL25niFspU+YbS7OaRJLA6GmrhbH7yKXBIo9gH0pCGur8K5br5wBlx6OF0
gYxewfw6McMqvsDLccv6q7tNGldL033XzJe4JGlb1Wh1TX/2Htv84sd1MtvPZ2c+MgZCVBOxYFGC
sFzD8WwbGoMvYmKZAahAOH63FWhDblzUYUZIVzFUT+bv80D6dKVNiEiZDm7l+PCgZb/kCNWgfJ0H
Qwsi2rjZUxqVOhHFFy3DspxCF7C7ANcMeK8WNYv88TwCVqNiarhCcKSoSWu2XM4aU9Cb71r4MELi
1VjoQe/apdcAIVpEYtiSzJ46zEyA/8g4KNRgh4kjJp2macBFypxix4TD7i6ItBgpIdq3W7zFwpWj
oRvUo5XTLM4msW6aoD27lV5ar4JMZPd4DrhZkHenLplOlw4uUNZO6XygN+6DdkFBz6nUPBbuKmC6
Svv5rEvF7Bg4XKE+BOiKD5Ey0jlaIDkB2pJDwuxnpyzr9Ppl9gqUmBrnQNomrcc5B7VYDsWlzuQh
sPB5DjodN8IxEztDiPq4YCKvpUOzOiPjOiyvsTPC0pR9KWlJyOX5yoWFVohDvzXQUyV81LWksurC
MR/TH3r6cLk4uLAjBq3wRX9niQkO/1aLft02yuJLbdGZFo3zXkAX40UQDGoaGFmTEHpolDeVvP6w
DZLbLb06ToLktyEzQJWc4vzzP97P85h9//30kPDMwfQS5sZnuSfLT7UWtqWLyk+L+opbajDLw8QH
3h9z5qdCYWPYlX9y5iBhvbG/u5Zx619XisfbL0Kla0sm+SGXdi4QKuTZFccBmTiNn1vE81fni2RO
MFJktb4wrfKif5SBJNQBdyrM/60ZoOZCay/pi9QH19qFY8Qn3jX5giWqJgRVqsio3MsSau8SNj/A
SXnWCuNU4l8l4ELNx1uvY0lvdYNcviPSsltW1fQgveoUJXNZu8FEhqxhSKMaCByfgk7i0AkRZIlB
rq+H5EeYnzsOXA5Jzsrm9KV6k4SPm1ckEspBIFMvvHKxZo5S8EI8yanPoafZtZszxBpqxxpP+4TZ
YrgrL+XpkuBuHCDacK/splHwns7G+7/YNvQpglsABbCVmToNj8NkGXqkJ78P66FQ7k5a7O5uAWB7
wAfyeY0rYpPEljRJeFAgBs2BR4eahizR7a8qQ9yhQsR83KHz2coAWO+ipMwM51zKRpqHMFVpTWXs
/TuquGhN4HhhTjiLIgTtD7MLRYfQNIVKRQkLRftRyXj+aGMaajGu7iPBFrunh8Jt8KDjR/TLnkAh
qTheJfPXKNbFVK1bkrGIenFAMzmx6D0Ix8qX7Jg+E/WD37YMF+VwpkobY9dJu2EcC/yMUWt8QU+Y
di4EBFKEFZ2SYZGHwTmmJx20PgZb40E2tK/70uAoKjcA5njiTab4Lc3u6xdieWbLcdo9cP0jhHyW
OFaWfNAwKz0VtBPhnYc55SaKb/dBvMdJ7dAyw1m4NM58Epdai+39b8mW2K1jTnSQKFiNUYJv51la
xRv9PXsN2pVOKJkJONx5Ba7qfMcu9C6Zuh6bcpUCYqpwaMa1UYYXXAf5pv+UltpPABWs2ZAQVsIp
pH48IBrxasCl3oOBmRnAG861BGD0nu/ZWzESuA2FZYdtQrara55dP8Uwp1z6mDFcmdLovnKzsH1p
N5DD04yjvNaJ4ylZAJQJ0aeoUjKWa4hKvsZYRyJ4bCnj0LMBighGzgH1AC6AVqN3LPhNNz1nlzUm
UUC5jNcJAMytXysXTCs+VgG8Aa74qejL3UjSGjgdd6O2O80EtyEacy5Xi+z0O8dAJFk4qAuFjYtS
vHCTYgFYpBVMTCHxwtBOkEAmFNyY8GpEzIfFDOUKWbDHf8379coRsNjOsQRlbDItSORbx6MQrXpv
+P5Rb6VSlZ9VwkCBcuA50YInwPu5ej6feaoX5yCDjUvKN7byyTb2f5oLWzwvDmcLULMRFSfzmgv8
K+ZXniE01VNz9W7eIrHN17QFTjtSlhN3x5UZ6LQfTy0biieNAKNWhaGtguC91eN4e0MQlbk66ZU8
xgqf4qZPGhARB/pD3W7m4n5TwqlwfxJojyToYZGO5WLEQRxyq4iV21N763Ajk/7m9sGigFCpPcg0
c2r+pIgoa/eVX7Io8neDeCqs1F/q1BBkYSwwAiGxTUYtjh7IgkZ79s8VHwxXTDyumBpNkX72mswl
etY0T+/RhEvAW/g42lv6AFUgegBNjO7O8YLhRzG7deOrZlxhcBo4OvPyfwdMgmFzXuSqwS3I9mOH
70ERIa21S9M4bwPvDaukS2juyBYhKrXUF02gVZQ2iuP9p8tHmpq+l4Iqa+nEgXAbX6Fx041nt0K8
QAWvyxBDEOqKUllo3jUasKwipngE+XpLhmk2ZNxOmk3w1IUTn5Ir1KkTcxL2cH4Z4j4KClUMEfbS
iodlG8z8Dj1jtPrIK8L/mQUtFxQKE/8I1glQoIsaSZVrvT3bMeW+4T8KStaWAU3ZGofVIIrJPCCH
X15varUn128GUlHNzcQ7Y+epBMgeMPdfHaC9qRw1Xhju8jgmAifLZtXza0mm5BAbHEO+lrf4pPbB
LSdbVDRHFPXDgcJ4acCqJke0sIcVgbndBdvmWEuxzK8Ebc9uA65XemG4QBbCHBw2tdwSZOeb20U6
jZLnMDRoGgh7lvADEu8OYhj9ld1xF/UaCqv10r6LmEZhQ9vzlxlPT+rq8wuWuezPqAd7pZDLt7gR
DYEWloduV3ej2an9kg/OlV4BASkh/pi93EIG/17oeTtk1qynmFMsa/w/RlGn3fpmnQ6eD1DqcVjk
Vzoy0lxoJ97T80NrWJMkEbLwAgOlMrO3r13Fs4AqBo5iqtLUIO6g7idDX1VGqqopszUkS+7l8sbC
4nFFfEJa4KM66XHy9O78NPMeH+yjqUHwB5aXu4A2mh9Qc3RDL0Qgd2pZYQnwQKNa/bfpL/1vzFz+
h6+OHIx0IgIoAFXed8G9/B4/sgypUzhRosMInuW0VeSKgWuMfsp2ZiOmIVvadCvrM/cskyDG/Nxz
2NHiXPlLcpUkuFuBe6tD8BwBoSdPvS1O6M8SkjyT3fAAlJLgzJG7iJhcwiyOlYg5Vsk9u0lpodr5
bEShw5qHZ81kGzq5jscn9tXYip8NrXCwPdzx3dpAEQ8qqJud4yNFNZMJ57L3U1VIUWI3Dwn4J/Vv
C7ykUL9zpy6XbGYLhBX0mKHRJR93dtwKasVszHf8pEXtokqo3zikGx466tkv+kemm2ZHQek3cf/v
bV/BdyuWowQVavR/XjgsZbmrg4WTR5PIHRe6UcblQkB/57cN1TRwNAP0BCNXNuHZ//dj1RTN5BPn
TS6m7MtMo3Ph9cRoGZBk2g420c0fXOFMz8lgCGaeOKqxhfLj53wlg05VfaTaR5K4QZ86UAwoEeaX
VbDHtFmWqE/T3LlbLLfbOHbXc/Z4PQVup6zYSrYU+0QGAwMfhHvg3B9HlS5UDegNbGxejKq+jC2U
rVQmEGbk9pfHgCIf5ie5qYFdX/pcA1xnkErhPdTZ2QTDYzv51XH/F8UT9zG5yFNhQLbjr1PPZS+e
Vty1zZTMSSfVIiYEtZf4TpMTtvH7f53B3p/8fNYNqtsmNhsAF0vWGCSBSpQ3zCgEJnOOp4coXFDj
nPYrBHAd8PcC+HXo7JhW9qbYlK+/J3rlwv9BBazZgGh6ewkE8iomus70AHahgv3yleaEB7heytgl
DccuHiGQnKYWcaWMNBf1adq+n2BpQX6qzfBGq/OX3+pH+rDN8nh6rncvrNgTItH34CbUfsK5/r27
HwYGtCUbxk52VWXbOkkhwbWu+XXFfpHC2l6o+h0Kf0ABGjgT/EEkDvbFiw+pzr/8K4soMPghlHGp
1LSJhYcTTHd/ZBMk73pZ1vXm0UWKfOWlsbnrnFORKRDiAtKzuPMkQLRPpGvhS7FVfJwnH9i9NO7S
yVTflP+uKQxNq0hrHrIau49R2Kt819DnmEjhP7qhfzcKDktN8FghROcFaGsUTsDDC8/1hJrl/1Wx
tT9S6IDSFvxESE6jK8S6rBwKPQsTieiCSrctSqVx+cSCfTnMUtl7hskQbOmP/+G6jjSYH7Rnwli6
VBp8ahmcuoINbOEdxPvT1VWRxWXq7sIxpdfRD6h5BmLicGcDUxgorXkfLKh4XX+6pTSEnU0sGXD/
p2RZHhMwsAvm0E28qC7LFUQs+X/ZGHWKhMrJqoXlJRAy5bscqUPPo/onLJch0mVrEoRg2iqIA34Q
QRsxwcDKHAYk/W+E6ULuUYuwXDBZd66xYi7XAawviG8bpK4a3EzUbuTFZASSleSmOf1jWU2wrzeN
4jM5l8mUBzhiDPXm9tLD9UbvkkipsaupObhR8n2Xd1nDDlfL2FngR6lbjHvhYo5LEI2Ka5Qcwo9X
h6n/lMMn2cMQDAIyTjmu+vYlorsnxQb4hV4A+cJZdVqzTQ2P78NOTf3nf9s/D1owobrZ3vT5StcG
x2VwuSc7dNIOvGqp8iIvjdHz8MBpF/lbNDakDWUPik5zkYUb9JrtGy9YWA9ZMiKLyLn1AdTTufMW
yhWY77pflEnS10q3UuTA/DBvp4o5P86zHihRaZdSt462FNFNKnloJ9cI8b3FtuGex0Tx8y5JJJaU
4/5gy6vLzUMtneDM/HVwv2f7V1Bm57rAJ02Ekw6dZF7fXr20iJhZvf/8O2aumyU84/Io0nPTN6iW
PiqFc3UMCqaRjAHmNaSH9lNLpNTcg5Il2JCW1D0Zsl7ZCMcGdmBrMuo18DSFm7Vv0TpT4cneqcYe
xI791J7mukDo2vKrlSEjo/OByOGSUlsvZ1vJ9n8DIqxyULiKInyDczNElltjrMYD/UvKV2LebRSz
KmKQT1Sj9Ic/BNIgrM4dL3L5US77AwyLI/ZYVVaW9f1Ldx4O9LQxXRX/QZ3PRUFGG0ekESxydCbL
8lVeaIy9m/pi4mkT9nWfATWebgYhi0UN02WozEFs683T39K9q1mGVBdw+3X2DCeU+vsZ2lVXxo9K
Gto5Uxbw+25+XpGBUPCzhM2hNZhNXa4HWtY25T3P6f5u9YEfnG/D82E06+BT/u1m4gh1Z+v/EV0o
iHgGL7+iWYmOkk1o2WJKUdXCSqRmvQYPw0yNhBWn6DkQMfFgPQpt7h2kzejxjjLrMQPCsICEqpkO
TGU4ZFIC05tLAtlIo1REiZp16T7hYbOWQCFwbDEdxourtf4UGhlqlNqW4Vv8MgZuL+YYn+3BJ2HE
/E1yRBeNdy0oR0vewwwNQFpv8DSrzCamfmn35/8kigkNaxr5ZvVYtEEm+mqM29SyHrTOfDy2bLI1
X9HwNPlGRSrtL8VtuxNGsrFDfKBwvW6d2oY9zenRW0u3tzwD/0ptJy6MeYCvK51YjBxNyOLpiW1P
Ylqt8hI6qVXGTBPtdK8dfPefB2iObXs0wfUhNU84Xwke9y5ofFUU2yJbTMBRo4Y1NSNJYUJs+yrG
OHtEYlkWCph2QUqMaYF7+Y4KCCw4uFgE5oCgAO9yay30A3riKmJw+7ym3WGK6ownuJuopUdNRSoT
GZ7fQDP+dWGwwCWuPXHhxpA1fN7SZAuVUG1jHjuDqQVLoqYH7RSVy7fAOltw9sbzXNmUHu8XTUR2
xVeUGgOocC97T9u2IJV9JCtgoZvEknp4dkywVL7IKVDbKDAMRq6v98rPj4XkRtLJLzxq0ew2OvAM
J3g44tWunofbylGH3tw7jvoznq/TClHxir9PmRc73fQoP3YK4ZMtQsB7ZiZa6bPEWTkJn1H91iYj
Lr6B4WdufLcmMIfQQ1eC3p5xsthmFgmtXIV9Y4jDUEcSKaUFjTY9hH2+XotG+Sw9p0mwJ+g9Xab6
8hK8CdQcq6oRn/1bV/UAP6cdUMj8HlIuGUvTXDGfxIgpeFy0jmLotptN+l5dgTiQFsIXAgBcxshY
akQfcFRNEl4nRb5T3mmEwZiUzPkk8zsilZLC0SLeNh9tvAdTN8EyfJTbzW85g3rvrFJB7OYbFzhv
hVGUAC8maIL4szDD2vwT2cVfqoJ8HJqbvxknvOYYsCc6SvrTBuipEyCCyauSD5idxDB/w7j197vW
4soak+ouMCB9WEf7xYQJsP9JOW1ky51GQX+NxsE/beX3p+To+ARmyKJKkxRPQ5o/B46EdhfZQo+G
dcBK+K3AmU4oKeH39vsW6JP5nYrmXj6jCIZCS5f26upd6pN9wuu+LgKelHWMB6gWwpkRYFjRKZKG
DW/XUoHhVBbL4AsckjCoBRkEyYE8/ZfbOzkfc6oGnBDnAs54Yxt7oA2INCwRlyq+fBTpVgFdN9r/
kS/mwErOTWkvyEQTkbviE/0rHyOZHcsYCyL82zXmeKKeYIyz6dBfnvapAzj/3qJFbtFRaiZCOXYv
MowtNlgrQA6DQB54gEvpun0tJc9jAO6zJ1N7t2WfulqDWxVfWdVl+gHh0lRVrRU3I1jXZFPiz0A3
QuD0r0K/LlQue6WpX76ADiJPqb8bgRIx6a8sbBnlC8JilxieMbBDypDX+zIbWqPyxTz73EumE+hV
QAbpkk7POn8Mz/pQKC6vKrwvRXkemQX6ypFf70/8k37/H2jybEiTZX/TYV6w1enkgp5y/tUR0Cf5
bQa9QAvHYVGgeznkbzGvDtlufsBNo2bye/LzGKN06O6S9WfJ+1OK/PRVIuvI5Ie0iqeGrL4VonX+
Tu9pUXABQI90bO55xerq2ZiHtC6//992g06J0oUhYsBUo9o1giAgMIC00rs2u7JEHgdyHTCmtSVk
Mf2GEa3xRvX2LkulToNUcpGECgDVxR0Ts/4UqRrP3WUre7pyKlUcSsoQztUOcc/EmnExxSfuNdw2
CMaCM+mD6zSn3+2DbcQoPrAAxtgptCAyjWgY4hVKkYp1bWu4ZiKdaLFofNCgeW4i1vdzNKF7eNJ8
x/K5OWAEHVWFiXo94DsJI8ttwb/Yr9dz6UH2Ez7iWUPm+ZU8pU1TA1zRCbPWgKBZUPg4ifvHPh2e
NwthG7UH14OxDxzjGGm0Ch9YxjzZE94UwyWLlC94j5edAaeGZ+s3NIfIIefP345xxCOeS3d+rpC1
sWBM8iEcne9CgN1Sf0eB8iJKmZv+cZ51A1f4nbKqPFIG2Kf1/2VZ+vuJMvf8W8XTDpxFgkmrNUeX
clXcpl1xTPki9RSkY9UE/J9itnU4/IfhbJ38hv31p1xy7zzTvJqeXxZAm8+xDmzn65sgRHd8CaYQ
9iOmBaB1qOPGXI0QdmkxyouStXTydRMnhQEE556TvrBvj3Pvcki9zGc5xSJDAN0YtrK0Ii0bunkT
Uu9wWekgTOopu8IpxHpfTkEaIoaL6iUdGaGx7STnj653VHXSXzs4lN9niE+bO3C87CXQ/lb9wLmg
fctt9ZOppKC42JSSy7CZ+7Ply6kAtHjy2u+Ica8x1JGi2rqkfvh0rf2DTEUeNW2k2sBQinPbKpXM
nI4/WykOc+mNuSbL3fSZvfw7V+kvsz5UYQqIS7gbummWWSlWbS6DvnS3Vz+uQx5VHcVmUGYg5c+U
Y+sCJYCXZhSnZhKarJOAxIgYMW9lDkEAtakTf+JhyBjuNSvNwsX1sOYQz3z+DlAzb5DdFVR2zqas
j4Dh5jxVlBWe3hUNPeOFBeA+F2DAxbn+cR7Vuqd5FvN9ZFzPYrCZKZic/b5+AgtRUbJrbYZVGEsK
eppixt8bmcRQXUTGS2Mg0GpJQZyFtJ7eD4AWHxyl87mDr7Tiv6VlR74aMUJrM9tfBYVSUq3QaPSR
WQeNVSdUGmuvLvxvbkA/7HG+jhEVu3c7zkcTZLorgezYP+TDxQX9r9O4b7snTaHI16fRXv9djD7P
TxtYchnVKRPSVpHmJOL1IjLKOqrOjxqlH2fMS1XrspPA3J1h0JySXF1W0f1FUQzqdRc9aSgLShFd
QfreY5CAG7mQjW0QXy7S1uxllzvx0V7r6vSbVU7Mls210CzJVCYtAFsG6qyHnpYh3mdQilWNHwqP
j3v9Uvo5sbbCQcFXnCDgHmxSr2a4RFZ8+3ERviojYlnYF5IcpNvOvskYmBoMJrZ+Qnxf/QEs8QNX
Q81xb4a73BG5SVpNdhlWiUNzniIUcByXDWfO/oZ8gbiAiUfveU9HRCR2BVR7ktqKMpobnjmOcvs4
WV/QIppXhrx2bAhUZmI+x3C1sZ2LnHFa4p/7v1VcZYw4plDTl5x6/OW8Rm1S4oqEFuyVzAivqtG3
CMHiobYDT6sxdilqDl0vhpQtWRnLUcjZrF+gNAbGPrAVA3+Q3uufHq4X6oH+3AF6mkM5yhmeaVpK
wljwWJVzvR525rO3nycH2l/dGnpx2B2i9/ItojvLAsiIDBV1iTvVEDU+6tHBzm4Bcw0fih6ijASi
QaDLc07BQzhtnmXshLyC9hMxSwKUtb3dlDNDbR+EYELvg0vJ3blmM4HuEh83jTaJ00q0DmBLryBV
hMsaWbGes+6twza9sa11E+JsRCSHPQpk0soxXI2bIWFgqufjaoBVlhWUzlecT5RADs4o5S0+DnJT
DWJ5mVYRRx5UMhZPnwGyzSYJacbXl3dTWXgp5ObnvvPnrjW9HUHsqY0G3lbCgsQmccgM7mE06hmQ
yVWHiXdH8sXKXX/FNIfR05sJ9nJp37qjKi1Fq0kOi5hhTHuO5+ggDJA49Y4JG8jnlxiY5z1h40CT
AaId/3XBLxEpCQs/r1ZP7Ml/S+we3qGKegtz80k0YRiEb/bEvI1TPXPVziVHt5xui4x2TgoFM7TS
RJLgkUXMuMeNRpovAzkaN3NYSL3a0jxWHG5pGsIcLNEgrSF/FY84ugpgwb6Hg0DneDuGldxZhGDh
ycsKmgayvDfReh45N+5rBtihNi+h9hAdIXi/9LR/tSfIwnC3bUeu5Ya+D8FH5UP/1DC54BHdhxFB
mBWUu7dv8PH9RvwUDSspcBiOQfy/4dgvebG3jzv1oY0ZOglzYsQIfsreNgGhm5lPQrnnDBQ5w3Ou
6nmraEdcQUD//n7aJstlDgskN/dta+L6i1XLDpluFPTGJx8W5o+hFXnPiyorBUcD6psT5CYm0JST
wZY+Ru9wQKUvpDamNXhqrbvOKaPPVpoFpZJ4AIxejR+rSTiEXi2bx4R+lcmPbl8zwYs/NiCmzbd+
490U4SGAMHg2DXPg3518dJh5VEfW5QbZD1YuGQt9k/2eYt3hO3nXlTKZxN686m2WCDYvomBIF8NZ
CFjFsgcVhXsQ6KG2d5Mka9f9/7oj87DfQfW4VcVyPd53lcvxjCiSxngnLg6PEBDqLXRdZGdSz95k
vKmpcNEcdIt4WctoKdzr/MKYiHZOIfHIj/pHfpj3J2srLZQ77wQgbIdLUpO0XozvEm85mjwzC+ki
nddqXMerwjQ9X9kT/Nfm1IJduUvGAhxrfg6mNvAujTkqTPydNbRbsUpoAWVMg3s8A7vmUei635Hf
G7Ugg4Tl0Ei46tc/YqJg+LmqTo2dgzDJfoppZ4/HEtpMidbLVWoUZPGADfQOadas6kqmOLpviQHA
5X+hsnXMGByMgMhfIQ9xdKS9WnotAVD71iAPdBmVMh1VUz7jd16UahYv94MiUbdHigrUJjpjZf/2
hSA+5JdG+ApaF9d+HQce+4KdhH7Xf1Vjvj7XuoODbrKgum3mN2dqMGT9/XTusUzlkWKeRGu+zmOI
KXK6u9qV5XxuNEFIeDQpr0607SKP2AtaZt6Nq4+6uWgJBbvD+fTxebkuekCLPe1JNtVpr8mIBhxH
Z9Km88kQaXoXq2r6P/a+HgZ8TkxasNc/n03u3Y1Y4F+VmnCCfyAYwLKH+nwHhHAgFHz5wl7omBhU
nq44YhaN39W72v+CfkCpWLI7Fd2NlSJ21XohY4cvvsOTcQg8KB/bOgVjLv5lP2HxCLzKGph0Ol+e
/AlsRV3cIa9pmGsYr/Czi9+xz1WtmtMRJFlENqShJsg47lFK1+TMZNb8ctG/JdK82RKOol9ISXCD
d7pwEwBm0hw2U47k9Q4NJG4TTeowHECJynX73T6nK+/N8q62BOyDa20R9Bkl7ZNrvkV3BWwmsYAr
4bo3Mbbr/TV3gpiV0PuKLTqmUV1FVX5WyXcVgFSj8k1XpbIKiHY/bRk1dvSKkp86HWzavpI7A+7e
uS5ALfyDloytq6kNEiYCtABViKGCkMAhkMbOo1C8b9qyY5lmr63vQ3kR59vkYKm05JaEVA6VAFmP
Zw0JUSlZ0kecQzrVM/dkexQc+3pofbcDbrsh27Ridz3mXq/KTonWy4XKO8PmsMfr0hjF5XpveLcL
i/eNHwqXwFDW3ux+gqLIq/ENOlDxvOdAIYESAnyTUEqcA7Dv4vUspwjBV+2tlMBQj5rLISx5hl0w
T9iinZIvgTQJzOhDhSEgfrGVoKO0fLLhF6A5ebZdwD2b4DEdIE3FyIPy+uNm68FXxhT1S+EPwWzx
c43nCLrmfKtjHTbuh9P13SLSp4a7uvhqTKViHnCC+S2uZHPE/iAhNSUh1MrOG16LhgjoA3Wmm5rG
XgsZ4+wHVBshv2b6I3AAc6G7r9NyXamQn7JInlImxezQH3tKTKVMpGJiEx5WPK40eFaiNHYkwfM4
03AMdhXoCJa+clQSwAHhm/eVnWT2qHPy7LgKfXNYmY8q3M+ksJjCXrmzy25o9Z86dZC0rQcZIve4
JUW3hQ1kOqsWCBSeOJGfiFL1sz4Ld7cdO2xUxhxGURpU7JMn+/5XVrjZ4a6aRBYXD4o2rXhDGpkv
Uhbzas4k+6gI59hpG3wepm9zQ3/ynKUN0F85P8679RBsOeV5hgdHcJ6u6L/aI5zLq3jPkqzH1KbC
BZwx4VYDTt8DojNU38usGC4kEdKR4mXfCmTF2YS21ZgRzV9OyPIqGdquKmyIvJy343dzyySY7+SM
CI9kKHNysQvPvbwihCMZ6lbhl0R3wuji9yaran1NRoHGu2MNyO/eEf++6RLdWL0qHID3C4JzBYkh
3PqzdlY11VOz2IqsDVR5wnAviezPXOgSp+5ieGa24s93i5bXJJxUCA4i6yH0w+EKOMjwPe1lk6k0
Ag+23+7j9Oe2WuZXnSgVd6zr1p2w2vTmdeCV+qHAaeq/6za1pCMea47S7F1GwUwTnptYH2nd/Dlm
VALWap8fL5GEQIXdQ8bcGrjB3Bx0hF3dWoyFwOlgKJ8fVOEa2P+njif8C3IJ9+Ql+9l6BvhK0/jF
qqtj37OExWIgO8WgklgAoM2QkmdzXY6dTsO1yUJc5UW12UWY5Y4ZH9068Vh1OQxfZstggHVLzzcO
GJi7NVvXhWmqmLXozFLFs7j+Zukj6xkQae/HLYJE7DmWdcEEcRS3xb+v0awxs/vT2FNyNSBX713i
6FRwOJ1+Jt8V6aSafYri4olqcscddfl++VXtlxQ4+nL+Ee01/VtuYQvQtoCCfhHmFTeJkf5R3jeA
CtmbF7NVUzE+wP7fhtvBixcdAkvdlQ1ZT6dI3ccUdgs2XCdqNHbkELULDX+dHERlQXF3et4c9yIK
C8Sfbd2yUS32gXWdDv2VpmhUGeVcsdma/b7IKYjHGvdIFrVSXYWD8US3OQTnmITCpBSbbpZ6RE+2
C1iGt6NkSNJEVsa05eVuksV8w13UzDNTMfgP7K9PZUspxFBJ6eYXGyaofaRNcNX/O2V8dsPiswy3
q4wsKnWye/ZvVnkmqsdYHP83yzmitVd+9M+aoQVrnsdv7C9va7WWXEvHCEQZrPYanOpf+uHAI3gj
gkfqDrhYBMxJhRfXSr3MKxvIJRgdHok/KysHn5Grl+KCTk6Nq89D5erd7Oo8Fti3F119tITjCAhl
JJ6LXQlYYkomF5T8h9ul6lVPqToA9aAID7wbuTVVPs9MbZzvyoSSeMSeNVZPBEwd5j0EC7NCSt0g
0eFb28jrONddN8x0tyRp83hwc6FyrT54J3RuUjuBzQuqiZW1ehwfAvlBIAUaeVWoMZvRsLx80eNy
/jCyy41XzWECjsjEqu1DeUNlJdPinZYVOgN+7Oz39YD7vrLTThaigoOvhsg+tQBqMAwBvyI4Ne32
fko+OLYQzyRlOMIKdOlywW1ZivsD3TFsDU9lmMqc36Hwb9KIzWMJ2jeeNu6P3a/xvHXyWu2VxFye
XWjEjrryOoL8YfpdfnzbPeFomHRaQoEp/RnNXWAlAJEJP4CUZruBRUXj/I6gOZxhZUHLtI1xZwCZ
CXh64EgWnu8e9TsV/rFAh7USEUHY6MbP9LYXeUd4WBDhf5alN1mZSpgAj5c1ebYa70URLIJLwkhq
V8EarShL9IOrM+mk007mlriRpzMDHxK8nBE96DnFSt36lzUfsiYjAQW3zbGyEVH5D9W8oSOdHKF5
cxKYJTeFjq8WCIKlPqO0XYeqxWF3HeMRJDmMZ+U4/puup5taH4yCJjgM9PS+CFXcfCEzJd/b1+Zf
AGFeYCPdf/ICJRVya0075fCMZ0szJo+0bMgmvmXXsEYa/RlVOuWuZY47qMWK03UFb+51CLfUZ7Ul
XK9wA5P9DVkE+R3LVuxwsalZ6DV/wu6iVz9+YHDZNeN+PRFphtC4BZEk6SKDs6qW8OpiXyPKmm5E
teJwQ1BzrRbV4A58AgI12o7VTmNfntEiITyd6Zutge5l0mp0Ljr30o1E9pii9Q1vSpajZmqHsGt3
U3kwizwCmpnDhrrcUZTt7umabKPgrFMLSWgNw4PpH+ZhqxtCW8O6uLyahTzO3PeLSdRGPT6kiZph
w1faSH34lRGZiG7gVOK3OSTDe+3f7T4P3AAo1Kb3gKr97dyhKIzs/+v8y0Tk64qDQiQP6N6f+X3b
xCphCpF6vaFAk/7HT6Ghwl0hcRa00q96QnE3v+8I8GOyvhW5ATLH79GzgFwldVD4Wkp7INEn2CWL
DTqpBvLw375rcjQq52LBDNO0uvEgAwE/+mQnsUPn3InY9UsdJhMx5DTNAoXgcy4v0+mYeUyJ4G3p
DbaQ3qlT2VenX6BScU9Aa6MRz7EyAibCRDD9Wx5dhYu33DV0SZpFS7dGA3tMzu9SF4z+y/c4M3+k
0A5/jVjsetDLLtbMtyAjG7/a4/zgLnVta6Omo+UzTBjqrk+dQVtgRbTlKVbs+0zPL1SgQKUtEIpn
KSVmVY3kxx4zvIe0XC9umHL53sMgG6Zf7yJT98HY+KiE1kbc+vGxFC5vDlC+xwFu+dgpBcex6ghS
B2jUEwNjszzJgeGXdTIIWXPsgE5nwUGySwhtkVIp4ol17J0QBYEOInAgnfEjr7cjpddMnsFnCYLT
7jXyIhn7M9tNfHfSFANyt6172K+pET2i1YmX2JfCYZZ/1numkcPt4E0FQS+ywlsTR3/+DX3zq3RY
n5NLYXE0JG98Npe9uat4fH5RwW9DGJOr8K/bhLoATPF/mjXXd7scrmDINlVwPDBljWlb2yWVtb7X
q8HTqiLev/8o+paNDajr+YXkev/GvIfmcWV8Z5QBDYLAvI4ZmnjDZt6DT972zHWOEQTSiS28rg/l
HHAbxqW5LOQqkLzvpjlfW7SWe3P7cPVUUnpgw5jFjf7pTf9DNADtxPc6GNdtMEfzJDMaz+qnYJLQ
F4hKRYywuT+dI84paqDxAde3gMpCvgUmQtbu21jVhWMZ9iYdpa1Gml0SLWsWs9+23iu7HRbL2b8g
8rSQ8d1aUlews7f08+UR24tEkHiJfSiGLkXzd/MKgr3oIEZNavaMmwdi11TY4t6WgK/pcirOIg0p
XPaNZbq0yS2dYgfYLretj3hUG/Idbafy2MYlfA633O0kqgmsYSlv+nzIwnzQo1EjBaAN7zV0Pj+S
dkcoNcFVZgP4zeIjfaUQ8rBfm6PsSRRii/QOTXm5Dd8ZG1eA9dvYubByrMdOSL/zMkJqEphYzB6G
Mc6WpeH+T/OMZuRWkrihuogXU+9znCh0UI5xtFUeIZR/MyZxjfb2zg4TcO/xurq3q9izw2GceB9b
GzE3Hv5zEuSoDY8+HX9G5Locmt7GWyycjo4ziU2ySieHaKM/i+oukU6bO/HGh7nMd5KlQ2K6ktbI
vRUcF406zGmsYApgJIO34rq9dGFZsKlGVoHpKSoK8tmUBJMoSO/KZowkzCgtQMWOljbUNi/F6S+R
YslNaoliWMaRHf+pMTLa++PVwH+tkOM6lfP8ah3SmmaaKaTV2ZCnbZ5ghtiKSkmyQj7fOcaDvD8K
rwO2vBGEyzwDNu1hEWUrlJPVdAKHMgub8lG4prz3IKdZ+2INScvcAxXK8TB99nijAxbaad1SQfBO
mQqgdOS/CD1oDyxfSuUdI+EZy9f41xCqunhhRM7dfYlU7vdkQ/KPa+I9OXkTARNCwKgKjFTFBYax
sMXo9Ym+XhbyvOR6lWwS+AJEEbOBKxm2Kuidp8b5NpHYKhyEkgLjvvanIzeEzu2yjwN34qbXhaqz
KO/txH3nN2C+uWIc3JjOt57qBA53nWL0PYOevVU0+2kWVSeCOzVLHwSJpI5rBYYI7StQAb76gAUE
9WXVvBFXPYppxWHiTCDwGD/k61lxOQEe1qJQi0Vv1VL4QrLaY41e7WkKC6DuAQwxUmA80PX/65Co
iTXQipaPG4CX/j4h6g0OvLqG6QpyklPC7XvEZAPwZU4HfTUdQ5Cq8rpvwVjQtWw5ZcX7PjPMCSoI
a7BTH7Yb+2AQNPZ3ayukb0s70qArlgtn8uJ8YEY3iJtZwRPJD2QsXa6piZInFwfotAvHqyzSIiBX
ASDYQd5zTKYYxfdzOp/EUM82fcf9kDWbLsFwk10rAW5G1Jb83l74ODJPQx8gOz5OP6OdFzuvmmi2
Yxv/f9l1lViRzs46ZsH+9vUvz683fCIChdIG0P7i9JaEjq9g/pJiEafvUDLe8tfL//ENPamL+zQT
cSnotwjsrliVG2QL4Ekfz/IC+eH485q2NE7SCYrIbSBzemxf9aMJwfIoHXaywyfCoa5MZA1dL90/
Gl+xAP2lbqFxa99rmz3Gm/2sYYUlK/FxQClGRSh4FvR4HkctRUCjJ6HqFQ/aeqDR0/o73KuyvUL6
ZVu9yuT/4BxbYuw3KNf2XCSP0E62MoUxXDbjEGVvB6G5KIX2ojjcXuOXX3suJv6tGHWI6QMJWA8K
Wraz9NbTcJhfs/Teaw8VD2OGu9waG7VOpJA/z2rr0w/6tgR0GWzmtSXaZVFTBrWxDUO9PzrTlwh+
DA4OyNAzMO2l6s/tspRE2qcU9DXCjIayKaSnZGUQNWHbsh7WSepvzOc9ZuBuongDc05amFQTa1x3
pDCMptxgUnPvrIS2hom8bdpfNmu+nhZfPJMSueRDggk9wguwbMN+JKxzkSdogbSeTjxpnRsw7lZ2
okn52N33WGaXhC0eCU9/CU13+sMGm/fhDwuGxA+/23WV3bXFXo2GB5rs7GQLIybZ/2nSPdfN5OR6
3XkzcLPOLJtvv//P232Ht+GTlcdaMc74oQ4FwApGhTYAv2gpgI95HxKPZeqWDGnMUn4x3+0F3fqI
39ts2vbuaG9CGkrb/WcVMuzMxxcwtYoKmANSyRik2sS8j17btI0YWStyduegHeaSIWOA3ytie8EK
ZHjjp49UXoxXbuo0GGds+ngQGHwFVmOidIhKvo+XD9vue8rg4zU0yVns4+/PdblRhV6LtMG7mfek
kpOEnRE/iGA4Yyjuwmh4u6upRf2pkrOCJUlt3vZmNpnmPV7GtXT9h+pF1fR+iDpoy/gUNqzR8+zh
pz1qkS7IO7fKD57Vdhm52HNmSVDU/obR3YMDbgp7iRJ6QMDSVFmQSB34U2knUJUNIQaHoNscZEiw
jxrWdUv3pAIoPZAI8B49oTwVCAivQB++Fy0WeO+IOJ5PSS7H+rnyfjeATUhg3nBGWr/tltAPjcTS
1fB6XiE3BGqqy1OhPQsCSH3KKacCHKC9BdNkTgi9/wfyLU8IIeFNVXRtsfO2xZorgY1+LxtuMY5Q
l2FcBLdFLm5aYFD923VJPT3XgfShBI2IR8HTFXUrVDj1LJvGEzLdLXZa024YDc6VFZCJMFtZp8J3
tRP6hhDOoTpReSO7fNvYKJMGQMMbeJ+Zv2f8MAT3oxLcESy2cgf3uORIYQqdF9nGy4PmL6UEPrpo
3yminkAtD1eHPlNyBJN+FzWQSbb5gJw3PiuP32Y63mCQAyWOXeKDd2DDKNv8qRyYRW5y6y/99s58
YYlnpZVjbmk+3HuACXiy3NnqOrCpjau/EF8j7hRhWSQRhaAaj40r6/km2mHlltVlzXJVp3DasNL3
1zYtvHT7aqZBM4tN7Dw5hPZ9ifSBY9V8F4I3a/vZ9gr8gLqY9/UWpjaQ50zNL6EOLPYPQqHTebv0
s6Q+/k80/0JQ1cSGGRjjhNFHbVDo5skN//ZujzN1ofO8kXMVBqPzvLKdln8bvWDegT7+I7MGUxhA
7t156v1gojFM3EWE8fOk+8UXViU6xx6DMUSP/pxvq6ewqKuyyOgRqnMKfOLGCRdD6Yh+0gAJ0T99
fRu69Ti7vB4EKlxTKIO5MGcI10pKRoGcu63ZxhsL3zcPdQVSPKfV8VwvGxy0z2afhvNRZS7fUmmL
oxCKTmwXtJbp7zOgArIBmSPTt9S4ZmkYvZsd5/O5SgoYP2anMq/3e/VG7OD6TtCP6XTKq7Bcn+qq
WrLvDsVL3D0OxPtwhoUFo4V77K8BDESiQiJuIGQxQSZkRVCTZeJiWFjApN8LgGZWGaKqwGOflzWB
BXKCQXEkD9tu+jJW8UPAq/eavXzoDmOQ6HqtAhs6ONLOA+78O+JByGBO1iF6WbeHbGjIWyBMkeoi
AxX0bHfdPNTVNf5HMyophT/5ZHyJtupNlQBB5+iC6M9t6rw7JsY6kUSUMLT+7YklJ2ydnsW6TVuw
+5/qO6xKXLop9hE7ujL2u2sepWlSWymIUUx84gx5CDAQSLBaUWkWuzwrwmT4dHY7Yrj19cKUudzH
5YOK5qiBGaarWtDhsgOuJlz8lprGFAXDLCcSRTLDfZfRIHqBYk4NVO4pU9wppFlxrZaAMVe00h2u
CHP2mw896SqiEBCccGTSpTfqCXO0HH4+GDqJ0ShRm+t8W93XJ9gjRJzbAP5bahFBq50WW6AxFPt4
LB/usbgmertTFwN2NjXj2mjOWN9Lk/ESazm2/Hsir3a/W+YL1NZtPTM2dit5xgBcNKq9jG7U/JWg
Lo3XrOPVcfGtsJ9Ne28qGuCryiKW4iwaHIlh+NCUkOdC9rqhILjJvqUVJgIRIapbxgRQZI4/C7+h
3H9hiuRaFxGPhBjE16L7WEhgdUyMpYlMH79XuRfVExfKYzqUanvVVJnqFA3silvfT7SVYppsk/8y
VAaJlKXcAKpG/OgKnfToEPmsbE8ZzQFpAxyDz2oB6Nrxd6eTM6I3DDKKNd3j/6gdpjDq2D2aG2cc
w2Rtu/FoMHaWzZONux5nO1fOpiY/tDaVfXp90t8ABO2T2M7GWcClOuOG9HiqCfqfCFfIRRT8gTVh
9Uz0gEJIUBpOYKAaQv12ffydJO8YmD6ymN7vo3ti1YQw+iYiQytj2m9KBs2e1GSmTumZ3nSHqqZ4
Y4bmnOO7Ra2UdsnxisRwV0PZWgdtDtZKc/YgpPoh7yGGVCfqUQmW+QZsNF7N5NPfERexzg+kkdRw
niI0oAWO1ofSW1JDF3SrZCTAbpFOj3tLYEDT6rPSwtV1ioYXIH133LE8MYNlV280rrFMrzTAW7rK
7gNxJMUh+YFgTneM4C2HnPK247I3sJ1ZeUCFXDsKmxCPlCfTnWTHtmxyx8tAZra5GBuZe2E1tSmB
SnZFq5ByQzFucZtm2bD0nTC9ghAcJAZRsqxp7T1J2OpG07fIJLx+JFuUe7m11XsvhWhH1QeAoCE6
CPuP/BcPT+VoftmwAMOfviCJethLtEB76gB1aKmLEvW/ykCFOTZPn/5OJ/uy3YP58SXzMwSL/bh3
NbetM8lpl7yOrCJNJof5Y0cW4WroF8VCplptwmuQEpLQPmBRqgxCUGScdl7xaTFuftL/CS8up5TB
Ws9RYQFh8iDcic/IWcpyn1wVqaYX/CSTJ315Pvfj8uYcl2qxiQOqRmIWOcHDRd/fJ0UJTh7v9wqB
8w07LKH5pr6vmQlq1nGyY0vobZ07xI+LI+Nlo2YEvoTWfJEFn0kH9tvmg6hQHhlKLrjPczfYlIdH
ZxUNkcwTREilZ6GdyBlBk7iRJYOA5XgEMem34s2IekqpmCL7oadpAw7fizXM2rG6nVssiMXJrr2X
6C63IDoZW9APSTIqu6cOVmh7zwgShmBRZpj4yDQ8cBEymzIkZ01hS8aKCxGrKFPKIF6lGfi7j2Fq
Jcbn8TFGD4si+00ONg+QdHcixaMkpLZxMOHXxNnFv8Ly2N3uKoCUgRBsPb9ZTMNN5QSJAUzLeBHd
UrrXH8d64Zq5hRTqf5rF1NK3pZP2ifnVrQGb8FjKu0QCVjR8uiyaOAn35fZCiHDtQBTXtRmEs5Tr
H0DF7FSzA9k4ST6qZ5MJDkgJXlKJvPC7TH6QLjlpNE47NoQUxTPtFNSTXIX1ByYP1liyBtOcGAK9
ThmCuNKRXDSmlWo3IdY63MNvDi0JhIhkEnsTVCjui0Ym+NVfaX0C4i2jDG7YmxEroUQbPQfGTBCH
5o85t2nk77YKX4zONKkK9I6h1BTtavYNY8I9cikU6H5kU4aOye8OC/BgKoeFcq4NNnZbINaVufsY
/T5nLXyvkvZC5dPuebzc8KISJjs0lvI6WAVmUNgWFuDtUpB5TShEX9XhvMB4oSeaB2nadQ9X1V5D
b2RIa7DjwV5eP6jpDn5Xr9Cg96tTrGO2WOlArAKXCzTjwWWau1s6IhALqVgPaRXLchlUcB9drsGL
tjRM+sOCsqbMONCPO0Xp8xbsgvyZq2i37XEiPqkvnoWoAtQVffC5frLxaBF4DWzB5y5wPyZakKNs
tIRgkd+dCDsiQmM0NI6lh7dyoeDuI6z7mqzawIJZVfeniZ0LHCS8AGqgRosIO2D+W10IxO+cqvw8
X1NhbAF0O2pPFzp8SYLZ7lR4ZWnK/rD3bOkbDBPUP9xdTAU3Satc/F6+QcU/XD+uc3KYEMcIV1Sv
JQYZsUh7ql6DHSkdnOE0bWnndmOH1znconxHZWOQK+DxusugObeekeziYB9P96MMY3vHKvx7rqN6
DZ00EuxWo3CqW3dWflPImjvy5L5R2m97H+3QPjxfDIMJNKdsudplJtPvkyBnmh6rE4HjIEFkLsrD
vSKDyxxz5UsrdQ7ExxwPmuvQ64V4ld44ko9kxvN83sZVDRo3HbTWZQwn4MNvpuXy+xGDp1fZqylM
8Uj1cxKGd6D6ZQCcUTNJimO0S6GaxUhFd5ILXOqR6Ek8Vk5dYeHHbdmjc/eGnKG4ot1c1ydolxDG
wIx0P93QsUBUI2eL1C1HE5U2AfWuI8XLO6Ddi36iWCzNhsNN5mnk40U7FpjWytu0GNkIYJzBDRQ/
rieqAkQbKwi4BKEHMsnZjNn/iXAtBAlrf+TU8lo7fLzAtRB8qOkZ+BXBa08iVft1P563GP1sfiJI
CifCUTglvUu5oBdGA5c75m1BTMA+LuIZFbEMZS44dPiu7toLD8vj+XWUNeznc9p0yWcj+M4Gahxz
qeAxYEarbbzsHp8czE6nOpw8M29rqhRbz9PuEdYfHVvKTDC5QiQLhF3/emcCrMOhhuW1Vp6SJsmN
3WqCIeJQiC57ekOv5BS8TaY21xVskigxXptNVPXm8A1v+z8kWTCrJWeB33/Fm2Sz3Vqmj6Rml6Y4
zS3iMVr629LNNs+r3FUck5KrhmactJmwMkHsP+Lcl4rIlTkAqws0CRFl+vsSTinemmCP+CRTp9+p
OQ2WgI+14buZylECGYIY5hDXUw7l9pUj9/xfr+NKPdww4ZGgWtiWf96apOUInNic3faufYfCUr9U
ZrPpfLErPPgVf2pC0IGuypI556AKMRZfwLd3EPTZKdqe2DyZD2jzpOL5FROJ9glk+csj00MfLEUg
JSfAoiiHSVzfRD8f0gNinD5VBsJRBVNuIYKOO9Ukfw3HCvjZaO4jHD5lEuODHQMaG7PFXkTGzTFI
QEGIMT5wfqWwmo5CAHdXTrFAojOfKV8sOYuc/gbmdCA+K3DLN+17IwbNe1EI+RL93vKpTdPigZYi
STnJrijFx9HPTWwW+uLRLnc2ytEYOLsg/0o/p0KA2JfYwqg4bi8eBy6CriI0pGTM7uttEcKblbJ3
KPUKEwcfl2aK75B+sFzFD7OonujP+NHuQLyAkraWDVZh81HwAtJ1Kspob7UycUjPZFS9FACxDdAI
UtP815MajW0/dIj1rFbdmGD7E0guBRAUeyOrN0saW2Mr/6kJ8Lz8zpCg3jCU9a/bCbBTrOdyEwkC
XaI89tjoewgfxcwI+X26yD2E652UfISF+s6sd4odhHd+6eCsX8qTBmzpS61MLur2qJoWxbdxArJ9
cbNwvDGvFlHW5yT3lEDQKwv9tLXhtYaAvpGd6vMRUgy5qvK3Tfqt/pg6V4GvzWQMJ7HuGA7UD7l/
tBlTmSM5jOb/WcrBlNsAmkLcjMu5aRL9n3wWfveBJ3Se3tYAkL3l4gwMP2Juvphz7h3AFNZHFf4b
PyLLp2Hnj69l2KWoeiGSkrOSzFT6tIBV63hWcHZ3cdOqsVG3aDx4EtRd4GhmoFfWIqVs0zd56VJQ
EBdZNq3lAsH1dJAgA2/0NMB4YdPNbt9xv4WypfPznUmLDW79oIgWE9pTAdwUp42Be5cq+2uVXcWo
9ItxMG9xjmuQZs7njwpjT9ZrFBhEOJkFd2GIuD/BbFgS/PXTeFqHpCWni3wEWgJiA7diIg1/OTvm
BuG4ajqA7nxCBENa8L9LXVLAyWiA5Vr4qVvv22Y8w2yzFLbqIyF5DjTsMS2lpvyQai4dMj2NFYCf
yOUB0Gak7BHIE/TG+uUpvvIw4NMlzItIybWDaR+Ozi4G+UYKKXYDoqYQtOBiWT7YNuZ4m76KIki9
v4m++ckRx9MwQs5eHbcLsr7jMevWyOx+4oITSNbGIt7XBlJL4clZTTrrvDvg92x9RX7twRDWOoL/
7OjJ525HpTuB79vinqCOVNefufYuprH2fy0yLfn6twSmW/jgRlV4eSuv+bf5G6uyj7tKSh4VId1v
d+8JtjT87glFd4+XAWghHSJA57rGvudt1VBxBjNRBYD5iLAedAogwjPcbIA8pfX9gPXoAX9YkOUQ
abaV6bpvoZo6pqzUtFKBrl1/x1Kdr6Y2gedT8NV924ecJDy1vx7e7idx2xIIAn694Tao7GzdwAua
SufZx9kuZ3Gj6qvdyyms48Yn7MZXce6ZWfd3Kf9Nn9pOGIfaalQmW/m6YcDhKWL+2zSSfoF2XQhu
67ap6kpXtcagLod2pdqwmHIoamHTAKW20iiOdrC6g9za18ntnVzyJXqsCzijpjD24oxzE7+Afd96
eMpv4OwB0LVxldGz0mtMTeYOTuh/0ZyvRkT7U0bnUGOUDQ600YBpCgUlvxcWB+axF2j0rlfxEjIG
D3ObdILn8S+o8wARqYY6JlnJjhk+AKe6VgZAd8OEJqitcKBp8pq5/bKve0g2kVnLmt+UEA3kdVHL
C9NuEVIAG/nqpY3QwAlNrrOBXVmiuc5WhmtecBYtGMJQJxhTfexZxGSBAzAiJWppDl/CZ+R8gqn0
n0jB+nOTpt7sVteaSC2HjYDgat0Dr9VkX05npDVfDa2yGc1MmrHb3VUi2EXAG0EIefgMsle+m0SE
4GeJEdoF384MMnigoi4uv73hk6/rlHSGRcoAhuvsX/5F4DxHsKRlTAkQbopnBQcnVL1aSHzxEFQ8
E53zTsMSDYTUmLtBYmCYjwfs8GQe74ilfgX5Sqkm/vbOFfrr2m41RVo7hAaX4Vm6sEPb37VsC48i
NcCa/oVLHkkm+qA/WSm6lEqKf/qCybTSUHR4cf2E+An4S0b0gbnpiUwym4gqjQXrQgT6UXCVnGBE
wPXG/xBbzmIeLVEf3Rjti7xX6l3FChTidrkETH9fUoqaffrSE2jn4U/wkGum5XLic32Y/+EuAn3n
f5KHSBkeWv6gMkY2vTlYjtBM2W3Pv1vS2gqe2eUcb/aXTmtu/qoOi9RlY4l/vMYpIbaZ3PzLABQe
lrr042OE4K5MEpXm9nerReQpfknph3nHKrtg53rl9NEeUyPXbM9qXLovb4MO1nhjCgpHVgmwtQPW
NvVepMrg1urxYRAFsskdFP9CXtRPOc4bPtNxhIRHZO8Vdy2UW+pqSbqzXTWPL/goX5G1zjVGwPgz
RtDYF4y+IgwTN3EBRZxYwsvRnnmyPZURyuajkED3aEf5Obqg7mTNNOhlY9HCXPEUATbiFGCihW+2
CndmFc5j7DD5E4PF2Rr0DVTovBfdBIUGZfnpHXJiFrHcaDe3CJsWi0N+PN1jCJuRPgPR9LmMq0Bn
wiFkkuajyKtboQwAy1KVrVSkD8Q5+xwtXT66jh+T9cWB7vi2glntkCzIlPS0aC0FSRXnPul2AxBw
UHVfAQ5vIW0jbm9UOdiJ2L9K1R/rwyxnYlS5sTknQhc0LPnvATez6cy3/A10EZpZjfoM7d2liWoG
nbTYHusWdij5CkVAETc5ikLCpaYtbXpiWpZbWA6HR5MgIgEkpUYKbxBuIDo5ihEo4FPcv21FfDUM
k+3ibWOWzNjNvagbCbJI0VHJkrDEf1i3jNHHLm8ATJdNhefNP8lKXr7yPdUv80ljMEbxsghFEJpt
jyDVFzWfnIV/gYz7WnjO+FigZJVr2cggUKS7ZhZMbqoGkMEaZYupkQd8OKULebNjSRKBpUOXujQx
z9id3gmkb/Sb0y4ekCLoCUC6TyKXDbegzvwysHcbO6ygTT+yePcPXLyEzlSLA0zO79GL5KGA8Mo6
MvvODCkX5Nylda6ycdpagvwJ6HeA0KJ1GuMAsZM8btb9WMp06ousVV7E4OfHzB4hQDgWz4WGdjst
gAfoLVvvprR+fieq7Nj5siTt1ddXo9GUGV8nBsfyohaIliKAnwSp0xxaEglrMvJYJHAUleXh8v0D
8KgBDK04DwKMnACaFAtNbNFQOtcbqYa2T1y+cvvjikb/25YY7ZE4CpncwcV7jWIU4QX7ASZFKLsp
sEqRlAez7UqY0hquNQdd+sw7qGSgOJNf3Kc1p6ntQ6MpbSGtkNGRJOjQT3PXeOTihrXGROWe1COP
fVlE6M/5J90yhCQMB2sglel24+oU3YbtlSZd3UHlfrJQVwZuHoVEe0D2FpTsaEg68Ql8oR8b/tmG
fnRVanxx+UT4+4T2rRVCmAsttDfc7ag5rMvLLvLYHu1P/7bngUwFrepk5DrQObUQF4hPpKsgBTCO
OGpyQiVkqqI4/qv5tT/A1gS2aox8HBl/HOqT3s24aA10WGjWqSGkoBrpy+EZAaGSHKghd6710NL8
fqDx/Kax5qOIp94IRj7kZolpnQYhkqVlR8bSn5VR7ykUZLeYUbKHgcXq7gbiH9VwAMbbau6Jm/YA
PhqST6Bkg77YVn6nF6HEysYVsQupadGXoUmRI4AkZyQyYSQ7DyplvGg8Lg0Hcd6OWvcmZ+gMxsHt
aPgNu+REYZgdhog18pnUcyQ0NxDrHW6EHmgrIKlA85/wNPKKg0dMT3rsvMeDbNdzVdD4HIS+vJEo
Ki/uMdSOy897SdfR420dVWur1cmbVUFXREitkdxg2ZhPtw6tsj+M4maxA+0LdsZ6reGRptCOzNrB
49yaEfncIYUozwMZ/VKCECSghnqffrhnq86kbox3oQNorbb8Zwon3DwpScmtACmkkwSALwRZRJie
fIZRSoMl58FX8H/SMJd9PuWPhIipe18C5tEsugXO0TnG2mvsQN95J87PEzg0ncDUsqzGEShr6eBS
ZjFFXpNs1IsP9KWy50av1BCiF7wb4yDsrqUNJfLAx8BOYHmB9vhKokbOSTdRt4aix9fxPaz7rtvJ
jFnMgHuwh5EL26N+FyVeaZrF7BU+nOaTABs+CbLRUQkrm1lMgWQe6WskNT5JaU9VCWNDrJphSfkS
w6of6syXLJy2I5lJhPBOv+OEN0nkmBoIXL2JRUY9d3OJsqs1voWNiFYdMU6LRvxnHmoumGjh/TIr
uR6r9gtYPsny6hoDMbPKfsZe75iqEnHvB+PuPUJroNfsO+HQ0B0cvMAJ1YgzDf6MhSW9E7fSyMw5
HUYwGnGCwF7JxsaRHF5bTvroNAbgrIrK7BhL6GkTXs8oF/4BHSfCC4v/rGNP0unhJwcY/CGZx0vB
Dm+9JPm2jpOC7IZtXmwybeSVbKYOCzeMVZ9S6vR1nBKS5PIGPkRrMYyihjZa6YNAznespM+YcMwJ
AG+Uy3t7loidWiI26bLFwq4RpuzhqGBRBFE0FRU1Mdtmm/AG3XJd017bjcC0x4f1pCk02hqkI6w/
WPV2+uXab+yqVJVCK0qUp+vK2wxCJzu7Yx1LHf6O1ZeNIGOQ4OMJaN7dmzSd0tSLSiGMClf/EcIP
tPcIEy6n5Ga6Jxam/vlk2kYitj/MxEJK2TTtgMLXOng/KQfhGhZjqHpt9dnms5/QewG2reEZzufh
JUy8LHfpjvf2qhTbYC0WfTHqfHRzROIsmvyilx9zcBweoDyNTpRQqGHiZuQEFTRawLD9p9h+Cnba
s6gjQCgGMpB0ONkT2HKotLpf4/LIuA8yKDa+pHXwmuVfKduZwpHlE9DS1yEfMwmcEcLBF8L3+MOo
DrYj/33IZtXAcQAI+fiBniPqyBw935DTpN3SDD2k4MzHOnt1r7DjLhRz1lq+bM682wnzDh/9cFUG
EV6sK795oEjN8kxNA2LmeGryCHouTxbarzzPs1j1JuJLo6bSE7NXcOjW+tY0MAGVqY6ToJLqbY1t
JwSFCRIZ3r/5TSr9Qtvnq9t8yRRmkl9QJJ5hhioIV6TqLntK61hmSUfYJasVeEnsKE7PsATr83J2
6D4GNrKLj34wf8OMlyDUEmawhyCNaRKaZTw12RIIXHOPGi/io+kHV17rUU8XV1C6MFzpOeR+0NUg
y48J1AKj0X98f86Yvoqr/S7IAhsCOr2MCROKRNvHuMIFxumcBYXwZsRfYFq6OYIYBWPygXHdzW9+
zBkgLX8QoLHgM64TiKOJHu12JyGXAbEbJ75lGlCtLlNrx/LqfI16rAisUGApnTWe+4+T2Z0ZqC1Q
/eVknPldxUajYnWcPjdn328U/60SR39v/vBoaPA+iWZn8onqN9TA/2/8lO3hiN0Dk1LzVWO1kJx/
ntXUNyxGo8ybkvIAhJ4P6Trkfi6BHKKTtPOwjeXT0+NNe64uv9orXxj2Bc+hQ8HkygiS7GNjkYMP
NHd1pG3NulXljUjaU4OvDHx1ZnXTriVkm94yH5BZcxHEzkMs6jU/yXBL3HwCpMjucfd/MFw03lrl
Lf1Hwgl+W5mSdMu2GnI8foTC1XemboYQdR47+8HL4d4BZ5XNXDBOSQVJLyTRPZvrV3HZ0J6xmLfW
z41L3MhkUi6bqretrQ2vWc9ol5hMYZ9wzHmqAdCQuqwSocOg4h1O05k6U5ho+bzTiJoxXFSkcF4T
zzhW7Enrq3wZnuroP46XNO5Mb2OB81a6+StG/+1NtdkJk7yDiAx7Tbs2UtpOsEbbKurLiQlmiPHo
wOEh8a9t1pUKkbstr71rOwVCLkj1Of6Vt+CLkVZ+UpLvWVqE4F/bFUFKH/xHBPOw4sxhmXBr3J0l
wWd5RSVAXWcV/DZ0KenIAXzxIKpgzR23SVuO+TBreARU5dmyc4QumQtXCs2qXm0t11DSRI7oZeOE
0CZLV3GHU+JNvfFCsivHnLrL9Byp1aUvGD1EN8UIG6mYTZ8zsEAI/T8pQQyxs8K8KsO0Dj7RMUF+
KIII6AEm7qAyb9obB5f+LCKgDTaVf6M/EvE5oBjLMdN+0TiZU2egRdbtTQ4I1tJQRf9yh9UdH8/m
6yYgwB2jO5h5fjTmi7zMqWQy4xzNeWJnn5jzdqi6jddyfLhaRxbNasGKZf4NAdyd3OZ6B1n4c42j
R9iNLMlAbFF4PT7ErI2cKyF6e94zkvMXw55JSrmVjM/cXVqsEs7CH6DLyx+v/PjcI6y84t0m/yqZ
Ehl89CU1nighMONnhTU6eQ53FhkpsFUa1rLcgkPC1w8k/Cby+j1pmasJOoBmjwTzO1CDqBBakvkR
uBsuV7YTvvPvLzKzYkc1QkDTTEF9Cu1nUvD5wWMom7xxCktiyIh7ciExLbtUFrYGRPzy+2H4QAlX
evOJ1ViVmokAdcD/gP81NFo45eyxv4/7ibbIRILziYJYMoE9SFSrIbU010l85NmyckCrE8qXcFFF
rpJkXwnvfl5KrSR0VYzwvTVmZnMLcvTEMUyDkSgvkKvJ3Uq2eRSv9rIRbREMAzqNVSjUhwCfhMfb
opw81lx5GH/jK+9TunzI5EMHWhl62AiU9wqAOhWt8zlDp8I16XjdcEm2UGRDh14Y6lh8KIh4dQuj
maX7kW4iKbWJ2nmYTUj0pN3yokpamumqneeEqk36Hn7Eixr9qa20iv788mafdcbUTVzspwfglYl6
EpnzNtQKtrES+u1TdwzRd3Mc0cHHcgmJQn5+lUC2nJLVvTj+oIj6BszZM7jVcxlqgaUKFAfj7EG9
rjE78pTZe8fT8i57e8EI0OktEra2ArqV/DBs2p/I6nkU2Kc1AF0ijhcO1s4v6Vf0NrIqf7niGvB3
NpirN/H6x41Hc2SbVGBjzJkiy3IGRHSg32tDzh38K/z79QqM2hamBjUVoHIWB3nDdAG0jHgl/j13
e5fGINrTY9JoJFl1/TiX1o1DGBKa8NQa7vs8w6kSZ62ie6WhX1hswun2RbdajUU+5Czs81cAfH1R
/B/0tFB821sVbwIlqYhpdQJZnPIVAPJaY9WS5FuZgUGceJROvLJlDc9SkrYNX98EkoOByaCvV796
mgDoxRSol7MEA5TVtfD4noB+8sg56DdUPBC8+7TjlMM/GdhJDZpYRdrHkHTXzS6HIzL9/TvQywbI
S83GsYtpWURuuyqDEba4ruJThdnwkdxXBNNejSxhlOpzeCwxu3TfsZwbN61CzZuaMfu30KSo87PE
LQbWO4G9hpnC9GP/mU0GrioAzdND9ITsM7yOF84ecPuv5y94SVkbN6prdTrtVlJyH2P/IgPJXAoy
iaCsajomn6RWu3IHd1QRQcIPcQA4lTbUgFFdFhf80b5GNExK/P3hwHHD+9j8O2ouZnFJnxR0QFg2
Ti8kSiLBkyJITDuruW6xVpn5AKPbG9gKuLvSiGflRvZ1mYk/kFw8PAPbotnB5u6NRNtOWemSsTz/
IDAYjBm4tXKPtUnvPw5iFwozunfsNZYxJVHDGwIZ9j6lnpVx6npYiOnYk6izJktp/S3AHyW+CGbg
ca/CbK5pJIfI5vlIdDsY3G4HHslnxV+G3WENf3NnzyNnKQJKkbjAcBIOv/VegqeZ18ThENGn4hXc
Zgf3VxPpAKLy930L+c0n5BPmDIbg/OoMCIdVYzFy0G5Q4PpIFr5xD0WN+rHTDiYw4dWJARxROKdp
wEYY1P88w9tSaMD5vkrcLWt8kB4YVTTPAqCoCtR0jyUfKQUdaW7IbDRXHVs23pnk5U2xLb/3j+CS
vQbV+d0teAh5IgrTxQnT5P1/fpY9lISTpiqxt8vMh7yoy2ihu9KyD7hO63u0cELOIpcV4je/wX7R
1PQpvFiBxjWW4ZUSdmC/26FHF15rYuOKxJDbfDpkxc3s+B01twucSz8ONTXDyuljA8rHRredPcJ3
KLhBK6iYcS24AwwClM4YrlFVSfnS2wvq5ecY76QuwjAWyMNiQZxMEfqwlHGuFNFTvyCiasVN7okS
6aNJCnHMaav+IIeX8Gu4FisoO2xRxp/AOPeTqCvX3b3aiv/jzCuBqnLh5y8Mx7kwSAEzDYeatms8
HRNZyMJ7huekNnH2JVYYZ8MqOfQQqF/+bFasXcqBYkzIGwHIipE1SZ+k/gtRUjQTs/mjow0vxgMG
BAJKS4LNnMejaxSL9tx6gzXQOfTvwX4qQH87ffb0aLR9DHlfjWWeYqoptF0zV8l7+pntnKIRsTLL
X9UQ45WbP80bvbYtT7XjeqO1D8goKEpZpLCVMdufS/xo3HtY7Zfiwse5M5JBaQqoBIaW/jSNijbF
TXOEFkRsrtZw9uEq20UlRqSypi1oK7q0sBL8dXXINq6Oj0u94Tesr5Lm3RwW7ZaUJnwdUWZjzah+
tCi8Ps42dn+jQ7I9czAL9gKyjYHV/ogK+A6bWCBFQOFEzzctO3iBOf57XYkVSp18SbgoYCTD0Qr0
c1jx7OLIumLxRpiQEygAsXPjoVGKN9vXffcAKAlXGgkgJ4L0J920Twb0dmWSEfu62xPY13ybryk9
TuWI2epQ8AzF03uMwIoUjCfG4pgMHkT4ZWKISYtMo5HeC1PTp30GuvxiHcUXMQ86COImpW4v+mH8
gLQXpRBx/6Ivej8fOLQe4qo8FhvBjn9iT0RL0FfeOVfk3zsFb61pGuRO/2O2t3s3nfe9tpR5SibB
GhMR8vw8D8L9mWCGiEurPg3J+7uRKwSM3ysQy63XdbUwIv4QZH6lzw9wNWXN/sQQ33jeY1WNxxT/
V//SEpSi90W3lA6481dtlofgFDDhT5aZuk4lDvm8EidFPLy3suIZhV3tvuRXDT2c+CQwebjbUvy0
ewXgxRX1U8dCfOKUXS57h5YtrGdD44nsdQsoJzlYP3pM9KjV9ICfXu7StDvqv6sZcr9XPmEsAef+
UHJ+/L2CKLAM1M+qGbk2EXkaTc5KrbgDtARM1WCgMHBYQMWrg/yGs4wX97dImuPelIxlTrp5lktG
6lzf0BuOx5hGBWw6o+x2LvkEPgTOQ0lHyiC9TtbbaIqe5ezP8qyolynMo5w1NiCR19X3nawPssMH
Pc+NLWaefGUld1J2ALEd5TjDTw/ffr+BjmKDFnf3S0tk0ixZ1s2V9h4n4EJmVXwTKGhOtInLX0fx
r2W9fjB8zNI+JIArUY7NmFqME0ht3W0wzGdY1J85gtRxy1UJijt0H8CKgLESbkmZWYnDuUXFw6aa
oFv3+Z40C8PUVm7cdubPPCkz1dLbHZUKKpfIGfZI6gn8XqWiJwI1APzxs2spbBH1OgzlYw5NQ1tU
8CGRqyk+mCTJ7/T6cjiN6CtF3ainuzNoFrnrIbRhTnyESNmmmBXzOgbauzWC/pYwNLi96lmSCjD4
xan0EmE7+/5kqWqzMrLrcBmEDvsxm9RMsbsNjibXgnL6u5PWdsxMBt3Cxe1zI0Wg0JwiExubCqsX
ifCjv7p/zukTs8YM+8g7h0VRb+1EuwmdPS3Oq9lDEzDtOr2mwhd8kqxQRSiiuH2GA+OMEKIz5G3Q
kakZWEGvwsZIxQ3ATPE6aNFiz9ZGP4ap8GTJymQ0qR2riJpz6FLVem0jQ31ZxItgupHVKyhiH1gO
YZDc0ujTrA6E90bJMmpnrFQWYbl+GniXKCA0OHQpHOh4P6ERkiYH+db81u3Xz8pQCovNaxLrn95j
nq+vhYNwEiVHlsq5w7imw0F+mdHTjosnNY+jk4s7ubEcwzolaWjLhc7Hq6wdtCBTh65lWkHMTXCb
Ga507r3ozvIoWYllk4yo7xjgLGAgLiCZE8RnngRWLF+wsLv4OOudI2GhnOsvMYMOuNAzwaL1A3uE
2BBr8nkl9XocZ29WX8pQ5CgK4H+K6brCXFrjTt784s99gr8Uc40RYWG9hEdpcImLIRxPv+m2fagN
MXNIp5LsyNFNtaLbezklEfYwLcODDSoRyKNNjTVYf4+80UlzT1tZ2QgcH0Us2uzJLTmw1rph6leH
uFxEra/CyoClECNLDc8Sq8EyZOggjxSWzAwaJhvmqqxBo9NmTenU0gwSjS/qhleBJTJlcR88toys
H2WP8zxlgrxLY/kVHvYHtrc/oTQXq9rnKBrIpQHKfD6cyAOvXb706rscbA733QIcOuOHs1k7klyW
ARk6M6DY/NqaGllYOjvs/zG+dMfQopQok1zTUyExhqSIaLFr230LzJZXpxvPLdkPtG55WCxZ8gde
oftISAoSfEV1HWPaz6v8LJBcQUkdGGBnnpS9h+lj3KSj76J1hw2RxK5yqDFfj6Ovixk9A7979ATd
tu/6qc6dWqBQ2IJ2Npe3SEcXe8e1lgwEoOm6j90cL5LJY3kg8irXUSoNAp0ZfQlliBohsZMfNU8z
Bz3qisYVxLQeRU522N3z0XFsSEiqWtbMdz1pzqv/kKmBU5s60jvdPg2DtQvkFug3bWjnc114sKQp
jzPlxmvXoo/vn4RUlQ+Tx7ZJ8WcSLd5DVZYxvC5qqyAEIoJczUvcribtJrpGxAmrK7kpYledCFKl
3LXEE7Z5d/ovjr2oPvzyw6eJOdOF5TPL6BUGYLWRRHxtHObwyCNBI5wCY1pNj2ZkfFtgAf15f1uJ
/BW+CywOlXcXxA92eRGZ6+wu0JrwIU/22/yHkcM949jm/aICwGfgR3zn0vggNN1iTPJz0fqC/c6C
yObOciXLUUJtjUxlMCUx+SUSfUb42Ycd4eQAusJOefni8lu0anjQ0ash78xvp94ytCsvLD4sroWz
FtbxHMcJdp1IrvUalsdcvSIh1MNo15dOfdi5ar2H5wFpvlHuJgZZokadee0Tu7bsESUtS1fvaayP
LkE+NVS+H35DozId6EUf8h+3JOmz1gpaixBKsdllJdU05Ac0/1ZSJa78obwkWiozhUBgW2mAjkpf
RH4pIv/XLzDucUPj2FTmzVAJDP00fPVLxxOmofb31aMbPuwCCM3It4ipEiBbtJuAqZbhLEj6JWhr
cwwq0+cn4U5UdgBshv+no9oGE/X4xPAsSNLOYkImQ7jOrD0gs1CWhs3r4S/HrKT5eV0gL4xbK8E3
08nWlSE+qEBTg9puNIGEFGUfUozhq4HGQHrihoqBU+W9n9LbOeUCIImEF8E9R+64PbxzBHOnp0JD
CXcyovK00q2ZkNkeItxTQNtaeeQJMb3gPDlhY4AkWIpiGqSVYS1WVEPcsxZixMHBkxJQ31+aDGrF
hLQsS+4cPvhRU6GiWAvAJlNhk1NzxesiPZZXEiEVwEIob8IZb+Mffk+Nf3GbLIke8NPgb4vn71cW
Kkx7DDPtwZM35mV/XaIXwXXM464seKz/q3FuDb3UInsEBds3vJ616id0Vi9IRVFlwmNPwnr/iAfF
zJm0hQPWBNitwEcWTu5x6koe6GAs3gpW7xAv9J+rwquFyld9nBV+R/FkLNi69av1cZIvI6fWnK1g
vmt6JEF+qMdz+BqpKVgzBYhWim19cMN0D/+trKjxljffqMx1e5DBy0ZYAPstwVJviWqvzR4SHh0Y
Gc2B8eufl/YT4edSG5iuEfQkyyL6aGK7RkKmd+EA4bYj5bHRnHwUM3oAsvjetUksaMh2g7K4xYtC
4zZixGXoX39CX9QbfodcfCjcZA9CKrCzCWcGSuKelmdLd4mpof4jT7gzTNCSQ2VQk0eKLrXY90tT
X6GeYUjPCmnd+w22LU1tsBecBBVIllSt3YIglwTazEi5odEOyXvm/DzRGVNBe4CQeOtJmsvB+Afl
ruhaRUhC3cEeN01aVpIbnMcIhhKP8xIvGHtk7axI4VxeR0lSZjJWF7EdeVyaG+mLPAnJz3rmW2Jh
Wv1P2fLrY9Sjd20YKnoSsgidPT9TbSpnHUI8whZSALOI0MwrYDc6wh6AtUInb6m6XvD71jkGOwhV
I/3jPiz6oTdU1m6GuOiRFvy7MmRQMDKD7ObbJQQXwfrWVAZdGp2sOcnmCtWk38bSlxAihz9iyqPF
/ag1+Ei4ovX9Ak92IwVfr7Hovf+gixfi8mkGyeGWZDhmiZ0YIliOBfNr6YtmoJVRZzdeAAU2SBwK
a49R7JH4U5VEKxBuHZ2mUny15CvudNgFUwkNLaeQgkR4OoORlsykWQ5zDW04lEYOidQckzzHBUrp
KvIxdkVt7N8eSV9P/avyngXu9X//2R+2WPwjWhuFn9QWNXTbIk2BmhFBS4lNZjDE+9usVT66Fr+h
6Aej86icfXg2CooCuVY1ESIKVZ9eFkqAQ3UicVp79nTZpeSKwUYqVffh3XFBAKqfYCLNKpASkx5V
Wwnv+++d/Miio1OUYI+CY16rltsb8lmpMeOwbxeq2olb5g9/YPUu8xImhYPNqmszqMJU1NdCm8a9
ezZ4iXh3wUwfDoClKD/6CpORWzQT8+YrMeQgn/uzqoM3R4+64tfCfw5n7k6Pw77gX9sh8ZLNIAcg
fwXSVavF2edcBCUaQWdCZ2HmqS69uTne39cMOK/IE6dx+cMfIhX4vrcOakka9HIRV/tf798GFvla
tgIiQll29sxcCkdDH26mbM//jwuuhgnbjr/hMXOL3A2NqvK6zKBktVCEmNQqp+nR1SRU6YA+cRlR
aPabpv7fNx+G+GpNdOzW4NcjG609jWGgZgngOFB0qJbh8oeNrM1YhHBZYhFosrvX2L+lN0UYplmC
eJd3BRKEa6FoS7O+GO1YDahO15ICWZJoYDk1FlmRnZT5ZOjGCbUHvmBmuYpfAlkR5JOLEkvrXLqp
k89kwTBHKb94o54obCVdKVHVkk+gWcees9pf7VG7sc1o4U+QDDgmnUMycLgp7QMJnBUw1czhpYcI
yCcfp5MmxCtW0QHcDdJm8kZSl3Ey0i6NQm6AdKCvqbWVJpRbLxHJWmGdI2M758Gq+qmUdlD6wqOI
m6Z3SncsLdUHmA035A+5JM+hk/0KcqBfHGmpAooAI9R27WzSmGV2wjsVSlcSyAIlMX3K/2kAmihJ
qXdaeatP6xqrsgZt/IMpD8QDPt/Jatq18jWRktfYXzn3rvr4dA73nihf9fMO3QBQeG7PPPq+HehQ
Oisu1F6KcnCNjWx1ilxA2RHnBejru96wBSXEEr38lP8FGV20Gc4+pyjV0nSfMi/SWdzWnoPtoOOg
YsKW89VMaurn5keUG24gPt4UoF2oZ5qGiQrIZUO7jPRdpUu9DhvHt/rQd91if5ih2QvmhFxyhqRU
Jniyt4+evEmrDNsBqyq240jm34IIDlmYO2XQg4Q9BjGblRDqsbgUBCbHWVE9/zuSAB8Zwmg73Opk
9IYQFLMYH2a+S/sFOVmn07lyvzvGN86NKLoUacBbstitpVOlAdDamDfZUeoHfJppjW/te6fxuaV9
tKW1nSOF1/1AMPH5hHNZhRGVNOTwPnk+HvbyJLRaK14gMz2DIziLwq8lpG6Tf6JVZhbohdFPMaHu
ry/0ILtYv6PTosAUvX/AwniliL2ScHoALaBtJafTKYVmQibGKkGsq9HpKK/zTnbnXZgmDkfM/Xr8
cr/zpm76kNcA0gACQKITAgfuOEgxD2LUZ+jRhrSUJ8JN5540eZuU/r7zk0mIXEaS/8GkhlDYC6uM
+cCzk5addmecf637Wc+WBwO5Co6WtKIa3PhjDhbRXmWvonc51x7Wg1gJIJNfwL5FMouLjF/BKBPE
PAsQXAE4VZ2/0rbEgQOzf4y98D44i3Dme+wODVn+HxdmY4lc3DWaFcbFrziw5gviLEGzd5a3Q6ao
ItU8rY2CcXEI8HkCbv1bob+lt9FliWd7DmEB0iDKXzOBKeeorPKHmso0ZaSNRHUVuXGvhs/0otqk
fLcDgIIrYCaKVYm097PWNjiT/ibCXMO5FJ26Zz3VP95BAXTxHMjE7G588LDTzrktXUY52lmhN/si
qFnusCUrD3wIX7JVbCT+ks+7fJzZVM8PuVOC44t9Qk+U6o34u4sdv1iIt//a3Xjf77e9NuleKVf1
hdcNsfPO5ggMzIkbmNz0v6WOPqw8Aeza6M8pf8PdO/fCGRYf+lqxMkazu2orx+a981xH1octMt23
ZnfxGXWx6/fFE2tdGTyMUpb8We3v7CpuJrA543Rz2JTX9HvID67oSM4I3CxKt755aMDPTi9EFusf
EflEfUlzqnEDlayLULpciIN/jpv9PgyyL1Ns6R2AS9g/9bjPB7g2bFqnX0AyO+/vCvmNvC1LLVnU
cSsoBgz6I/1fecykd2NhR91LjHwKNsoAbMtKtDgL5buy9Bf4mZD+EODdygv9r/kTPhpcQyCCzvY0
ZlOS9+5ulGMJktlFoNPsSwggWTEJRh5HHV1LO/8JD3EmvDHXrgUSzODXMT7UsNMfzadXWGgYi0FA
3fWHBBM23FlpQLmx1SdZCn6bmKpjaDvju33BEQcRXtwhpWoUJyX84ImRjCD+2ZuqNm5TB8VEMfFP
mdfWPayf7Egfg+kV5Ekcv56rWdgHMubeWkPmvfPWlFso6eFsbFpfpfTtqKx09r/R0AIqN5mrQNxr
MXXcV/3DduBLQXDU4+XnOMkFXY6oUJJ52jSJmNpEBXBdwhOc2cmmzhxj5WqXQ9VzF7LTVuHgEdDY
RopVmJEoZaHQiZxVm/DnhvCpWXwTIQCefmD2pKHDqCvXzdpQDAJ+ZndSfGh4GgCIKXyFjO94DHyF
JNNatb26xXEUsjhaQ1Flr3ICRoYYhxURe6AscahbjNJbrjWGZmU9+RyoyYLAPxHES+hEJ3zpgMyR
26bGfiUOtSQbfXzafXPkYmz3pZTGidJDiyR/um0zQtBLQfapjXcLlZQ/XOjQLB0b3DY4L7sbFB7c
S6b0sjSSj4GseSUoTEbWLLg/+7lnUBfvb2N9OWf1KBUeiE6NbBpjC6Jm5Cz+rEX2n7/qNpId9pGB
/aM0Py62lQ3S5cv608Mj3URa96QAk+02BGAuTQSbn5XidqizEdbNsyDy6sJLLYfmDLLKEt12LyAy
/lCys/QnkAJxxxCBgLkWFkG2vOjBbSr4ElOnurnQ3FMenTrh9IpQFaB13b7uJrf9IHtxIkhK+QLu
CBeRrhKsjO6CS6EgXOvfjUQORRFVEsShX2Q6fxTYknppCp7jLDqiRoVqOtyM34x/wmepbDFv2Rvz
kZWF5Sn+1OKWpFjyNsCOrNfE47KS3tOVYeSnmNJWi7jCOPzyuZs57+/lIiFSKaEDz/ICPufyi7P2
x9lY2xjqrOPII300+Bp8eNwGtrgimlDKIN83Yh3Ob6H9lRBRMpzZKTdlkMyrIl7AOilDVcSnYHSJ
aktFyXJPyyAj8QYcruHD9ICxKSl8Y8WYBX4xDWKk2L1FHY0CUQWhDOKzFzsSnE4rLHjN8LDEASe9
qQSyWkWRYtdSQL7eElmYTC5oTwBmQXLNJivX/dTkx6tsewYEjAdg4i91tAtPgUuowmYtHsFAV7Mq
76xgqSlnZp6Y7oaL6svAD1lIpm4vZZ9bghINlN9bj5jTZk5FK/Uzc3+zLkF/zgIj2ZddozcyiXV0
vqSSG8KeUk5YHgxoXfMk8xn7iO2lNOFUBEzUYIOO+5nO4PCUM9j6aQot7J2+/yU06aTU1grhzmKO
tAH8uAr9wP5hTLooMm4zlNvQh1bsuLmIZbSQRbsu7fKFA+rU+FD2JHCA0GDdgjwy338WdgzjS3ee
PhgZj0jEWtMP6lS9bmzzd+hwODxpycS1N+pqaUuOiDZJtjeMbhBDHm+lxAwuKU83Zf4hSdk9BY3S
0Du7hnUdAUFauqRR4FUfO8CyQNr63E0sd9KHYkphjPYKiJCzTfWoKHydXY4PsvQocC+sBOLDKAHD
8FR2a8ufPcqyc6/YTwBnYxEijOSulafdvYpNd8xZQ4W3Movv18AxyJnVqHdDWgUz8tg6ij93X1Cu
q5qEnjRzP4KOxCM4a/vBifkgH/D4FvcOs8bTNW9kRE2zG0qtNn0uHEPjSe3BcF4g0GOfwZ4Fekw2
C31aKIyw4MNeS6zxDGTxV5J8CVxckY3NH9xaMktDrK8F+jVHXnObuGV67w6s4TNCmSRUVTbtIlyf
Uw3P5zS1KroCrCEtEdQjDo5XToTnHi/LG7hOBTE5g8c3xnm0hdoyrQBQvIyaWEAvRpY0kTO3llLk
PihGYbCzB/ydTJemlklswwqKh7aQR0PY34g1zkRAcT3ItCpn4LOMeffO1FenQdLIN8ySm1lXK/xX
ySAPPCrVmaO1tpeiU1WTJiDW+dlaQfyk8KR5GoTZGiZnZoZGO2aDLxR5wOKl3Qg4INnzucpD3lPP
EId1yIF0J5F4GhREZdsOrWBzAc9KnTZYpJlxpqqfAarRK+RJy6LUii8ndhGdvLO5967KXMgVutE1
rWcPJiY4y57bWnLuFlLX0tjZMED9/G7Zo3IYx3mq2IPR16BYtOxMENHYdUmZ+EZxMR2wvy8rj7zf
r+6K7VdKzWpWdWpeNOu16DzX8AYFV/o4jBlmuMoWEEl6H3BqH7kuVYfJYlH6X2aAYfIipyl4XKB9
UWXfn9/bft2SQbNJ4pWOhYUKm3EplON3UlXibkRyRk19syli8gmboR0sEbLAZC4GJTNXU6y1l6r8
KEc/1jlRBAI85DUIVegFsZ81EzVpahtcL5GU82XH+j037ZlKfxt6XYumUnvJw6lF7oaxV7fTFR0g
7iASb6lPufd8gcdDdvOW2CxXdV624K29iA3OYKqP1++photmVfzZgLV1uM7pQFi9wK0B59Uq8JS/
yeaizve6J5K0u2gfBlKoefKy4zBExzb4LJCfmhZueOQzmOU4tfGA2PqsNz4BYD8FeDnbbuvPD1kE
vVr4lpdHX+cRID0+Iq20bbA/ZlfTNeGN+Nil1boQtZffQWHK+IR0zeADi8F1PLKAkakcW86Uu5rb
LRqzsY3s4Fg/wxEw4D9EJCMQWxBNyVzKWmuQsZKa+nOVbhYev6DT8eO2EFo0uCeEAA6pr6+O344o
Sua5+W7/I5FYBPKlEV8FhVJ7B7gV6ufXgkzEuoJKjGvxIMJT9H4gC4bGp4byS8QsFiROyxbXue6a
eQr1PG0HNHBogyAi7XN7YbXdkVpmV7CekH37BgeBeY0llHofqrRW28BERDlKAJyeF87+xq7cltrw
AoTHurG9Gi0Qy/5fUDZW5x+rEKdSm9Xj8eFOMd0ikNp7DYAj6b3iuJnc4s9V82IOoV/cRd6U4vjH
VL5I1jkgvQhwCVkmLRfA3dYjx+Cp0bA5eARACHsnhZPr8vZudhWn5xt5TuaqLXh45eYy+ug+Xlju
+5aE1ZxONSM5TTl5mdafyuV20FKF+XqLS/bk4sfy9fqon3ZmkJH368HDctG3TOSv38w99C15WjZK
ZnWBU0p1M15a37NM3WqTtrZw+9K1q6jsuPjWFjned2UoO2rFLIqm+9I3wCJLA/4/Q5fcx34EkpwB
Z/2ugqlB/5Z2pEvzRpZgFFtvs1YljgyZO9HaxJOX1t1wg+dEhqN1jSNdO1SbxPJ0i9Ep9qaT2KC/
ayKbjNTl6TvlIzVp04GdeIweyPqqm3qzWN7rivZ37auMK1lRChKTf8RI/XDlnrxs/QDm6oK1gyPK
Pv4kF1w6M6CvoQjn8irku2wEoiTHEAbPUbP8jdyp5UdBIq7bDMgw5wafExYya1cisVfJMPMotsFQ
eWVa6pwkpkc+Cc9+BBU/roTfPBMojJFT4+5bbynQJIrhlFIoOZ8VA4v6hIRJwMBDA/udrb6tdLL+
RDutw+2+Z86nevrhEds9TTv3ugps3BwATFK8qOzS5lmTyXeBb6FLh/BsVdWRjRh4zvqNymkcTNq4
N1Skq5v28WE3krO1gvlzMVaOQNrxQb0D9upK9TLrAvrzQez5EJ/hTXM9sZzl4OR2d79DZ5ximL7F
vXVUhPFK5lyZdserpMfECAeuLqaiSDa9PeLRPgvdzIgVkGfeRW5gD54+iAfNA76FEm6VlhDF9MfB
2hInggBWD15kyhv11JwhByAjLAQgnJj+ACw4TFS5Vgzjh7o6xlHLX2Eyy2MMQEyDJpzKSftSRhJ8
7jFLvoFYlRHytYxuGyb/oAGC7uGUZyywLUaG52V4WJtD50D+ahyeYqF9Dsn4ptPTRua596EovKiG
KO4MC8D0j7OGp1XwJ6qst0NJoUk4WzGVN7VQ4AgrrM2JyhL3cKeTpzFsCF2mEZA34nWKIPWSp9Ew
Ovu3anoUoTmmeSaoJYvPhG5T2ptZB58MTpoPLPdMmoBOlsdgmqfTKonOi6jYlGDXRLv7tXIx832c
bxNEPz1c7yjil4Hkne9IYvhnnwIeqk+UcVU8POi4QyuQdQbxnc/fkLPTwQvTOU32MWXb7cSBz/Qn
a2M+fho5/cLBuwNryLVyPocdll93b8/c8jSLtySZYrJ8crSOV0X9l1p4eG9I8pFztqGTmY5WqGIQ
EVHcxUf1/whbR2eEBYLYWwLVWtgNV5zTlUk1YjPMEc4XyG/Dm+Cm1lrOaYrPDV9Tr0F0k/vpKGeP
VQ25uGKjEGiAT8wAOwHPX3WbnK9Ah6B5nVFiyeg/xtl/1x3//wY/V0cM5yCDZrJ/KCPwg4nyq2HG
6g0M4L6vCr9obM6HDU2q2TVZjpcv5qAbqMdwMXGiMStBM7goWLGzSrZooDDaCp18wf6Ovh3TziCy
lEI8WfxqVUOzLG5n9GeBStJuX7MT9woxWLaEaQAt31v5X6XOkikhQo7k7QV/20nlskjeCbF9foxE
hH26wVqeLr53gjR2jeZreoV3h3V5qmgdeFNNLhud9WubYbU3I/mjDOI1imyW96rHjpfn1gawh+ut
un2SoS3IVCLkssEbEp7SrIII3dBbbyI4z/IxDe7DMrtrl0nc9EjZz4DjmjnwRxMm1GS04ZZ+Y9H5
eLU0KjnP2pnQx8GN85dndsk7FyeTPIO3lE6i/9MPgcXhpRRxnslgynY75Sxp7KZO0fO9NGY5DOwD
Sb4DODr8dsYFfiKYhPhCphW26GbwOd8x+NXqJvOzCJKkYjTBQZsKbUfN9ZZT6pp37wyfUaeQ2X9u
Wtg1bLXlP204xYJeg4RET/khs+MWNAcYRcQJGY5QP+BnqJ55GHhqfu8DCJlrgaDEM93ITFmpry2J
Je6mLmiF8kmlqY4MvZ+yuGIk5+Kc107CR027OI/cD6I8aoOhkCo3jNlyGzJxzFrlkqfBsvAUYGH0
WG7d/E+6HgwTzpVXRLshbiU6BbeqhxyOP7k48okyiyrv2m3PddGE74Nudpp5rvZyonSZVxpFTp4g
30Pig+Xp/zUPUNMPPro9RMwlwXZraxd2K0txvu9/9ipKVOrmCHEmdUsbQ8cBy8DoDYkcdSHJ/SMv
0RiLM9LRWRZhT3G3A65EUd5PaVinIL8rho+Bq2lGkbfVrWGGh3Xinpb54wYmXELGwgmh6j45NjrZ
XVMaoNzlaLx+QdopK2nwR3cXZSq+gJhVwU9zfPeMabUVDs+pMAphFuk10mgzrv/5oEYivEZJ0UJ1
/UKdJyiI0HEGj/a9cpPNUSHp8wrMgPm2O7pDS37sbwfJsXFHRJBWe35OU9AflRmzvmIUVT42YTPD
F339VxhDAF8tdg2DwNYvnTT9PeA8VVjnRqLjL2JHwwYfGLVsul7FbVi5XdYl3W1lz6jvfcebIJj8
KRCwJ3HJE6+Qjjr0qE63Sgf5PXA8xyh8l0xf5CEoUTKYduFnBbrG6No2qQ7WAMQAUhIt9CJa+NdU
RkZD208JQTm7NycfBPk9DHBZhM7wDatR+r+Fykj8NRArb0iTvXFNPIju4QvH5PucesqVZAw1feG5
NAq+pE8Xa1V4nWsxCxALuINDif5VrNJyv2M3Ysf11QOBYTUREZ9tpGo6FAU3JTJmFxD2j2WqYGUT
908UReIrpuWJlEsFdR0qVZ+9XOGfbmo4yww+L5DWTF3bKXlnzishV8NC2a8sb9dpLURLXu3KeF3j
eycpXFbNP0TZop/UVlehIX0XZxUNfIlTAQa9BHtLZXrEee5ffB/sDI/52L4ZYU/VYaM/OyLkMRb8
NUZPRlv6MAk7b5yTHWQ1F/neI0SIyjXOBDkvT9+Taxukf+LCG61yzx+dIf892cwNddzZs94J3OXP
u8XYPPP1BgnSDgni4zhGRMh9/CxL9i4qHtH74NcAPcsjD+ZWrc1MVmu324hD3Q0fEzlhfKJzYxMJ
d74peFeu3IRSp+LsCu28K4cwSr9fy66a0e4RAJKHUzmVAu3fbrrspfwROmDfU5541AKBIhNxcnYr
GrQ4HF20mAJCS6VBB1TaAHEPbZfplOtx/HOTp9oySwTthNnXBTUQwe00C7RbOHVrvVyCp5i2Eufy
iywv2PeuRs4gZwdld7rS8OSK8aZnhJ/wPCYnnrBsGuYZND0wSIlsLs4sbEau7mhjeuH7epJaNpfd
LdSNsyWxyEpmYoJJ9/Kd0AJTByyGe+UmUVyCpvFBSIig9zGIgYycEu77CfsvjNWiECV43YJ2lxW3
6BxOoFH++c3t+p9zr7I0Qd/oG60AA99ybzrlGvrXuGCqrfIYpz7CEUBy6dpda++B+IBHJU4vaba7
F32s/VzAglv+IYjWrHUiDsNTDvuzu2ofFIVAE7+viaspMkcTKlv6oayONZlzckWCSBb14qrasmtA
+fyyJnHAGJx59RH8atc1uod5PAv7c3Kelteytq+EdWnKNlSV5C4dAGFpxuMXfyquSfCSYWbKe8TJ
CiMnCNM3lbPrMvTiHaK9giQBj6VDRL+PbP/9Q/PLqjAtvPzM+G0z2ydgTU8xgiUM0DJJgVErLAai
g6h0bJKWJOapAwM3pqpNryYsQiUgtrttE1oDPGPBUDRHT3kA5UAL28nmHxHHG2w1oXtc5Qcl7ip5
vO/KJnUnvi7dKfqW1RFp2eE+0V7WeaU+7fTDZh8LuFl2zH3hHqXNKWHeDBXrNtybrrt+i4+D9tX2
zg1r81RwLJLWRFBjNdaeVML+vKt8zwP4PtA6Qrr3NkE2c+FhjvalO1gmAJDuSsK2SysSzAgbqQcM
LDA29CZ7r75U2SmR7pV6qjn+DAOl2YnEDqFuQdvYwQf72CJAVGLGJLcqyQft31MMs9vtubujKEpF
Zd3QLL2AXr8bOSPyEpmDcl/YHrz4GfDtWuw+L8OfBpIVJK0BJxfuL7vri/oje+9jFejaxmmL7BMg
JZPO6e/7L+u7zsOWcB8C6urcatJ/Bz3j2aiCPk+XFCln0nl+8pMcZMHiQhbkGhxneEyDHJmgex4y
nAm99MYol76++Zkj7l7xMfpz0uTfRyUBVm4ZvA8ArgrzpITqHzv5+8yCab0/HAqc4lrTFQsu9qcY
QKMUSX7FS3lhOUYaYO4hOhWhNDsoNV5zfH9Loss+vgD3gqgoRO8mlUesKKhIRVHfDrJVBfue8614
UTktNGwiLVMnGyvO9uSTH/zqysiAE2gxaUGFUl0F6wbzWpr1+hcKIC7bqboxFClYQVLefa8xbxtU
j9hrxX45rxF8eyGacVvnTQ0OE6H6CWHGW6P6rDG53fhHvvW0aQoRiDIY4aBrKzVk+gYnjEMNX/2v
kJu690ZsuQOCWAL8DEJUGCuNNh2ehU3SIOPUVVD5ui+kEljBYT9pplO1L+aWvxJ0dPu9Y9ovYtoU
FCRywRa/Q3XFkZgF/pRnfr1CpayETI8SJq9XjV93H6zJFq8yyrQQLwe/pmqjbcPtirx7vNbWKjPL
/Dr/jLAK4SOF6JmeHQtmUYc4qYFrdBO1en2IfuxvPxb1KxSjd1/INlg60BioB95fPMegA3nFVEZD
lX8dw/U/iIm4/xTmT1JFPhVd+7axEfOZ34k7mBzN5P084BPrmdXn0RXqRqwejdBytksyHHM7N7at
wjhwzwUz4VQXqu/S9ycXW+SY8EYIKYbzUxBCCjokhqGIm8IHw5DJPe4KFKK9EC9+UUW89t3XSW4O
/Q5B9EdeU4x/LQZj6s0mhOR6R2NuRV7SgRDRv8WMehBKiBbd8V09k6PKqlhpxSZYffoLK9fRTwyj
BJdTPClipd8Cx3XuPAPvfiMw/RVCMfJE8Hrx4rLvER9kAX0VCIC/vDwFjSeWRmAxmQ3P29QA1mIt
U8709NgJ0O8wcHqYITruu/LIHlckIjTfZ6CgjD3YRBY2EqJZfhlnMRc0kB6fZmWMAorvn5QATNGF
/Co7Bz8W7Nv0mVWkNY2g5wH1w1WRsZ6SN2O4EIVKVqfGJ1Z2a3uOrJ4xCj3QyLi9mWkf19AQGT/Q
NxqXBUSZ8Dhviee4Cfs5fept9IOBIt+ePauiyAwjmrr8yUCmBnfoyxe7H9H67BZVBSbIsN908Cza
k0mz5XQwV1m6GAFJaeAydLuH3HMPLdr6gkKxjtZLEtOXEzfOGZXJ14lZWzolS8/mEyR+mCt1Lp5H
Pu5cMRimGSHA4c423QrEF/VT7zbDCYEMxcLfdrqvpjHdST07r1SEN1qv+sPro9NaExT3GdoB7Rv8
l3GhuoiZGbpIUbrOaqkjNosG+q2ii15eDOXFOY+vXA/H/Onz58FM7njZ0bidDPGeffs7SuYEDhNF
Km5Y9UVWn3ShIwczwT1VBUdke5fBieoypGl67xtTzzy0k5UXfPxb4W/KYNLl+8qgw58ufaANzr4O
OVVmavSelcqZhfaFMppZUCxPJ3qt/yiVpv0IuNrOQMH3uwIHxmHKAcYxE/sJ5saCwCKvFtoloCBX
fOyJGgGuKRm+CDxonGT6MNtBE2h9/2mBaWHBYAbArLIZTCI6BF2CNPx94F2YEwlGQWt4460ZEBFX
IGT9PBas5WDSRAK9lzDl6/SkLm4KXvQX5VoxEIdg2iyS3ImslmbWNLtsFkF80wZ9SDy9YS8rc63F
6pNbYJNqJHXl/bciDEMn84vUVdTRlnz+4chBBlCyF4W2L2AkZ7vNYzDNKvT0W77I7fIVvEydKgAZ
tKNkVVgpsXMu1PohhWhqhbCdyMi78BAowuqUchpqd1+ONzFHsPIRhN3xNTOJOhZtFvyUvrCal/6R
ybp+siMq3i863SOtR8fb9KJvidyeVebMaa5Nt2keTEW0MpcM5x/BnUQqTJ9KdWFqHxCh23hio5uT
oIAvSvA8UMXgqGA8pYWgJIl2isY3Bq4dwJ4KgYgfgUE32esw4e5bNDtsKrOS0ILsel6CVjWihb7d
nLKoCN3O8ulNRApd7onlLIPzGg/VWg6y9AXPb07j63YtE7oJb3bvGZAdWH+iPAHDsm6kDmevnYYT
MOkXKmYE/pIpZx0ZfsnK0gLRPa6qt+rL0HsE65Y0ajgd12ORbWu70m6nZQ5ZGPiS2VwC21iTApjB
OwpHmmEy9XBgkXaphS+CjMA3H9WTpU0MUa2+Tv9lA5d3ACZasfBY/Dxq1WUat5nscaq30J6Bu+HC
2L/+mfk/9WywqCHc2j3kVbIGRaooQCZnRanVru0L1YVt5rqKizNmo6MbnnKaeOCzFbbxG/V981NV
JphDNru01V8XctJFOopz16LyGY9tI1sjS0qLqHyN29+Bm0iUCKiNmgJagvN+9ShVIxz83Ie4haSX
x0T2kv3y6ldKaEm+w0ES5Rt8aCKXRSW38J5ZpzEGkq+apkIqN/BMR9nt1076IvHgVgi1GZhcXWJf
2dT+0RoAPhxER3FRgPQbyV31FxOHqiZUXMXOdLuxoxyqPWtbxip3M+MN3n6+ewmESO8Vxd/2hihx
k2ZklXRckRGU8E7shUwB0RkKU27OarnTyj8c+f+cgWK0yNbfBtUR6W3LGRRcI7jViY2PiLZb+/of
CxF7st5xVUNBD+6qYUdh6jkOWfdh2D34Hp4jc6fOE2F75USVq2vH1VSdeSRq6KLu6yFM8/LxXq6f
rkh8ctjphJnK7AxVrb03nXPlPyRMjvbDQaJKUSkHlPIV0QPFkgRpbvkx8FLA94leEMZQ7pM2NieH
rJTY7bph03lGMkOlE73QUt4i64Q76DiHbS+dYUxi7nNzFf39JybV13XA8gdknXOFM0rCg+RroAdl
nJmsl/wf+HElo48gjKnxaXZN1q8VKkdx93uIHmqevTkoD6R+NkldK63i1XxGiOyfetT2VsqTlsaQ
VoLCnEpCvRj5ZVGp2303lIBsqjTvuEuGDWhLSuDXZ3hGV6/MQwniKrULNzyXCA1So0BWwkT0y/xq
RVu04OkJnZO013PbgLsD7vRPjpHv1zk4Gdw2JF76Oko8bFEmrFMHsQtt8BYGgMUdqxprTQbYLfMT
djBep+5iSsjycH5HrCVie3O7+Xp0GXy7B1HEDiaSLSK2s5ZB9bqaZ6j1qBLY5TOWdv9gfkAMiLNS
azQA8Fm1kiMjxPxsNCZzCVh/AA/eKFc2ulZdfFv1EEqJ8buiM0kDNU1eET3Me8y9QCBOLnpSSzQu
D54NP4IAWylHbXXzMKqywEUDWRAB7tALFCKQU4QyMbcvJMcWoxxu7KcpGJWRCY+PeopHcmq355RF
B7RRnVIDrSZ8zyHkftMljYixdJrYduHl4v6w8vmX4imFtpNqW796eCrDnCLJzr9KXvBaHp69K1EZ
gFXarnx/ylYdnyoR9BOhpoNdBnhukiYAjyv+LFTcv9Y9dLSNg3BS3T+WkhDou4mDk+u6psaKcXqm
pJaaccngPzXnKBeNh5l+nHS65CH3a0NuSVOtouPovhSpVTZxeXf/jNp77ig59pEV7VncdZqJEFGT
evILqICxdJAiD1ngGC1AjDPvVgZMvVn+PQBB6ZdFWQ6h+bF21vV83wMrbCNBBDHAwndLNgwixtDY
TV9DAWphnIhrRu3Xu5xOR0+tKv5NnioHiQgQDyXlTXWNNeN+1U0Um+ikc6ofJ+Eh2NDTubfd7/c0
pVBSsZTEF6XlrGpddNBjEl2sFbcN3vgmDuAW7dGC70LRSk6qPgSvocrItjHS7NCISYE1EJQEvNlM
KbHQidcFFGmHkNODJouoRylqboSwhJKVZSAn5Q/L1PyvHD+GJ2O3lOkeMq+FIWkrY3mzhJqlbw1V
iZFJ9Zw7XdrboiuSLHFE0TJ90etx4GhTk442GgNHsmz9muNN4wH1MsCLpi0ty79HAEDPzrWcMVL+
CCyS5ymCyMO4QTxqR+zsjV5uh80MOzWl6go4bBajvQOHO4cYd9Yf4BQxiqZS4Hm6wAd7IulCYvjZ
iH7c8z4gysh4taTkV+iBRMPnJf/ZUs9rWv2wCTMYFYexStJ/3yG8MubiwXgQxOJ96ulPRlwp2Ean
olklyiHRlJquoPbNHeQglisg7xU+Ozs3LeRbZug6N1RHKuD+ocVUxueLvO5xBpTkO4jDbS9NvbaR
b0QYjgqwYGnzbiM+rJgz47n1tec0rMb5Ajv8oGLY0poq1t8ATLXZkLIF02FUKFaSe8z21yMOLsiP
Z1NGN3038mECPJnuOfpR7LONpzjP5p2N5FR6hvjaYksrYO8MpMHxnV82/x8pZZls/oRxIV8aymGz
5iBzDlWMu506zEIP/POVeKncK+ejoGuCOULbMoPM7lyPW093meOLWAuXLRTwtQDRwMGkU4am8DEu
mGXrnR4C0kwjOBfYkZ+8oOI++Swy+D834tW61/hUJEOudD2UleH8VjIrG91IfRl6OaPnrcLeMO+i
eIyVeNsWZ9vmjAtGN2Wfmc5DLbhv0cBRlHIsfHSMyS7CuRAzzJXVtA5tiZuC61/BVDO2700FXyPm
BuxQiwqiI0m85MBiMM5wdxrBuoPnFPN2IjTstcMFULhYsYNYNUZFNr0DXfTCi2j5j57wzqwtOI1F
bISkP/Ys8mThYeQrbT8tI0YDsx9ex9ksYEi/TdNJa2sIQkCX9/BUq6X4Kk9Tz154wHwMT2h9iL0K
J4G0JM4A3foIlOwPQukuEfNx8O150tD1E7W27WqnegMd24hF52Ir0gL3N8MwIeoREY2d/4+sUpe+
P9b1lzpcLi1+xcm0ojqGpZimrPrE9JnPWmxq1tmiJOXagW9m3ef77GKBjKmZ9wDfJE+9Kc3Qe5Kq
qHxH1yho5rYQOVztE0t/CJlK6hY9KYpQ7E3ZAziQUQujkcUwDVettJOo6/gzxF2UyTLwoDQjHxne
5p6mvejIJzgcG2LZc0oUNrLef5ejCdYt6QpPa4B0DZtEM8K5m7FDjU5Ug0hF9nG6NwGlC56Ng2NI
yZcNWWb5qJCfaV+0Bky6rPpQjGsmxxkyK3ialByHVVOZE81ZlF0VEi/ruTMKobGFRH/jaCix8CLR
Zvrc8usHXaOxjaR979+t9/eLa0YPmTH4k7KF8zSstY6XV+KYTm0yHJZ89e9AknBSBZPlX84sj4Ih
aVn6i+ZvSsbjJiK/0qN4/A/gka2Cry0EZc70ehCtq0DTeGLPmLkgT6JBHBWiNyHFevk3ACIESVho
bmY1ZE951kqbItTfvdzlIR+XERgUDNoeeQp9/4UShnx9LlAsFcovWY6CA+i/Yk0R0Qgml/cwmQE9
cyLqcEl0DwRX6lAUj3b0DB28LIEQr5Z7OTS3rQ2Xto61a7LYwQEhUhcr3Lho5l9qXakw6i+cD1qU
mcI3lJxQ0kqWoENtofkDIxoGaL2pe3KI4AJ7kr1vKmRwwpSSmB1Th5C3hgrPEDBfVpBa8MJ7Th2e
+9hnEMDbqWX3Hpvyp696ZYT4ujaXL4KJkPtLcONnQ+y9sXO7Y/7LQg/OGClgUEmnfrObRu+4Fi7B
I/DqEBIZheM8Mdj8oPxqJ6k7reNC2cGkuwWZ6oNHtfF4E9JA2WAiVkuRv8ru8r80tNSdJyZEe8gq
Y1hbe9Dv6jhe/EPeGojKzFvnEeRFXTgq+Ve7ulJWpFbzivllaaK8yhszWiCjd7nNSI+0/kepN7OV
Lxlh6fmzGXBv6tk3VKMsDGHs7+LKQYsKVwE3HR4RZ7DjW6Gigj7d4plAAwAwB/SAPNWXZjAJBaa6
cjAaQo+SrpjRO5+q2o+hCct3RuEIrVyHFVhJ4JYlokU+NJgh3/KEYBp48MVddYWT10X/Zv/3pMkm
+wmKDB/MLJgebw3SPbAN8bQ2pcnR79Rea283HajIqyY8AdCEPb+tiAprkHie9AkjT++JPwnrXY8T
lpJKwJF49pEgO1GOpJQsTZ2yqDALov36n1GLTk+2SbEK9a+D1tiG0pzdY3CQpb52Oz2GLpQHnA/x
60hZkVQ4hk7Fo9uBugkkZVL2N3n8pgjVFT01Ys5gbJIRxKSOTvLx7ADE8bdmDHFJb6It/ZS1igUS
HcO0oywbpygGuTlVGpeXKw2yuozEljTQJYnEAVRxA8pEs7yfYUZ6ChUrzJvKUBPozJCUs2Mfx//L
dpsXoTxMJsu0QaVkNgl4aoR0Up30izoDwugR8vaRwOy0+OMVZs/AHhMr0DiLusa6sWZCZMCPjMZs
ymAbtCwvk8cODyxivvf1dMtB02yRKBUdBr9f2j9s5BmlSlbs8E+2saISsHkiLMlNHJfVLNiNBplM
I/aITUWm/y5wrgCgsewdGaPktkNZm9uZcsnSv2bDwONTpQP+5ScGMK9UHF7mSRnI8tNM4C5Lvv7t
YsczhN8ulgM5FkOYCCEzbsIKHtYJlulOKu2dIMF9RrB8129VX/Dv5DFRhQUjsLoNdTU38b/zTyJc
M4DtfOKt5eewEBHjmbcaB7vib9XVZmgdobQC7KLbeMRYQlkKyAW6dMF0CRSVXboS3/exZr4EeliQ
Y59DCsempTnk08DMITBBmLtfPwutbYkMpT41PMF2UOaRhjZ1JasB6WhjXUl3tOUMkVEWhWeTGfnQ
ui1sxxhxzhxY6c4YZDaSs5Gcb4OSyd7kj2DHa9sVpeeivaRXWa6qsnv1pesVF62fZTxU0/xmaTw8
T/d3nx9E1S8ucJrW3FNfUvlq6NQ3lexpqyyEmtwC/bWrI6R1GBWEKIGll/cM1XZ4fQjQ5/7rPSNY
Pcv+sddN/Fw8hXWIfWMKJWP8ubp5Z9uT9OST75UYbZJq8XUM1zGGHcJtez8Pk5FRZTXqYUPjCXG4
lj1RNnlHE30RPNOtmDzhrw07DCu29kz6C7T0u5z+ifH655b75kK9WtAqdUiwLxcaxLZ+nO3Z0HvQ
lMN8wL+KZC01UlvLNR8Hy1g+Hbub/LQ9sLxNXXIGqB2ZZftw59BW7fAAHEQBr6SBV0kUFog8bol5
mYO8jnIuoG9onTiVqDTxVd5m4CUJmzg0IzuypGe1h8IllruUxyWLSBx/DziCnQ9Y5MmmxFsrOcf+
SH7LwG0QrFtVC8Gl7cZeKVmybLZelvIsxUPtyoBXZNITVjMqwEx0WufBtKmkh+zWywVmfZYEDOya
/xkY4Rps+EiSE5Y8dVndkl9FKTkXH9gb6uKk3JisKUEuTxI0oknI1KGByEAsS6eaZktpMHTXuWfZ
atQyxu5U56zXRoTm8bErJNwDbvNLPSGm3ozzJ6KiSoR5QWHO8Kw1S4FLZOT0oM4l9WjZn7aXdp51
VOpvDQhwTygMw6lRTMct2pJqf6C1qpI2c2EulVx9lMQSr3Rsqq+voDwpdAQbBOiuIMWuaQWJCxRg
+BtDMNHTkZREUbGAwPSP3cXN7CPMS0YF1JAlT++eCka5nlHETE+xCJo1GYLLZlkW0tS8Pzxx1mAn
/v0IG0/1h0kPDkeqD1Ch4CiJe9d65z7aWMGsR/kjq10vnXlRVbCCA0RGgrsJARK3IS2jFhLP0aiF
cMS2MaMRM6Vftj3KV5t4RDOhKsNu9VZLIu77/St1m5FDnt2RJuqwXWpFChJcsv1wZ9yrq81xR4lD
GyVv//91kOhAzBHaPXIOwZMPMT/xuLkbanlbCr81kLZYq/HrQSOBLTYSeFGs8W3HGGofmkIO5tnN
NkYzsI8uQDYsLfgojo4NyTG+oRyEq35omUgO+dJMCy3O8IVUbAb9SvNB0Jz461IVuSfjjsIe+5I8
dBWWrWmHfqtJETIA2E35lTa1dI9N2gt7CbinL49RH49kw3mz6bT5KpoVoXtIGuS8x2ZNyO1jTeW2
RJlailjJWsvB7965TxcGzXQoI8JEBpydQIO+I/ZqrFJ6300nJre+Z5Njw9EAkKWDDpYGa8MOWF+Z
DJTiIMDX3sUhgqTSrecxtl9gFsfGiXN/TuvsSoAUVlkRFGBL0TJ7jcyl6KCzXoTaZ/Hp26L411tc
Ky5HBWeA6CuEKL1Fa9FYaPesGdWjf4L0RljJKusmydyUmKo55/mQX8o+Vzq1x4D6yFH98ruTDgYr
qBKKgN3xA8QRhpRcc6j6CNPoEhp73ToalIfHGIBZjU5IEeSbQZusFn0URCODovjH8Rwk5Qvoqvdz
VmdWi1Hb/PMqg1+ezDcwHlSCK3aM24hUUkXOb7Lqw3wW4kFJTb/3fQP0HnJZmeO7qalBGo6n3olP
C2RVQoTZGnPZ88caD3Z2Y6U4VH5cS9f50tu8dgBuPrCaGDCUrOwmM1lfcShdj4blyAxSJIPqbIrF
QO8f9V3TWj04s2+KsEWNyCMezbfDpiRfSMeczHrB74U/vyKwkRIkrpZxaiAfTT2zyjmXjQEszp3W
qqflIo1EqsA+84EkshOmu6k/4UV+k8lPf5nNaw/AyFo749chZeyVb3M6d1be99kuB/Vu+K1ZLrcG
7dqcsRf7aS6sMzITuEkZ1eFu9jFboskbQ7GlrDCJjWa50O01zHT9NGnDXZERTAGRIvhO+OwJ1YZZ
92ToZyXEl/YxrLNbB2SNyfIcWc3JL/UL/3R/8cI6CAFZ5FobcdZNqOCo2Y4lWNe+eRC3kmjBqT+B
YFoisZqx4lx9sv8Gk9NURs+5yLvkrWcmdsPaGYeSEm9KEDPZ1cuDprMdUFJ4e9KX2koUWmovGYo9
1BQFIAk2bNt1DyJCfdp+8b+hHuIXZpmJrqTBusoyAWXV9Sjp4YihBZQc1yKORGDnzC2AFo0m1Y+u
Qvec2VP+FzrxhFGa00uSkciNEFc0P+1vQ+6xWuhOIukYdTrhrzk2QMGyjTMlFBsDe19Rf07BOanI
fYxv6GcnGwiErZHrbPPfQEBcUf+xQsjcfpcjxbTYZ1Amxa+9IRWNI9Ls9P+ZN4ZVrKz7Eo/J1OWt
2gZ65sCo4hifZg0zEU3cMQXOals9vw3LTx2A40k0u1frE+MFU0mHdOwJFQ8LdDiFgNvT0wKT9a8U
xPhYDwMyBVY+skYInO97r10oLmGbtCdjO+FyBBwRN9Kc1WlatluEyhqlEJOd8NRf6Yvd4Nw5nbKq
LgOi0/gvkse3EPEKI6oJRCjvqkk4xcqmpQFO13RTXj6pG+tiqFrM60uHM3foRwUTWOjloavKCoKm
MHXVR+eyawitHcO72d2Mna7Zz8ayeDSNyf5PrOToFd4sPZVZ8okhGVkeVqVxN6vi1FhA6Rk1f020
c6y+YfnhML6y/ktyH5jqRJyU5k5c7DHwOOx8CKhrw9ylz2Z5EMO1O48EL1DCCsTG5EEeXqqnZ3NW
o3bOzGP8jrw+0L9Rz6CLTxSan3ub3FgIn3UTBCHojTwkRnbqhnG54U1VE0IS1XALaGk2yOmQK4E8
xURG0XcddEQw8o9e5DA4ZOKmIHghDaINQju3WmQpdRwvPwwSOUMzHMMULNaRcXNJuYBuA9MuGOH/
j97SWxY/2Ted4indvgeXSP1i4J7dk5ov9fvpUi+Y9DF/khdTmh8OKfpR2iS984TcYK0bdx/m73lF
CllgaCFlPz9XdI8wXsIn22UxNMSqXK3KNKGqtbLQNkXQuGOfQnc6Wt4UkzJG3EEH4SBm1QiWhcx5
MMQiG9YDYuMiSO+nKibf/tsKhYsZ8Fy/lUvxmA165VvyAGAkyrYwkYLVNxTnCJzE3luqwW5Oq+qW
0tIg3K41VfDWh0enhS3pENWbfBSWca/yXrj8KByTW8E1ss7kRWLgnp6n4RYN42xe51iXxZ8hT1+o
+X3kFWHyPnv76D4O1Mq1/XSrF5KuFYJP03vg6cTEH0otZ5CIPF5ZTm3QecO+DxIZnXJYjZU+iCGs
1ebAJpyqDTfHM1FcpGHT9uSLeoWC3rSZhggo1UXeUI/7UgsfWqWD3+WGC5QSTIsoLW0tAHs0hgfw
W8VziG8lE73syjzoBkM2TWwKWIGIVToL14Wk3suSdYoxEb4sMEQJ7Z/fABDvW8EtSbDFKjktonzt
1EM7fbwtLh0UMCiBmtkLi4J7CE3OigZ46P86wz+etCIN5WGKGQMvqp86EQuV2r6n6q+NI6lDPITx
tDz64CRS83o4IvG3iBpn3HUlbkqpnDigusot/ixUqe9bnR2VIFSOdZ6ouUGPLfX7Oj2R+cJRbkm0
1n2GykWfEhVP9VoNSHfZI2nP3sRwEfVwutM8XJSW67TnX+4ZFwzHuRa21YUbEfNaFWpnn0K6ZJHZ
TsfPT5cHXXXhfoq2fLV02lSm0rDZTCIM4ZYCApwqJoW3vAv4wOnFovjug/NBo36cjTnwXhmYigBN
V4+z8IvJPraoJtVKqkbofHgXh55YQvUJUNSftrgp93EscSiVgkZ/zuKMyGEW/0NKIYqaBYe7jwAA
7TeNrkMhLTb++eW+nU/JlcI+I/Jg4AyBy+b5qvaw9HGkPijrHyWcYYL4pdnjGcBH3AuL+bkpgHX9
476X0+xwO5g8ZBgsxhB9Xk+BJpIcyo9ajUGCNqwY2kTG/Wwp7XeJe6zkJtdptJjvyouaoBs2Xzue
KVnqyb1dmM4l3t12mgNOcPuCMNkgMJ8eP7yIVfilaYlYrKA7dIYyfkjrTUcOnECc7kNJPrvq+FRD
Yqo/2YlnXOb4AsU3yz9bZpJOc8dvfVayeWQsvsIzX53GMl0Yexux5bqK2XVFMnCG2JzfhVVnzPx+
ZqvKaP8942WBp7551z/1K12QKTtQpdNaCJ7Zvopa+2Gu5XE/MYNX1xebjnDtJSXiKPaY4JtXfwy/
F+A1zcuWPjVLbjMLrL2O8JExuSrF31+HKR7oxY44QhaaNOsrAz5iuHsB+QXX+hm9Coh0zxP7rt0B
7jOo3k2j32AuETJ39F1wiOfcYom8nPxSH0V2T8Inu5id6ZQ55kDygj+wtf8LZiLOm1wIBAQtwIlI
Nja3AzsPYkF8xkY7OVraBa4hdn4+LAA8C+7qiM6d3udysORKQeG9k4s+cgUpVZ5tZm0O+HA5ldBs
x5Gl8eIbZPnFM1Pg3F9i4Dij793tBgKMQmrNaf0guSnlxWonIaV+GE2YLlXz9K2lPEkokJF1n/ZA
V5OkWcMKfcThpiQV5dYk5uiky6QxcoHD9P2kL7q0H/LpCGOsSJpwkltSS06XHGHMtfnhZsDJ4HDs
lymVBBzvkSUZupQkfCkakYkuaZwxvFinzCv8QoyiWgTyN0V8wbBaGiLNYEfqyN/qu24wLJJIO9L1
azNUN2LGNpB/CUghrNFSlPS7ZWHBlNFeVMns88Y3vncRfDfhSn44vEEFz6nmD0gqfCUdp2Tv8m/i
NKa7THN9IzGjm0iHWXG6XDtQRBg4MA5CxxlN2qVIt0T2k1a2BRE2C5uWUhX/qf0YEz4XoAwzjRN7
Oo8cC0Z3O1bjlNtX4Gz9/FlAhnFdPlblWt4wxIYKzU2YvWpBb6OYD7CXX7dcaBEWXN/7dms24v8N
lIo+Rv3BHdiUv1kzLXyq2HVc8GLSLuKk1bsxlNB8QQ+OxPAuYfOxY55oWkp94pMxBLunneJqapr9
NkOUYQ9wE+tOAbSruLXp0qKcEUqmoM7+juTGfAej/Z2Tn9g8tiyfSD8BljRnIawVe68HjuU2p6j5
qjtS+/72QX3mXcPhTcI2HEAM/ZkCceTkYefzI9s36Ofs2SIWFGUr8Z/OBPxt8twvIEjtK76SrbiQ
oHQhfsi6onGKdCrli7akifPK3bI03D3De4LrQiy+m3c2XWz1C/f/r9TRSlnyPqqjqUbwO09OFSP1
sVxkSGjJBv8aAwvR2gyAy8UeQeoqs63yLZfV6pnj9+wIFZylipqPDR+ukq9D/oiiVHQJYDQs7y26
PLqgiB0OVBhOhx/YBNy5L1C6VdbOmJcJqTNtljm6nVpqrSNCWoxY8CKlEsPW0PUovOUB9g22EwsY
fiDfC1MAoDU9QiwWLGB3kjxbjpuUuD4rnnw6ZhpR5mzNn9kWfvwxQ60jNG6fhp9Wza/YsJugo7Au
h+a7MCbAJMD50c2Stw2vS7KdgyWwP1UJdLvxEJNT5oTrGlpM1z2SfXiqhkiVLDgMiJNtJLRDeSeJ
gqJx6up3S/c8EDIbDNcc9i0ns71Isy3r6q5cWxUrEXtApDLqPeoMD9kcNnNIs97/b7BiP4Rt29mI
9Ku+iShyc4zCu9Ch5ev502LMWw84qiKCgJPiY48Nu6/gqVFtDHfXJgCxUyp93TD5uJiUMxTF1gKH
upuQwUF+STm3r+6WBnqEUJomulQDH9n7wDMH2fxO5+1grUptpxifjjHAKgb+7sLaUYQLwPx5XYP6
86Jhm7B47Z8wE5beMdJOqLpOuwFUWfQpOPvM5uZGHSqewBVaSWWo5NT3/9UoaVaS7/kZwl3invQF
BXHuVw4n+CQ0WNFjwrH6IbIPMdTZdkavhXRjsbPRaDU44IRgobSjDamc9nHPf3mJfSWlI9go+Oy9
cNBk133HtMKn+Cr80MrDKRZYKZnCipRfNi1SdOIHEGyI6PL5Z2Jb2Sb81KQVub3U1qP9K6WCOue8
iLfxmS3DgQiCrAv2+kSNQWUkhCbnwrsNgOxwMLt4YVSxFtZa0Gq7Zdg9inCgrmJW0jpOBcNNQBVu
DCyDfTpIPuDTK5F42XDWGyQgqArbKuJNYVW8SoOycaW5W8ZJDJ61JqbpokXWnBW+my2ivnwj6wC8
M+rZhEgdmW3BzXTm77YV0Au84i7SujVH+XkfVwJ0jnyNMoVo8kDEy0pbNfnu92qDPyyGjzq3B6/A
1GUQJ3WXY1UTEjB7EkHYlkAIsCNaBqc9nEd0u0HbirlavdzvTkKYC4/uPMZWOyia0RvYj8KUltq8
AfjO72udFoXoK+mRJ8PTieACS4yTaRXN9imDDzNgGQo95HFeeVh78HvAUoxO6hs+TzFkSC9WsHCj
11MjdLAIkE/+sh6ceYQmX5ARUbc1XT2rU6dE5CPo+4Q5lZcYfXm+ugaO7m+0/pxV2GZ6RYInivpq
kuMW13TKgugxyvPizi/7dVCZ5SDXTpiX9fsqcvlUPcEFqqkxvOY/cDJXfonXCnGrX17/YfLCMlFx
zUMB+VbwUh2V2z/GK2ESkp8dSLixvCHzSRP4zTTQ5xVkDKHRGuMJFaCWBP8KKo/A2yH7D0UQ2+Pj
IQv00o4MueI53YbRU7EJ2rp4CofYwVFAS7I45whnD+mnnIkjnQfuaUVcgZ8tg/fkP0g+O0iU5wma
9CdDQ0LEdTDyeWSJprYzzOVFVQHdotOZHFs/OVU+upEDk5p6GeUP+Vffiq1uiwNsQtJjbTavQujl
T14U0wAgmP4INqS4KHFYwMS34qBesMafPOrrB7ELbdmg62+OS0btEiclyNAO8XcKfNfP+peMhQha
cf2F0g9fQml2SM++PhrSf96q1xarDIepD+VAnpqLKJ9wrmfmYbUp8ZaQr4+S+gZa556Ivg/67t9C
nK/EcCX3K6SSnKQggu78R+VU0gLGtU7I6c0ujsdU+ygFhhGj4iXoDsn2ym/7G2cvyCVIELTudesb
+9JrSk02sGjXAxn9NRCve9a++QAOiG4t9eGgcXNg4kITHBTwUo8otO6xr7rItQQchwtjbsgHNMsb
cPFUG9jolaDb7E/NK7h1BeqMlG8mV5JLEG+k9ooa/tzzuiKls5yxX1yTMsx9dSgWMQeafr33YZxu
Q29Evj2x6G0MeHRdfg2YBOl3XLkg0NX/XzA/EEJ0ia47JgkajMTmOztt+ypDvGUDHgfB/oyhhZMZ
Hv/oTeDnQw6MfXlCrd7aCw0o0PZGMIwk/k6StRyWDS+U64TU5Dhh4jawSxUxOm747OKXJKDmIpda
cbcmAJt13ZwTSU9NCmKcuQCTlynEtS34bO68ZDYbARfyre1ryQN9cFnQkknyD4q2ioF2Bgn/rATG
/Dvx+eeiXev1FvdHmnfzv7WEWb2f2bJJ3CqpCLYeKip7TaUIhlHHzMdqlxhO7+8uqSP1AJJU7GGy
jRcYfBZeAPm4sFQFEJ7XDf4Am0D9oENP1s3G6l+/wsd3EzzlrjkI5jG6MGXWQMOSBXL8N+jdN1nM
JlDhApMzAto+qqPp4rHZlFVZmXURBPN/kv+5hr8UVVmdvfqL7LW7+VM8d75KVMvckz+d1bTS6yqY
F882lZor/w4g7vEgbSCepwksIxJD/rGDzmOaBEup6bww9QzDVKhnglI/eJJ/xEonTJrCvmhWRtQh
JW7ZTxHolYKtRSrcBdtaPtZ9wa5JP+44MUjWqM/DfvNUjQn2pM0dh/PJUmpX588n76uFUvNudUjS
6kaNGbfWt4G5AZyuZXW2zGQS25UOmvjpL2aXDW2o/C+YHv0w9utEBOFtzfvK35Q3rgzUNDM4uR2A
gbYrBLmwQnBpmpB9nCuDs8UjmNowRIJuvY0tCUgu5S3WJDNO2f6iXmtMLy0HJmGqHJESwd9SWHAN
RhAP8Ge/Y8h1aKOpJSFvsvgMN9p+PpFtd14zj34y2uB3LLBRg5iYtR3kte5QWJV5duGe3r1htioE
ZlJXKoYBX2NVWHqpD1GWYZ1Bmk7USU4Yt9IcXei3mPqOwWV25YvwJF6UF2KLq1EkybwU6N/IOWPF
hl1fL42wEF9KkLdUaqOJQA3o7ZOGNMS9wO0bh3OPEm4V42RgJyd1xtffOvoor7BfDi4TB90l1Qui
KVKQsgEcL/HotlRGwFLhPk8IRcZLhbGm4h0Q3hFQKYqFnuIL8L8c0eK9qiqgDfMy7kcVaITI8Tet
6xLH/mG36NKmCKtsF0AFgWT9Q2Ih/SAvyhEfS/0QLLGJHzE2E02hxzXhBl1swFP8fBaSgBCq2SfG
qJASINU+zJihORz8M6ehjg/wmLZatqoIfeIWXAeDXqU+aOIPxaQ+IMmlhwAhOxWTarj8LDbdBPjG
flV/E3C8xad2OOBRHDHQDNvpN05iLSTnRMbt/d0zcJidYCuS6clXgVQTmV0X5mmMqutDmqR8gFwt
zpWqxCeTD2JKJt89Jt5F5b2y31uAcYP4OMKSVINMfK67qkJJEVp7Lcwg54q9VNmDOVQefozJbAhF
A0Tfo5s6WYZtM/MoxOqDLl/XuiDJVmlF5QbDcd25BPBPERyoWTCfDnv0wFGSTx4nHrmb5DsQBDnh
ntngP1WDdl0Ih3moaFlTcskuANM0Fz9zzV+QfmbmaUevn5CWVzC/wWYDuTKCkfcnv/pymiQMqfJ3
ZF/xdeZao8LjBhn2ki1rnnkWLb2StLXY8dSbvu3MMfezutSlIYp7mq7/ArUrmsdZ5g3nRL1AdE0t
VgHFbGUIjxOVPqkkbOYamYfqFTTGwKzfRbPYMnGZvkgCIn+T/DgPEfibaTA0Jl8AY4bWCjni5Vd3
t9tNW876LtWb1Rx6kGsoyowtzdEgafGXTAO8qqAUBaTG4t6DVzRJUQv+OnfmYqgYGMQPKU3XNPl6
H1Y8FpPKdeocf/afwDJw/h2TOzz3WfejgujXgaG0WA/yIT7QBDoo5DiOhxhhpJNjREyoVedlK88/
ByIB754kQN+NnnleLvzwLkycUb/wTv3PgcfXNf4ahyCI7FE+9mCRztIGKgE1FBGbAE6VLpXrFcUK
/YdHn/RSLOPavwNnd90MZMqL6Q/KxGjrVEVq/uhH+PO6zn1ORYD6W0DfGI2zcaCDsuC/lW8r5BlQ
i7kT7XXP1lPY0qDC09RPAjbFYNgsZu3PmG+IluSyZXxJfHBu8qXx5VHCFxEdPAxnTsRWxQkvfvhI
vZR48B3bSHzkQFVoz2SctfmJA2IzJskpxG2iIqYpgeQq03vmy0yJMTDlpZ/7JNzH9qXcEDRC3EWg
nhFSzBVMb+7iOXoiPu4bKQI+CZv5sl6ddCd1vQpYudprptk85M9SWlOI2R/UuAk5XBC0mzkotyai
ppfYvxOWOkLcdptbBfV0b2AMXY2r4tTIyemky0rZOA35MlHIzYTxkpZVThJxJMmwuHZC8a7FGSbL
MHOE70O3LuABkOIiLrzGiBKXdRWNreXQnxDFJ7F3/yYMnInGkExHCH09Y7JrbL1lo1D9/wjjqcu5
CrRPmTOZwKo59uHmL/zNXcJ+Gr12uC24YrZPoktCadKFaPBpVlX3mjoCPtUZyFshdZXpirKxVsjG
F1ozijjbx5xbHcOCmJ15d2N02GOXmuAicczjkLlCp462dbDux4UWG2QfGlX4LvR8WNIKu1c5X066
tDPcTud9VUTWwtxkJk8UKb6UATlxGPMV3GNeGxKlGDkv81EbAbo0dL/dRe5m/RTLq5/+FA2Xh/2/
abaaPzYu6PS9ixJpEGprSZQczv7uymZD388PRbQWPqZEOP7bnEh4udHJUNonOCCaNxhw2qQeFHim
CtvHDk+l9aMmTEvVSDq1AnLpe5jN/vsDRELrgybIw120ZbT+2NaAqdyCCgPGgZLuEe5iJa4NzE2L
etsy5njoeuB6Au3QXqz4uttxyqisRZhho9JmacMwt8uWwL3OWCdsIbNdMduMsicLJ7MmZg52CLU4
xnUpkM1C6Ahv//B7zwLqvHu9niuenlzao1dtFmse73YQ/XEXgPo5mQ9XZmzMqzakP5rS+8cx9eBX
1w9gimaPf0GnHvIh0nCCTX939+pUAscqqAGee0hw0i60nBWrPWtoydei8eg1rEudpZ05+EJYxlXX
8WFZjiKXFwo5g8kzzjw2t0Op2UhvrKsnbARdSKK22r6mltK3bDop1zHoRNnXWPos3ZIO1dNdm26Q
WdQHCgBDilyob+pfmaGl1knMl/c6/rcOFr/X8Bb/nqTePC8AhS/6xgk3Fp7TicBDwxIVL83ATx1P
JV7YYF50XU5VTs7T1tlNDfERZzUTztT5+ePuGTag7TlzsjyhEltmHqH12isiRPJ/Vi6ciimVqXiM
dY9E8x/34+7tm7UMuosREKtUpNRyrlj8h9hEu8EJnYWijx6IqDLK8MfrU6YYAipnqTFQVONiyj3x
GAK39NVEzui+C55p0fPnluaSwNvdLh3Vte7Qm19cYBQu9vyoltFcGrV+wSMkTicI1GDvUevElNit
gqVsHAZcpty114DhE3HA9AGGTkpVxvXhSJpC0VtIUBsq6SRmDVjonq8zCtOtqkOHLtKv8LoQeZ0f
XgU9iNeMBG+aKi0Sr3oR7t82ox7B6Tnn2f2/yx4rn0HDufI1sAzW7fkr7b6F1j09l0A7xo+QR5lw
KK1i5WHDcLjodB8xALNK5Qg4BwDc0CLYV2pFX2yOlXKgueQbrCw361L8DDYwjjGpczlQd+VsIOd+
+V+40LzsZep8i097iLhhTDn+V34GdbOMlJ1y3RiRb/2qiV0cgMtzLNMogNyUUcF7I0r2RY3Q1lhw
vI0Z9gI4udFiwMpbTKsWeaXNo+7ns/cT8Pa7uybrSTlr4daTx7h9V/WSolone1UCsug5V4rDlOd8
NCIwf8ugsGGpQR+U4ge/VXXt6DEleocv+hDv0OJ4GBbFdrZa5ADLHWe114iSBmQnP0W4UIxKTra7
d+kGvJWGUYvj65KjUWqngNRcurQBoZY7G8Fy7Z0gcVyjW8whBXeb8lyqDu/A9rRW4n2gDuhSVtSR
ZlpF9DOIkgE94OaXxVN3c+BSg1L9GmIna6lSoCC6IIeBTN/LUKGDVsA/J79Hao7BM4qyUrax7eKn
ma8+ZcD/ikBZY4IT7QT9f3BmGbQJ+rBu0bKMIrxrsYCyV9sAs8CE3tMwfQi8RmtssnOWZfa9ZE8W
vZZ/V/nepRek/FZLN31G7T4FupImCvlIDjz8qPRKf9BVwCzegyyLZn/3LzWpmT1h4UlnOySOY6Hd
lWnFYPp3qJxuKj03g0pRA0dmXtLXxmS+3qIuo2ZGn3qO7cQwhf3csCB5JwqwIjXf1Y6FWYAPFgxB
de81eQqijclPqqeToryM9MB7YUF2tbN6yHEU/Ao6oJVeh0kzzzHhy0XRflroBXfwvd643rb4ti5J
Duh9Jgt3qX5EVt7/CCArMUCZPbgvaFAKy7y9G+wyBUiwlCOPqMVJsHnPv9ZYO8cZ53I/Rwxlz204
fvtH1fXS48yMNdtfoPBWJZlruWzqtx3QHZx6BUQc8MCknZVOu182oPC1azWLBiU+dz2xDuLJUAdE
3/V7jGdNQJkNBhwewOePDFQKKmCpmbBbGoxOUYpdOAzcSboDrU2Hbd9jXUauEyjpIK8qJ2eTyfum
0myWpD/9j35tuD9SK6c3G7uNAKgAyRhZgL68i1W60dpe6lG5nEtn/TuX9yKQcaBqFH7D+CPymaGe
BVIvkkehZkcmJP/KSkzjtsHp4HOJWJjJqYjQy5nnxqdlVoS8Z0yZULdrwfY9PhmKw6pxkSKkzgwg
2Cuobn9S3bIUBcMbrQ3fUwuxa3B7Ca7FAuwUHi/6keK3OtirmI04OLhB5c/3UZZDMWR8guRP4RMO
+sPJp6CScoL2tn8FiGRgKnE+k9ahoN1+R7I0MijExDL/frSCXGnieL08OHzVvFmtRBpRgxjtiOrK
pNJsb5CQk6Au2gpmqyhVLasjenur9uziaDtVkreVtyGleMoSlTRpPOUo4xQ7zgJDreuIHJVAF3b9
7qLyZsaRpwNHheDiyKhrlI2dgnGdY7/VC/hvQTZgYKIgfPGSkGZZFEALmGLw9uYEnG77iYC3mi54
Y/XfImV/Yd8G9ylQMu+BynvaJVCpd/LzRlamrXEmdqUuxcLOIfkjgYGih0Itcsne3Rn+YU5r9ejR
VaCm0709OgmMTfClFXwhaprTvRUzlnyqN38xOCOLAENNu465rumz71JVYhdqLpBX5s4LIRxp7DLW
GZlvRDout4Te/7jHeyuMFg3mRuPdz14eg8ztZzSenbX+sCiMKrfNfKn1oDGf/ZekJKlSFKCR+dcX
/hHzENDREkDHeWavcozhLCdMDMfZGSS8801JNjQtOo/8T/5r6d5cVBIy9oXszbZBWXuf5J+6zuD8
svpO52QUcriXRP4TbSdm8aU02kLQ2VIs7Ywk7jwdBKQ/dlM6D7jguhYPwHa+TTAdLLnDKAh7JxcV
poXgFP3zk7R2vUGtj0w/zHncfFyUDTvYhm1GAaSzuP/TNaLrMqkVbirUGGDNpfFRPd709834bEkT
6ZpC3UckIM/B60ZMdRzZFW97D/X4jxcyUeuCayeGoFkttEfIO/dccp4tWVVeQlO5VYUq/J0v95tb
qYTvCmcZrEf6ruxkHUt3tflAQjqSPPCczC2/POjUrV7xU0+WCINgRgCzRqGNRq9nV65e+7A/vZza
cgRkuolUTbtE40yxvfIikmfNeQFQgsUwxdIjczlaMrGxWur66Gr082iZzhUK0EeniNSjP62O9qs0
z7SCNV6LMhOyhDqLd9F9dc+B7Jyyr2NAmv9emUnXOjEns51lqDuHzQZHLGLak+wLuAvK+1Nbx9ue
ia8x4CkY/eGHhc+d7/Bx6KYvnstKa90bCeTm0Bgc9XSU0rOTi3fK1z1rEzQNF342hffIs2/44408
qRacENfVek0+VPpLIG1ATY9f/MZBzs2Jjmcp5MLaKCxraivZvhGFjKFFE5QCcBEYFC2UPyq/RMzc
YaQZuNSZA6k7GwJ2oeG1zwliW7q1JmPFb13Ht1G6uDXEwHB4fU/L4qNieNp7yf2AY/yR4TNdqzp1
dZGNNWNJq8mQbv3pUycoZTXqwrUo1o2cC598n7mRT79PCRm7BlZUU5VX8MuY7zhtzl7yjAWYiMGK
nKmdeIYdtnqxMib4iVdMUnbx42/Km41oMRTEHFK+Qy8SJFfClXjmIYgIjg/mEhUmD/EATh0RWqEm
06206RuyNXPXp1HCtY6/+UXMIieY+NycuEPs1+2MxCDMZew9s8jtBkSK3WS08+/cHwcNo69FBxc6
vMa5wPAAvKFH3DQtrpf8QxxykNZ77AtsXv5rpNb8evm4nCZA4ZsRWQeMw44y+sAT0RrfxNvaPhdT
HnPKX8YDRYNokoz2X5lUN0Hv7SMdwaqXqwcO13TSKT0ksMbi3A9sTRjUbGIvbvXOmiZgxx7ca2HG
XA85bt+ot3yHDbiet8IjODhUbHgiscd2bLz8HTQGEN7rTMdpyTjAWMfNtWnigfdrdpktDcFnvwQE
Oy0W0GbjN/3nRE1ARhhpmmSKDP3Pq6iXaQgeaQUt8lT/lH/o6ExR0bd6/ABBt/02eW/AKrsyoI/B
xML3Sz0KA2OZqOtQA1EKcn35TSsxBiUgIshjgEg1GtBAdpOPHm3nhK9SjtsGqKvRSkx6RwzlV0zv
xqS/rw7iYr3bI5JlNrE3nRBGrwlG2zhMHkujJV2FuDMHsGoZFgiEzAmOgWgm2dFWXHvuBYHdEKD3
dMGM8D1ONTphAiavpmkkzomMMkrJZsqzlZSYQmOCfB/uWMydBzj7sy/m5f//dMA20dElikq7gNCp
H1cjqHZ0MbTA5+Z6AKHDdpQ0E1BJ8fMJmBsYeqiVoYAaLJ+7TxsXRXSIFZ+n3CgBkxHDVBcH4Vs7
qv5o44gmvwbTWgrSW913BNQXp3u+aP3CGiNN16m8bYsvZiIYeqMFKbuX2JyYMkVsu0KDsKQCyVMd
1HOBoeFiAxu9gNKfquYwNj9X0LHBuawasBkdJbFekmW88MqNtHzb81F+NBurWKLrYS61CtGwz3EO
F2eSe+AeKZICIxz1SNstbQg54rduKTx3GPsa0W/HL/giq86MrseC+n8vNPnHa5iKqfDLl7tkq06e
qaqFbS+xkG2Cn2da4luT9hjQRqAixbI1yd9KLbXtzMV4iK12IWbHUo/Y4vW4Bfg66+z5zr2iq9QZ
3UiU8RDX1rR4lMVY9a0K28iEpioDMbn8McrN0Ekfd3zHfbPyo5/ixM0Xbc5kzYAr3IFvABdvO2Tl
r9zzDMa3rpD9lpkXCCnIatljZCERY5pfclQHUbuODXXE2ad+HdHZt6h8NFHRo5+NUW12SX9AImPY
p5PXhYYwurcEUztZ7UC2te/qeonfnokcD/I4p9pWU8GllcXK+S9LkG5hybvvwGbnenm1ih2mqm3i
/GmLdis2zwR6/60O03b0E0yNP2qFiaENofgkNhRCA/3t461ldU5KJvXDqRX+/aB6GyxwqLVJDxCx
VsYLabStovGFk2Wc3ZuJKLYmdvxYxn/XhB0g8m+U/9o+FO+RCCMH01Upcci2Io3Z5lebh7k/Y1xM
42iWR/HTkbv2XB+GMPiGqq5dAxLgxT0sg343rXbajKf+ZR2F6nnJe6PyGnQysHu5cU4HUw7qaO7o
Cz+8PaZ+uHOJIZkMEUCirrsYxHlo/D0H+FtE3JEeFoV4r88PdsluX/3daI1xtTIooLLCA8snb+a+
jjc4FIJRo4wW+/2B9mbC2AbgZErwLNezt474VPmrsCifsCNRmQyatFHkjAQ3cmxCe+3ug3xwUBFk
WsfT+ZeTkRN6EaeLpx76JckhW+YSB7+k+0C8OzsGk/KCoZbthnZ49pDV3+It3ipdXP0F7MMBZ158
SomXzwF7qqSmvOha9Us0h7nQViRC+U1+tKwaj84r/YbZYZ8YahCC9r7OFsaOiwjicFmq7RVx+W0o
92L9QU8uRo+3POHWo+OS+UkKVrZbPiy7/tli+LIdFh1QUh0Sp3Z37r+IKVrzo6sWfrDsKTOpSK9y
VB/fcjmP1dF0tfRQfAQwiTQ6FJtBRA04MjzALr2EY17XhxMK/n7nRNgAaVF3vjXxZP18CH/T+RpR
4mo/tzYSdHiOGw7wjQu1ivNwunCVlOOtL+Bq6djxERUCJE7J5zPzhFTVUW87v8Jed2w68znh1Ae8
Hadp4UkubNJyqfOWZyuroUF7foCDz3pFojj+yRiSwiOZJIjlZKLoyf9dyfqXDGjWDMhujAnhJzE8
ftm3E447as2ZnkKnwmJ6Z9b41qJMo9GLLY6/n01lrW1Rhk67tohtVb45cATk+8TTqm6Y80HxLVC6
zTb204ppAbYhGP/sRPmiLdeo2IzWaq18GJa2o6wmq10XRp+lzuLwt3ERaC1YPfqbnO9UoZWCXplA
L8rJf9o9TFKzlLQWfoBWahWMlbCD1ENfLdfReSHvsETHnwN4VdDEsJJ5mPF/bM4OmwWj+7Q6a9W3
r89H6XLY2BaLyB87BS8i+mWEFBvXwjfBS7xlFpx2r+sDsjDfYLMyaCroJKBnxrhkxqCtAsPoP6tB
N6Qiczvdl5MnEHdTfBdoe1SdYW4+uILxRhfRF9VN97jbK9//e2Z4pGTmchn+XfwJvI9xIyoV7MDi
LNIU+4d74LJkaxPQWo2o7PfQ5qopI/C+LlB7DqN4032ac4jTtYEm0EOB11KzZgr/PtOGKcqdfDix
h2Yr5MtLG9g8k4PPHEDN7w2wAjTv+fdAkJP9SVjT1mYHfGblQspho9nLHc3OB0+taUeY5f7ZaEhA
M9faM9RPc0Kn2tWlJ02s5nssI5qpw0Q+MkErmUvX8QC7iYgCUzamg9h41ASr6bWlp8VnyeQVIP2+
/QhkkB4m6VMqBmj+ZT3FzKe4XEz+vEPkN5ZP0/TKF9UwrVu9TIfcEALaaHm1Pnrxb8LxKLDvqxOk
26LmLx2mVfImx+YhLpl1TfFH1KtX0d9PAHSYVkKvqHUdjdOC4Fz9sqtRJ2JJrEqaa+l7IZKwaByl
ryh3eGX1JKEVLe4M9v0OGmJH42Xx1/dASkIKWu4jUj0Ctp62bSISMbeQM7xE84kL3O66mXWZxNBZ
IzIv8Uv2EqHL9SabpQsQBfPoKv1OfLgjPl4Gp70XkowNI+kflWYA1Uww+VLpX+GNlDSuqYkwI+tn
f8HV9fR1lzQLBfcF23JfUlXIx3hv9F+6yNJ0/x+GaD/J0DBfEbDhX9cP/RrATnssDGYhhYnMyTOW
m176gvZs3QFEjlwv3qlbKs+wNRrIIIEPMrZMre7Ln9i9ih7t4i6uKY+ZmFFadMO0orTnawMWJgRl
j24xx2/r6scMiyRgE76Rc4YHeF92x6R+oKJJfiKPx+fpbwsLSojcoL21Pdex/LpXGTMLFNCcLJ5p
qrjIW+VUlZWKl8pL63ZoVRA7OLGlqvB7Fo3Ju9+p31Nn5mrlWUIfKsGkibBdPcVWdAP3lb+n3rni
ppTxr+KDzk3lfNxbvwd0bZnUPWo1yJ85rpHHvulxtJ5vSwrGQ+YxoZP6oDCYehsDdVMZK+Xd3ilp
0nmG0YYbIMXLaqgpLv0bg0GUbUHStGBIPf3ppj89uiri6Uil2AawgX+lC+FlTQtk5+DDUqcWxj4/
HRpznYyXntQtzTusBRm6cL0x7c/ymFIPDNhy7jexzYBBhklAHQsSZowLUG4/LDUPib7sYAqGnmzi
YHZj5TP4HO80SBfplBUka1UDPjHvAGslzfpSv/09RBqsszqzRzoTbIjOJDf/zCpoq8o13SROUTy2
3C1rMZXrFYPw5fZ3c8E1Q+gXEKsap9P1l5kqttuLabZR5OUFuxIH0YmGb5Yf+abqOA/RHsSIrzQV
Z8xBjaWGfWpwoEEOYuXFSWC3l+nkfgMNXtZdb8eaqoSpGGStEMk7QcRC1203gvp1wVqduIKnZTml
mgbKher9LDj6lAJrPAIJ/hYtajxktxQhD1kNxMVJeewsuM32Zee7MrN5sWMygDESnqy5WO/JrQup
HQiscpXTR9/qQozapaL3zv4BhLewAwr3xPbZsLbY0Bg9ViuXmLmkJWMrflklkOyZGQBDikPaGSHI
7xSUkSybbg6xU54MKbcVvniC3ZQoPP+aY4mfk25ymZMInZHk41tLlRyqxdCPm5xMlbjW+53NA7O6
NKkKvPb08zgMWnG9RfcVVN7HXzY57xlfr1Sg6uoOYTcwOrBC1zZ7ZUyUdXGrFLjQQ2y/zljujN6s
10SOmShxGgT4QYCMpwriRXihVjGAASav+qKRP1vG0kcHRpeYeUYFflWmoloJjgkpwSEvfp4aCVcH
vClScQOQxPCjpSB+/1/+5s0GcZYcUORXPQ+DUvo/vk6Doz/6/THWrPVlvdI351X76f/4WpJrs5IH
+X6UsSDMm0Rbiuhwp1yWTAT/H6evDtKsi47MPygjVAoZ5SL6oBUJaza4bOa5oonv5ZxPzAnmcj3f
w47RvOvQWWMCtZkJE/y2Y6q8Y4jEyczLhj8KDtZcQ3RW+lfB3cfWUsCPYxqLkU62xghzEhvQ9fQu
QijN+5wpAoqGdwuZGUVLcFhFIOg8EZe09VCVk53zs0qS0Rb3/BT5Gl9DpNJGNNTXFN14CeeRlKU+
2geyAGepTZEVwTVcM4KJypmHthmEleXFsDtEStKgZu4hEfUWy74JSHPMH6wR/fMQxeUXw7fxxjcN
PDXDbr4LfOQ9biisdfgWTUw1shHE1+3ZSEpk70QrsotO/nkHsJyb1lNnI1xA7llEKqFF6R4Ej9rA
w0D1WDhXkIKEuLax8QBowrazWWMVzqXtDhslQCqQAI6lLE3Y0585FuqFz2JSB9jhQsccpWkMxJLh
fXB3bexBqw9XbDHx7of1z3lBrcqkvz3NpJQDN3Yxn4pAGYLL7PFX5FCGL2nXHyZJhyZiZNSpGd8p
0bt4qlAEAqxPWrTrqvwutn/Ln5Z7tBzS2jyAkd7L/puyezGgqsRAEtbpUhYnumsSADTAbXhvX3A3
W7LEhZ3wDQMg2SbvF6y/0pecwCXfwzp/fzrBbSSSqSXjPlP/x3i29PXnDu6Oxrp01F8o7QjVxjwg
f54NDxw6YjNtyUWXMN8zGxM6/72Zhrliorl7cfUiggVE8pE9X+Yu94NeFHxOepvgWS2QLD+S3ns1
HHak32n252ZDrh8jzCEBY6K6wTnNO9t3QaVZ0k+Jdsd0268HHxIg6BIRAjyXZNLU6El8gDM+oNCs
+BoqjLJLD/1+un+Ape4vQGTuqSYgIR4x6qTm2IVJLVzSsslI2BQYqSgN7vX7NGnTH2Rr2FCcX/5y
zvoMgCOVVgk+fuq4Gsu0SIvoIyCuedATluQz2PGAXxUSdzi7UKP9NJHVncheLEK8vHklkJJj8bhO
xkTE0KuR0zKpw61ANbJV8b6KQvXGgbr2LKrgEnH+sYtuvydRhmmiBLHhwAxhkDtnT4vev02Q8KTf
sX5NkBubXXNDj8bPTE/M7PC7IJ4Dak/z3bLNIL7UnM09IGkiKNDnsNvflRtX/IVsCZCJ7VMUZ+ey
3sUPFita9/GK5KbL/s9MXW5sf2EUuJiZ9ex67Ib6B3nQk2ybJcmOsu6HwXLUxZFbZJZeSxN2YPTO
qo0Xr2bMVMSagnvSQ27jcHI/nw80OZfu93VMaOll4gdV0+krUOirLUg9AMJEKWM/eQR8kxzvH1UN
PUgGQpyoqMORkhN4xIN5TC0tA08QFzJOnjjt1CXoEP4LdIuElpS8ZiA8+99YiJJHO3hqzW1kMhP6
7tXA/qmyAmDscv5WOFgxyqXCV8H/fOmgRwkkTpYFn/zmq5Q5DRCnvElskKhW31F8CULgUyJOhw3F
P2QRX8kSpGI4Z+c61aDGPJw0xkx5kAYSZmlucJsQFiS2Wx0jozLh3wUr14/1VkthEuK407DQcgqz
C/B1KHuKFlxUB1nmdej2uEUEi1tkINiMKdPx+zY8g1BBl81notmntdAm9ZC7Kt+KKmMYpSxvm1Oq
jUrHMa6me9uFagVMWOas1J2pMWIsjd3LJgKXXP3RRBcUeqa+a7mJ0BjsLpfKrZhiL7RY+wLJ3/kj
fqMTb4pP7/DRjzqPliIOclkLzL2RRORXmjpyG6AE6SvUaqFydRM9Bs4x1xBCiDvNTydrpF8Z9Rnc
Ph1PoSwaLLxU6hIHi9GvXV7lzfl2ulwNoHTwJdkDCL81eX9xGWIZrjNrL+BNsdqhFrWNxMIjqE+U
fKgtE9Z/LtB72v/gLDmE5Ch5qmEgjjMTGtr7bXVXNPqFifWKC5DIxVxqcWK8v8TgbxQQm70odRMn
36sOr8uMcl0O558Kt5SRo2eEyJxpWmIkYTrFZoprFCdoGtbk1f5nQzSHKCMqnCTXH9glCCxwbtRO
7AL+Waku2hh0fXbKWKBAiKWY4w62tfF0tmOd2BwUQR3yWUA2QkAQm3sqf9IAsrcT4NLrvu19sv4D
FnMNFBnY+ce8dpwVCTTWrAG72uUgWR208/RCKwyWzK0GtNyVdpx/QWHXkxL/4JYAQYl18hUoILml
2zI6J7Vfixi1stnwBIyzmeBK63mh3k4eE56goeC6wsA/yfh6e9T8j3F1mtBcEy/G/8JebdrUniAs
G4SanEqz6iNxpVmuRB8dsfA14QhWcSJz4bDtOc6UTyyf2CtenWpxaRi0HlWlMfYYAtwR+tn7CoNW
7lNmnxZZshuzoh6wcnvq+VVKz0rSjQ6nJ3NSEVvKFOag41IdECFBw4tWl/26m6SSWPiiQZRhRNFb
shcFLhLLyatZHUeyX0hXVyiIzuixpM8Ceu+yak8cIeOWH5EWnu4aNzLY0J2J+PD60Z6ynkjfqoTO
D4sKfyALR4MpbKOAqqDAxnVWJ8TniK1rKpRmTjdOsrJ3qty1uGhc7efDA8/FyYOLIh3fGu5dO+Ku
HRRYqBHoJhops7sAGNhdudgYI/7OZOH6iLX6KJvA1hhRH6caCKd1kuF3NtoHTwvQWx3abn6Xk4pn
/Abh0ynDAHxbZ6jBjatTSuIwYXEKxgmjlx/K6qHIsUVP8itJDJ82n18uLVKbB7MfSd2YRXqm6isp
1ATEPrP+creWra5nDIjUE3cPK2XnGZj6z9I42wxesa5Nz0hHXn3fPwL8sagWVAYz+NZSgT9yUFHw
O10+AMNgPnup7FepmcUCjwTGsrzpzjsNRqrLir7gdKgNnmBLggNMbhklZrBX3kmu/IfLAZh7R4lp
KrYoMPxfgI/tt2IcdnUuo2jJqhS+v5Gd2rPDX7RvidrqVBMrropGPXX+W0186ICEDNkGU+pqlqJ5
Z11TStv6mAYvmLfFrFgfcKyRXOHK0FxiwCL3mkg2G+XRaQFAMh8DKMxkHzyYRiMYNkd91IUsRjEF
vDQFkAbw5xwgS0npIW5T+VKbIyJde5O+lISp0juNOzJSLLuq+oKqclbC06qnDN3OuQrTKgX+tITE
s3BTokGP/2apN6GSbWSjafcBbqhF6+/He3ed7KbYlFhh3j4mYNj/osS1FwWAMJ+blD8MmLn5fvWX
SvAyckB41yHj8DGH82X/DUY4hvqndCf71fUuTncGECsP1EiXfFfaFXaiSrBB82kToZPZJtBvWkd1
rY504zjNPGFEtFmFop/nDh2t0vyZEo2dEG7epdTFMgaBuk/EWolbETwp2pkX+kD0Hw1Dt8COzao4
BMKsChJkgc193qUBtKHo7N9gJ6x7KpIE5PK4bqMeQRQODdJuMUb6zfT+/jLByPuzCxcYv4sYfk0A
GDMFhZ/3rAdvyhr0eht9vEvPnL4EJgNnva00MfgbAbBWjUDBT81Ry81JFJTpYP6ZCmEZPqsALd+I
84NksJY0bbST7Dn56LHrijaFsw3lkFVOsIxtBCNAWaHarJGmUS+HcB8pbMSRLxpq3c7lgPZdpU2i
33IdttzewjtZrxMeDs15ufsP2v/9okORVIWyNCA7dle6OIfGp3VpHozmRLQCXnC/a2m8ZogDznhS
6GuOjKUIAes3T7+zibnWwkHpw1/u6QyN4782yA/eDoDXOPu4271K/CuUoqGApS6/DJJmFQjI60WO
oKb10k0WtnrTV2WJtNoGjPWqGdPJgb4AHpJOhD3oXl5B2MxUwyavhnXqRnRnnAZULvabPoellPYq
KXeGNcqDBPu7/cOAqcfytAyzghzELAMvb4wq91JNMsyqgAOKouZSt4YhWrAV7EFit12StlTL5TNn
YA+owIEPbZupf0ylnI4fHZDtDrnRXGsUhLRYgp9hyWT1T6jLlLjkYIRaVYcj8M2emA5s2+apAnBB
ueGdLzujzF1/iNIe/4wktB9Z6RNXzSDlLk8imO5S+jHpGhRYStYRzaF5k6HC7OXQi5Oh5g0fHy0g
f48Mt0aT2eZQF9SUP8yWXuZD611X/hfKidbPLjpaTg0Io6iGpxibCjp6GDiBRujJv06lAWmvmPfk
eqG8xWWayhHqlejyQLF2rX2jOHh8XtypJ780rVmgDdlu266QaA3axJ9SUOg3aPZ6inOg6iJXOrup
Ud8+aMl4pFt7JLWe4smvOSMHiQjS+x/6v47jxfdR4TA9HxTAYfOVWWCYH/77kCsYv/Bi8RCMALfU
6+YEY7kUrO92LmXKElHnO+EnrX5HOXsSPvCWj1bxVEFzn/uYkv9bITlim4vG/sOp1fq+Qu+CSmMQ
dc3cmBkeZlH7s4wu+cU3z3HUBpCJ0GW3xR493yQhNyOPtmKNBSgSr9f+2yNoBqAxJfi0h6TKRjRq
wemmRIy2T2g75TC3LiYLWsyIyaFFYGmyf9hD5uOvwMf2b25ur0fRTXjrrt9Vyq+kd28NSIhGSQ1K
wqVAh7z+L/JkNJyAiMBW1lt3STVj9N8J7TfjNmZUSr44m1sB0pA++cgWxCUnYJ0WcTkKrp7iJKhW
i/hc7p9hSFI7463QOIYSmhCn8nzwF1X1Yuo94MOJwhSL9mihsbvR2GZATn6B5VCWdLVJYvRR55K6
YnzL9z9oxnkw3e1bBIPJkzsaWqc+rrRdsWFK7UfsnSsCGo1AWaAyvPMsiP9Dt+WKOhkezF1/DjOE
pBxel+7HAmug3ZQ1FwTtSbi3PsSoh/IG9HwjL40j/zL8U/zsBBoUAxDicB//wlZr0LXK3976Ereh
/rTjxFuawHlSJtHb+nN+qAcPDkfHpopmbePw36+RB6wwXo9+1G4a+O23nszOp+z8Yl9YQMGJwbRS
vPNAw7FKkXQBPb0OET42eDqYjKjyYcQhJtW5hRd5ARLr1+MAYAaHpGDdvz7u87CGDfFQOSa+Q8C3
xXJd0uuOWOEpSB53p1LX1dBCyV77MuxAAORrLFuzJKvv5k2YvaVDCJ62IzJ2/3xmNA/clDTPRPFb
QXXzUw+yd/sBBTbhiXxDtNiFa1uejNye8Wu+FuHehzgCt2ykFDkibjc3jdQs5hrnPcbHpaSa5Iti
oag+kQsInrHSDwSObwuZ5AfyGAX3KhQ/ZoOW/qDomxq1LXSFZf81kypK1g1mGy3jeXe9ix3YJNxv
eALERjCkYr/qrZT8SZhrDyocxlrKbUcMuznIQvCERdxR6sO8NjvE4mTdCcU6DpI132g8dRyqRf7C
GWTxnqrIGdY4sKZKYm7m6cbMpfDUuia+YhdBkDyql9ow0TkGyg5Q0dvmRg9bIvQ2Q1MQPRAhqhbt
l/jL+6h/pPpdJleS5SSm2kcW24xIGmBjZNVXFsEnuAnYfk3ImEQ3NMH7bGG06hv26JvnYddto+B2
FHGxMecgGDlCgjDRzh9E4RxGi6ye/JlWb06isKpm8oS5ihL2fSSQAuFxGIHxhjkxSGEeRtRisSiZ
WWAbTr3SALtVSz4shXZqQ+V1gKZuKu/0Llcbmm9EQigwIpB+nOwCLAvWfSIxcpaNdlZwPYnKkgHj
g0GUj3fhBUnrAJ+tHf93bKC3nK/H+PIZynWHvSHx9jf94ot0emzfHH3u9jXwvuoPCgBQtvfOXfYQ
ghtD4TPqp+oDMcgPvWaNEvULhzLf1D5ci+x36giJ+IcUV0MxRyfA9geJ/ShjwuZbef8AmXCNrBbs
Pn+2UmdlOAD3Mz3AUpMWmOg+ceAg9FERRbha8YXNyq1Z2weLQXXlV897qjh2gMcCm+S+wGFkXKWO
0RuRqt/AeUtYSNuBIqRZH7fDXb8IZRbXHMXiHXYxLXMUXTtcLYtDcXw0+U0onFdcDJwCY+2W+7vv
o+XhDaZQRkMPHARLNGLqrLQp7sR9aFLFcyVOGx7scob0tnhLW/4YL/tdbka43mDhPRbUyC86kUdY
mmyFgXXp2tV6JV9GRK1GOalLc/ktZTCJxL4TDpO9ooovNNjO42uV10qPK7jNOHG581HuTvJO3WjN
THi5nA9dmMnNKSlimmUp5N4jcZq72njmbaI5+yGvr8Vp801BuGRuByDDcONoT6S/XkTEWGWlKzFm
rT2DR+PT2TsaGubgMk//VUpe4NwKDv7kyz6OkmiOAoY8Br6oj0j/EJ75Sfpj7IeIS2Wgrrqgb1fc
KO5zQ+q96q0jHqvM1Ma3T2HaaLL+eUI09o5C0UIQGOvz5vPfl4TC1Yz5BBJVswSB4ZqrvOtqgPjB
lYgukDuAVKsfbiw7OWjSy/nnTpScnSdG9K/DJQAB3NVzhzVr+BvFPweqgXWcl22BfSSXO8WtRJrZ
jZlHPmVm6MNzaWdMLHds72sLRRYMVt7O+c7PRIMZqsmGEfTUpp3Q1S9u847OHDIjbjm+0kRIFE7Q
ezkNlQ6vA104IxxCoJohqqtszMqu+KMVnIpKtZoq4TNLQbM3y+bP6+BgppBTmEamE311Fesu6VvT
2+6Qy5g5NKaOiy3GFxjL+eartUI5sShqxzwnmXnXCgIFFDwwVf/Di93NHRxMzbS8vyjVPpNc6w8L
FZbxzMw3maB6Gyx8SwbfVBe9IMAstaMR8fHxRlU5IjS3qC5J9aKtJFZnhG1e0kiGbGywYFh0mN9F
yvxcWK//965gfSmkPqTlZzGCyVT11ATZV54FwBK8RpMNn4yMAqNTmAxQaHxpeFJ7R/PrBl194Xc9
iZxA+IzTxpAghHn9/pdD3msMwzwZsTR1AST+DEBUphSetzn8YILLDlr/24Hw37fecTr2ApkKverS
W9awR6p0zRMfYe9TUumOxb61Gn1wgKJfxad2JKvP9GxETM5Ymv13IrrqCHLmlRLVK/fOlqTBCqVU
gglZCpNAgqIm0d9SNvTHqoW1ZEvSlUKhNuDxKieJWCMLRIFKaIZkYpq3MLttG0IeqxE9t1DXTm8S
zecPNBsDafIZNiGCsT64ntbKxc0CmGaon8cpb8DRMW07qWnbOmE1DNkWxavMQhb8BzgiWXscMQqU
9Ny/yJm4NSASTaCo2cAnMl5gyaKo8aPyo1S+rBk/GEFqcM7dLNClmaOnv7gtoDODIy3LTyhwHxiP
rNEQCVs/N5xyXtVGJ9k1L5hL0NsTpHBqxrqSsr61gE7IIl237opQVbNColtC0wKv2X24lG7/Q/jU
/bLoRkUR+K9WSZlxbvV9Qw11fwbBLyVFmTDUefNJDI7rKln/YYPS8uDFu/JNOwIvxU4Qh7IfVmnM
uv/SNCujJxqamDCndi6CSmJs0JolBY3JgH+jHExLLB13MScwguz+BRM+K4Eb2BIMJaMf474+qFbV
RwFys7RR/GBp+5n5nn9L1B/ynWbUxMVJv4/OC69lLVY2+wD6hFV135oiiTKREh+criD2XYyeQ3+Z
R8dFRZ0miRs+0Fc90jLTsTpp9RoyP1+OJt0PFalRa3zLPtYBkCwDwv5Skuj4I3JMN6+BYQdj9dHi
BTi8eZgrhJo7XR78r0VoNX6qZaGBYVUDp4HLSDExO+bQDHgClHsNwATFG6CoLYzKJwKnBQpXi/MM
joQ9I3ZKiSdDIyo6tkN9rctNPLU1HEA6KMCCiDuBOtFwQg79hnLw8biJq+y3jdvVM+lO2AtEIiFr
jGLishyUe2VL4kPHTXN17RxcA7UC8PAETMYpaVphetFNe74oJL487FVb3gbBohEDA1YZzv48EiMA
jnUod+v+7BdZuI9XMFzcFJ9WoUBy6PGAxNvqghAwInJycCZlG87QokhujZBC4A3eElkAr6kGBy/H
3Fybm2RzRB+Mr+dIn0ANBCdrSs191hy/nl2nf3/K8T6+6ac4V4RgXBKaou7xeqtE4/g7DoKH1Qpf
huj5B7HgkEj6UA8rdkAcsavBg/MCg7sXUv07Xq2ogHEWTHzNIPr6iw7cRME9hiWmdy2Yilml42ZN
q6aadzePBgJHblovWXH809UTQY/+H/lvijAoOyjUTeeDvivOEVsZC3RyPcOAnGZwwCOuROAPoNY3
IzZNc9Q9m/5gMmMcA9CnhiOc6vfcDsEiJKJkMYQLqJ+laXW9h8obcdrTELC650iGC5iX7R/ZHfvG
kpa5kY09iWRJZd7kBVouqNWd8C0HnksLS4riKXJfyk6qxtGuFdAJ6z0BscTQmH9T79DKr9NURYHZ
Ke/DsGRY+p40Bihb5iEfu9Rq3RNOkzJffrqNUg36htDFoe0jUVpcj9kr4f19tIdIhShe0Yaybsjs
NLByOODkg6bjt+SDMZOWv017xCETQwOoWPyDpZdTFM9S1VQafj681epnhJLXVguUxboXAbxKrgBk
M23cpiEx/ryW3QGeI/jG+vSm0DahN0jQTrFZFjIvOt/6NYvdj7oGNlB31Lpa3Ri27ZJCX+EllIDx
6sCUFobzsyp5lg9NuWFzcYLkQA/6K/Cm6dWWyOuZSVlXRGz3JfEo5L3cVYV1lubj4KlUrjrpfBSu
LxuABUM6ri3rvHHVyWbOnPcQFOtvi8yvsKhnvaQL6cwk3eiDHap9kzwHRZLGhhn/C6nTuF1o5OQ/
v/3h2NuGXAbWZ4ETOv5sirrma/HuhL1xcNkcdtCr7RAZACoTIuwuag7QzKNUvCsO4RK6xeZ5hPUq
TeToQ+Ocr22uldJNjrXRRMTuMwHgwp6j9/7Eoa7yyPFQljbHcED0WzJB9D6CV38mR1d0LuSuWI2w
SeXmXW3yDFoZFVrfZo9u7nC37gKAKx+Sjl/mOc/8dxvawfi8ikdJFQPGoVdvs/aG5EebIE3sUAl+
tHEaBKgKO8GEg4QYw8pOBXjlY0dK1OsQo+4hVuyOrUUC7+oGCNDLgEH05Mj8tMOkTBvJu7tZxgkO
sKLnXbskeEv5QKgqxLRR8FrRB6Kdnhi9caUqpnbZ3YEgv+mHkLcj9YByW38oymDbdHSPZmFT0uGL
VbasAchS0UKxJ7dKRJ09vDwVW34HpIwx7nLWzdyGenoZl3EbOtuLWltaD6Gk9r+vckJaLcQ4uCb1
fbeKz+BEJW6tqbSfqp/BcZyaP2c5yMk1Ig1CHf/xWLh86Z9EaYWfMZLw/X5F396mFE88AD62FQjj
HEJiOF63Sg7luHxp5Yg/QfLLkZigdnbuZJ+U5O/3owEzFMSE9QiFCigo4NXZqQbyQP326InSEhJU
mGZr69sBSe1x8HCZpacBuFSv42EoKIsdkvHWSFhLclb2xBMSOQ5SIha6gzFh5CZ6uq5S3NyyA55R
5NSBzummcxrHBlPSfzwpSnedTKX0DW+XC9YW8BT+b+KlPjC2WE5godHVgJvmmtvak7aGl6mOaLRJ
d0kpeURuedT/aIav2hceNLeVPoHZ2xvTSRlJiGR6MQUAr8ShY7h/R6o3C/FPT/FLUmFfOT0QPzTC
42gPBJlUOT5gIsA65JHsx3PI/JOfWyEi5HdC/cKKpLRzxktC3brqCphXxlXv6LJwtgb62B7vvUcf
iGAtkEwXKmgZOjAfgB5fA5VsEU85GgZLD9eawaj08+iiV+9Q5IPhWCBSfGWukzt0TqmOEi4BfRVr
JPosmY4uHlujch+AkJU6wouIzYSnVwA5Y9JMmnaWT6bR4ts8Wt+NKFCEHVl4Hjkr2HSmA89BsMwh
lIjykxSIg0fYIdVKvqQxa+wSGId4m5oa3RIde8oaiBADX8OJGTTcFMGM/TpbhLhug3nK2b2c0AMh
ZH7ugTs3mbP6QREXo7FzBDAk3CZHGta749W0QcKeqGRqL2FCRUEncysPruSFBJ5mQZqDUrRkEMGU
8okCP5w/exTUtXeDMLBsZAVJYlyQ8rnPsLwSkIDOHMJma1XlutKUMDdpsFQt+4W3jVm1gpmLyw9V
RA4JTHu+hWGRR8xs8egiFb9qYlZg+fnAnKMsKRXPXcplm6rjVEnABVqocDZdSbpQLWDeCCjPL70J
STpl42fs55+SmqurVIdgH570HLw4egKkHgr8YuyYIieDta/myKTf5NoNmeCoVdZhjmZq4qloB7Ho
kIyHG3kf/LB4vZFOlaESAgNyQ0LKJwJ+hJDlZ4X52FpKbzaucHn2eC8E2g5hauK6PekLRRMBxNnL
tNNGwdUoHkaytoxgWAYB+D8nh0O6SY3U1AZowbJIFYA1UEcqZhpaj2quJfRsWBaSqpFH4T2uy1PZ
fRRaILcgZtqdEp+Tm/te7DLNRdag4mMnBmsWNEQWG1bo/3wrkAkj+QkrWvam+Rs/Miy8kDSoS1hw
m6Awm/5NSLIaovtz52n/eq350Mhko/OoBLFGGocq9jw247t1dfR0CCA1Og3uGF62sUC6tphIVjK5
p/YBgFXl6sQVn6TDXQTKTCA2sPUMT60XFXCjqA9Ssv+s6/GMiGJLXYU16ora6H96vkuaVVP9CwT4
Ob7TUvospedhyyeOsn+oMrm//DHi6g1MPXYDgDeEvQ5HvFLZ+p3Up2Zfi29DDPUm4puSXR4nrG+9
4UAoNcreRvB9uoU3t+aYJl0n5n1TJF9vs2rbmYm8wBUFSfWW1aJQg2gG0JaM5ViM3SvkqxURN8+L
SejQ29nMnXLL6kR4fe0mdNkoU0krYJIfjaX6VqKPuloLt5fPu/sObzqC/Q+x1mLPrXW4gaU37GD1
T+BwVhJl9JlMK8SK3Zh6lRP+i2blJ88B8m/BiVLOjL9kYulMIzhzYZ/ZxpwvNrHv0yyWymyxm9v7
M1klbcxmFddCUONUzm/xNrFtB4NIHCQWR0YtxV68rkjySn2/ZIT7Mr7YKPgvjS6TveOstIHRXobP
Uf84i4c2k4tKm4tEVRFF6X3a4GKqkTcj14MC3vVrbtSVRb/6u3M/tlJFZVtccCQAUrs7va3kTSfv
XmNozhxZhn+9YH7P/JrKayvI6C2y3zOCdTjuvyLkfxldrnCUsuIUBk+zhp4IgOxOGt+TYRt6KBSY
+YWFDoXzJeICYFSTdte9h8jReLyLcJ6kPranYy+6bw92V98KDf3F/gx2UhuCl+ZZvJ4BwVFg9MEf
W6BR0yzAYNWyHLFeqPtUGwfWowpChv41kVp4z/yRzxh6cZ1GqsQ0InMVIupkmUfxPU9f7ihkY9Ql
FEmyZeua1+2dH/Rb5foHlMECcbFIZYeA1m6veQom9txJGFy59V8o3NvHN8OJXyIzyDhnnQmK/whz
ymUvoE4JAk7whFBwMQIYcQVtEflwTeFHS1MWVeztgBn1zHUkjAxxu68QQ2ZdKTl2sdw3bE8SRwFR
tIXe6OilC2MFhHw1B3yJgMze3wSXJ0UI9l19Mgwy+6x8H9R0gnF+7HDluKeiR84m4tCi9BFxvG4d
SeWKSmOjz6T9+Old8lpvFJLcjkIsaLhsUxIITXuMcI4fEY4+7L3j+dRvkQHfISmE+TvPLFOearx2
DywUouLGi8tGTzznPXTg+t/5EzIk0/J23dq/jzjZq99oE+c4P+Xa5Ka6i94TSjos7UjC4o8w2P4Q
wINcAmaQFmzKyad3sLa8qod0LmZR248kXmqRd9BEkU2JlYxvMhR5b3c/wKmCbt9N/TjFyCERXyze
G7YDSEmqWaH73g5SXFIWzL3bDCXjJ/IN+3Vr5+gqF3quY4j8shfshRO6kHFWvYknmClBIFIHuNio
lwPO95czmGygkTUvhDakc9VedQv8tB6gYWRj6X0P8jKWvAMymmvk6qY477XNY0RrQCwwRkBP0Do3
s0owuITeuiyR9+EAQUJf7XiuGG7G60R94mavOAF0CpuhslTJ96HYvRhQ6FZMrJtMWnEjgyY5W0/u
2uUpPFLCFqVgG6hmHarORtSMjeooYPj9z7uhQcZ5HhwvuP/OjVnqge0CRttjejk0iBMUAd9RLjTo
MAyVVNjjCortAyp60PYgv/n6Q7gWgGpkO5CKbdcsyJkLyaaKU+WjZrqVjPPnpZRdW9yE81foFMQ4
Imuy+WxjT17gIpZdAxIsNaebVGivyU7An3IeddMdhlPb/Oug9yw4h6+YKOWDU0/S/9ZZ9eV7SQdR
ZOMVJHtChFFByBvbViK9xeDe7eIKBWOmh7Hhbym3AUOkl/1eiF4BsJ8YP4lJvZfNV8XakHAtiKV8
ayHXDCMn6p4XLOWBHnw6tM2TAUu4HuYAEvdlWjE35vWCCNsD70AMfxUHkxgpnzV7pN8PbaqjLvre
K04Ai3fAJCCdvedbthYzLc82zEUGO9VrYGeJVRIqsmg+m/FbGu5LRY0HVhDxj9pKUpaTS1LbLrLl
VffIWCmVLG5gTFd9yqM4Vtk7jTLVsQPDToq0npBfKzNqpQ5CkAUYFy0hH+xWOFYPXilNwirxpitT
qm/9lhY/v52L4lOwJgU5AMirgAVMVoUoWLPhIVSyc+yo/YKtVjTOALe6D5KqlM0ZZg+hohGd09Qf
1JR7xbSMU/DXji985DYitspxTdeYpnI6u57gOFJRfUKGdplmZgCZ1F/hEqpqtBI6edSyGjOLCX8y
nVh7Zs1sz0a/6be0tU2PCEVZ3sjPgY+a/BBRuDhs+M2eZC/Ya3TYcvydOG5BfTIivZWCSTyBMRYh
1GlXiApFpUrCm/LbeQK6vjhYDqcD7CyjjqyW8h2wwIeqVqko1qCHMjKzKHa+MY/36SowMJEYCXNr
KGqkTJjpQ4gms/Nuz9dFl7mXYCe+IO+/FAtPOg1c2Y+KzI4ztybhfjB97Ktg5giuXEsc7Egp7zTs
m2XVxJBpM1lCOqAQJwDIDugIB5AfS8MTq1jY2aCXK2Os4x2kj6zVmnCHZ91OdWKJdh/O5BvBS3tE
chxOVns4bwsz0ynE5v6h75MkE3lu3jh0AEEOiq2irF9n6czL/6M5VDfkaFjYLU/2WqfUpvL+eHOe
ZjP6FCCe8WMuyt7n+8EOD7wujwxA+vwWtp6SD9FL2VgZo12PrI/mmNLQZrqMdwW72FPey0901LTD
/1nwk/OVHs7k1+5efOXp+2+rpocnnCgL7nP4a+YCvFkC9p+l+HQYRK6Reku58oGx8P1z8yOhIdYc
SuR4HANWbPJQbtIqzv3pKAwqK8x5yItypJDzpieUHVP9FeaPpIw0PzwUmG8+vdSvqstSYrq/iMsi
Ge46azELXCua8F7D8oQzzb6PHfp6RIiJUld3dlNIC6qGl9UK8itDFzDpqdoJYCVQdiRAKy1kpMEW
6ymcagk60rkB6xOU6xqfDJs/KZTuy0xP+32AU2cTPxII28e10bfXO+F5m3CFe3a2AZm/22nHAs+Y
gSZGoMjgLeiAT15hM5fTbcLb0ylzoWUdCjMMQkoQS76Ij/0g0otK6quHyVCKMuULytFuKxnLE1XN
sZJFLolOAtG6E/2UOYikNkoU8t0vCkh7T7RwllXfHVOZzJ1Y9D4P1z6V1RX3ET+2IzMShqbcMk8H
KQOLeQbgNGnHCJIHv1RLGIj1Og/rujNYAbZu+FTkXPB0vZTeRfuzxRkm21T2Pr43W/9GGmNu+BSD
w5HjpUD39Lvv4Qv8w2dY/6DYj0YK9EWTN3mQoKnoyRG4TQDuKB1BCYna+zPo9SXoMSsy33p4cwnz
aJxdrDnQxIW/4qWLG5G0U6JBUayF0bruqzZrEsUMZKzTuCSD1oEt0W2qgpWcWPdUbJgv684MZjFp
aQTYyWmbCneYXEa0/HZI+psYamNPPtX2/manYKZKzRgR6n0QbvBgHgx+BzudHiSXkyRq2X4z54xC
LLSAeNc/978bNwk2RousHcWIw7b089sqmB81vxB4/v3qBdpa5lCr/puTGTWV2sKikD8FKTPFGSqt
Tl5DgfR4k0V8/Iw0D+IN5JfNUMEygSTtBNOoXmLQyTd52ucoUmtnqj5vqsWIYJPbUoPux+LIMigU
19p8XE/L8SKLMM3GhbawdfgqMEmPmbufoSU7B0Rpd2nC+ZsKZczE29hKN8LUcPMqHxTiyo2/GeLY
3uuwQwnRvqRMRspwJrqxXa2M7nCmQv41sCPWQnCvZufotgT0N+Ez0Sy784NjbEsSiLEP2RZLaaBs
dsnik9xF8PJleiYgZWKW/szJMUqJOaZocRLJ+O0JbtH9HT3MJpGdW+J3ThtCBZeqekQhWFDEeqZT
GlqhoYWV6LIij218U51zQ1IWmhlx5fKir68WVFtwVMg2GnYzcoEf0AiuvN2Zl+DtzeUiV9lWB//G
+7vOsWRcs6ss4N9U2HVI4wBu7wsZwgrA1tE3zpoQpQSzyELVsCMdr4vSYvL/m2vABgq8iR9jr9J7
zCKCY86JnZlehAJkGocVR0rHd+IInU4SHRmlmDlu2ujnLMrvz2FKoy1Nv+HuHwFqzLhJw8RXgd4n
A+F5hUjTUwVGKohv7torRCwwngXG/Y8hdm+mffRVq6EhkEkIEUzuZyse0ytxlXtb9ZbdLLscsH5m
g5Tk7KubK9GWkyLYpY2OevhUrLPHgSi189wUvDzPV0KLCFCeAzx+sk6uU73n7zgt7fMzgYDkpvsk
4JgKkF7MDi4EFbc0DQD8bOYp20cQ+4Hfq89Pwl/FvXlXribDVesqZ5thO3Fnyot+UavVsLdboxwz
xfps5bEEyIc28OXLVVuSD4/BbQ2eTTE5gCAdPYfH9eWf+XcDqy4JRwM6S5PcNkbj7McApmzYJvHO
gyyDgk6OmnkqZf2+qOEORMlJis7BI8m8hAmFRbZoJWddfWKdGB4uLR/mPorSo5Qr1QvTtBv4JWEr
Odz0kK5gXVS7HIRSp8GIEuKzMZSqZVGLZt4+xFNpZUbM6SJlEBjGbn2b66r6blqtry91xY62mUTk
tHUnSrwl+Ka2Z3zJTVyzErEQPdifhJYKfPGXW7IzDFYRFYrDBg6wglrr44v5jJ2A6DykrPYbECRw
ny01rQfgq1hBjngfLfub3nt8pGFA+nxVxyH009p3/ZX+x5zk8+DkxBM16WRAsVkdziJETcXGOysD
Jfc/DMVFMSN7kR5uZM7DJoG5AxaugTQRYhSK8cHvopLk0sSbxBpNLwuiKTsj12eZDRCFi3KeSNDW
5aBbHWNRyFcIKMbbXj5AZcYNWA7rL9oSwVQ5WD/X2J5wXOMm1ITTzm2k3ejK2dnGZ+K5MHWcwTm9
3TgYDpdg7xFnv1KeZKMN1TQU0nxDofPYQWipS/fUMTiWGOenzOXNY9KzC6Xaoyq5a+NVSxinED4a
7qRFmKvlP5O727vd0bYpfviWOPPRiyd91Qyiq7FsGwkWHW+KjOWTkxwASzJ8ZBc+TCmhephzmO0a
OSY5p9VUS3kZ/w+XWax08epKVs99nK6WsUpVt6/WebOf8wDSxo0fCuIDo95vq8L6b/1ZZJXn2oOF
BQI41pLDZ9lrfJmmsgbO0xdc0w9pMHQLyazx6AyM8x64cAjsGNMCap2nUGdFPFb5ibe628DriL3N
GkuzGjJcpavNqnOJv5KNOcVMGLJROPjH2WEZ0tL3VYBGRdpVIXdfvtMvkvSwApysNbX9r8G9MCEG
KAPzl2DSkkcHNyPiDqzDON60p+maKskCbBzXoq6GX6xiHT6cXJB3mPxmwoc7alz6xWbd1lpYMoAJ
QpmgOOfkcK5xvlZuy2URYIv8j6GpbDVgH3CiaItD3MGvXyT1XXHqaWUsb4cRTsNBne3pWWF+ssi1
hD4FB5lMgkymrc+XfG/p0ykc1nRuvQe5l2bpcQEUSOv3Yyh0nOfdbWtmKtuurwgztGXGJ773D934
DaAZeFAhN9hEoeVZ2nOcHp/dv1eDuV6ueZa836M2BOz3H5a847r7o1cf94ty7CTLrVnHWr2gqEZv
U2e+E4HliD6Gm7bffpFWC14hkB5kN8qA9jopIT+/E6n2kcJgPb1dohUE8PtZeb/D/EpazsWQRJ7u
2Ix9zoOHpLItFa7hpRuhedWvXB2QT4UmvJC+FmuGRHZDsCftdka+ppgLzP/M7T2zlrig3okqwx2M
4P93XyuY462MoL/sdew5w/wngu0FM+WeEJ5jCCwWDqJ7ydTJ81M51WtiW3OZiYdqgi8Vwb7vr2mG
bKroueTcrGKDW9NPyazZQXRjwTuDKA8ebKTaqfDWQ/FMF7ya5SQ6+gGZ9waFv0HWIu5Z0M2NBwqg
BxVmHvNKeTsbNkywvQQGXZ5LvjZAdW9zCzxYCFOj+PNzqtKstpeOty7DFMDuOrY3eV2GHY0gA2E+
RlGZoc+jmAZpPW4c/6yUKmU5er1ZTdXxg4tuLJTjP4jy0AfdNz/+xXCTRm6rQc7KlXf5xteN8HnV
AwwEYRM9SGmlSzqw7FJECe2wiNLqf2SopQ9Ec1S94HcJWrBnK4ENkTeYNh0KwjnBxijSVyJqgIeu
8VDCVCTxSA665LDG+oK/C8SK8FX8S/RdZQ61tF6AiL92QxQ/EQGorFm7XJzP8B6VBImUoHsLUe0I
eJ9eSJHL3AIpuvxjSco6K4spF5vGnb9uhB1+zBae6vHXBzV+uTQsHJk7JkByrAuAos9mtNpn4YUA
IeXbZnB4HOd0o51/yuvQVVLp0mG/pePY6FKngwO4gGitwcmb4OmdKVJ3+B9Pq69FIWf2pFlPlTm9
qVPHk+hDFh24SnGhJ/zCBHK7XrA8+g9daBwyY3YdbFQTCdPiP4Ig6OrMNkPSnBqdTvW5cJSPp9Vh
w1nJzOQdA3Yx7PirBj2Wr9tlh3goTE9QEMmKaByKT04tKe+Jqxi3Yc0cdmW2bXZwRRE7OXSiK7nK
FrpKd4Z9pMXzA0qNs8gG5BBEQQWFIg0DxJy8nhlTwDBeNgb0aeH8QZAr8qtYA0K444yer+E9vl8S
KEnhRbifT93D40rTHEFzUhfZHeFz5havSuEtbX8hgTVFVAp73b9wBkA3jI7dZBP4c4ZbgOv52pqk
q3tCQspjxhlnUK/HTLGLHVOVHsx5gJbunkJ0ywmG6trjOxAPGRuwqU0PzrRTJtj23d0A9O36Rf7O
g9nQCcIYabETOAyGO8bS9vPO+Pelsoywy+w024ps/rS+oPhqK+91edg87N1PDp+dBC3izvlSQBWD
RYeyp1uxftid47Rv7UZXt3jb4h87dcdew6r41QGBGIaojc+u4cdo3DmTWpt3r2UuYGURG9Flqksq
zehRXnVfZf0VVal0bpEZwu2svtyVl69whOc9y6IQbdqi0o+26bsenrLhfwsFEV/uRoWhweRDkUBl
UcNSYtIEtzS1ZR5MoNddvXSfyrQGrzMN20MLeB+u4XM59tuzs8ZttjMij50bYm+zXUmq2eU/YuMu
ffDFja/YLr1mV8zuFlFTiYrrlMTUrgyyLcBCaEhpEBFz9YDEGOSzmywudk5sIbYb+aDYLLa2oAbt
q8zo42IxqbgMCBnXIZ8l7gg97+A4tb0Qoj915CsK58DAo6nel1ED9ZonI6KtT+mVoAuZHxFD4cOZ
4tAYmH6eWE/qFBVVEhFW/ctJav2BfhnCliDDLN6+8h1dveYktSRdkTZG94m9GfxUE4nAvz8eR6TN
KGhH4W1E//XrSQaYOA7HgFeZ98G53djXOC6AmzxoIamPUFde05iUZ+uuSvkQKLVEwo3eBtgruoqU
LNh2htWdKGDmieLiIUByTjI6DvS/muXjLzno+4vmdZqMvVtZhwYabIaDMSnkXjfHWmXBEzIjoR8j
XtlaoMgjo7m5dgI1g3KdSw49NfHVsuv7c8QV3ehfwHcXPJafxru6s1+xlOE02QAXesRA4q+X6Sbq
8L/f315i0B55qf3iXDNQS3EYBCIsbzS6UiReC6yG6PeHuYPBsyyVF+FzM307jcC8XBWlPtyYDgQT
uOyEnthGNpH6uTIuH+UwnbpCxegKiW8tiptbWNGM8Ije4fNf8dfzDoNeOAHUPXp/FUZHQQf5n+/a
3nGdd6PGT+LYzgioai+BdB7HpISyMkE/Vzw7JLqfSI7OgdNjGJh7/XNBymVim6GFGoZaNFPMlOF2
uDW8qIbB4diMUmxyCqrmn0EgHTXyI6JohJ93akFweFuiclYXoBvnHQjI+HtA/CUftthB0Gfdfpc+
6mIDQmUJBAXQWXtG4IyTuA+za40zMeDvqlld+z797QlkuA+jOqNEs+qG849CL4WvrfLcRihgYY5y
odnSaykavP2Srih2cXYIzqsMuOKSrvIlENsdpvWe8OLH5RlahcZ65r3oraBVK+WMnciUlytetf1C
0bgTcRMAOQbw/T2Aenld+ykE6Oiu/ax7MZZt6Np9zWH4NIzD8IwYC+9h80+I+Ryz0KQP18xAbecz
RpIJv9TA9Xu0DFj6dxaw+I+XS/eELBwgW5yuqhU86aFVdORYSBeSpOHOiELVW/+I2ThKhL0Nmizo
QpvyoalV2cj9MAy89On3rSffk+25wWkG8IhMyl/4uKwBYEwCWSuN2JZf6w5Ht2SEVyu+yxCNl5e1
aDKKAMY2JxsIg4xD1u1b7c2FqgayMztkrsXJcxR6Yj23c81OXRjtkfZNKaX8aLtS9BpbKEBuN6hO
PS3cVsniXn6kl4wYU7RlQPxGApUW95sNuHA+cdV1hKLMJ2Ja4LPxPPM4m/ER63A97ht4oa8iM6kG
KDAWhT6sqKq6e1ep6hD2tCbuX7ysNg8aB1ZcxObzteM4aVyooiaIPSRR7AEPWTADqnb8tEAkgJwj
eTKcHjw5+Jo1pV9+b9buhTzy7lG7Ko5xWOXBVAK3DyRq4TSjz43tD6gC8Pmf8vBZAL/pnj58RS4R
P5eBn732dJRQqxGWehQCLcx1IT1rZjVlfjQ/hHAjCeEUtTS2ihjnTReJN3C5czIvx01EIWOZqkaC
0zOImgjjDp3d0p0I7vdBeSlVkS1IwgonbgcQoQ1bgWoQHy1mETUxpCmdHV10k2fGMf9LmutcO0po
0Cykxl/wQ4yblc76xo42ayk92djoufdD8s8ku64d2k6HEo9oY+jdhzr7+rV2S6BcezInTcNZNP6N
tuaf0FymVna9pG+BR5i4FxUp8qLRFzLqa7+xEgxPwzsFIaO5CebsKSF9May6f1w1wRm7z/MZX9Bn
cB+w0eu1NvMOaCdHpV1mjNYcJZbLRSI6LUWHkZfPg7ye+ortfiC5WYsgeSpxyMneJ7PZ6xuKzfOT
BbQlXFVrju8E9Hb9648HpIp7m+pZgHaBhomhYC402oFjIRSs3/5Xxb7+W/uoqM2TPPyAS2dH9Ddg
Gxg8H7iNI83Bp658UTXqdasa1hVCOMd8XkETt+aufubgrGUu0/rDTfcCXViSVZGbQVa47SOiv5pl
qDYFejagj787vT7Ml0STqsdGB3UhbNns7yfeX1r2AKGgf4tu3knZGbhg3qD/W5gxJ4em3mKW6Oxk
xyReuCX5PE0YO0nCMI1j4FH7MXpMU6K7Q2jg3WIrymYQzginMxLWvMkAPBIeaVDRw4FXT8LvdEpO
vO8EDzMMXRvL8pyYTTFH3vtKYaVdNlZ6lYMtr5CM3GB7OMET/t9FtwuXNR32Knlqr2L4cxj3OCJ6
qk90jbtL2JljlIPVCTZZuHWVJ7DN0LE3NMPM/1XZ8NQF0Ulnq248kzi3Y0UmaGa8yqRQQKHpRP9z
bsMVmGnT/5u/Xtz9+bOLvyG88lBgQeVfFEGfNCIXQnBlycmq6UC3HmRi9nYtxKX1f1GFlkaiCCLy
1JNpr7XfnUtQ06GMNQcDxy4syPq8tA3yaxaz8c5NZxhyYo1/UENs1Y/XHzdewwORCK8v+yiAOK0+
N4kURRFDzin7g3w82Qmd0Au5oG3lgIY2BLyUO0mEMDQlvKBcvFPdDnisIXNYk3YpmIcUCi8b/oaL
spd1bvrlqPRRp3dmgN14BQ7OYQR+xXp2E7likDccN2HNsn7daR7Ro2a+XYTZOwQRyHRWOKn87j8p
pNYCZsNeOKfdh5rPgLeTOf+Q+SKZ9SvylyGjeDRQd4fVkcF3yq77OTYuLw7+MQDNJPu4/fXLYrK/
zfXyMBUhO3fLG8WQRXQeagTGqZCwv4FkyuVkw1zwxgWC7yKFQQ1Dp9yyyiXy1OYAhjD4dxxuP9AO
uoHZFOP6RH/3+7wy2aJgae6Ot9V5UURJD/yafVqOZgpfEHrMVYNMkx27UVNNf8qz6hoxiqu42JDP
urlXQ9Nsk0ocCVG5Zq7BrQ1J89U0I+0A6qhJ7YK6gD65tAMVpPXXEOFVSrsV+zUolIU+R+9gwEQC
IehBtTh42/LreQn7N93wQM6ScA4Ww66D7hUjwUfML+GHnKEWZNQrL12/3nBf57Qyc3AyjIOJvnoL
JEbMsnPn8EEh+QwNMq2w+UgUpyyGY5XaKNkDgHeIFvQqVU/asdPBLZSlyxtDiGI9P+x38epGHG3v
sg0igTdEdcGjb652I7PLa6wCb/BNelgT1PpIROLz7dd9VSxotbS6kUXirgxvSraXyxtduQFQgv69
GuaUHQwxQnBUEB7Fzp/f4lM+uEbCx+eEQqdPTyAXANr4ybfOjZqsRHi6e7Ueb3SCdczXXU038Wak
YH4luynDrcq/beJRVP6/hHcOV4ydbDLXN6Hco+1fs+8jvVVyPU1dwphojxPGsopHvuMseEs7CS8v
ojOz8waI5SSbtfo+BBEhSzQNRFEXkp5myd05ZylFAUPFf1Sb8M7iVeJ713V9WSpKexJG7TPwJu0N
XfrfXKk18Ve/+bCIF9pYSr7pS3OM3SLAqDBBXaj8su6kIvn+SRahkJFsX5mz9GuAuAtSt41DS2Tc
p4H/HzLNX8UZiysZQU9YBZDNpssSQECn17Av8ogrc50lLWqvDZ/vsNQn+gnhvtrtQmH1zErble8y
rQIg2pg+W+750tUCS9DN+pMGoPBQNpPCmnyk0EZpVV7Q8JCiunngD8tlZJeh9XxbW9fLOE//ZRNP
gHKYMBSpeYeKkSeXrGYQzqu+ne1Wbmgbrbt3EigZZD7+T7RhaYh87Gt8Apn7txFmTYHcwYYNBbRA
ejbC46NUMWl5HpRyFkndSXupiXl3WuXQuXn32vCHX0+cdY2IW/Oy1sizacLfXUW7q7RJ2mzPSCVh
bPjVEC5T3V9r0wrfcyIuTez2IXzJ6TbcNTNbEGPxJ7Vi8opUWLSCzPjz8a3ij4JzBCrvqgl6pOkq
DIfXzUtry6yrQwgy4lc1wJhDP9mf31u+o82O/RJlu8H8XM13LSKUxAGar1svqaHOVlOax+ZUqPoN
y3hauFwInfE80nquFy6gaQIthS+LlpGg3RFzJ4iSO5BFr2HIo0ghmsDNlGnJ6Eh1vi7BIPkZBLH6
ownz/Fm7laYeoU48SVdIZw6NieILp485IdGZHaRgleRRhXBBEL+kVaEnBenztCTzOHovxFTaB97K
deUxb9nFc9MupuxD/bnNCyjc4F+N/4U6k4WwSfspSIWH0asXWLlV9d9/qwatPAONQOpijq5VfWmu
0OLJfc0WZEgGTZ8IhSMQLUVppss0D7ta/DqWWb6ySjSJ/0cDjNpJhbZ11I28sPCb1yrTXoQ6PEy7
IQH07bHfLycBG9JvaYPwZaqR+nFYqHE6EbptN43kbTiM3y3URgyjQHb5NZSq0xifKCImxozWNf2B
/G0IcuivbGwBZq19dYWxpcqZ9RDlAF2CqlETVzuEFtDyF0EbVvJTWygAJ+vpt/pLWVE4qbvvAuZ3
uhHDFmWzvKYwKZHhUy5DSx+mZ9+VWQBqo0V38WuLoWpQNMCiQMq+6sJg9ZNJiBhZTv8+bzmkznLu
nGykfqToKeLsTju5E6sJyZPjtAfcm5NngI2T1ts4MBM1KcjpfSL5CFLW6NnTdPIQal0kxpn2G01R
VSTn2ARBVFb3LXY4ieQn0N/nbTD9CPHXKW3GbzNsXb6vLSznn8zbvfy8HRvL2GO7Hhh28cFq6IlZ
ZTv0wsD/7iK6I1G2O7hVO1q5DimqOygS+gCpJYlc2uNaMrkubcCsOYFr7n/7qhTwqgq+uKSRIZK1
xB2O+s9ZYxSaCcKAdLcDj6rai5T4Ec0X339LydB2HyXnkgGvu7b5QepMV/+PwrJUval/3ZQejg2l
7m3EBIyq7ui6TEE250te/YtgxpZz5T2FCfqQx9nIi6XQZKumceB4+/ht4HM5Ln4PKMgezKubJ4dO
luHGW+KsB3zLqMPAB43mKbac0SUbjwz1rOUnk1au9H16EfyoQiFPOD1E7Fnp7wuKumDssZVUXeEj
VdLiyl3xKHRnSn5ZGoBoOZhx77WBWh6N57sbC1p+1/2Cwf5ZLPaR69IVQyk9NmCYxiej2qVDtqMk
h7rs4jn117FGArEslMGM8OpfElVY1ATUdS/cBhP9gmt9EZH16dyhtsItViThcputZBPGbw/Pp5tL
6irA6ypFvs4ZmynOY5qTvzv9J25vgHDtRYK0KclmrN2zne2Vh/APXTU6XiDBmb7O/7Wzji45OM3o
t9Q2OYnRcBLB+06UIXVOkQacRVYIOcxAHpxwbHLTbUGWfwnuz76RnWrQOvvKB2zgIylDZV2GSTRt
lVHiAm9HJP3bk3NiwnowJw3TLuDfRyTqTeZoSBVakpNZLb7OS2oWqb6ckU7BFqnwHKkkn9e1oinU
fWPA+csYOtj7LAEvChhv7Jnv9KYNNKN8NCpULyru3TVbd1+ZfauXF/qDnEj2TauVHcyte6t+UORy
OEYS1Jd+5fdhSbDYg28L1LT1WudAV+14HHzmCxz3Qs7qVqeG8CvXmNlflCpCc+l9vfe7/13h2K+m
6SNQZ79fvzzZvXc/QC4AeyYXVQm3dg4I/jP0gmo40IEwxxyDLgZcfuZVKP8jamEiHyUyKH4EeH9D
ZS9j94qavhP/7gIzTpCGPE3aHtxVsbo+rmlj8gIJTAfrLBu4wNoNvGf9cgAr3ncnZpoy9g8Av0wX
JVum8ACfcvv4yOmPn0HuHvn5o4nTN+E76Ty7UH+YdppFM6PWZGex0tCHr8W6FkCm7hk2IE2goDn/
7SBZfdeNtbQmJgUgveyLAKSTutn9slBfqk6YlwFpmxEf41/vlgc9QU8Cs9AUd0TIOGA2h8dkSGdt
zp/Embd5p9wGo4HuVDiDM3So6sbeQutqC3KhwZg+PHSQ4UaCX2Ifum9VEnn7zShKsPsL4Q6hyTM/
9p5H4y7BZFO3axosDWqoAhvwh/d8qNnJubPwzi41fsXV6uGAjk+m2o2c+1W+QI3JnMnzdNogkUoE
wq0pQMOxBqgEeaTMkzxjIbWACgE3jPweFTJrItwRO42Fgp9bMS1jTmqgDYbjsOYnbKVnIxQJxjXU
lLQhumVDm9Dw7+JiBu1x/GXtPLBB1utLYY73gZ4QEQlEj808rnrNDHturLKPr3HlebjnDFnbWZZo
4bP2LPpu1mrACCyPkcqx/OcfwloIB49FyYidkYUB28ybj4bLHbsl22VFPSVBx3K7d24cRZaXZU9S
me/fm/gg8GZ0yC293uiWWAjCVF3UPJcakZi5mnFLSIRMffCNFlBdE0rFeZTtRl96kR+KuUILIK7a
LtZIqKnE1bIXzb/w0xn4WvZbr4h75314G2vIcPy/+MCAkeiPMjHrjX1plbGpMbjyrrQDhN3foH7r
VPpDeTyBZOKLoXtQwS4f42uqaKbYWGXYYKfpxEkemRB0yXVE1nlebxdFetKXeD06IgEEom1OJfiS
0cBZpsdKsUecryMQrOXZboEFZSZjkaGr6XZtLWfAZoh7WAX3TbGE+rn/0HGrU0RamJ/E9oEvVwDW
WiUt7BSAy2JwcEzSZpoY0re53fjwTN47DF5aOfnjRYPy4ay3Wd9p8RWxctjmh4bjbxrnu5uzoggU
DeMSLuLgwO4U9VvvWMrSFd1qPvmQDF9h1Gw+Xw0iuP0tSYRjySfU/Jq6BjGeQB4B8PqoW6Td+1Xi
GnGjOfaO6oiCfYBAWshWDbcBfnSG339b2AoSfY1KLU+ZaKVksQeaXRRaaxg4l0tVBkaQlr0BKPXt
AiGXKJwF3Ki4LdImwYyAw28IkXKfPrUPcn9Qizax4zdy0LKZ0fy7sMRTm28IkxWfTB5RqXzQ9Gaa
Tea1+ndZlz2D+n5fuIdrOPDuck120Knkp5fCpIgylxV2x1vM25CE54MwkiC9dhQeBJ6zwjWp0Qbd
vvLGVkJtAIpmxsfEloAUMQhcHY1+J2rcL8jilU9JxkKWGfTMTeve3YFcHyg51K/sggKg5GtTgNrW
fohxBedgSkqH2IVT6p8Tfle8KTiGeIscw/Spl1wuentrhGMyrmTfI5QBU1Za0ndomlicnPoNDgct
Y/Zjqhm/2LO0q2Ip8HpIJkmBM5yEI/pEjXFcVTWAntNJb+eWtQMWr8Znkamyf2tdBnvTMyUWIwFx
SEi6X1a18pjg7mbZy32gXGh4NJPHpZDJrXmchK0b49NlPtzH0s3CtxKqPTGGBvWSXiCyJsDPOEOM
i99JNBBDICZaIZA2YAzhzfPNfhok1by74lcTZoGVRcSqp84sHfcMVFGrZ7nQ++GNtAySPbLk5tiy
hl633vf5ku3GdLBQ12TmEMnRAVNINU+WU3N4z2DFD0v0v4mL+yDE7dMBvODzVTwI+2EKsjaoBU3S
fNTegEWbrilJr8Q+9fMGoXlSjPHbMZX5xpXNy+FwnVvWKtNE8BmHm4+s9zHL6e04XX6axLYrMTir
yT3gNJM0MIJL5uk/WdCSlmvtYC0DEa4Bbmvzl1RLU3e0MrW6TUTdpO2YzD9vl0r/eAsZXRMXKt64
Zi2UAjqZybQi0rIpI0tTZr/JtbNDMsDS0VmsJ0zch61GkakKT3/Z1ZEyl03nTv8IbEhSbRk5RyyQ
cO0Czt6Zhdcg4fTgL5uHO4jzS2pqDhF0zAkKK7Iwa62HuFG0LixsIhYmnLtJAMHonofkii0vt8QO
Zz5gzgI3zUIL5MQVq9Mryzp5IWcJM3ZRODlx+laap37gxQMTFA8j9A4RxteVuofeC4jGh7kwJJhR
FqxL7eemeReUvvXvJSmykF5bcIrUqEY6Gt8wm+5+05+KQYHNPQr+YJ7k+EP4ra0uteWPAJ1QJl++
FmOSWgLgxcFoADDa+y+E3IuaCAwLe5yPPAINy2l4vVBLTAZp7SrOQmaEV1MwfBOfRl+i2m3mYM6g
ydC4MYyA39cyKwiwyT0Hxdnuc9E4O3et5uJ7+vVZYVgh/6flQZHi28Hq2xlekp54pJFZvORMXYX0
OZzHY5vHa2gDfY4ZU4f6RTQBdqPst2q8dQeyZ2MJ/Jdf1RGXxSnhH5krskJCJaCVoQMLvS/m1UXc
JAjXOrcsM1/uapCZsFxAiSGkPV282W5VwMAHwTx080NBiK6xZcme4GfO7/JLhQLbdcYeHBITnjYm
mGJBGHIKis5ytuRx8DBOfSiXr0OofAoL/7qeSu72wGaEKw0HXrksee9OZ/ZM12OiZ/ZnNuoMDe9G
XF+XvpCGKqOqlpZ0e8mAPJH8t8uX2wwUEX1OBmOl7E1yRfncklD8HYrNCCYYITsJePFXIPitqJxf
DgJHBihWZmw6IXkqMkC+4hNGH6lmTVrHgPKHgEu3zFE3ggWvzR401lbqzXfAtiy9ZfmBLHwBN1pZ
cuPwB50g6clQa/N6mRMI44i0SwWId4ayHAgS6/4k03BSe9igZSO+ezVpiCRNJk9yBsh9lIfM6dm/
oPthh6F9DzzlzKI0MFwSrwkGAKIsoX0eZ6YQGqJfckgXRnfTFflM/Xnmfwbx3cE/NcZ8j9jjWCFb
4bHqLB2Vym0JWAA9OMoXaF5o7+y9VqBCBXphCkbe/fvWFNsUike9Uyxfd6FDwFWfY0ZXQaZaWIiN
A13Ody9VQdOK5VVr8hPV4jHnXSZTTCD+GbLAX34PhHE9VZk8NoKFSGtJguLrCwHhVeB6dXEQqE8W
o5l0qz4I/JA1o/TsjB1D1T+drE2l8qiODz6qchGAhVMOVP6w7o73+UR/Z/pdLQUBWwjqeL1lpFt0
Gh78SmUjsLSbuSDYEtlQtzxGtYKW2PBJ1g5ASz3hg40ln4GsAKh8EUCmPXBsRcVSARMh352D352c
irI0Tji4o/pXVpbx9+CApJ+ToxrP8+h4gXCer+jSAHx72EW502FaDaALGPOCqJvDMzUV8dejj4uz
P2371HqHyI3M9c7LfWFSk2jIHLZg/GhxXPUO1TtlUcHUlLTsN8s21qjq6cm7U2sS0aW0AJam4rmv
0hWRARkKWbgQLZIwDetA3AZxgDHtbOOlpcNykK46eJ4iuuGBy7UwqJqY4CWxRWeecOn2GWhvfdKc
AkZPB4YTY1+PNh3ffMy8SrWohDJTUxWTxQ0971JgJo9pPFwU2ofbFX95vDSqvtc04CzbXAuxyDWX
3HhLqjXPFI6tszd6DN0onOUs2m/peX71wNVmmnaMVnEEGM6MNvBVOaxUqvTGK/p/OY/l7/yrl4hW
69qldx+ubhl8EAVHJSDtk6bT9mN0BJ3IofEpSgak9th/HwXfbr9Pw6juaM/cEuBDPZEw9jLHaRlt
705Cp5YfBff0J7bE0Y/vg4+mspgZWGC2J2Yh05AjfqJHznBeEFkS6q3Od+uA5M2QmuPyTJeSOLBq
L1HbmW0B0YBNT/8XxJyjcIGLcoOexUIV1Gxo6nTnl9kP0LecdBSurEncqzG+vSK/zUyHvWsr3f7R
/5mn+OUtDRMxQ3IyzBZINw0sk8mixX4pB+2y/4FlXgYLpZ9gcDyj9Zi1haU6ESZxD92tWem4iR/R
oeKBcxp8do2avr5T3+J2AFg5yk7TCBHqEddKf8rXGGzhie/uMl7cPL1K8VA7BTs7nJRrJTNEywE1
Ra+MuYWv5+rEvj6nNFQwNNzk3u76pGcA6NU7bDPr3o4l4UvAuJRmeKrMhIXjK1ChiuvfAQUrZwib
O6GYKT0ooWA++/eEX1+CDxMmWtYESwiGwKovxE7hp5Z05M/p/OXCt3gHPOWNuY3GGrKaOdYnXWEG
xL/5BGnZz3HSodEs5n6McEq+YmPQtlF9vA8j66GWkqHhTF3tu+lMCD4ChOTXnDsZBehHC/HQNteu
ePdqI6CLmS9JwdCWKwyv/0y9c/8UsVrMyd4fD+8sWgCcBvJaOcPbimJzB6r3Et3ntsrcBlWqZw2W
qe23uFFTpJUWi845QThHiTMfF8dMyz8Rt6R3mA4dZLapnvAqR1k4WBG2WeO6mYLRmxbqWw5gM/gh
PdueRPoC6/bBBDNX2NV86ZrodDp/msAFrx3zqjrdol3JCi6Vd8ErvtSZ/X3wn8llfpkjDyQzFu9D
u9+KvJegHI2b+MBbONxUn0JQVNI6VROSTEU33X+I36xb3Ot2TYz10NW5MLsXWsFniVJ8+POSOJK5
craKIuxoAJOWa6WbxqDijQdQjTcsztcFlOHit0pMQfLJzsQH9zyGGlS3kbmHmU+NQUrAnuO5TvJu
aFjjpQfE26TpmHUES4OcOiGMlGxHiGehYnQ/tOzDEqNpV6FPuuth2slTIp9Kmw9h+DvBoqcN4F5S
gdg5RKcJ77HIJkrri5OlskrQLW0MBzz3sETcYr5EzZXuP8qdj3J1EnDu3z8+h7hUB/LSaVmd28bh
XhdHeQpr04CqJIDxUGoxPR/BeFKTsPGI/7+z91inZwhWpfRa6BlnNr80CYRgJUmJoKx56OkovXhY
XYEsoB7ILdlUdjr5DCWf70+97EPwL+N9VOd1+SVU4NHY45y1POkgkPi88o1wDdO98rFgah/ASoKw
biFaxGH7hCNLvmuWpV6iN17OQSQQnRZAirSGe+svLhun/nq8PTT7p3U+P5yoPHEwcT4krCL9JETK
mY3bvAYgESgp4Vt9jgwhBo8hjgcuXcjBuUvEoEf49zmTrbNj3gDFCgLD+WAR8wFmOWN38+gSACxL
3ovvNhCoq6eUe6twLsk71cpnNGC6b7WZWqf21j/DR1cWu2leOEm1Q3lmeV+8ZG3He4lGfhTI7GlE
nTKxX0Cy2KZEkd4tNDFXlnZ/9iAyjugdFnzKT1kDrQ0lHsVek3PSrCPFrDTnIA4u/7KAwIccnbZJ
Rvq6jZdX9qwM7CLWttfwbf8LAMpqWqSz97zxSuHRqOzbiQwZEdUvbuDe0Ry0HCJ1auQemz0uwiTh
LuCeJi6bNlr5Sx5O2TcOeZFX9wqTsCOV4x4pNSkVenVNbODkfl6aRoDoESajv5hq/SmvqtvAkE1s
Yw4Mu2ZgGqBpBX/cklXjwJNcdTuFg1Olk9+AQtaH5JLpP7vvWNJCUxeCtfAd5LDRQFnAflyZNAcD
6t3uOJvoRo90tP/skW950b3LfN2J5f/F2atIaAJ3n3uArWlo5QkU9Bg7fBZHg60MwJwaCBefTK5A
GA73JNAIPRuzaUNwW0P4lBQgyWq8Wse2ezN64vu+iwo6gGXlYb/l2ZdJ7gwt6YeezSsh3Wf4RME4
0ZEcgDD/Mg37USpkPeNCIU9FaywTuCK2VMZCDiUlqN0bNXZjvTOgICY7CdkbA9PJiqnKA5kLLEPo
k4qkJVipZq2sJ2uUsj/Cqa3g6Pfn9I234CJ9h9Rob/dIhhReWXx3aEY4wiyKjaKOwJL5EuN4nOn4
Y9rbTyR10aSOazTZ9xuVInB29VR5e+XHw4A2WIgatxIqHDVNX70QfNsU+lzivBJV78DA3QF97EeX
Z4/ELEWXjOtngTOzHXLN84gJYGRoYU5cEaFuCIZR5X6JOQcbma8KMnC2Rav0oJueE60uUaBkx24T
HgSkR3v2MH91Wpn8ZvA0HAF/InUz4Is31T0ckyghmzpB+2IEb1PaCA7O6tkECYdKody/DNLlar+Z
yrogZdEfEh9HIiwUIfDcI1jSCXGNW4uhCO/dUd5V6CtY+pgBCLVyHL1c3KU6Kj1MKpwZbt5qsW2n
VdzIOYeehnCHeCjZu9X7Tt032ekMS6MNg5xiGFTLfujvqqr1NJGPYf1lIgtsknZpWuGVuZ6C4ZEn
dPwfdIyPRUFVuwn9pVSuMPQITNo0wlOFACehFInfmdc6dP2768BWFWgi0WbE+tScdXXR+SL0cdak
lv1tJR9pih3E6PM2jdsjbiJ1+pozgFIAFfFDI2DM7SiS3mBJ8u60dhR0fpW28YXxRVIe76/gHUR9
l+59VDhuH2Ya/7ZBpoT3rdNzV9D0B2g7Uet62f2FZDPvZuJBU4oSpgbg7zJoKi2Ot1UVNzHmfXJJ
n8oGRlczRi6w/enrX6fXEqoT+xo9xffBgKO63gSyLO8cUHgobA5kPGylNOLWUrfT7WHxAg/2TWQD
D6a6SRhBfKBCGexbxiUraJg5J06UO9/8jtilxwUPGZqqj0ZHBdNOOYVEn6SmvRywIMG4B5QQN8/D
LvoThK200+hWOBbtwnaXBpTVpfcNbjFY2rd5F8fjXH0haEmiutaCQNqCa2vf6SrE8mNCJM0F4QXX
K/REZUYUISdJwJjkZ0us5vOrIblrcyuZiF/nGq+PplRrFI8n1FRmGw9EvM/AEiHM3guPvn0S/jip
WQp6ePj3dsrfCuCb41KR6HqZCQ1H+0h2iqw4/5eYVjif84+0Wj03dF4KrIPLJsvaNxCDdlAJlYmg
XJUMXoVBCiXrexfCYF8pIdD2g77jR6k8oFSGh+Cyv4oQnX5G1XCrD4fPztKXrfN0L9s7CCEOXDVV
bqoffSKSfPtXvJ1kU33lQrKw5mksz9stYcXxsnHXNbO3cvFPbtSnwOpEWXoq+LJJaSX1ny1wPTKY
LXIWDT/Fi4zqiJ+3SGK3W6IPLx7K5z9QjGebgkn8LjQwr25o1Uw+I3m9Wq1+nsxEDUwcWBqYKhYY
4Sx4UxhB7kaRXtnpgdEOGlT/4HCUN+jWjpR9QVbwIlij6nEn7j/3pD4Xhib9WDiLKTAhugUBY8bD
6/ZrlLveVLL2RZmhDGSInucN0mW4lmjJ10lrfSpX0ACL/M4/bM4+0dpzQ8YAmK9NJe5JzwvP/Os+
Hl3hVIlvPECLExoGX6V9aRfA85wTcq0GMLRnip84Ar/yYqfcz6nHIlkCMJJaFLYiTsPoZRIpBqgt
hH1DlMTnagJA3DNCzwayVCESbQibC862xicxEhSkgelXeJu4fe/M/vpiGZIVSvtDiqJ4zaja0pH/
50tpTWKCzhb/bYXL6bgtTfh7mf82PAmA7x0/F8iBCeniurb/B6BUARD0jXm1NyE4jzbtPKv3T/lD
NsaTOD/wgGnJ19Egqf2zYKALlWr2i/bSeNbzcpFgdlZdftAN2deMkNAcAI5LkLmxK2EHI8MzLDgO
kakuINvlZZmF1pECAjwO0E7ifzQNsqK4gXLewB4mDRu1lw+3Q0GoPiEmeY5QNvazi19pCRNIHOSr
kuswXVJD4+veTQ0TsN2lVnGi41xzZruVbpWdGAsojIGSFSAvvbZJym7bk9zOq2/lwJ8wmpWTnkCz
oL4Hc+k34RUSL96z7VNFEvdi+F5ebM4ElB1i/ArJBtpPmUyN5/vS9NGK+NvZIhjUC3rKQCv3GeLp
3zSm0SGFsg9y0ufLijJd0xTiERpiFlKnWiuu4hakxmewWxfsvjscyQc294q+LgLQY5XHYFPzmi8Q
PPPUjel3T5FhmKZBllVhUnnZ+ATmFaf38gOPrHA8qE7dKUQq3qI96XbWry+rrY7Qo049nvrQA5W4
DZu3/wysW/Mh+LQ4ySIykPHXQoq0yk+kZZq9YoPqB4aeBiDl69AcNepR75HtUauHoMYqo/BMlaBx
rFUC9JmbrBAPCwe9QyU0fzo4dww427bvltlASvCLYpBWiNXXye4cBhf1hxoGNuOT0zlSmPzIELIP
aovw/lr0iD1vMJ117W5llr05gCYzUA1ySh/efgYLrN3TqrVSnwCD92CadVWKRMgA7x9XVs8KS31c
ZltYYedzUf7K86yyQ4NnMH8jGxpBdtOJ6S+kp4nRQXTmataw1mvGfY3jq1knVessNSrWBT7/2D7Z
XDI96+YvNDiZueMKLoPbT5tha0RlooA+h2l4Hp+DhTHCxYKCoES/sjvKusYJxL3PIvsvqEJsUg61
c9vSwRj99r3BaUBil1jI5l0FLEcKzI9cxju35yG1YyYrna0kFiMudb0uVLKwW+u83PSAQ+yC2CsN
4HJdFy9+tIOb+P6WaBmYY77nW4ytVFemoYEBU6i06c6acp6K+EXlL7h+6xntjVQBiRBnF7tzS5Ap
GVl6l5DUks0ObQsBGId2R4aKD/x/83VoavWSvI+cGm4BFdDl/1O4NmONzFI/i3H3NV9xk6EZDLyO
EA4RQfBM314vQWmq463GsUPaIQQqrEZnP4BslGT00zQRNiQYi3njsVpjnWy4urUM6uATlrwZh9pQ
zDfNcEZzR+fapTkd1F8uYNjJCbnL9bYAkgjHIAb4S43b5xZdrFX7w2IlzywYNGVKRkz7SQshNBy8
RgdtZk03x4YZQ9759uvSOwyOSVe4G22wnlMxipVTPG9tIP3J3k1TJAICDNcJvIWQ7ut6woBdDZex
DhjJp/hSSk1nF+nWddbhZz653Wgn7ay/ojOfXlb+vinLw3hrccXIWA+gJfYKnbWm7kJSCjbuLgmv
9/zWTmyufO/NaLN3PGZrLEVs0+i1JyPKhZFCZKFuvJEo5651f1eT/I92+lcz7tzcDdkGC444uT1p
Q4tl7qw/Qn62BchNMdph15283gI0juNYkxL5ue3n+UEUb3NcV0m2O57F6BJv+a09naxIxLfI+3h1
t+61kwTURfajIX7PrB7qu1FagxD9T7DK9ivRmxU6TKu+uV6MU0UtHbw9Z6WQ3QK56L/Exy01d6HC
WBvTRQItFjHCd+T+3ENAgsDlZX5i7JMMF38bQeNRkhOAyCLWobwxvPtRy33YoYPEr0bgRt97cyI4
Z1RMZeRsL5pqSkh3+uoKOuLzv7ZtPYbUH2/V95rn/vumKj2a/Qmx/SCchfc/mSaS9rdeo6C2zpED
ZdVgMZuGBe/DWOIWUrJJavS4Om63gLihC/RNul1v6R5OXakxLYKqcG+EQvXq9vihf8vRZvXa7AYe
0byKfcDFtDNU9Og9Ewnpr+fspkUX6nRd/fOk4/ZWJ80Z+BHgv3LqKsCd438qWv/yT26nocxRb4+4
gtd08QWz5bEL/Dqu2tWs2u5ecQAOHDn2/SdtvYPe3A3Azo1UUaW3UCBIJTqVmNT+bc7JqdCFtT+5
RnCKDWvp9GsgsUiMhXxNTcyFvA5keR4RlvzvF4Qs4ibOg/o4WOimb22iyWPAo2lCPING5BxUQAGA
NfaoQhjDnE46ZS9wXF1jXOVwZCtcasQgrLRYhfCoeYUGPSa93S4fzg21fE729ahv1FNJQdtivxeR
5l8qkdqPnFMbc561L4fXm1O1DOwyjixsTeil2F5yz/m17SIxDJQ/Oa5N5KC67ePBexqXVLFYs1Xm
0LitVCgNIp6AIJZ8lYkoQTpnTJy7pSmIpL06Zs+ivLCt88kl8M/P25r2pmthGVJGMSrYJy4NfEbJ
HumWpjzkBZUJ+wVYOse/h00us3fVhXt8Lkizg6N38fvWRcZheoTDUx0KyPNdxq6LeIihPCiRzKX8
TuiRGnmvzlt9a09uWrJVqxuxKI+j2uuxa8kyOTB1CTZlMuHFMjr0JF1H14u3hJCZz6j8roC4TISw
mYQybTmf+bwKR/2aeO0FxP/aQ67OkEZGLz23SEp7485R0Z/lPJd+OpdCNAJpv6bB+Z+xBSQh9iPv
JP6oGXAyRIRPCKh883flppJNtNief69aK8GROtVD4+ohgT9uSIRhENuLP3wOz9fwFzr4MveenvoD
U8t3MlINQyX0pKbbs4113nJQyCmqyw9uPie9mzSX4VQ8Pv5olvagoGvOUoVDXeG/1IJrYz2xNQwY
nHtuP2gD+5Hb9Ml6OM990r0qhk/Q8DHHPqL77S8tS3sCGBfM/jYhByhzTM0Oc+UXR6FCQziTGdtC
KvJlAm1gvNK6G1prJZ0VhTNBMiulobEhQq508dLcggtZ2H6uCmMV4q3A16TUns9fpUvIjlzasR19
EJYdlNlfqaFF479TtrM6C1rvyeZ7rWYG5ovDWVeuahEuwTau1uZSUngR2F+bSH8Y+uvwQdItmHLv
eRw5HHgIuVvZOOM7Ol7oOMxrQWTacbF2Tuw324qXSgcf8gabAPcVU4AhhAyYbVNKK6/I/235tPWR
d2a5NVZtmANLqP6Gvrj2UAcDLvLH2JNmlUcO7EdrGrDulRVfM3ggctCkB/G6t0ahUPzKXEKhwr8K
A5XPt41EqZAHSqx1LbRqRA4HaL3Y0+tFG1PJ/QZsOOBTEqVVCUvxcKgjovxyZ1/Wvso/s1aDsXUl
5rSW0ynELVbX80a1X0C2pJh8z8XxRQ1gMmVi3fpTynrow2pv2dZPXOquSqsxuvxxbUUL1PuBy1yR
is1aMzfbXrQGdgSEtDkBlol3CLk4vx8HG+mDLql5giQdU1KFWFPRNFBSw96GAfGWI2uZGDltCEH3
2mgZuOjyx1SGlHJJ/A7AR97MMvxVd3lMKnENJ/erhxFW+ghmMZ7T+DfF13jGb2wpS1MAX9KEARnq
DQrkvBMQgT7XX+piGbl+QX0YqeFkMGqUj+TdLvtPSJ6YUMPI/bcxwDC6rljUwaok0yYGVMGhIKFD
DVIGifVSBtoT4n5vqx6j6Xwv8WUQOZXxi0RkwTZtuDPn1coKHF6Bji0i5/eCP151KpJT4YlZAYV+
yHn22aPc2x0HLEYKBtqNjxrIvBGsb/Y3AO//kY2b4T9OcN76SmopF9kcODRDhxnrzB8cSH4OSg3b
56YNRytRS/5pv1wvbb6eG6+mibfE7MEMSLO07nlQJhXfpFDUYIfcOdjZGFAYJ3VryXFQXciAa47k
uLl438Drl0AdbT0TmcVCqszctInLb62t8zfGohv4DXs/jp9TQgOblPyXrCHoah7QastEuAZAjowV
x3MWPckMR4nP3P4N6D50o8ZCXppe9+fGpFaKmNmWn8CH0ldBj9QB2007E1/h9YqypLtOdZGWgzev
JvGNqjFu9NU7Bmh96aI+Z5xn88OZQ5XV2i/+ZqfjiRYdhqsGvUHakDp8cekBSfloG/bm8c77cl8Z
OEO9mG7g9BGPX0VC2QuWWqPqMx7h9uaheOI4CHviO4VW7teF+eWsJVOpnnilMdPDqjACo27bb+WB
WWEV7ZoNYryIUDpB8E0HpYFwC/DRFu/rAN8i2NRgSdkP3/LKUnd7xSfu/98i3W7S91DZ8qM8/isA
Mi2yCiLWNKlEK0bARB6cH3xCLQiBowP29wqMrTeuzlpUtBIYNb3IqApcjR+BfUEYhHw7eWrTDp1o
DVNwuIfeOcz6inUFCgQuA9dbUnjF5mXF+unjcuAtleuJdH8uES9voCMxyhth6j0CE2VpQwEmfnWA
LvJi8fIgh0TNbAFLNugKvnxKm5Jo1srvdr547V/ERVYMw7SP9GKnptZtLrtU8CFSwhUG1H1Cz3Uj
94w/xZXM1cxXD8rYyA7q5kYlwVlGISM1mIqbRfol+A0Da4dlNovIyWPWzoo/TdwIZ3G9qOFXCvoV
lUYQLLH90afKlnWFYI+G1L8hv08ziVXcQSU1pH5FDflNY07a5rPwqtQBwEiz1zbvyIrhR28y+z/m
477ZrW2EJpf/XF7I8WkzuXPFeAwSpy7EPWt9QMYC4+dxk94/CsUFmV6wH+xTu0XK0hXDokOG/A1i
c55HZ77fyKdYecEBKFwHO1pX41N526ztNARz8+MPhhFEMhKLes06NQHQs9Q5v0I39mJ9l7FEeWlI
mgE87N7NcK39c6BMjHknb7KGrzHS4wpLGL3/jq+LCSF9B6M+FKuzu+/nRZgceAam9kRjdFHyDPGb
HzZXH3Fm3UjnFq5CqBQJMuUwTEsIKCnRFKXnNCacuUPVJgnZVHVA6G2jLJjpGPYPr0zGt2Em33ZB
O4yJXILOvHI3NjG6VQOBCUjQi5vkvlxHOrcyuS4NnrBgFRWZ31cYMc7TFHLnlBYTIWDyje0olyH9
mM+JgggjOtshWSmb9YvcYNu92DOAV8wbGquRuehXra0zFIwtYj6+VZHZfhbMF3AvoTRkJ7ZXf5qd
sXpXl6KrSrQ8wyCM4DFMFbOSIrZmdo+xjxGQk26V3K4hT9oeEqa0jm1euBFC8HnxmSfzvg4y7b2w
lxI29/6JjXJ+dQin3lASMRjgf2q+JQX7L+T2j3mnoPbWga+Yza+BCI0NElXKuvhvmrIaXOK1cMZo
sdTY9cl8C83dNWqQyJD0ilWjit3S5sVqVmIYgx9KoHGSjVL2+x8DNa3MLxQXPPGrpEGXyNmSWaJm
dT58kHZNTTsUOkTUh+PR5YHjqcAJGrdn0NyFtFBxTdTDIhfs6D4TyuORBtq1OK9E7Pe9T3XL4TFD
v5mSoCKg3sboxfIKc6QJSa05DjBEl7I7WbIOXdR53U57DcJh/M/1WIL7kee2jZiH7BFfRJWM8Am1
Qc/cYmaSsHPP6wBms/B2WFl9hZP+lkUQ6nFPMqYzRqsZi5SJiMO59kl6V2+50PEdtEZFgSclJHOO
gB1Fc+8WqfehL8dMBP7vBAGWgB5I1xgRPM6ETb1THK/bwXyaDNb+R77ZscKzWv7vG7ezX3juzRBT
+6DFnAptIYMFZPz4Am5rzUpZJof1YG1JVJqv25Zo/tPDrOY2Q6SVQzs5veVI6R5+gaKrHtQ0/+fW
2JLc8QD+XP5r/2ZJMvqBAE9fNCdV/rptPIq02g4QAoP+iixq5Pe+TxiN45DCghjMlC23PZDUkRQ2
hOjTPwzbUIOmtPyM/EitpknKj5PgOJ3Kjg+FI/vHo5ana9lpp63nybIe4IbgC7xNkD+DHpCZgN2t
pOqHA5v35BD49c2nPjdjLoIe2/MHLxxFAB3Ef5/k5olnoXcA2/ZNx946UoZSFUGgCEBNoL54yKxL
4CDevOk7zJKXMeLL278o+LwgKpuCuZaL9u4q9/n6JHQvIcMvZw1B82R+3ulwn1bNGJd35724CWFA
MIRNOMDZhtbHYPwaijn0OYcZDBjp4na3sqn34bnQ/ohxnpyBLrE+mUG1JRpha7RGeuYprlOl+Rqu
XdeaGTl6tipP7IvSsb8MiBzWCNB578L6nKA6ptySmiHvzPzEBUn7y8qaRpXSzHmrq9/SL/yEBVei
tWg8mDwSLAuZdJ3I4S8hDk5XCCU6+78DpRu6/fZMupm8rA1DA95G8Hh5TZmOOpe5TXqgxUlBLnX8
v57s19vzEYaHgdDvb298w1HjAuq2Txs60T+NtRrAJRUb0ieM1Jdb3UWpIPQGULCEBRgiE9nzO7z7
dXwQErc2AGDgdlnLUnePiFu/XyvR0cnbIA3aGDAJkM5Py/Uxg27siJzLoWyijGBCxK+Wo0fLFnHN
d0DIPFSSKEwlTfIxMitwf6G2Bwq5mbMm1Pk8IUphy+K7uvIKaXSQCt+UCp0q2zq+Ke7iwM0VFypY
GhT+XhXwSWowQMA9VFjcp+mD95sBTCThOYYgEJUGhsziVe5Jiihy5yh6A1IDFnrHAL+xshqruO1D
qUjUoMglZSWXg/Lue2nO84ssnkTXByIfjQz2xy2dmfxYP8dzuvb+rLl4Bmf+hD0HYKhWkjyZIzhX
uv3jZ9BSp56J4mwXMoCvzzBu7+gRDPeKMkA0ujbrCqQs3VZi1vhY4HvldjkywwC0AymsSICEwmE6
+bMs+qh1BD3jD8CPM+b14dFwpbhlH2bvX++ag5hPEbD5EdgYAka5PpzU6chdXW+JafjoobXG+0Ru
xBFY1pHZQs8OejYFgFd5Ptk/kKa5WU+D0Tqy43k0Asdpqg2aUmsEvjWBgxKxvEjWs5XAy03ldT+t
DcRxo44jquTlWvl9+AfEiXNlfj2DX34emKe9z0KvHSqjIE3uh/4ceG9UsX8TH0WPiS6v2+kVF8YD
WyKJhpl5HhyfxLpeWWeB81X9mZ5pTf9nGagPDt1wRgIhooDLRbU0AcvEO/ipdKLtQNd/qU2XqG07
npaBtKi7dNmqH9OY9fzcuagh9zZ9n0wn+MdCtmaBqnZRjgFL43Nj5Za2LsI8cAb/Ql4Px+PET75E
LZHtopNb2Jct7oYR0DM0Th5EzY1SgUaG4I40KJgT0peg2liae250cmPDL4FqMX1Xf+O1dP0kUbD2
/F0DSyGISYq4Wa9dtjpSYhYsgT2TP+EBIdHE3r3yqrsBb09k7412JJARx/928mAx8sS3oD+2xw1+
jCRuSMWiSKx/1lptnNedWJ8eDtVYLV1uPVLQ320v4GowQTi6Fb6H0wzYDTnHAGoT1uyMtfsXGaEc
euqgynFk68JP8awBOaAeaL0kIcKdnMsahmis2g9O7eIHhn/Pt0tV5X9cxEz4dT7nhTg0PNYbCPrL
eH3xzdh3n8sNHpEVTDPBrvUvFBNZfs3RgnhGPLa4sxxAXuEwf0Wym7oQKJyDQ3Gi+CEDQqDPG0XL
13/MLW5rOEdrvi7Gj1PBKHlyQd38dl+eK9iLTtWI6SPy62RcfrYPaBjOhdijCg9bymNefu1GJRkP
WSkHGDRNYp0oW9xQkp57NBkTfk5XhS7o5eOK1/x9qnu5p1OFfw8kKGOAJps1Jaol67Gy9P8uJ7Po
R9HAlIz20ZQ0m6gEFbfO8nDCqf+lDKFcrFaAwPsphvPxvFVtxuSYevh9vA67X0d3rbnuorZBCx6A
T25gn9mdWjKFWB0nLXgZYDvexwmhgm9rkB/E4aqt2QmIbu9Oftj1dcsbDCFHGhmeZoHs4fgCC7q7
LU6ki7+8i5ZOPLe+HLBinh6E29EBFb6fUKL26LjXinD6ri6KGxn8iULpn+/g5EUiEvI7eqF/XhxP
a5aNerd0fdwEruRnHkNbKqESJQaMeE5h4IdFtUzi0NJZ/KDIL8f649jrdaE82kBnB0xJaXRFmbZ3
FJxP4JG7X3o44kmnl6LN9rDswat0TPxpGFeZhzx4zSoG0tmyju5iRLDv5MLxYlBmDny8EX1GMZyn
fU/Tb9b8jsqMGVlz27SojaRRAsEmgGwkeRLoPUqfJ57iyDlQpLxtD80a1oPHdXeO4+iWFZLaMx0u
naUFfd8QwFsgIHNsB9b87bGBql4C1cb9xINuHuluPxwKegUD498srzXI9qhE+cfGmD5RXmYWvqys
j+gh3F8sJAYLqA3ULUg+sui4+7ZhCbQEi3E1LtlSI/GVLYFBPA03jolWp0S1YBHa2It6/jLt0nJm
+GrVuSALMkkqwsbTMNekV1HsBg2t7LFJS8nOJqs1P3V3x4aMInKX1y93uCvkeB4KxHu0BZEYzd25
eiusgBugcZq9ISHgXboypRsHXVcv+uyuZEVR5pqpwwAkC8QGzaZPrfiO97xnt+zv4l/1eOFA2SUm
EHhfjAFLlNsm7IGQmYJnXbdqVnlazY4kQy8bxPEFpqQ0xxkUU4reHr/jvU9PdpL03LfibIuWXAuE
jHyMh2a+VPFBmF8Zcv6aVIsHDXkeSloKkn9DFibdjAjzW9HwFPpxdsuxCtOCKVbBK4fh4XAQG7FO
XiIyL27Mun/bqyxKolhRPejcGR+KzpuzPMuAqBg4z9zbSXwcBLbgJHwufzXEXhl/fQMFqisPFLdK
ctiKPp49PfIGEnv2B1g5ylcqbrwUP4HnnW18zx7UuAF+DIccPRQcaauQn+tXveeJGroJtuGJ4X0M
tu0BpOSFX7yYtM5oqOwd+EMreO8DKl7IS2lqzspXSvfd8WLRg3JxjvsD+e86gEbGw8VNd2thbcXt
TZIEdxU58hOd72wuqHqPdwuYX6ODqskakiekFhi700rPfldI9UklV12sMpN40qigrJLjDwSNESVu
EP0gfE6TnBA6qiY6nbOeWeKlJ8paMRYCjN8gbq1pEx6G4O3VJYNl+yp1XhFh2IkOJvUVgA2Jkg6k
z7BGuVYP+d2FFxlS+yjYD/ipcDPChaeysCh4KevL4o4amB9O9XihozqG63AzhzfbJ7gkPzOFnU97
NzLYC+XrsKMci3B8GN+S6Xku7/Wdt/ql9F/YcLfKwnnv8j6N7TSUANvSE/2Y/3ln+5fEl5fGMzrd
XCJauTjrGqWO9rQaz9cfJOrAUfzX/sRNW3PhwatMYawMkZ7Ew/Gapo67KOgCqR7d5Y9YIiyXJsmZ
8fFNFZIDepObbjX5xVeEIyJ6LxG551wty01aiB1l4w5Z1/CUBVf0+5gDFO06G2/EQD/RolRQ93at
LURNORJxlKIUP0plf5ZzuGDGqN82zjg+KtH0DGvxhLxz6SQWNUrXiQUSDdGOlfk8lnulHJBfv+Wz
uFivICzlGSwk8p0sUiwN4nrFdEhfrL9eEPKvIYOCqY6bp0uQFN+pNi/X7AdG+3JdpHMcSoj00xz5
GqqU/gSt5HTisAnpkz5yfXb2iFUfQFm8HzvH9GPGsJ7P+pW+W/LjJUfuGNNnNIZB/vBDb292dJHl
dy/n6Ae+sq+3CEne316wAMRGsB6kTzBCX/k2VHZlrznWqF9FFJnJjuIwszAGoT4f6H9koZ212awE
2j9dHQU2v4GvFARisbEIzHvvMg76CDCTze00yjG7v5hHjL9gWcS0iW1/jnTBNoCYcqkWFRtHf0OH
saY/g/PUdaOve39pInZ+w5oRYeMw1jymzUSzzlpW5owcstdLsgzZknYf/9TL4DDRZ51QRbD/aREi
Nr52eJCZ0KEjipqCnOAlSLoR9VJWWKdKalUmBI5CpZWoeaCpyft2bAGLcPHHHHRJY6thXuilePfV
VcOJHhn3WKiY9N8p2UvtzbmTmJC0cvPe/TOXYbCzLv9cQmJnSiG1Bn3rNzruh+iad6S4F3knHEXw
hhWl5IWzqGtLWwUj3mG1zMksBApuiFRq/eHYox7zGqRstYtZAyyt6x8vrc/XZd1PoNsPDMicBQx8
PcfB9d526cfm3T8IhHGp0HPIZe7+Fs8mTBN0Tb9AFvOwsXvSYA8cQdc9NqIeMgXaDfvm7HyQJrb7
t5aGWby5suToXfjMVwIYgPoCi5nv+tg22e8diMiU2PfgyUAMbTjW8x/neSRrEQPm7DR7M1P+2MlL
0xQkqzyIOJFm/jaNYX0q0Je2VDDd23tr/KQwOsGmjNRzYiXMfjB28HS88uQI7zX6kkPsvSUQcQZ3
2H10Nf5TFdmtro685qvG2rMMVc/aa+b3oyeN5pbGbNB0PyYyhYpjKV3cSGyXjCusKiLA2nSPhIhc
trR3d8BYPIoP/NBkZd9ORaLpLf823F5gndEhNngKfXQdwMd0ygLl9NdhJyiQNhuXCRITnnzA26Sh
VZI98qDLb3gA0W3a2m5Np+YQeGkYMLW8YCzN+bcVlCyvKNfpjdhSYW+Gy2Ys9gm8lDDB55L10fW3
QHWN59qwcjViUW8k7fophdjYpY6ppn/2MSNROUZAYTAPR4JO0DkbVFv0AC5DlwmoST3x5oo7dxQh
7/YTrEM4x5G8SLwbXppfMflX3Q3HU8VWH2V9IOwrqgCn/8GDm4fPAIhca8nVbQRseSLE1YF5eJNR
K4GykilS+gaeAnfOczY0WpzOj/11r/eeC6OzcB7kNrnbvDwpG/rNrn3t6+/hV0RrPJxFlvGSqXfk
Q8qY2LSz5NcfAUdgvnJH7nj7KHw8ASjdPDXG+BVchQHGbiEZKIG2eOCKbo2MrJPmwOkMaeAgdZ6/
npeQNsDwlosZbKQiYr/C7Cy9gwZpZIjsanxzvWks24Xoqh4MtqkvgcEtlpA57HeaLBrmZ/4ceIE5
0//qBRyYI0OTJ5x6NxBNGW6lkutypaDugnsg4fyf8DWp4BesMAXOGOr6xwKp6dnkecAejuLvnwab
I5cYdslrl9v8FbFQ0gX3V3xDpLNuxOgpSyxnMDvq6Hkm5Hcq+nWb//3HfBGjOhByC3/faC9ADMrp
mR7SrL+P08UQSiLjsE6K+w80y4pK8LZAssQrT/IWtGmFQkUF8waH1TU6Xd65JYLjv6qfM4j9iY3b
gy8kah0k5OOUSUlbTeSYJFPnKMKAaNfEZV/9gcx7uj02+8SWT2eZXVWOk0DwpTiGiFHirkEoIwEB
TqBfGdBLcgOubJbrY76ykK2EqdPsz7rb4lix9f7Qn9W7PdQUBSo0HXXYWIdJn0xL+e7JOA2J5rM0
y7ea0gYDw+bfCjgghAmFjFeqt8cx00WiDLjeTCajGkSd7ictFPorl8BnE+octxHzee71SCXuZRM0
o7q/ztIm6aEM4gQH1h/7tJOtkwuxpRSlyGDgBIMiOJyc/8o2TZgnaPMQ0iHxlHCmW67RDOa3CwWP
mgb4AT3zkbBZ2kFcnHSnNPqH/O2ZD4IG4V3sPpVdUYtU9vvc9INS0SqCaQ1ofoyY+MBdiopneixZ
ssi5PGFZiRnyN2RpSMVXgIUqqd1aZ/3xqRIw2K94hspDon5gVEs1J7h0eQXF05YOiQrUfx0rVn93
2ntxLEnkM/zd/1LXG07QZQBgeOAIIs8gBAnmCQaTZPcahopXGBXrXw4/ikFM2IXupSDfBFC9viqJ
vY6DjS2AYKgT0qlbMz9oqnH8/3iseDrcmHPRxdFBmIYMREzCK3oANmZ+SFmgBh/lq0X/P1+H07HF
+3ockKSIwk14jvqeeB0qv8U41HnrQyNXWccSdmvR4qnIkbH+X9E8DjJDpFmDFIudAJMH9Djyl5cd
UZx/jT1IW466g1dZJYkDOizr+Gw5cKgtNHjlQH2UgqhSwtLzeNl8sDacPA9/edv5eNF67IDySntj
s9R7v8n/o64I2jCKCF6PuQX1VvGTXoL6SUKqRb6nynLCyAoGgh70JHRcfxQbpMc6mbrwq0T56bo6
hzFT2n1CBQvwiS8YtbUrrF0J+YBncAgOCSWQ612ifdsosqNwESdEDnQWEq37yjCXBjMk0eWfdmW6
+PuBtoAau/9XMqIFKjhc1gu04ue7krFZiCx7+Uv8HiTDDEU0bklsSCT56aK7FfZGl213YzWmiKBO
xxLS1lZGnkF5IWR+QfMMnbkh29iGy2MTYsq6kdoPXSQu2Hjk9gH8oZFdAgJoVykALUBplhlaAONC
zZBIIhiFI0p1vduVwB7rqm1aQ89eOFh2HrtDeYtJ9q9KHk/9wequo5fm71Zm+NmjezwpAAgOG0rx
eBhEWJBgZsujpz1G5pjbXipml6gPOHSaYQMtVtS+XBK/nPfWyGq4ilIdGC8FxQ8AxfSOA1RMU0LE
3fh2nndYEoTnTcJHdRAeoMf7iBWFq0vJZ0qS7cK9+ZBEQrSn4cWUlFsvS7ixoMizj4oxwcVhvWG7
Kxi8kNjKQ+s0qfWFt5t1PhbAG5p2wCa3yaBcGg3U3ucQNgfepMHvPR4JrBQKFfXCX1fmL/9QtmG3
a2YB4d/httf4x1AexAUfWygHHS3SbGq5hlnRxNxZCsw2zSFHS7+O9BuCKDz/EmQM1q+u0sDtkVgi
7QxsMmOkrWZ3ucaBG24v+nwuSmgZcRTqLk+lY0IdErxEpfTxfXJprbq7WrnK62n4auQRoxsD0nxt
22jhRj8ZosH0i0aSjAmwJzA9VrpvK5fBZpNSJitOo0lwWDYVvemDNzFZGFvaf6DqB4egFeilHc7u
ZuYPFAsSBkY+RE9Gx5JMW+s0y8qxbJT2dP4jTfyshuMhLHF9evkdEWnrKzG577eWZHF+UwKdb6Ge
FlDixfnXUSO67YG9Z05crTR5qNRK1ddV5FlK5OpT4ZfiLOVUVeS4DXiA9L2nV9GI46TJiIE3BQQ7
WHgIt68e21rYYRj3u/7VgEbsc5pyKfjobhIHe6MH4CVSZMFz5e2yWQA3tqPTxdbjPIWQjeayYLNh
LyIm8SQP06FTMMBCEWBW6f7n6kg4t2FKMqJJY4Y0xC/idVoi8pYwhjJYeqmSgu4Avl6gOfY5ZsUK
Mu4tqFk6D9XM2L6wKycLJbQWtM/lInm8yHpAh1aZd3txrVA/xFn4pg3UMkXflP0ZU4e7r9X+hXHy
zNak/vqUzSY4Tjq30KsSHUgaeaeZ/yx9NzF1vOs392M+GHUgvn2s3DY5aQlXAgiJi4pA59hTEHYT
vGDETZmtNbLdd4TDzfRyuUW70L9RT4DrtyKO0YPnIyqxZRDCgPK9q+YNRIaNcFW33D5pTWDazMfF
ndi/BCxUPQXvXcKW0WkOt2Z/25bygYGWTbcVz9J7myUaZ3abtAcliE21d7w56rzFDxcVR9s1VA4R
GAngVz8jncqgsC++NmlJwbrNSRy0hQPpD4+nqQBiyRy+Uhtcs6V7ulbnsfjha1lb7oiIjXPI9aUe
IrgaMA0P8to+k37/d4btYi6QfXXMIYb9y3XaST1MOkxvRqu8DE3Pb5I8jQhmhkiWg01LZ8Q1EX+A
l9AbX2mDk1WALAW7XjQfAniRGeSdrPaEJYeTMEFKRQ4JPphFz51PCwPYJpNv0Dye3rgkRecA1KId
yBqltoW4mQ5jHGeHNSCfw/aWRUG6zLPdGO+KLgQErnSYd1oC8hpae43p4GUYt4CGNpDdVtu1NbNF
U0deZ3Gw75hQCHXLb7vsMWmkZLwmMzPTKRuH6Jil+z/hwKNY4jzBk+8U9IA38/EI6cDL7H4mQh5l
WzqniWn5MhO5rwgjvoOguR2q25uinsLmLMWZ1/CRAgOp6woK17Cp+96RQjwAh4g3ReSZmdOMI7tG
zhAt1Z/cr5scvZPDmJpW9+tnf3QuBaNZrPL8SPeSSk4X9SSiwJBtUxBhsYzBmzsp6/OU0mCQZJze
k5kAVbXTfkhE/Wz+Zn3Tgrryt8r8h6yZYlQZ77G7c/km6lSi1ubjGQJbs4H0rRbjud2IdMCnmWvU
BMpZxmx5tqUrveM51Y3LQ4/IsflENpLf6/i5fChx18I19mjdYYarQvNZiHMaLTEXXayQ2Es0cwOz
Wt/Ey5S/gYI1taEtN+VISgpYaYBWOqHxBQdY5PsoTP/hVl9SBRGNkq46MCaL8oZeVaCX/+UZL7aZ
pV+dBOUM28/Y+vpl5DqQTmiBQp6XokBEb/CvHqTzkWIkNMYKlb6kSwLAHQ3QeA3g8ryA7f+UUnwd
flP80cNmPLSD9Ba8ObcOHwkmilM0pTyuKrjyL2sGNhktvipGVirpW23Tyfiqe9LdnXf3TXKD0IOn
6YX0wVmjTmKE16Vn61FR6Eo2o6HOTtoIQPcunro/Yy/p/GQOIBah5yfa4Vqm9KS1MphiDFlu9Hth
tI4A7MNIROxQP4bzX+cZyeTPHfOa2YybmZrEjQfpHvdamz4mBUJ9JLRKUd+7WzlE7vWEvHlw6ZOV
PCqYaAQSFEhz0tfpj+KYq0lTS1rgXluIqrHI2d5uPrr9iFIxeEgQbdLC87EJqATYnrGiZb3wFaWM
FAtrlX5/Nu5Ywi+xnwmLQ9MiKollAfUhuA2WZGQgmJEporFsTA20pLn4WaEKFNjCJDui/5QexoQq
UEwfeslBeuZB4ti2h1w+jB2gp63R4O8FizCBnEg2bel6YBbp8WlJMpbo/U3cc6lE7fQpfh0OQpvz
jkxT4jkpOJ6AFjIvv6d6cZXoJSOVb2zT7gFFHxvRNeZx39u6kK2ECRIPme6fTLdIU2x03CaSbDSE
sQ+KLq9XmnlTnj38NNRoPrhzgqc3Fo/8UKvPo9Rd98LocQ4GOgZ4OaDxYYBe754uThcI7Emla1U/
nXUZ7/PRkBo8OuIm3aVwlamBR0jtIzXS/RkDjppslgsUOziIuFe0wBXfhXjaEon95/1/EvGt/P7G
p90qYn2uZFmMpmJuPBKA0qhKpHPuYCueb3Eo5IJvTzm4aJYBjcSS5UxnbxW+RuFASUMJ2XF790qx
i1wQqHBAn2wRdhuSAn/RJNjDXGkhi11rLJeUSlM+R9Yc7haBjlISdcHSr1nFmT15Y5AoWlG0AMIB
SenQnukVKmEdlK7b/x978sJoig4nNuEUph7ea/enfSm7BNPvOO53YuxqKDq8xhZzRWr3aXwwujWt
K4eEeXZraMfX5kXtLy0bumVa250MRY4BI4pS2A2g5zsVjh4zemynBwqrUnF51+iqjnm5qnNwPiN2
Xd8zr1QA5oOIhQC3L/QaJgz3RCtKlqbWyO4uoOyXS30koRTN6RnbmkU0xWOsIk+8YBBFNP4ynh28
9iFoQq0ax4eDzapBXQ+czHJpYdpOQmuV4RtJAO+FQrMx/hKEfKGxuvnfxaYsUljEAJ3GMGIVYifx
aEPS/D+ARTQux8n6GqixiSGlXHIOZbordco8Y2S/FSBA762Zx4t4gvkCttiyG8/tZINjNXS4MuN7
9tFrKB8CUryg01CSMSDcGjlQb47/UmAf+pe+j0S9OtodK92njHzxrjkOxb9KNYsQsrYgs8XBxX8N
rBjkzo5MiB0JDI8LCobpqJ0rOKgI0YR1yOG/p+hh18cAmbB02xafJO8BXmT3x0ZfvR80Egbg9a9a
8L6eKNIJmO/KE81sHLtSH+WQRtOp4r7oMm2TzhtXVux6Zkpyl4PaJQb/0hdlDz/O2Z4PamGJNXIZ
M6EaJMgsrqpZ9Hx4fgDCClYFSXeUr3aeFl9dq6c196wIHxFAexgShmBtCbE82T1VxYbl2Is2dmz5
ckOkodwlZhVqocyUZ56qqlSptWiFptY88aXxrYCItdxrZYUIqaHNd2Y/F32A3Z3/jEJ1a2S+HWHL
mLYn0GDPk5rmR7lD17SkjsjNz47lH270NepNlMSI5/Qk55EcBwsPtI1Fekcsl8YdZ+umQ6ZeKYN7
/j9BYiwT9elird8JyWcRAc3R1EqvaN7XH7qZpPvtguZ9E62gWu+XpxXMYtY7xRa24u2RmrIX4NWY
qxkJyPLO/UViiXurf0E2DEnaWcL5j3elyCOgJkKq6LSAHV8AU0hftnfoybwsSjwrAV/qjev63bCz
MVHZnuesMxCqRBuP+CWchkTeZfNcHZIqIZ61ZX3o7CHhKn1ycvyBR/WaNUZxMvrMja9K8lFA6zJA
tHTujaxAjRI8dm6wF+oh8KTGUJg5eWOutBCDKn15A0MeKehnJTtcb3fEteEPUYO/CvXjqRgmhjh+
6jaK8lylvNpyQ8QFTNGLH+okfPS0UgUQ0LXKzSrLEtAZzGC+RDlg4UTQeO4EQQzx1hrmKxrl5c5t
sy2rZPG/cfF0rBKM/Wkt/QuMDCLxkHjfR2NRWf5dNpHuVcz3+GxA++Dz88Fv2VXCK80t2KBe6mOA
wtwbiuwgpSBgW7hY+DAWCNsAONlyQIQG0K+/PcZDr/enuPkYTziT2+TQIk5hECmmY9D/X8fMF3xd
MmHfe9dChcvnwU21w3/uMPoj5Xkw5uebR6a13IJXEPUaWf6CPiUytjEEFnoYf2DSr0MGcPb/oEzG
Lc2K722iFvYBl2D9pBxvXV12OajjibWq34Tw/Xl+AFC1uqY+oCOPX7qN5anH9vdNct5cz2nXPeyU
ipdSsfV8a5JxbbC0wliHKhhOiReAWU1dK/rjH/2mV8CvuykAVlQxh53XMko0UEv/1Cp9drkjjAkF
bVSJb1QQybmOR290eHWZUFgimjIkX6jmNcmJlHwGLkq2A2umwD+5hXt21xujmldRlMskdcgoPSPR
a7fnPP1kKU+OS16UKT/UDJwakjaxmvj8pp+ZOmVDF1+KSMI7lVedv+okj/CFMMipYXmkzxl/nV6f
wSsF63YGpf/17Tglx5v8xTs0F0W/cl2G2SBHFp44wf+BVomfhWSSG+isEiznBcJL+eMpw19MDc8b
svrf8XESNNpJdnVCgQa9KZaBr1rmNj1YSzTXJ4K7ELJGXuRa3r+g4Kb5lbKqgffSVPv02M31YbjZ
5uAQvTSbmvmDoXrFawN0eaD4EXjNl8/RjRkgWyzLonykYOzHs6PsbO1IBEOE0uZ2ojugKmdQxwi3
+6TDZMlG9yKHli3C2edxpGxwGGHcnQ8FLmI3lntaGkWWpm+VNVFJF1GPg+FwWljaTpLdIxo5cJ3l
+WA6FS+imjq4PSeXvLqQ6MoE0TQFd4MhQGcOjRcx52FhwNpF/EmunGxvglnGOfnLgebxiPJmNbzx
LLgqtr8jnKHB1LVOKnSKvzX+D/E9dABUREKjzqTIaThlHhVfF1lRQOpA7X/MWvf7Z4bjWGWYL/B8
1PvlkMfY3hDhrd92xxl12q5KCBK49boIg2LUqojwTiGUx7rmbzosaslaYGpaD01YL6bGZkezNOLT
H+7zwJoq/QI455FqmFVrO0nQouz8r4t0E0UpL/kCdNDvBOonMoDanfig4tBmS97kV2fj4UFAXtOe
Hi1Tq4WozzDJm5dezVJrN+XgMiwpPW5dwQvjzk9AYnDj3l1p/1LFTrIVZYbcQrkAHrCFTltPuGii
okL+JY5na87kC4UwPfFXasQlXamj95sFg/94nxfOiOhS5rP4yIKCvLT/EGfHkjD9K8GyfI1dJsRR
c+M+L6sqF82pIKABsXoZwJwaHyypauHvxUo2FxvYA50zAXbF0prG5QSBEe/N0qGGJ6McEtkzWhHg
iheQrMjzIXGY+uz6cDuUa92h7/EuZDPBt0BvI3jfT5H+1eCPHtibkNk0VTH/FxxVlxDtF7UCMHb5
sEkuT+21vFzAkjOfMIW01Zj1nl/VbEQ2esLgfu8jXmHDOS29kUpPOjw2X0LMQbidsnOxyizqUuN4
Tbm5OxuYImOD96SXnWRpK5NS/HkGWz3zVw3HlrsBlO8PEuUAHkpacSjMSEArDZZsGVsgdT0XUdue
OORWtc1TkFrraHkH32FTuaGl3saff9UveVzK9Q0CwER4lxjUvPPh2/Rp85CXpiXz3IZwNlwqEnLK
APxKPHY+5SHwlo3QqLU7ilNHSWf2NNm9UMEHOSoXv3sdm8VFmZH5ZXW1vTl30uG9kWeVFyAEb27l
b6etPgMgvNGk7oL3D2CjgnaprSKVm0r7ESEHF+26hc+9JK8afk9z1Yhbooxs3UxFiLIkYM+aN6eS
7e7etj2fUPUm5VyPwSs1iMJ4nx92l3i4d+HO82AbwrHxJPwPxrBIjCabcupTnDFLZs38Uy8wvcDs
wZi8ipeQ6JulUQ3GnYsxEs7zEFwAM1d9LXiB7svcrmY7SVnJbzq3TKZ6dRvcCSTNucamWXb0Zq/O
gZepoqmqAQ80xe4USVzD7NgD5Si1pmu2BRyQnvFJezVXUPGPisodiqg9SzWSw1t4dJ266RdXmTzB
EVyeb/cvEhSa7NdjL1TQ49m1xOm2ehsCsMipktzxEgVZI6YQjKWL/zKFrrO6Q5kiPaa6VGKTVpZr
wyqx9WY6QOPs5FLhePkBkTpd5/uC7N3Q4Ld+AUUcnATbI7IOExF9snoSToZSR8Wwa9Y+rV5HRjod
0DMlgFJJXi0ielaKPZ5FprszPYkv8d1BFwhpeVe54TXUSX4v+PYP4u8MpgtVRC32cFZr6QXUXj9W
QciAmCkYBvT8M2bSOtvZ/MbunXdKa980uauxFdYJhOCyz2eFRIQ3Xt7b/fxr+teYEcRBMC5GF1AM
sulOiUghgFAi8i9xaBuXUwu0vCJx8xwNP9ruJv8UnjRSMwzv3YI8pR4jxjz9HuEKs1fWg6PtzpX6
jZPbkm/GwAUBKjkxxJlGJeia2PJ3E+diTS8qPmj9uUO4GykSCwZiIXFrNDzlN/Kc49mHnBlNAfdM
XdYxQJs9p1GucURGhjgPEjYjsNvSNHTtZ6zX33aKF88c2YAubp2hydjvph9tX7bPzoQB5rsptVS1
l5VaUHayTAW+2D1XZRe/2VOn6bs1PXjScqUSQEBnNam9M7HjgjZIAp09CDb5ZecIhrRu7wnLYAVq
X+fOAG37+mhFOq3myRNATxSRaX89vg6U/DhFnsHrAi9DoZyjvlRm0q1h9wdO/YmgMJ95zt3k5jix
KeM6lPLrzdgFaH8OeU42fDbpiWQ4oNKA02/WlzI2c58IoLmY2Nzaek2q1skjTxPzM4W1h08Nf8la
oK0n48qUEiPe58qWlRfebHxrUqWYIpjpmwzpkIDMsnWRT530MYAGHboEyfNRhdBZRvFsBA+6CmiC
X95MyS7B50FJwjUJ+VZRo7gFcU1pgGcKyYWaz0HcgokLjWQJ8Y+da1p9AnfgqtbdRq8ZmGRFMBKr
vbKwKgDDuDjLvVaHqDzzFYtDJKaWQmGkgxzmMg3ggpg6/V/3bHJqdZ4Tb1E6HmCUmwxczcEOfWuO
BRs2KF+umeP6ajUw/5MEp4IIBPbb9IM6cKIHrEEaF5kFKRfUrRFCaqqpf32dmKq6e9lKuAXKBXAS
UDg5yMajzSWif3AwBn1vlQpGGc4ax0+tux4hjnE7phmehSucQHo4JwK3PKJU+5xQJUdYOmKGA//i
98GwKDFO36E4g2d01kt1063mVCJ91fVbKJcYPtfcQYjlwjESnR/w2PqkrLL2rA6bKhD583TrvWfy
JlJPfIqK24cGQDC2yujpv0XVW1oGG8w+KPuzhoVJL006SEFkK6j/SR+BBzoJeaIgBaSUC1bljrDf
H4Fkr6zedoCyypwZ8fXdWchf6aIqZWJPO1PQfhjtHpHbdPjNQnhNfdFOpC/ut4/s23yt9HKX5wIG
BqBGHzo3FZNQhXOTpygdKMYXcQh/xHEmv44c6XKRA3o1CXovya3xqWHNQjZokXKtOzGYqsi8HqUm
PH7eQkqjvy5ejJrKqwVoiy9PICW5x2G06FVblk0+c9cup3P22Zx07AOov0KNctGQLLjAPF2HaaZV
lEGIPzkwzJcPCQNIqtDvHZJE62DQBsXJY2SOEkKM1rIKaVkrdtV0iUByqfcWY9jwwvtAiJgMv+me
XN0bQE9FVpD6mVGMnDz4skqlhOdjeun0DlHcCMPXrof4koDg6VOtJkTTiWYhnWkqeSwoeRjM9pPn
WOjDkl9rKXWcpa2eTF9NjhdgkceVqQ6GWQpVaM2/fXoPU7nFYkaZNMAi3ruVkMLI2PXIzDJNcg+b
gH6VGvopC9AtVX9Hs1tG2hyva9qTa6UltZmsDCuyWXntlfvRZl2hcUTgsJuTrfC4texe2sIo1EVk
kTV+y4KSZqwwUcaW3qhdfaX1f+9d5MqLOBTA/lxg6eLwPNga0QTg56h+F5lgOH1T19URllLB8Akz
1pNBKgxuVKX5L5j0HWJfQ075w9pq7aQzGUOcr8+D4yTt+ge/WsT+/wGh0xZpbh58ShOC7oG+Wcu2
0Nvn/rG1jJc4jm5JEb4tEwprWv9dbzLaHLgkXCPfh/iNDXzFIIYhOogF/Ak7Cp7VJ3cM3/rhIvPC
NvNarJLPvdfKyCaPogguBPQacDeRdqXMJoaCVe+KIfB+SwmpWB/MGSF0dOT3Nl0CSOtDumuYxJ2c
km4HyFRcL9Vq9G5n1Ta3il7dSRmPm9Paj6o4Gj5AWsqyabl1TvbL74i0Ef3xuGBDJxanNbkVOmGk
CAWlTVW+befyF+JuQ5hk8TsxWkSCFSoI8YVex++nshS05H/2fZ5efT97mnZLmGM8x0kW9jt9DVNy
IJspoMSJu2cxVTmftjraNvNDcrEIPjJrjavqxh9ugzCZNwN5caRblu5k7uvbxikxHIBCJn74FBwP
QzIH5J8/AmiTwRc07hJnUpFARv9f2P2xlOh999emoX4a/2qpBxldOSN1J0IFsVz2G8ZMDdBMjyHH
EwZWfLr3rMYXO66kVKnt+IiPQZVQZl8hP3EVSwFyCVPACrHlyOcVy/3fbinobCov7kavEp4IdPMW
KxAi2FN5l5086MHVgWqCZpzkQI3RR5zm+sgXh6zcEkq27mVuXjzBvk62Wrna1Rr0myLN3UzDeTr9
9yp+hsJQ6C/Rze+9OLt8JYgO9Hs8CAzDNrkO136XOnMoK8MJXQv2X18g1qBQRLdieUIgEJ7BI8DY
B9/7x227zRyosr8v7txPghqpySycTzeWTf428IzGJfQmr6hUVPgtyiCaSxJjAYLCcEM2V3NXhSMT
bLMB5YnK7LytUEXzrU3eNV8jthTqAR2hFKCGyj8sEuN8RuXMkzxqfpykOMTr1+32xZabDDJH3758
7dG9IRWxkmQyOs3hf/QvtHlQ8+AHqEuyV8NstCa1PPeNahiPCef/3e5gS5+2h0bbwkgfI8qkiwue
vbAQzYlrtTZZlLJuv7p+gl3UwpHM2breRxz0wljV48k9EirX+aU+ZBeue1hEAnVTsyPvLFduEOcY
0YJSFyn0zsLgJzAYtUsQoUulpsw4O3jz/zE2HaolNVaubPHPF7EntxOSNufmmtoFvjjcCtwqk2di
1//ehcscwMsc+0Y3QfQySj+mrBL+vBb535fteS69ZK9AA1+7w4WYa06qhEss7rds/sofGglxeHFf
887frKHy+738RXifUAi6iXIzhfA7tboGbF5IZtbtHhAuHCWPZeH5YlMVBCeKAYW8Ebe6FmdNL11+
UU4NRzG1hNz+VxsI5jayD4vtdLeIVOQOQn4M35MYS7LoDn0hGDt1WO0ZnVzlTAadGfHQftxeMu9n
8nElh1ysLymh84LOqQ695dovC1OfDniecl1oXa5nAFbgIldntXrzZk3MmWo02ZzFKW50OrfYCTSC
NdF/wFHPL7/i3kqeHQXH3se4zfBJCThjUCoNmAQAgqc6zckIkmtmZCscL5uGOC5QcGFJuDMu5WE0
fH7Bfo6w2Vh2nSE8khPH9sCqAzNPvpoTczQHnL1Mh2v2Us8Ec/AXqGaie05M3sWjFX8+qEtBDP4z
Hd+bV53UNEFeGxjsKtzuk4SCvvkHjVafBf27mAZzaYeyNe56OI2aHloFOFRKdHLqb/KtXohpl/vS
fK977DCpfaBHUSHoCmV+t+feKxAuE6T0JNtsiFHZ1UdwVrzD+z6D3oqf055qPXEBjU9U8F1dzwjo
DUumdEHB6A8WK/hJXrnZU3Ejtdd4iAqLvPSXve2/JPCur2PecPg3trIX0vq4BHC0/EUS4XbDXy2v
7IhU09XlU+Ktv3LLcBUgWiYHYefV/UjTZX8l8XFpatSxveUFvSzqH/crV9TedIgeZPgbgfgCY5Zz
sEvFMCEqCc2W2s6hx00fUh7x5R7W/x9I0/XjnMA3xRBzUr4IuxFo2aibKA11EygmdHGCzEz1aE8l
xuZDU67JUzym1QrC1Im5sK2K3363RX332qCH3LYaCUqb3mpzcw/Ag1Eu29InFmvU2fI2Z45EW9+t
iKNOziOFvK1RfwIqtLxgk1fCOTowE/st37Fqkjuk6huIzP18OHMFOq8BvhqFBHajOSY/Pw2i2AfL
Ixnc8amEdmZqEE+X6pdQEUoWU75TF+68t/4gH8fIc9X2WKqEv6VTk+aoMXfW4DO4G7mjCWu06MRM
o+2pFJcaxCsGLvS6lIZX8+Ejjf6aL+Fw1sUsUY2KGLsa/tMyx0zIW8TFWFtHW+TdzWq5Z1iXo5ce
/vWLSJIQDNbCVZOvCUR5Elr1r65AlPJTeeODHmEwk12Y2JeoGgrlVBSlwidZlBni7rTREpT+ZxEI
up/Y2BaFu/apJLIMa7+aNl2G6z2EbZKUOBM3yTi8dXSHZuHOvdSJ1UdXUgbR4wkzumjuJhjbI0Ww
56py0OyWIJbAuBRBlAtQDpIH58NopAj2VUF0XLNTnFMXLlw8sMMcYkLy1xBl4eg/ylWlHifQdRK0
5d5aAq70xgDSnohovDBqi37eBSX8xJChoS8OvshlO7xKwMbDbe55lP0nsxXgRCVg+K3UcbVGOzhc
dgK7ZKESwV7o24mHpQtQA9fJB0vNe5uvmmUK8QrcLS0yUf9kA/BjSRYwCtDrQDEfCH0sDjC7QfNA
D2QrC8HqeKkH/VVOlUblVCRRtg4K4P41A2kJ5tCGpjXHRz3qDjIOo9bg8mGsGpC9asx/ayt5rz+J
bvIpBsw7vvftQOmJIOW1ajAPaNZVUOKcuMyS1inLd8Myn0RDbGgQTR5fWpOBZPf5nRs7kOWqwyc/
3t+fdc9/QvNfb2w6THFnXXUtuRe35REqI/vZevreiDvSl5lu94P8FOfNT2TOLeokUj8rN03JBlyJ
BrXt0XpNL9DzXW/J+kpDeIy6quF0Vu90eTOp/i7zQtnhxoZafxv92YSWuTI8bYgbZtOuZBWienn2
LH68SRo2qKTq+Pm8GAOpPT3J7bH9ftnuoGar4CaKQq8/LexnLCNKbb4MqlfP51VM2UHoAYKWg/GI
dVlM/DS6ZiZbAZ28GRaRwZ8vFQO5Dsx0nBB1QgUpwmO7+5RZ8tdLuAD1Mo49SNWbW6b+lLETk+3S
kqWByrzTefxJTbZjNRcUcJxxFvMD27u2xIIP3qTdc5UXkjS07vdbBzKNHcvqR6GiY2XOWcIe/w6q
CTRNQN2UMRYDTa6DrV9Mn24sUZVOF0RbI7b01PCkVzDHKgh4BZqm9eDNM8y9ez9TvUMBbwoPrD+B
iDQXQCPLAjC5zCrhCdfdAdQ7ja//TxJJ+iV7a7GVp15FYamSaYwR89gqatZDyCrkDzQrMNt7T+ko
3aK48ebRFr3MlKtet82Ax6hbu8zuooVj3fH4Go/J420UuAcC+AWrc9yGjuhIo3LGhKfhcbiF+doR
ssHs/+caOl1jv5ShISo7aGjHs9oZyvauiDmOQCXgLBJapmF+nBNosKUV5psiheeomsUCFAXRiZVh
2d316btvy6CbmVPWcpwItfjOr1Fapz3Y6oOSFO+thx7xuWzkoSVv5g4n7pabjeNHA5c4BpBthZLV
vQ7ixp3Yxy2k4n2X6d1CBC4wLN66JRfgzlCl7juHsyrkOx9GWY5XFXV9b7qjHv+YqRQLYs8wk+on
UplpwsTyCbzair7CHmxwrdFEfBChTb3L7TUAekxy7mmNYdO7drXvvI3jfyAM71fqFu3EVMIjk5jv
jLSg4ItenY/bMn29PHvBOU3vZk+0r1LNELc1BMcCtPD+cYL+eKBMgJKNKBhUVR9bM2G2qwDW6+Ne
jZXqeag6VOYUgFFtYHxu08SCRNc14zztBEW5UF9vnw1oZ44nEsN9IUYDYXcNBD4DURqTd57kE0Pw
PpctYDp8v4n0k974l+YyNVqTGYrzwrfTbs0s3pij1hRkaeDoZy/0DFt6GdnhLNroWWBC9Osq2fvX
Jo/C2m51CamGQ7MD2jAgVyk9MgTJamW3B/smZF7BVSzjPSRB6h+shZf58mJHmFmWRuGhlbOLDW50
sGmVIq0XL2gQXwNezg6sKqabuxpB32+XFWCWw2dYwbVXAy8MmFgpdALb296cJXw7Zu/l2H24NqKf
BOWRQbjH+x1FUEl67uhWL3uhbp5NQajaCIF00GNV7daWs3VOPQrJGgXJYr32TY6h+o5M9Pq0KzHg
QTpXzyqGwbTS/0rR9N7WnhAyZ0rpw0xej7Bfo/94PLQDcsPIXyzGVWzRhNARoBsc+MkNBTpKY2Ms
MPLrJ3pI1hnq2oFbR7nfEfYblNN2x/v+vXw0QLrvJ+B99qJoV+IsjEQzf9wPl5RrwvdD1W0focl7
iVQ9vF7kcrdXYC89g4VVzaLOt8X1UrCCcxfbdJ/+nMwdyls/VBezizsTOgB/lORrkmx7c7DirJas
2Li91pJ82Lqetx8IDP+RfUrCH+IlvKKXc9BoW1XtpfrnxaA+cSIwYYctesYIMQZ7HUM5SEn9/QbT
8uNaR7tvvT798UmKYCpqovmC2+fJlORz6fHqzpdaCxhbv3G/7lbpDMeUgvYjFtcjIB/ESuJsMqK/
DQB1BgR6JcBuuBS13+gU+8ftYWlKe3kz6Ot1zAI0QRlMWe4QF3qKl3ZAjBVFCpD8Vz6pkVDJgjV4
enj7xtS1fh4ytkmmirCg9nm4OODUMn4bTKzf8c88wvVMldNaAK0PxWBJUa98w7pY6HWjF5kxUoy/
m6RzpEBYRtecKbCzvvmrbHCFmfWvM2ZNYpY0QnBUpCe/6utMeoY082LTDSd017eMCVKSYvpFZoQg
N7yr8/xumn7EaxbioYtk58s+A4xbA/+xqHFYwvW1Zjqu1qFKjDc2XFJihXgVcUncbmxiW71q/Jz5
kmw0C8l4EQlopWB+vTL7ZkjxlHQ6PG07yWrX4VgL+vFSX8Q+lhC5N69JFnP1MIvv+FFARRsV06Z3
8mDu/ZSylmgXkB+sCDy+t9rc+8VgPsGMzWoNXmn7zIByenfQlb4LBH4rfwT4g3ATIfzfuXy6/gzy
GdMHBSY7fX702HncJrHMzQ/HG6PFdOLLpdrO1cKgWQRF4kFxCi1gCHunHq6LxJnm59SLyLNlSPcU
ieK4+nhIypAZLH78ljBP70zrTxhdQQUaAxhngV+x0MpCWLkLcOKJWb3Wqx5gND+pbt9X5A/OFYAD
JrhJt2NneNasScBNt29gqupHr+MuSgHmCb0ljMFfdiCzk4USNEIrM8TV9ImnB4LWgDJClddjJhyQ
wnY+gzw+MtgsN/tb5eLMr2xQD8uKmnYtpJraqEnZ3EGRyRjcOcd4cJzNdGI5RdVud3a2YGWlmQGI
ezdIC4X66ln40mW77LfKNNhWwRqCmJXD9p+KVuunxsL2NdqSCr1f1mW/vd2JTG5sWCdj8NBo/DKQ
EqF7x88sC91ADPCBo16jVI2RZOu165RlUpCpnuiPV7+Kh3oBYg5gcpQdfUt1p0S88ipUmjNZsFLR
HB+6BKkoGUov6kvYHqK6bUaL9TE76uUKTcxuAQ2NaHVWKYKvfyD26fmDYkkCowZvQUZGWGRkWcHX
FiQBuCzKr8c0wmK14uAwMccH1o+l06YwRZbWdpOg1jE2i/U8x6nIdV2W/8kM2TOZ9yvXIM54oLN5
icWdZezjOyeQ92KD2d4Ue3mLAPZvtULIM9NqPtvzk9kdHTVkrjQY/tOklE+iZ/sIN0UGoocj/E2o
eQCU0MDjXz5gWYCe6LwPAZEjUBmfLueyhXfIJwQjAnU09kfi0J1m3YqbtvBHLu7VKrsae5hWYBUM
3+zPEZ82DTE4h+dIdd+8WdR0+XGCb6YXG99nQCq+PRDY6mQvEo/cfz1e+dt3McJ15BWJGsc8UyHG
lhmZ0Vo51pl6YAXsAkPbr5V7gh7YjjPbppyiEPP4hs2oV3XndS0B8UWefT1tEqYvPrwPFszli8ST
7bcjNAadcEautWuHHD2nb1CGLsdx1giZlgIuydHm0k1O9D61CSdhNubFt8n8PfjDyw4IutEH6AXA
BPAqeuLUrrIje9ZCKhOXcztfVTNyas5PFLIdqk2pNlfIQxVR+Sz8TZ/A0khWFRq09F1HDWYk1kpc
axkDrGZHhbSUxrNTjxCcBNQkIbXp4OIGPN3Yhsyx931hgqOK7EZ8y7oulLy5qwkisXsQyNBP7qMX
jrYn6OXU1S8fdJ+rU7Jw4ynsPtjsq6cfIIWLDuCmmVKwKdGcCh7kvslw05d95HaGxlvutvfQTw4p
EnLGZpkPTNYHKv1gkyznTGISn0jXx/YfcO/mIC0QKAe1WS+QuEKaEXX9sLRR8+H9QharkPorRNqL
n11k08OaZWC4jYe3kyPXPZQXpddbdeN9FUosjhP5ip+5ewQIpcFovRqmA2/TbOFQxe7vXCMM5Fmp
CCx0iSPdg3+RasoT0s0oifJqCe4uRJE6JyYD+kYetMF9IiwpYpLhOKv9lqpcPRfb0vCi/sUbyMPv
5sIZgIRYPndmVhiaU01xz3C0ZVHfovNEUVBp4pVbYG7czPqpVpxUHvsD0tee+lhdOuk3dY887kuD
zVquTMNQRx/ypfmvJkVCQxDIHZ7Cdm0U6uQ6uNxk3yOxPq5fiTY+8j4+7DfQeuch1eZ2xg6eMJAX
Any312lpyv2OgEMHzyCVLPpy8PFJ9BqCf673IzQPQqGLVZLw7wTbOhhNmhIe8c/N33/AvVWKYolr
ahkQtIyvddv9AakeXzipzjSa4ubdkaFB/s2HuCStjr+KJ6H0cCxZ1krkvxGuzgCwPgYEZugKz0TL
nCopfF1TTx/PqJBQJEPRi88R1Xw+ob3DGY7LelDl7v9ldIVQ964FdwYGZfWYh7ZrZHBAHHq+rgbT
RcQ9OhnG/sVTKEHpPWHgFy0jzP6l20I27AbY92EDGMzySG0bcJj1N0ur92bCRyW/4xt4M+FJ/kgU
HCKRE23VKQv3bV+tZzG4CmQkP0KuZev3KvygFqjqU0Wt5iIXvredmz71fjFfavSLvOjDoQWv/pmx
Ckzqg+MAooo/OC2zZAfKt/xpWxz5uXw7e48CuVFYGMd27OE7BJAdXy/AJ2XcNuEZ2FBvB5deQxlw
DvyYNTl6qxDU5Y6t+V61mV9c7jfeFQLymJSNPo6MoqJD3/QTdiw7vZHn+InlmHPZQQHM6fVCw2Kq
6fO/tFI5jCVthDi6QkEQQlYEXrLZx4TCRRv13LfQSavyCHv9Np/mtuZL/3dCSC5TQTf1hFC+SLsf
4DBVmpv78FZRRgv1ioqusIH8jhdvQfG5gnJ+mGCYIR2+zVB7FpPFRIa65abfz7fo1hJ/e8cX/Hz3
vmXA7VAEZHN8AUvGjMhgggzUUaq36O7/2gJVCdxruyTkNRvvaR9rplgC20lYkQuf5TnHpyv7MZVO
iz8D/eFslHXugZt+JH5M2pl9HNjOUgtYSI0o4hL1T5SLvjrggbbtZH08sEaHqc/L6Mtixv3HELPn
DC+M/4dso78xh2gXfWLkNiks3ny5/KgRjkgInE6TEc/ICk3vUF6/s/+CTQUS1RNSc+5ayJMEnFBH
01xENfCLmXPK4cjAPGK94ytPKfhJDrIR7kn37lepkSloKmHnJBZ87M82MaWuLrBaG7x7LENiS3qf
0qEkV1y0c+sf6fzKdz18Qq4neLWCO/kWy9WXfAWFVKj6FcBJ7qpXdcPce81OzG89MUlqDF7W4T+m
oqfk1dca4/0pCWEmisxBLHe3MyjjZ70upJ7nhsTmoShfUkXCzC2NielHc7YIoxOmUaCzNMZOnYwa
mBy9yfH8Wr5Bd/Y2u7yRAOjxlpGtkQBixhW/p/9cYG4ZwTsYJXVSBz1y8kJy8e4E92sv/CxxgUt8
XGuNUywHkcuCbjEaqhCcX4PSTXvSVQNTGUtgsav2PXary+pdO1lO+oQOjo+Eankd/yGB0/O/A7AS
ITB55KTBkaV5fANH62TfYcmwOOCNKKTjeLkZtZioFfyBfX5W6Q+AGNV9tvynuDw4e78dXpCRVBVq
csr0MCSrYB89+ouhKnVgH2cVrxTwU8etXSLF0ix9DnitoqycRQ30eDX+qexjG/4klARErRjdCpiv
2/yey4DqJ0MOjpcelKT+OSjdf93nbD+qnIKspNEF2DQ+iez0794vXimBRf7u+L+ujMyZMR1pixG8
KDC3HD2ABTu7X+xw8nKJIN8RQXxubSalW7TxyoJYKH3MJa+SWEKdXIqTvS6Dgqyk+wKZU+tdhKWG
3MNMc9HRRAuA5/BmvAZCKXfC/KQ0rVRoBJUoy0Boxue+5jpx5HRU7uTfccplkUKOETbfViQKM5zz
OySS6QulP/qUqXoRzit6XONooqJx2X8jiDI4AIBFunKxGY/+W8IphgSpRLhIcmMpCVD4Z0lm0dV+
+iluRlIPP4kGlpiZkR96crzKdPxCr13nHwDfUejrgZdg44nU4oE81ksIgjO/t9eEC/cSOXMygod3
mRWUdTRx4XzvdVtfVJw88kPAhC92jyxpqkvDsDnnXyRgYNQ+fglfKjQLdh9RMWK83NZ9OTAcKVRo
Djk6CYyINBKVdQ1Gvw4VSRio66uUguaPu5kL0Hk3v/59K/L1g1MmtF8oP2wamvkkD/4+Oc1Q0DN8
Cu6xm7s5Fetsq4ndREGcE/ppq5OwxxEbjfYa25NPDv+kP69q4aV6+dXysSB3RaU+qLoYgC7ajWOj
7MtOSRfBtWf4dhZvl9Flj4nOx7qeO8r4bYucnbzqX414hbinTy05ctC7fb5eV3vNEX9FWTqQxl8b
Ny72SuXHI9u//QsedFnjSgq4YkEPd6shUDRxoKBYRhbVd8mm+nl8rQZ4XWuJ/L/zeywCNpd7fWMm
3kHDQ8ooNlglDiH99WvbVYQf2Z7qoyfi3Xe+6MKXvGXyeoiSC5ftckAFM5hgO9DdFetkLd6p7jhl
VvLaUIEMYL/4nwH8K+XcRWkyUhsR2nWGz4NaGvMcTskgz8BO0dsXBojfJ2KwG94yzKfo5Pl8ZsuX
M6VcHW1cZLuJDiz4koZO8zz1i27ZZgVIi3zGOgvfYCo3XMK3dNPtf7kwYXmYYfCwO1NcDn9O6zue
pGfmDdtuG6G2FnBLH16SnSXmW3P5SGXBEtPo8fxlrdxfj+AR3ylboOqbJyOifwJ+5Y+SXXu4+Vrq
9lsTtV5W2iDXBWe1V86FkraF09Gioph4PC3XABBe9C1Iy8ODTiwRk5bIKKnXvcdlkof4l1DZCHxJ
+CtYbAF7P5OyqVaT2Kp2oF4O3UTJPX+MANO+vTBmIUWdeYT4Iq5lrIin/mAsZzZ11LqMpAjEB6ej
HttsU99pLCyG5z1ZNSjs/47i6yCzwXX/U2j8JJChR6kMFoMuTTBoaUiQ/HKgjIqa02Qhi87J2FDs
gZzb6I1/WAzKknIwK3qhJFJg95w/StYJZeXtsVE1I2WujfU2xu06D6rhHubK5LmoPBaaIalMAx0y
0twRy+Flr1iuEmwzAryzf5PZOAoT3Ik0sdt3wjOuNYXKe5nVzcqc7bSK+Z9DhRM+hr1778R7U8+g
Xctlqsay9IWxNVmmp8KYW0DGYIw821KNnqQh4Q9rAG5gKXNa7bFZ4pnJnmd2HbnagvXRkvG0FLOq
zOc8fnHJhAw10DWo5XhR8Syg6ff9cRdwsTKdUSxc/2pwDd5B6jMol8w3wX1crZm+prhj5+XQrABt
fouZNG/fk5hUDCzhdgZiKw2dVZKOGZwQD/jP/RHuQzueFMbNPXNqVo/BYrZ4neAUu5n1GP900K95
M9Ymh7BdH/Uh15WM0z1ur9TOIyNks3DYZUPwYwqUf3iFZPiSVkHnTyTSe19xZad60i8zO+CQPGmw
ZCjEMCBfL+93D42ZWBmSbMSkRvR4002ZcsbSi8PbConUAUSXlPMc/mXQ0OKfEK2r6mRdWqqT/ETh
nmNvkfFLXZDCzeKkpUnEFCXfD+Wt0EuwECZCjet04+/7K9dfRPEUT5f3c2S8iY6DGKYJeXs00jwo
fhgtrNKg67guUwqxwzmPEus61+J6ov2qae6iDhR7o6YSySOk/sb7xevKVkXNoIIpLScX1zE0H18A
+lYvdfZhUe/UdVGXqmWnDgwk+5uYV/qZc43jHapXbxVrMBVBOQsjo1IxcIuIDlJXfhecKFRzp+aL
xhVDk0E2CBUdTmJwLFEQGfaewBO9NvNajUq6Ge4vD3BPNfI+FV4LDuiWo1vPEu8u+A4x3/E2tsnO
dAqC12UbBcNEggrWBLFEuEZWlh1AmVeXz+fTazTXMVh1ux8TKNVpEt0MWJxrWSRF+2wUNZPYQIh1
gWd4PrIv1Uc6tCXw6PyzMkid7TnaXp3gGFw+Y0VhPEl3B/5yKlRSpKvMu0OTFOyFJgvDpZxUCyUI
+Eay7Ga8bdjET1ZO2x90pr/U8STf7olJ7ss2KcYyEzzGPnaPfADSdKpCcE8oxK3acOHsz7KKnIz9
ZM4McpurgU4fobpIjemoNYPaCbnzeNHD1lny8cyui48FM+hoinvTpksT+YvElw54kqYSG1KvGWGJ
Ne0MLdO/FvPiyZynHRsiwvYQa7Q1RCdqHYws8G/r5fAuYvf1BSU3Iomv5nrjHAxNWLlrQD1sOU9W
O1+WX9he1NS2tx+NMlfaoF+AZDQJaSHs1JjWNyJ6dE/m3/D6Z9fbcvhuMsg0i8KrGs16DPmQQWL0
9tfHjCNl3VbetQqSMbS2ECpp1bx+GBQ3Qiln1CxHIFTiYW3bh32cAfIjYM3F7L3e3J6A4IQZZQVQ
Evhym6Vj6FI0bBdklwGqKapTZsBtA34uevADFN1waFUOByEKDzT7t3Qm89VNTUCPm/bl5c7LMhB0
/MJse04OoVa2OL5aoq0D3dH/RZHFAYqaVRiDhHZWgkAZaGUPn0hnSZqdISMuRyWJ+g/DOB0V1bCe
7NUPB/DIn7DCEhmY5SUJH+l0GMUpncjm+NMw1SwXtjlnRbyyta4ZCo3d1J11/9nESGWj+zhWP+j9
yLI3dsYSAuWJkZ4CtTWSdNi+WAhz7O0WQBYRFDvbGQsuRxxMrwlfw7TqzrANBoJY+x6g4TDMBIuD
jS+LzwilY3WhRECCgu7m51539DzuA2JE0Z1IsoLJbZnC9+Lc1mXhtjcvmWcVrm6jMx8zDNAI8GQ6
rqYNmX54PCDIOswiz7AheQa6M6ykxqNRsWpiS5K7BDGyCC02HuPrnUbRvyIwAzTUYJrqRlg0P++M
v4diFuxn5E34xZooxmIC+RG5//ILPPF4E5wdKK8uBdgrW/jxefjmyix8/cr9RrJryF8351OG04SQ
SBjFJ3yZTUJqkuOLEEKWd/cds9H3agFScVyXbDiNBjAZC3M9fLZ5g0v8Q7bdCv4FfmZr7ccoXY2a
MuhblVtGK0q8Qd081qZRNsp+ulYn9JVgaVhbSjy82ThiMmcI3LThIypaoOjMmKa1pOs29iOpvVB0
mSb/023xcMGTsKY0AgrLpgaiuw1aNJayvEaY1MGfys3T1+CZO2DIZmS5Xh1wrOoebzrgpXuUjqiP
3tYEy7w9WyN2Abm+NLBi8zJGeTNLYarUwTDNgJD0nCPwC5b/HzKaTn4vyoKM2BVFbU7KLki/iKvB
OF8L5mHcXI7ChcNJDKZrx0ZC+awGPdBpRt7RrV2nQaAKnCnwQslUBrEaAwjE8lSubSBtWINjPzwX
SAzYuB2SuRrUrWEwhREdqxMPQTEEQCMeLmD+OdeTpA+gAusSeQI8KTdwCi451vnvMtmEdsGVHNjJ
Q8dSycswyuFrM9AtB3y1yDr8ZnX70hd+KgGu5qsB9HNCyzmkFbXaIMZ6WQxeJRNpkFEJkYRJy4jT
6WzB0xxDOeeMROeJTTnUsnKkGe3YnrXX9K1O9t0fOpSXwNhyV7XNEpR3saf0Q2VBr/tSQ5nsfP8R
bNcMcHheX4F2T/ENmjx39Ijj3xEh+L8W7Z/pbRgUDTsVCZuCuNiDC56bhA2EOlS7SoArbamfzr/x
F0Bb+4uZrzpKL8moxmB5EK29ob96TUaOIRWSsGEncc1xuKaPh5ph1grGApl+gQhe9bwWyKqk61AA
KIV8STWcsQHdc6/9FC3VALCqW5qxnYatbxRdQakYZjpzLS9otwvSWJiKx0GZ527yOPvakDtimJqQ
wBrAE6Hg3z+5McLwZTg085aDqh0NYVlgCjPIggYozWonYmiYCFwQXzAsgYgUbxc5EtzzFm5ZbehN
Fu5WPu2Ii2Smnex3yMi/3CPn0RQx8HBB/OPIQojPSxdTmuaY6Vw0hjrAYrWYdVmwU7OdxQcLf6VO
88slJX8+9UDeRWZKKwRoDh+ff7Z+VkCdWd5OIz+FWlirq6JBmedg2mmpClFjXt9NDjdqXOLUD6dD
hHM085M+nmP3x5+n8mUTZok/0iSgxoZjucCi8vJqToWMEeDc0slK0VAkVCXooB5LrMuXxwTBARmv
iM50P1m5LUrAmB11L69C3A+1TxnT3bqZ18v0cFygFgszH03IbGRwP5NuEyHcjghKK1udzVyL3iXV
D6S8MRyP984F55+c3dCT5VQYy3Wk5Y+ODNjBUK77IDmnTNHnErXqPQssaA6Zb8DUSR29eve95nLK
5bzTRsEVgFWTJ+DCUvU686Xzp+yEfJ4IiEiUKon2KdVEhTeRUW7lmXJC0Zo6CW1Rvzp3oBqwCKfC
kMI9qU2Zk5AJN0YySsGsnHOBUAFNagDMS9pVgIbVqY2STre8MHYgfE83BNpJJKF9k1JpwNBMIWc7
D+1OIxbh5sdhDaYJBckhPF/hXcpbHINwt7JQvKC66WiOSKlNYKVGRyuucR3D04JFGZJSv6c5uFjl
8SyAhC4PGpKR13q+U9n8rNC5bK0sdI5ACMKsdTcXwoWsr4KxOS7Zop60x2Zk7m1vcRxhfT33TDa+
6JXQCdFjEmWjjPhkvQGjOeq+GpfbxVddz/qwuWwIL9ASHsGgUaSwd/L3W2bB8IBEIY/+tEZ9DiXr
e6kXCJmeqYINboOlfkeHSYA+Xtn7LLTuLEs9aRfM2t7Dbl8iul5dezfH4166EdXfvMVYZn51dI67
eSE2nx8yf+J4W9eJNlRhDDqeWJ8b0IkXWBbxvPnpz+a2Pg0L9+QXjx6SPgEHVDI2HhkkZA0gZYXn
S46k4gZMV1IDe9Pc0Na0xjDD2hAUKYfK/VHn09s1kTlabUtVC2qtHjlAbOTRCAGc49KuD9WO7RXu
1EQUishHNX6afZfgtnbqDscy7LYZ5hspD4hYC4O0wsF+f3VeJ+0MnDKcOpmt0vIqxKCrlmxesty6
5aqvhYzIyZDgfZdBTc6PtuGNU4n44HKrWUs0qX6TS3ooulxyBsj58f3/oZ1VvGpnHXr8QqlDZ5gy
8SldeTyW8V/TWsnC8ZO7heuAMh3+F+l/hrSR/tyk+M6y/9lmX6LCHKoH7OJvO1wiHlfZu25nIyM4
n4aQhMsnoRBNE5qE0RmFCN2879pYLfDtTiZc6LuVgtI4Y+77QuV61OK3dAW0wp2hwxaDN40j8y0i
bIQGN+Ddi9LDHH71qJuxB3XckUJfhkuT81VhNsGpF/iE7jIRqdhkgz6nxCMPUE/Y7ayEu7DcERPd
gV//jF53kJGSg54I5Tj/c5DknvMf68GcS1bIFthnd2Y0L8GY0yf4KK6SI9eAKdGFfScuMTaIz5M7
RHMVqwJTpjNteqvmdLomn8LlIBGv9VZ2gtcmgIO0miVMppIIfDq0Sj1qVWw1vUw9xZvdH3kghmTN
KT573Lp2JQV5qyEIhLs6V8Cc7J5BuzqKK0BYZLrqV+5z8dMLRLht0oJCmkFPa/ENSxxq2zZsX3oH
ZY7jy99m3oEjKBNSBm7jgc4fV+fSPUPSOdLCuk5BVRiXgGwEmwuyLvBGEIyhDE3ZzkfjZPC2m/HR
CGHDENaJwSYdjhDkqW/zw/I/XoaoiOd16rH4iiuXQUZYoiWwjoNTy0+P7bXrvVmZcGr5BoevVXG1
hTweF9xo3vxpcH0G2t/7iCsuZ/ZyCztU2QFlmWzeCGXiQAjiWe8EEHVLahFPaIChfaMY8esv9SvJ
oJFCRq7PiEhmz8Zz6zrZo/479TuP9m0n0wkUyFsjcz0WORofbubAze3ERn9AW8kAgFnFzOPXEQnw
QGBEqcHDHrvq45ktS2FjE3X0yI9ceyR96BrMyF1U3iQIV4ByG2mf9ONKlDTdE0P1+tsJ0xWtjJrJ
zv0pydl6ZA8/04qvQbYPwmTY3gQ/g7B3lLxNKj+8KYYC5YPULE9R5Jf093okCWjgnL3lRqFWvoK/
8LzzJ3Py1DqfdkBLf5S9AYiNMJ6mYF8mLnTYpXcTP+TJLJxeDdzkHFzyAuuRgGHi5NvSAIkQWaSz
sbQSMzLLrA2VfI5Gxakh+ZvHoi0U0UplhAQrhLUv5MU2uy5iUSlh+UDHzF8OjAYUnUslP6negviS
gFMJCGeIbwVywiJDw3CelSXHowoeVqV9Juv2UdKZnXo1d/JYX1IUMe0WzUl+woGOimyJZIk5q0nj
/iY8ZUiEFvOlnRrbjF8c1IibVBgN2roLOrh5390QlHKg22OGktaJ8UlRgng1958xHiliy9PdpLGD
bcdBkarAoMIOtRJH0+R1kCyHNaShPEg1GWNC8kceKFMz1vavVhcYaxFsU1eKlV/Xf31zQ/961MJo
Yxs5dhltZvOLYxdo5RWd5DdFGoeHFkU5RZaSQ17qrlWT4KzZHK/7B/gthR/5NuJbGxtZx+bv9wKK
h5GqsQ1nqMDYM4YOhhaNl7fuw3iqSsN6s+DS4pemddk8461eaNBPfkMdurW2N929TlIAyCjMYF1r
GMievgtOlEqwPsJqHoL1z1T/h5M09+X4A88oM1g6Hy2LAoqDYBDaWGspUdG7aqVEd0+FNnPTBcWa
fN/sdlUoAKH2GU+IpFlZ4fgUlOBlhmj9p0s762vTiQKQB4TyWT7EcPtjoH2306urWs6z2SIU/Ets
0atBVBO9Dwncq+ZOISisWxucFyeMzskh/SZWczuNWLF4iRQZxzSPYmFiPMPth56T80y2sGs9biGl
okrkIEu+PVLAvidjbvwpXaxellwzAeE7JsA17PYhKQSyNF+0B0tN0840uKmrI0Pvk0Bsab1mMpTu
UkBxzfPN3ucpG7cx8jqnX99KzrKeZrZUBW267lBdMblz6eqk65BTL3WDdX713XUXcq+9B4YpqLD1
aFWgyIpRRJ6S3U91n3zGXe51t7LxGrG5MCAcOWDjPwax1D9WNhyJ6bHRPLmB3r2tfFSRUgcaqFcy
wEgEI6kyGoZqPMPpIr8uFOS3R1syA6hLzIufBQmxX+g7mKCYql3Oy6JZdmvc05JLIL6BAimwhXnM
pX8SeNA4Vy05PTO0J2OJHAOZqi1P+54q7DzioXeSl9i1jxEfxG953p1p/FZ/eEHOCKFXwQAc0SEy
ZE4i6OwNXTcZYG6XBdCgykBOj49BVVmOS4glUN/oIhOJMNb7OGvgzi/wf4v1MnRzuVWlxcBechDo
GwT1njMXLOOXO6prW5E691aWxGobXXGLKssGUWgp2ychVkKyaAMjcIexd9xUDkA5mLos7xvy7RzN
VhrG1qEY0bxge9evbFsuLTujlyK7eysFJpr0jc7NJsKoJ0vIlVWtcnQtqGM20FTDCCnK4AifVVCz
OESxKUnrHSQniygeYxrQUHfKjMtEY9QrNoCn7uTmkMt8jBYeklE8xkCzBkSqlN4aZzVJuVGqzqY3
GKVQHdnaVYbzDaJ9TSPCfuMuIuhP8ixhyI81qtWnWwf0/OfCkCBFNuJE/hYkjy2AL47zdQpLQst3
vJjrkNk+MgPzd7lUOdcGB1nlygCpMfkDadaNs/Hu0/HabJyGpkmTCnMhq4D3biW1CLBgPnvkaoSp
U9fQ5CiNfHzQfrgIkvv1B1vMe+c8UyUyLPeY6xnimXGvnXWrQqphPdac7g/LnLV8uMBcHDE8IHa9
AYiWNFkO0Zl2GkRr9ekDdsSxXxWnGErkEBWAW6VeMna6SywldCTk6pyPTH4YlIiiPSBPC5QdsKqs
IMZvidR3sluzzwpdAwhn2OYbAJ0SK2ZgMTB7QZT4EQV6ArMOzaclLAkJY9SXcNFmSW8PwC1BOGbf
CnlPw4FZ2KmTzGpDkvgIBrtjuhH0bE5IBW7WXNEkfGdEArhIMQBpGrnMDl6rLs51bHag5z9gwXs7
6n0pm6jdG1Z+pT7qGPTDORGMpOlqzR8LTL6YIaTjGGAGH1KZVUW39hWkSwm5swBy0qRfPb18ahOp
5iPpUBr1cSnoS2qGljLyaaOv4sygUJTueV1y4po/GenrFu9cLJT1TAi43weNHh7dWkGUSjzLDc1m
6+xYY7Cc4fWgfn5CaRcWkjocP62DrUnua/N1PGdny7QrA24i7MWBBISgE8/8CmOXLuBWX9j0J+Tn
2VOgb4cWxoJPwwyOIu2+oXEfd5DO/9tEg9dPFaEWWMPh3ZHqwfCj/+KWiB/l4hrNqtt8YaRETpdF
B9eMWKGmgurIdw4T6/YOraXVae5cTfsroVhkPwfIWXP49g/p/aXCJGcfpPqoCJGGn9XYOz+qzLcq
kmCYqwD/TtOpBXO17YoAQuI297H2Ju/QRD3Se41auN7N3j9OU0t6HrXWOHL4gxOaE5LFIC5lySER
kqdiYwUtDnKiFFeTwPHOsSWAd4yqFL9dfzvgoFBWTvpowUhngk3MvSbEN+ok6vB3n240SO9oc8cs
9foDH94DzlXe8Hhw3sDmqx5BJPzqtVJMIZoK40lLivPkwJ0SeUVihe3UKrLWdA7bqkhUvL5wYjJP
WpH+0EP3SNoDR5X0RrA3WpDCaZcHQqtS31cSdsWBp/tnu5XvInqZNTdvmongnjwTeAlF1O3IIg6U
ll8fo+s1gP+v8OuJVIJDCJ8O0ri1kxG35XaL4ejG51LvedqtCU7gZqcBbJcvzot3EVBZCn0a+XA2
73FZ/78ACJidg/TgfreAWe0ysRVraC+Q58taiODLY1MZgdgBiNPLvXas4nV/OxtLiki8tH1K1Mad
zHQbWw9dZe1Fy+yg6l4t6hRjxD58JB9jl4nYduDtlkIlKS638ipPDBN2FKZvRf/Iv8sWg4XCbvqp
P34v4EqZ6T6WtbW80oinlywhsYQL5xSS4NCbALZS9tiiuAiF9pMiHH/pwE7YrrDRek5JZJRhDsGI
+YvcewUjvdJLTgcgPPrBMMgxXeOHAX7p/Gd/43bTj4+eAtdYtzTy+697lt+LJHqp7FgDFtWMFY0C
kdzxyHPhjRYEd3uvx3o2spKUi/W5ben0ztw/5aMBq83wQ3e+14JpcSPWel2nCDX4keBTi2t+qxiZ
/pORFq7d4nLx+hbyFia0Qnz0htyPpozWUH3hBGwvQU+BYhcDUiRZo2sGOkInAfy9N7O+VLXeMibw
Ddi8M6/tAGPlm/d9F5u7+ht3gfCuvNv5yovYtlPb00BBc0BTRe7tTbmgwFXx+syjCvMyU3+UYn+u
BB+gjkENWO3w4HFM/HSSURYScleaM4Tp50HjtIf3swujEdIzz1t2OaUEMZEiHJ5/lbncfQnD3avN
VjOf0vR78+TRHaTEa8VPSxW+k8NupXbOcX7k0kuV/teYnAlY88m0eOP0HF47abmbRrzHngm8y8qv
68nJI9HtqQJMUGMEW7JyKNwCENKDmB4j82vlOrRJnyLGBNR6Z2xM/Dme9fMK1UoKeJjWp/iqmtNE
w/FvvMZygpR5AowKAnP0DWCB0DkwYGcZUhxSZkCUoKwQhZuMZDi3Wizy7I2kaiTG2JwS3sG4mJC/
FGFsue5O/8LRqfEJlDuk7MklwtXRbqfd/grrZ8dllxGd/PtT/9LvGn5B+nHqjjYGjEFBnKiMGgWX
GZTMGzgpdgXLn6Pux2+6DuUEtw1OMgk8wlsrgo0hzg4nRXZC9tBKoPW8UANfYaBvsQmB0K3yDNm8
L1/Ql4NAeMWwu85mvjSqgCkUCR9ICdclDHTjTWkwBaVI5FK3HBasbkFvKwlJ2OEn2PKilZdYhxaD
HZe9OL9Rpyidm6XGBYQF+w9bXBYGCSp+pfvPUkWT89mk+tFliS4k0h2psGRVEZAynS+ZQ0YIjJoh
HTFzHCJa3syHap9D8ahDa1aT75lthqXeO8Kdnrn445Mx99+oEvRURoxdbHvluc+uK2otwgv2Jwa9
HZvYbNL2qYjA7RNrrkVq1Pe87p/FDCqyl6ypkxY1GSlMK202ixPiZCKOxRGc8zYLauPJ1ucwJJsN
zSNYmIPIVI1kJAtx2O0kXHq6Bnj4aR/d1CFrnyAD7sp1IfQUKmDBNcgbNPYicQU0S8QyUrLHa2dZ
q8lQGjqamerUUbbteVQgxycIvPH8Zcgs2PjsK5aTdJgVbuCpHtC/D69qPp6ii1iznio2PEQcUlXQ
L62VjbFza6BNqFba+Jx/b8a/4NO/mggJSLZoZp+3lUu4iQ6gPm+01t4I7hKpvZJ4qo4EyBA3Tjr0
K8gS2aexSFWqs05GsMwZP+RZorultC6XIi9zpqW/SO94oEzLYA71Gl4wHCpmI67ZuJq9IjKTNMUF
CcH4WYWEBLsKKJ1QidUc1BcK9ZTBeHgO1FHdHvtyrDGYaXJIdgT4mpxrrkkrVEjmiJWb4OAEKGyQ
gJ6lTbRNXSqPwGHkgnhTMjphkph2qPooh8r32z4VCmgW4YrdFi3lXZiVGxMmtE/pyZq263ym0iuN
n7hizzDSSPPeudUFWgbec1K8XsX6Nt45uN2S/yd+8DmVoiYkuU5daJnS6Ff6CumW1Wi585c3zBF0
vs73+SMd8X2tcz7+LCXIFW8xHWB6jvO0WMxzLtKiMjU3KbnkHiokHOjIH69pORUMIVdbEsEazyOi
F1GlEnm62yMZPNxIV45L+W8rFR8syXRBlmaaUBCycDDnBLF4RM2xaxPId91OImknIBrMrywZHX2T
+59lwMHxytbT4HhrCkT/LPrFa5RQ8fJNitjgIsJ47tUEXbGR2vZFczz7LP1Xvcq5fHhxfuumrfmC
a2zZcAeyVgf1yoljExW57a7/lTISk4TyTm6tg1CF/TALru6XXpM+9tgg+sYniXb/jHXxCAKQfO2F
zPAdPZ15FIysEu5Mll10R44a6geBLFJJydGkhuwKPcHsnTT3wijqHvGQFQEHPadmC0H+OufSmc8H
mgxOG4hF1nGRFvGmXO0UHEyZ8gXN+/GAkTpeYeGb6zVg0LCyQ+0KbeblXEJlcP3816/IaHsD8RBs
QasrEVqyOx0wiNJkJFZYeXil0o8w+SsOLh+GomjD746sc549jLr0N/P5yyYIx/g+gpgzpV+ryaSt
gXRMFa8X1lvklnDu7K8tBzUmBzUHMMZu6nFKVvVjebtNcq0pg6zZDXEuIK2rfyMnP+S0rLbhQp/F
AFpr+UB42dSP2asSd/U8KhEqPfECA6m7bf8ZHsChMkzDmjqZ0BU8/eMYQTmli945+TQxrA1Ch/HC
kHScdN2zB7Tfn1UP278URE4oMh+nHXPGtYhnTrhsUwEojE4bJ4WvNsO5NP2+VRVFICyX2dU3mU/f
YTKx+CGC4U0JdMoZ618oCRr3fj65m4IKbKA4Xc2HNx+F6DcbZoPmdTECH3CeResHG+BddwIZY8o3
yI50+0p9O+Idzyph/T+lNLlJTsReMZ7qrqLaDNVTGOvrncS2877nWeQyDrmj4+g7ErsXxzvbJRHb
ep7UQbpCwZX/Y5mnsJhVREDzGRHhKxVB4ZaKcL3a8E1YBRD3iWSrmS97LQEND5Up3ZtQBdMScCAN
vALnzSh9/ANkgBFWQavMLsPALRRChUj9H2aRylrV67mydlt4BtsTti1x+rvrjxJcTc6IVxIUTcgw
0ei9VBT59OIcILrmtBfLmuhMUTsqS9C6hNIS4Yg11In9LnXhcKUruXK4EqEY4tjqt3rf/uRLiUhN
5lRANJwcTaSCgCAzQb1uUT189vfFwE1Xkh8ul1h01JtccSepKgWyatJVYJh+NZrMTUAjQmbc5yDf
xmfOLR1D1BhXv3PIVxKzZx//8Vd0kfeEQCq/jsiMuyZONw/G2Wr7rVqp+hjUiO7jWIjA+iOS+oz0
r2FjigRnz3L2hJBjKmXX6NGqCzlEg9yBEzcuaR3TNoPKvgck49aQIKhwUtUQGROZ2RTLSeHvl/Sm
ledrvwR9DKZy7YPGXIG4QAfmblSmJDuOChi9KroLpooZPW/QfDeabam8vZxZAU1krt2dCuzd18bD
8dL9goO2ZFfMUxXlRB0ggmc8REjqCK/GBfCbYrCbw9+w6cyJxyze+U3wqyfsZiTrLciGyhlHbRA9
wWYpV7GyY/3v1tEacXPL0CCw5P1+qpgX+e7EeTUdyd6HzoFtue7mp10BYQgaXGBOmfKeZNcPyvbx
lh/4WI0at/poolqzPc5WV3NPYMFqAFdtetk+9xgmkyt/DUwkIjqoqJb1A+IXN1N/YdVgXfKctacS
Sq9ORVIGCjjgOALknb0QGJS9Nbpjzzv2DbufJV3zQQbEZQbpwkh5tO1cNkPXQJnBrsPNoKXdwMlA
Ln+aGarfZp8/laBrHQNi673WAzkIWRGfVbAL/97rGqzsvgfIJ5roDa/kpbiGX1bPB9YRXYfTq5s+
uDHJOUlFos7DgU9foM6VyJlqcyFVW7J+eTCe+SptWcoRAmjvmgG9/AKBchb6zvUsUk6aZjgCCOLf
Qcqrm8JpKbTa50tp475bx8EBYmEQaE8W7jqPtcMq9/sR3ZTNz62aBj3dWMDbaC43NezBnHm+BVPN
GSRrfETS1knMdkUtqLYVRj6m8DbDhQAlH4Pl4kVYde9TnHEXf69PLAygCSaNnPIhGURe5licYgT2
qmbzW+5p/1Ru/azi38VywUDLLPPu3vU4u3YEFF+1DVztwSWdkVPZv1gcIJLZxR4n3aubM981A4bl
gwGcL3iAQgoBv/5Rwgi63vErYbToG7UvwyI9EImA4Enw226r1akmm9A9G6saDT+FIFesEWFfUUro
VDfVkJAZQDN3xZQ/YYs2+0t6J1a6yWiVpG/Q494rkU6bSbcKOvzVJk00OGzXW+CsGKJdKboyp+uu
IOHdJhxymGAnsgEif+Qg2iZkabg9sn5c+0AwyrbHMOn8ZJ7Y/dKM6YJdekrjESNv722OWMu8yKew
y/8/lmeLTDGMEaF4A40bbYtKM+uVx0NtcFqafmPZzJjsxcrrj69yWs1izaT9FjyVvA9kNjTfhe7t
oKtOFWYedXTABztWllLtlO/RUccFj6VTThW+lYHJ+zfBrUj7BkS8bhuif7jRZYzshfIsEUxmxHHJ
adXUkMINMAmIRI3BmfJNzvdL1efh87mhUwKC4uBybkEezDgkPd3HlkCZvq6rGLNNfm8116/Va60z
dzYATAbM4tLPxvlpYLfoIBf/+z2ki2KW/bEpfAayjglnjcjYr2Y51kgvabXusHKAy1OPtZij8Z/2
XR2eQqwfZJoybfOFkuQcvMrbB9EOEQCSesHR6V3evlYuPxK2aYq8RimYJi238PIICjVA+kpAI5n+
bizxOk+FDE7tlFntJ7PfagoOHChEXTd4tknHKj00/zXGyT73t1fI2+67dyiPqcfS9xj0khykkqr9
b8Gfx8zDdDcJIPFtSjiZ4TR4Fhksr8Zg43Kgetb3UoJ2tChX4VQKbykVbf7bxhWajpvSCnfFfNFv
Hm7EJFHMEnuiModdRND6ODh5ptr5FSxfhKEOykcnvQtsekRKFqqhbKwch/7R3f8Pfp8VQapB/MEV
9t2BimAmvJvzmcltQO0xpCvUTOR6zmQtEvyAosrHqoDL/pMTj+4AAU1WZgCkAgdlG//pIJp+0YPI
umtcBdD03FNWLbcDcM8uLSk8d1L/jwZLW/dHg3wUx0qGxJZUXfLNHZeQMtVooFIftfBKNEbfEwnS
pJ9GTLZS1l5VatX8avmJ5Rwf49+ZJzpwvAzsL0utXV1p5Dq1gFOA/8fomY423iZV68/AmRRkmPgW
33L0jzGhDGh5fLG5T79BJvBFlLYA2uUnkpjHq+NN/xsyUo0DfYU6QhZpoG1hYNLJoqpH6OyMpeIq
xVjN7np7i5On7NT/ZARKwWG4IbQywVQNVs6XHA6J9C61AXiLNmbartP8SoOe2dwTK89vtBsmPsjF
TGVqirbcE4sZ7VpgmZkY+bluE9gZzUzZ6bi3SqPU/lAd9K6dnB9ugv9ElkwVkC7h1h9TEH9kFjdt
CzcgW6QwYaJduNY39ZM4vOD15h2ZllNSbUGHdMB6L/+jshlRIgkZAR+SzN6yoZB/6dEzrYvnUzMo
vkKla4n1vrM/ywzGPpXF9mtyvN39P5S99DYOyeCCUKQH/wGob5xlgAvYifaxnOTPngkWJgJNreFc
YvvbJAnM7bG51Y6r5sdA7SU2yLhtFbGnRnxTdFCUPYLprkiqTLD92jr56Y/I4erS+zjL0/UigiKz
koWbMUV9OkqLnw9TsbVo2QGwVtrBCrN1GvOQzHPy5Pb/07iqYEe9/XzcrG4aKM/t0TjKLkNMYzqI
pGe+vGJ+7pVgJDiRuq7+fRtmmB5yJztubEBcoRMKcmcRuAYl78QjN64lU/2sI4xvj8mSYrWrFJiQ
mLjcb56YHufgT+93thyLrbIDY+x0C1iI+96FNvPJbvFEUDRol4uVtbNgP4qL/eGnFYYvx27PZ51Q
X2FjV1kwdyByyQksaEWppaM9oMvwMhyMn8oKhXKnbqNsReud1WatlgO98+I0H52fT/w2SFBaZxUc
x0LM1u/ftKQmdcKPhZF638fBs6Y689fKBTDeqF4WOZ3hLWXphg+VgXZXkfjJaNZ5EVmrxPBZy+Jq
JUInVUQygez2DJK7PcAAYeyResEcJYNEYEX9bvlFgQ46BbAVq9OOuWjb0ulIhxwx85lJxPvCRRv8
PVoojM8Dn74TQ0QF+OCAIFz8a/puh3d+0m8tTCZHFV4Weza9Z+yjA2jS6rZSohWYTRJJzgM9RnRx
l98db9AZOES6VYDe1cY0KhDxcSHENORNlpOpkRImL9/Hh9gRw91EkcABnju/ark7H8c4Il5Ma0He
npYiWJcd6o+8Kjh/rzRuW0Th3OaBWr2Sj8qXNald2lzybhhAzNzGaew5gp9F15xN/dIAAClI6pso
gaRn2PcY+HD+5dYtUZP8IJhf2ZeoUHHmmg500Ps6mFbAMl8Dw2NP6/aH6CGWx3lr9N9rSjuEr46H
4tR/u1YtXn9sifsk5iW2ZXOUqkvXQurzMLxuQMfyPRYSUvQZVF4xmwoERs2yLtHJcBu1MUb7J47f
qCNeCMmk+RLqIwxVn1lOivHuhLU9j7/Mn9hY6iQDNVEOhS3FY0ZyMocbSVlhAZprqcsVk9bkK00V
QB7c5obfrQ8YiTI8rgBpBx131YsvAE89lQFpgnYYuWFfMbD9ao+TKrNOMuN0ctg+DoelunU3mPEs
IxPLqPB/7+pVGAHH5eZP/Q4vaZTN4m4Fxt1WSAkugIwTJUwU092c5hR6ZlfT7bApZX0dAzxFdl4f
PjRnZHqUaTNv6KTbMcubxvqKwcGy8D2N1uyV+QmoDUBKjjtAKTQpXp559RsQb0vrIFbCTL4sJ+Wf
8RYKHw5YfiO1rUTny64MV8qwT6/0qvX7oZLoOLD/pB0BtuOiSeBMtTL0H3+r6WmKJzq3VnnqJNQ1
bXsMJwPFE9c3eScQwPoxudClj6MZ7Tebtw5e/s55YMIhQHCQTGg2qiHCvMJJpp87va2KtNorR07z
tmYB86yL74Dpgxkkr7tsV6kYVFFVMQLABDASQuawnwu0fB1vct64ZPU2ZHoN0ZeNadQugwZxFdKU
7tUm2ifD3bJrJRswffkEcCSeGwNUiR4rRLEjkb01rpI2EyVbeRppNmp90jPpah7YNM6ZtSREtLud
bFAA0Za1VxsAOz0YN/tly7DEeNrTKDcT9Dw8EUgGWO8R/7OkxXcM6tMZg47T9bbSaE/KuelmiQEf
Lu9iMAUHZwi9LBEQ9HcHLmKIxuhOrfyIQU5+MJ7VeBH9a+AqOyuactu6NhFMPMo+RjrWhL3O4cyT
iSD5nkHYXwxnPDJWHPgxfexUpc5SS/aIK/SU/dhOwxOpYSZHBVQw/tLOfKvPKy7OtIa3I+1Lrh0e
NBFuV78SNodQOr4TVitOhtjqIMg1loJ7Go/L4bm5R8S1p4+xezlp9afi8kNgxXIc6Q4OgTijetiL
XT3HPJoMEuW1LS4Nqu7Aoxw+022RyObinhdY/lo5D04kN5aGu2IGhP70WIONeZiuIsyUhNa5qpdk
coweinxwmVcpfuidIXU4OKiuIK6Az6WPlvAw4RzAsP/p0nv0/rwIbzdfoQjRCe8PjUuMtZo95AZE
h7YL/5XRGAmVBwyCWu8xY3t3LAIvJNec3OUkqRAYmDhCRgWVo0p5RGmCEzsPj+4NePl9m8veNva/
tw2D52vD2h18ohmduyXbLCxxnJugdAGas6MQFAH5cCbUhcVKc87H9iF0Wch0i3dGCJ575sz0VZIe
A9ORN4pQyaCObxbMxrt8A+ErlvRNaAZG2D8Ng/Q79F9nrklWZ739iIjgAlatFoQwROemQnrrsxYs
o9+pGMuLZn5AIwrud51S27YpfrZn62TC+FyRjm9Wtu6tWI3ABzbDPLiC4ZfDsYnNoC0QSlzK4e/g
WH983lMk0tIzzJnxqdy3X+TiAOIc4hFsh/gfaNHh8C4lG5UCRYUzVk5r3vYywKueKuCqEMYStf3A
VuTwqucxqq+HPgAvx/HPGCFgd3EMtaGntzSO/SpwpECdborDKQwfAq6q2P5fsJpYwGyoO7pD96K/
BeVc0gyIzrxEb9wf+aCkEpJHO4kusfDjbMHS9GrkAAij7nmKfhkqCZxNcDDOm9gnPBNABG8VQpN+
67WgEMmslF+8ENTPOA6BkYcn28JBtWgiJ/N1PZF1ZiB0zDK3eeNtPBMwlSnnqT4OTEikVsqd+NsE
9vWqtoOXI0HpwB4C+BAK3niYMgjROXLZmdDzcm48080VKOZdrdezUv6ln7TMAhy4PyIWWYLbXNxl
HVlYCFQPXFFz1mSqoa58HNv35EE8WSxmMM7JEPldfq6Q995B04aNvywGlGiHUWjI1Kh1Jz0gtmi7
6qHXqluUq6kyUBrbU/35lUYqzIE244JW8amB2fLzbYIYFnGRIy1XlRgKtpPmpkFygwSabEGxyqJu
DXBRFhdqSaFjyThqPMCIq0rCq8p/m17UVKRTZuFl3AnsWnlTJ0UXvO9xAdCrcYeJREqFys+Sbmtg
ercJO/Mwk1z1Mz4wpl0W6mJCJaMAzwCAsDBNPjQdPgoi+skpFslQDv0euPOV4OHC5rcloITE3nqc
76afrf26ot79BFgnGrdHs8p7VQbe7F0Gb6Z/9O55BSXY9Xlt1HuyfDkvll/u8kYMrwELJNGCPgO5
nZnhL3zsbGa7Znyw0R8heSGJObieQi0NMMIWu8azPMY7Vgy8rGsOUbp9Ds3A8dlH9gec5auqoVup
pD8eqVlKxMp20Lxba0mQtGeTGoKefKeF3q49pzS2BwJbjWRSmhHGREedG3VpB4qVCACi506kKw2v
IUr7FmOJ/moH8wVoPEYgxIydmVdM8KsoKDdkMitW/atDpky+NlmDCWm09mq1dn0jsxjWa5gNhiFt
uzYeDN17UbXwmkpNtt1vP3fyJtvx64m76qHhwziioiFVFXmPSgjZm0UUN9wMO8oC7H3snxwsgn/0
MnL2q0R/G7H4skjZFa6F6wulQsPoryRu87XTUVTDzZSWXJxeE6CwoUCASsWbibt+NljEXsW+dRwO
n5iGoAuUcgr8a452vTvkrueDiQ309Dk6/A7DQyvLWsY/jeIPTh1iUFgXMd+7XdNLidvwgFPdnsKQ
+OYTvY2lznpgJfHJcR36wC4SE1j3NxtdyCMwis0fYT+bUzVVuFHWkyuAbS5g5nqUDF3apZMo3aAb
qgy1+Mlm/zSHifo6y6pMVB59D6KpWi6tPgbM4MIXsyLrLzpk3x/OqmlAfO1biViYaoS1PFvPkcvw
pMaflQHwjtwI96YaHrpCiRwKCrU1B/fatEOPP5TQmk5gCZIpHqhHDiZ6lNikQcFRCV/SFjHXmz1u
vOxH9R0rowrFUULFAWyE1U/kJk9CtbzUpMDBmXS+cp4Uuj89eNdfryUc4iOv+fTKHqXqQHyiHn4X
EDhFhnTYSGk9dRsOPOSHPHWW2es9JmO0XbMP41q3peyuIWH9XBO2/wA/xQu73nY4EA5H3WH9pViu
ivLwXMFHHOPPnG/N5xXm+/d3jeneDhBM9vM2xyxLRVxZoWgMp9ooNL4ItVJ3LtZNYv8xMY2SjuxT
zoSvkjHAr563PGXjdoO6giQXPxjd+GjhvFabnfYa+StlD0aCyfChvHeMWtWWdSDJJ3WWdfyaSauA
U8XJUluAMVhCpjP8h/CfgJeaOiapfWc/xwzCND9XvjWcjmpEps8Qcm4KkIdA90WM7YMm5i3roMOr
P3S+wJNz/8cFKiTFOxWfgB3eHhBgQRuf+mm3kLkygf2razOKzmj63sI+hne4gN0Z3+8BdBWXAhdU
NiCvMV+JAGzUBc3376YonofTA1xtOqEEFiCmbZrOdE9OWTzUYL9Ua2fnvzdrnXYsWtJcpmnEd/Up
yvMDmyDXIKqSc1BgNL3XrmRAQ8XtmsdeS/gA1xe0Pqnj5AA8D/0Km40SSHBeb6BP32siSLjutWA6
zUdPWOqe5S8BWenFeYI+OxZLEis1gO+qZ2U9lwEJduz7sNM80lh7b6Df/G3X25U3j2K+/ruVHNA6
sR86bO//E124vzIHwnMJtyRAH2i/t7scGlIXbt+KbxeDSSbcwL9sqhLcxcE/lJO4cu23lbSnzzUQ
8U1Bklwg7qsEmULud/fpEwrbl8k9BUqlc0t4l+uKXCdx6hhJkxE8CGbi2/BsXUUU447j1WWFnZsm
0+WZcwBt2mNlylKy9UQ6OuBhr9/40dSSiGiZ7wOruXUB50qtpbOdLMNi20NVK++B47RVhpI4CUuw
843XjiM1FNzfA6VUOXkeFJmZXwnHPIUtmOV+kKuRuqoXtJcOb97OLc/6S/pv4hMuRK3+srrxqfaR
omovyMg9jEnabBVavj6xELBXlx9i66KEWbvwvtF9vJgqPZisrVavKm523dMXIygxhJBV3b69Hzg2
vEq4H3UhfZW8CwzlNcN4kSY5sE2XKzZcV3ICEMBwhVd7pX1XJXTMt1Rv8g2cXjgWQyCCpPBmhx2m
FQ3VNW9/0huUAP3tXpaMiKEttvWe5ASjM871Ns0+CkbE8Vv+5zlGeG1RIWLyrRuX40imlwXjzCfm
mfM0DJaL590M76pEJ9c0PVLDYcXkwshF/xCYEflP0KydvvEr/xfO6l5cCr4fJgxlKsAA96o58bLq
FTFjM9vws4I5EazuIohyFRA68xc4wUQtn8A7WPRi8dnsjLdQrvc5C6cgpwsOPrJ0tYWgETiBYdmW
tuFu6lSwQotPGkDFA57o3Vsq2fH7u9RPT9hA5MND2n2eIQtlLiPEqJWqvpEhl2bVg6kDbpvvFbvR
IEAUy4Bygd8acJYAiDzqS/FctiggaZ5of683PZlkYJdZSq2fHp1FMvHvel6rQNmu+PvOrxLkKf7c
OA5CVeSXAIvO/RdRgGD9w80UXxUSRORYRtM2Bgqc45Ww4izGHkdjpFX9cOUC80AvxJDFxaCJh25S
b2vyQO2TZAL860U0uIpCjjIPdK5UK2ne7qTbpY/IA9wnD62iaak02WGck2AMjQxr5Sezr0/wz+zj
M31AUIHm5Pm4X6y8FPWtncmJyuLvZFmTDxZLJSzX1kpgL4KyTtbnouwHZP5VQoBHRSxnx9x93+ql
18QUZs16T4xfJInqJYANxuyQrrK2jnyUhCG1dkezitAJ2L6KmyYUpD6vad5Kxj4ZMQXVveFwluKy
nLzSVUsF3UfB4sQg5qFc2Xn3hfR9VaHno5JDUHOHTe4QtFdWGdDkNcG0zj0hWNmndiQVZF4+q64P
b02o432+xlzi0aoGDXF6eFUn+u871tsW+Uw1S2vRRIrYgxHxN8drtan0WmpVIRVMSTwlLFtA99yY
/rA7cWxhggWU+UZyComdgtqa+7LQEMOZk6bgY0aLUkIRJv5MpjtDEuvY5jusvB258uP0XMNuaExF
N9mkZ6vFnjQYUJuVOKqx1vcmT5d3+f+bS4xuNVKewSnXYEEMGlHQerTc1c37/E1uJUGbx0TtCa8J
Na+7RG420Z+Cqsf97ZwE15W14AVdOasUxOAO7meUOxsJ83dOOseAdbF0ULtOHKSB7i/rZ+ATLhH2
+WzuDZDmVOi19jvv8/HaDm/oVyoHY7dgCLr/xZWlSqv5Erg4TJrM/W8vxQ39lsfuhMDj/6frqPXN
6hyqCacBnc/Q0j5z2SvMfS0e0zKDsmDYegmIUyo18U86KpBEYj69snWG3E+lD9UHXj8UQoDqBtiw
sOvK/OW4XttEc6UZRomj/VGH7WnCEN0ewdfCz7N9D9oin/b5NXDOjGbOefYfv9MJ5E//mtyxu2dm
wMwXLzNbdqYEQXaS/2xd7RjhIQIM7z0ql9RGWOs2Q5X4lx4xHTmiymKIBh6adyE3z70K7wVwr+pe
axtmNksF+F15qPPlvyCKgOn+sNhwYyKK8EJ0K/5M9zS7INdGqBdTd3gkcb7WuFU8WcfRWyg8r33F
XYlK2cM7p685PEzS7fXmuFdmgCg8DexVk6C/VWqU6pVjGogjjrPrjsiS5awRRy2pJSzqZL7x3Ney
RxfqXAcWm8m3AanlovV7JgKQHqX+Ny316K86LMG7IIg0jS6dBOJG+3X3SMj5FyZRXByxRHKr3lUN
p6T1tnYtW4jlR8G+Fv39xPTnsTpge1EDXi/Y1xYoalmydCnnoZymKs38KZ78+RpnV3JAEYRsSG/c
HKge0rQ9i3QyPvzNUnLrlXJCtSldpVsgho6JUKYF0wOxL7skaWGEo1k/XpzW635SEq9/OE84B2SY
lkLidQ+jpqdXZd0Busl/iu5PWGfzoUUQxPGuPKx7Dl3ObFf6mXqd7j3DpW/3i/R1gGCghIB4j2TU
Qjr9zTJqiUX62spjRp6uk9XBt3iW0IyfNBajcOpLNomj1zjex1X4LlcKnCYPBsBiY7OqM+x5v/nS
4ObxPaqk+HYdNvqSGq5Y88UXN9YdkUV8h9VlFWVyeizBu/eJHUZOY7FH+oMvutrgLMZVZYD3/t5L
DYAlviD1cHOuGG3LFsfix52MArEncjEAI0Cl99o1KgzT5S9Dnye+ki6TJqVKl5phA+e2UZLVO6Z7
qagBdlap6AOCw1CkkvG9JrtYDS4yXuz1/0Im7uNUxLCgoIwb0LpYTTL8wxqvIJJIjiMSqSuZmpmI
v8D8SzFZY/HgZsVZDYETsiuw2pbC3m22a6y8UwDISWRp1/vgootke+3Hvf+urwy4zgGDrQ6c3fcW
uNMwCLnU7m8qQ3rQci8FlJS/PJq9Tn7GPtBiQOQFLEZjrS09ZdQv2A4k6leJvd9EZCrBXNwvu7Hw
4tEMzZ0kFuO7Y5k5CvxVUz+870MWbRPcne14cEGJ8E76e/6mo/mwJxAqZu7v8SDjtSwxoIQBhPFa
ZlPUTdsmPeA/huRvWCdMz0yejGp1YZow2gMVI4Gjq5m9/Mp8itiD6Q5hqD14p2xI1IC0+TEXdtna
W6gg0QGSHed4kJnXCFBx01rXdvhfYyLJ/IvbM27Scp6XMmQinVyu4tYy8SFVQdzK1ni9yIvtzg6M
Xc3PH4oR+F9JFCNLe88S6pB/6qIRFYtxJ1WoaDLm9pUcf0s8wiD4Ec1yXcQZU7wCokn4BDaRbq0E
wkaJZ2fg5B9yHcpfSp4OJSdpvBLadPHkM49P6l/TeRqkv3AWnhxWS61f+haaqicUwHlekbKosUlP
Tf+eWGhPc78sRnDAlmb7/sBZI6bg79iAMh/9e3IJIbK/yjX+5YPfbqTaW0XXgBSlIHa7JAHaeom5
IJhwXxW2mzlpDiUn5scWG8wmyzNhpuGcBLuEZVmymosf8OI/bUskwv/GMSGRKepwPSX9oGmIJOdb
J9EMJj13JB/1lOdOux4gv8xpYHIkoPvF7WcpjeguDZhmuEF/SlSWXv9o0ncHAYyZRVBr61d+/GnQ
fygU5gYH8jRwfy1rFtdkwc+DMg8pWvf1V6gF1cPTII8bBMvAg3mAQzfFCTDbEplu7B6WRbSkuK+Q
Zsf4/eKW5Max26hmpsa1d4woVsFiW1KqQlHmSq3faBxOpB9oAptlm7HyR07tBVKZR1J5l1MQ3Zqu
lk6570H6X7QZuDnNme2Bmt5cQsIoXl2ab/LCKaJTgCIz7wcL51rZx7Z6InwqZB6JmKfVCdL3lpWO
84Ih9TOFNmMCnRrWUA+JqWJQV58Zqws1Nh7uedbEm1e24vZvd3pEEIcRQ893qvnB2QKE2w21S0lk
VEeIyyWi2ZXU1wnvhAnYpxNAD/wZnVhTORDivpAjv08q4J1Tg9NS4wfsEsKjwq8R1ZOThAl4zwJt
N1M+cv7q4wAKKK9cUxdHQwZe9k59dG2POOOif+SpH5U6LE8Ywv/VhJ0iUMDig4+JkjnxqNYFG8g4
DlbvNVOlLoXQ7DrgAoTlXepbbk6kRcUqSfUZq3n4LetN3gEBaSv+EHCVfTTmTzJWnSAR2RNmsysa
2AdBIReCIOVWSxWtY+B3/Ag1HxH32iQVKBdDBy0Pck4XXm91vuXLyUEqdTDJj6dkJtzGs4NGxCuo
e2tcilzVwaENuEuOSNcBRTZWGI0nEywBylgTKi0dvKEJdeCtwz+krZZHmhykMM95swlzLbpAOc5R
70Mq5MZ/zvxf6/111LeiCHuqP3DW127ydqBUT8P1voBGY7XixEy3OvyXj0AYObaqVXyZ4Ucsqt+7
CMHDx2Xg4cVWAAyD2y+pR4SHKl5evioxYQAoefUizrTLBBhXAttyolpAZaKE0/8XLSxt+JAnh52E
NPJiEW1s3Zq92aPzNe3aDGYWxsaxiHVSsqhjmpaXzz9Z4341lMfjRao5Khp3eaYiZX2jKFtTxzNt
/Fo87sOnjMvYnfwny58bktqgx76XSDdKOn8+1brjLpraNu3XozcidWHS8/UytBKV7UrhioqBZdR/
OpOVJ3z2wQjiEs7XOscQIn5di+JbzHPZGIm6EwCPU9QcLcT1KZbCX0RCYqm5VzLBX1qxBxQh/I9K
Tuo+4mFv3SV+7+Kei9DgU7ifi1VSfln6HdsqV2pevRxqiQV9GE5MDjDfd44fezdt4ua5gRg5lWb3
/dgtm+1Prhh1f+AVwriYgIMMvU9y+7kfSnwGU+MfBQZmk/VW0O+j3XveCmjPNQTUtkgcjJcyNCqi
I/yEZ5hhmvNbUlXxW+iDJO/ntnE+hOfDF4EIIj7RkyipkAEzn3tYIVKCfYtDPoSsv/rugYhtLHax
OCJ3ySSFcLoTRii66dtuO6YdTFBIsIkAMVlGARobFlxdjLW526ojGl7fFGa83QyrgaXIHQ5tnRuM
JifORmqImb895mwGFq0hD9xL31V9SxUZZtTbdQQO2r23Bdu9dUSt1Qg1Mfkun+2g5J784rjNRbWA
TqIjihD3Q7tPFeX2ncLY/4SPGvCkQ2bXsrhxrsr4crGtEBDYT9wupkgE7PbQtk2Xj+I+8Pu00CkE
4doR4dNgQK5UkjJs20wHF+QmeiRoUTwtHBBAAdCAu0mHImIkBs/lGQ+kuTV/C1xN+PgejfzlD9CQ
gSjn3nByPv1/TJRRl1fCgJbTKhpgahDXRkVh6hDWe+0vOBRdqUsOXm+o70Esizd2Udfc2MywGJS+
YPIbBKYcckDFmoO89vI8J9z2Ug1aCf/+qlEq8zwYggZzj8KMkQag7hHxd9oH/IMXzoMfZ7YutWj7
ILimv3IuDDdjl7zgaiR7a8xOKmwaTp5I7SqhPR7p0nIXIWGYpAF94G3XdTfsRoEVDpQVCUnj22IJ
4jAzvMsvhweXU7xCJbzUZRX0AzXx+cPBQWSLb2ruNFzbUzW6UwF+gUfE68qishuD8uRvvNSG/HHn
j9wTRIiWvMjqxNcTYwU0sNKd9/xxP5tOOOtAwBXv7ZUtydvBiIqujw+fwR+V6fHYY89EsCmMF+BY
YNkUhxCJTsWn9QI9K7ufvYNtrPINwPZCgUaQkPesKMH2yLFb+Gy00vQAl3GRsV1FWf9xTQBrccEL
abi9hfpdk/089+USJyy9aWnA2SdzdLlMOUyaMc5HjuuCLcoW645AQIWB6VilvZyFog+ql49J9LAc
LbH2v8YiI7lRMjC9zo199hP3cAswIk8Cl2JMhRXYTqj4dW5NJSqivYjqXE9SuZj5r8mBgpwhp2Zc
N2OO979sVPFOf7FKWalcYkxNnT0R9USkdrRwgdw9RYFr230zTY1y9lx5o/jpUb15M2QGUI31d09D
thiJrwFeejkl2mRQAr9xEhIEYwz0uZPXif3cGA2OO4FrJjQbML1UbtOaU+tPsEYJ2nWWIXbfbnRb
oXl/4NzAKQjh2NXZ/U/tn+RYoR6U00/iGFBo0YX/s4JN/MY3BT3tS+a8XVnIvKPocFNr4AjExp/g
b6qPZJWo3uANBrAltVyemOqEn7sGvNwDw561mu3JNN+VOL1NaL77Vu48JKIIeCU20f5KaOpHydNk
LEkdNrnyhrGEOAh/bJlMXM87BORlHerDt0B2JiMgmFd/bgdKFcXwVTmXHRnTypRFdj1720VXrf01
orA8ktEMB/+qfO0K/alGX/EzlCeS3focivdzBrXXIBlcrF6oR/HXqL5q8d2BA2K+rA05mJPuICuh
DYfm9hyjX4L5tConvrpTVhIn9NJ1MnNIBenUe3+OpFbKyBA/eqBzbG6NYwKPHbj72lOLeuvTxpQe
LBSXoXkPlG1I1BPfonDy/u6CnnXO0jdpUJ3xECny2Q57PLoqBJkhrnAr9uHu623gT5eR6d5yj3zi
wISq7dMu0l0dgm8zrUwPvpMqQqVwR7ZLQ1y0dHrbiw/1kiirs0PWnPH+66661LoFmzP5BCiJFY0U
ZCzLsCc1BSWzbTtt4YzjWRXz8di48HKfV0f82jCIjRZ3VfAksXRaffP8ddddBDfGXrgiVahoWy5W
4sYh+pPIuzgfVwayynnyFjrOSkAb/5fL2b5Rul14W7nhzkJvndotkS1QzldcVPuOoQemrZ0u/KcM
gjL3+5fPYxc4AGlnsaQJmeyBn3PLbTTaQH3u2j30t3umITOViqS0T5zG7Erc9Rj5/Fw6Vv+fwS/d
QGwTWagvIJcnfhOvaM+IGNIn88bifesviifwhi5WZ5al69XenRNpaczOtUOUFFrUrwwqI5AQ3OtX
3KL5ods9dPcfQph9SuPuoSX1XHtRhC+bYzsQi2wArsR2+OQm1jmuckKZ9f45L7ZWpzElBBD//Tyq
UIt3HDy0uA5otnalBtq3rQd6FIM//Gcrvkj0gn8SHrBSBL06rlHLxl4epccLbLvn8mqacpbC+p9A
rdFpaFroi/4Ef3q4oSxtufvtk96oR6ooiK5h/weMbVjX8jlvxmLJcNqo2TDyxMYzXGVxgkiAdS0J
zudfk1hhTLrA4ycOaH3BxQaUY7ga1mxMzRVlmDkZBG1/JVdSjZy9k/YCrV4QZDQVcXFjElsyRTVx
iOz8aNZIHjzE9HypyFCdr1wLuSFBJICjiPerV6CbztvZ0mtkjwVnqAbvmttqaUTFrRyoKn3vCsAw
wtWb0eWrXBKi8VX2U/wLs1YKbb/rNB3RoU21DnpUzlJmpFb6X0pMi5qA1nfeCB1YFPTEbjP8qAcX
dn+2biZRFPGu/LXXb9QXtKZeI+CsXhQ2eH4dmkmFRoodqKEIaFEpIClwtc8Eb9v5WgvY1Ip/UgTA
73El9HhqWeFt9xyHA68BTahXolAox8oIlgGAGEq0CGFc7icdEi8z+rimxLefGcL+Hwu+UWlMq1TM
3cx8yyGLu1mqY9XVIk/wa7mN9SA9fRA/VoUuntMCNEAswHhyBlkQolmm/hULZ6ZcHJK4gVquGqmp
oUCKexZ1vbhqx9xba0q/QzRnJZgatdvPChV7NbGW2niEA7moOGDcdJuchFod8f19D7ysekSc02Tq
2a2AFbpoFDX0ufqLHiE/jQBFUu5QcvIoP+RhTGrIA9JrTI6aVHYvMbFeYrZjEnt0M6GsYa6Y/7GD
ZL/nucPRoz6tpo/5xw6OT9SiLFjDwg89sxkDRMDoJowHtCsytMWf8ofszMGcVrd1eHwGAWXXu8Mw
Q3qHiMBxfhIZ7NTQfTN4jkULqIpfqKITdDggpJySOFxGzxFg7QRceKtmXDpL5CjldvJzqLM4a84Q
uAWqSr2aCv0TDJpb5BGZO+cZ8TMKTzwkRm+kSqOW0HxMeAh6xrTu3dXTRmQKsa8afrBFabad/lXJ
P0VEP7R1vrkJDtngBRKVIURlZFf4P3t/fNorvgO7kpFqxlRqiB1OtWMbKIyhjbtFHqwE6DukGdZb
hg5nhMXZOD207OXpJuJVGRPayY7CZmffbm2lVqnRmjcSm4M+pdCHJpqd7vYJs2mCsDqMw1ryw3Hk
kl+y9akTrM5TNXegKwMQPYUq6j2JnyzvYd0rLpop9PjQqSJVAcd1ClLYpT05jQp8dpPGpuwu7rCe
KUZFnt68lPuNwOuzh0xVG+JaLgAWRJjaaZXcidh3YMJwf/IHonaOYWm3SAr8aoaOjHCPKJff8s+y
3rr68tXnMI/neF+LE01DccXunF2eUvs+E00Qv0EmraAji4lKI2Uw4Tgg+BfwHKvwpit4yfdzduGM
VesKlkHsyeVQZ7BmpiaRxCeJirVsu2hfgE/DSnXUh1kkg115YwDPbOIoNcpuOQB7PhGBVvqQg6uL
3EzsQ6KDVEnjp9xBqu1uNSQ4ECm5JlJ92CrIPTelhgEYETsKmlzp3msA6SO+p0mki33f+ge2jCDC
go8+Ad8OEqD1mBrj24v/Yd2ZmWhB1yljGgjb9GfJWDzgUWN754G83us2hcjjPY8ceR33itXR2lqB
PWCcXoFAmqyqX8m9U9rj4q2X2oEqFOIon0bQRzaCo01QYhsjcvE9BTvYRkii335+r6z0AXEOGl5W
PH4ZT3VP+8B1Ohp4NcFvlf90UMZ6lpeezBqbu13i2wuo78sh1dSefrtsbebiejSsl4gL1mIGf3DU
FoJZmtEe1Ot+1lKYpK5W8mitWRE4OyB1f8WQ+m4+O595pBEi6Xqq2osnEvyYEqId6yUVi2kjnGsz
ZwhUQ+f06saEXQAnVamxlddGpixbQKjzSgRbrotgf0vn/sCzhNjWWpzXQx5ZFY5MSRuifLiXYmJw
Jf+kxIsrpq4gupWqx8tOGS475EYkul/X3RBSSDxuNCRNNJqiPeaoaBQtTSvy1Poxrq6RN40wHQfZ
VYU2FcrZBqhHrrWXw066qJ6AWUCtEjFKG+SKEfq2r3InbznKFlKzuhN/b7dnwVpsVRuWtijv+Pfa
l69Td/neIUjtfZtqRR/Qx6Gcud/2KK3FzzT0yt0ucGg+Z0R/Sj9jP8ZqEvEErTeI4Wkp5qS+QY49
By/eA1jMuZXftur9dQZUW26pK9IC1kfIDSiwTc1xCoFL2rMPZ3BCVmg8fCQVNPS7O4PKy4RSBrnC
jAA2YLNjjLDMx1Tntg0RGBSOotJwxPUriTwnQp8NS1NzGK3FUPAgei+2igkJrTfbcdqZZVFvJCSK
oDnY6Ov1JR617RegHAMhMgFaT9daf4Wpkz9nFFHSIIVSdcVi37mbzW7C0ZIk1Gyj5cvsY92PaG0v
PWChgaeV49zumVcARi0GRDZwxN04H4Sc9fklrdAyAiu5WUcGxI2QysX0QntAaR6Yx3TTUvU/IP5D
BFwdfBY8WnvWjw+tr4hjHrS8z5Vr12b9zZgI6fGx7YtpeuKIjUxeqAXLCwjtZGJXYcloKAZWDm9O
M+tSA76fTQspGse/LTHfGdDzLrXGFzHiuOLQz923G8NP/XxchvVc4lI4iUHG4l5WyWV8xrJ/tqZM
fKkWjnIPtEHtetMMIygzoVd8pR4D80tzwCLPmIn2i72q9gy0SgT2V0X6Th8FfLJS4hlmpJuLgEyb
gCpSs6WXh2MVbUkSkoA1F8hssrQJoC3owRKN0zUDpblUP/zx9lOL12sYSbGozumJiOmTRqoBL2rB
r4XYq01r+DFJcAqI33zwHmqdoojS+BI2WuxdLFKXdbV3rwtvqb4MZ21qI8DotnsggHibuaYfHBJA
DCAJOu7D+KVjJ+sC9VRG5VOb19pQFUbPg+RwsoG5FPwOreftkF+u132YjpLBtQPiOKMSahplcSGW
Jkz4+WZSrDAvd04soR4juRAVJDhRlWO90bamgPF46Mk2pI4gbtzBs7VCysvLKBoEGIGUTzIaDVLe
Qbkt2dSBMxY0vzf33HYIULwHeZ+DgFXhRMYYGWloCmCHgawhWBluq6Ig69kOpns3mqGeatwoK1e6
R0XCiImBfZLQkL4hZOj0MnXBlf2WSRi8WrV0ciIsir2tVAy+0eOTwscZ7MA4w1H75NtWsHb/kTZM
b9WqHsSvMdlHLlUY1T110TIofX+NtIF6MQY0BGj1zKAPdwh2H9AOnTHYX4cMxPb5eWY6ojrXUsVT
Ozx37UiewIxZZve3l64KT4qhZbwF5QPCv5Yu3xGta+fHnOhoMdIAAp9NmD13Au4wxuz4TgnDk0HU
9eITPRIJBWBWd/ibETCqXN/FDe99gcD3EDGQYhG+dVf2jOzewQiApz0bT0bL2LyltFRs+6pXc4BB
S4lh0Aes/4Gtan5ZeiRpbBQOpQEYt+GVU3IwXCPlebw+ZKVRTLxlxvvP5iADYQDm0reTj9mYUvBC
HhJSFyKaWWtDJAXNnrK/W6wJD/jq/zoZlygM13CuFK1d+LRraTGbYNAZEtq7PXQZumq8eV8v8veF
EVYtg8NUSKJGnb426LfJ71UUXdjxx8bQPJi0VngerJT5+6tI6ez/Bu+EiJ411pHuYqEnTIRQDl3t
J1D2JmY0wWto07kqfGasjS6e5eFM04vG5b+fG9GU6CFEV1kL8aS8VcKl3h+OAWW4M2iDqmUZlvDQ
k7M3n2t+mnbXP3V1iUTMpqVYF6eGbS9q8lwQ6OuZjvI0ZRk6ZAXCHX/OdItbDwtoF9rdhDpExk+/
IrKsYNKtzHTqUsFNCaTyMnDw3uebFWpjOmIPTCt5oSxdRcWdXtfOVLv3UJH+DDRl3NrrUuYbVDtD
56/CZ7kaVdC+Qnqt2PtUzv90GPTnw6GVBZEi170/MqziJYxaIU5Vox5sXVhsm9dB7OBO5q8PIval
mzy33EcgjmlV9eCE/s28pdD/Fo5Ivt6ZrIGT+SpDOIyyUohlJKzHfgrPJsEHuBkThZGo6IO4a/Sj
0isZfA9wKEWuu/hEJPhmZFzFOQ3xWtA74ki2V6uksgCbLfbbCqmK2MQaL61Ksdl6pm/J8BvUB003
ES//ZmXRKy29rJRq0JpVsxgeT9ILJZTu1PLB3IalwuSbLbzO2MytzPl/2C3L66PrY39hMKLXxI00
npWlYdaIiW+Z/qOw+z1aEpSKMxrykf0Uddfcv+pR82QuQpsEtbndnfz7Yo+zfJEsJT+6K/qiTZBl
cLrDC86y2kCBXi2ly/ddQzYxHB5bw5MDaG2BSBEwGJa0Qt2mhRVPnZVd1Igi5xWumHFCvebuwvtg
II6b+MQymWD574OgRoq/MoEkBY3mywsk6YcY3wjuEsimRjL2ZyMKz/MioTY1qLlAe3iS177l4RUt
48Zzzf9oFCsjhZoR022zbbzX3it2Xy5aJEBKDmQ3Cp67DBxskPqaN4HLS41CDQfctUgPpzUtGaFD
5soU72yd4lgFEi4Vbsx6wCIssZ9/9K2wU0JKvosOf7LU754oU6BWg09llYRo0hz8bTpnAavBoHE1
xmCAOT6P5Os7Kmw4+sZnC/OyEAHsqfDTiAUbTYBGnd8B0oQRFXn8AEIsFBU/ycBlb0Ugau+nYXvC
OxxtcZsW1WLcWNbbO3depUZPaIWzdpID0vTTrbvdBYryJHg4SNwAIkhQ7dnc5zwGge+3oggzBelo
xs1TsDJQyxQ8lwMnDBBNRnag9vP9iVCLa6ABqNzgln91kxctWPaRTciICvcX24oY36GZMkHT/a4+
0ENS5RzQPA+WARqHRhassy3Vb/AITjqelxvla2fRUs9sBRVkVC1KaupLDH7U6R5S+8J7oDVHRM+g
rLhWxgVFQo2jCUw6jcB5L4XpXMgEys30kweC1c6L6wm9A3JSQO832dsSiDtvXJJyH/wD0nyJ9bE0
vKJj2yMuv6QPmSo8CJzM/YbmGzjlKjW+s/x5nAeDobfmvKUbfwNMn697tbToc7p3Jbrgtg44ZowM
3IdQgf2FhCCOYv+KW6r4cRuzfYEH69ygiRAwNDWR0s5lUuvtqdEAPuxIdbCE2KzZVd78AbzLjBHD
7K4OomUt4bHZvn1nc9XyrIBrXLWDsoN/AZBN6lu1pPSwxadNGTXgMBGTxdJ+ug0mVtWOjWsNB5jB
lyFnR1IxlqpdJwSanSnk8jhlxOooQGZm5vA+0NNq/5ahL1GbSe2uw3nYr+kfyVva2HU2H+QHDUld
0ohjc7AMLNQsauveU4L/SSoE5nCejaYo57E9/kYqEFMJl3GQBR4eWLLkeGKmmspOOsYO/DFLqP1D
GsdLa6GL0C/PWEmBWa6K8wvuZRSZLS3BJWlPy49dUYb2PjMymkCwrXczZ/ENLHftqahZV4bpFAiZ
bXH/vj6vzbPvxZ1AqnLclYJmNkBV4YQ50opkaU5ZHhZVha5VWv0bgBv9HqmWdrq2UD/Vi5txiFEa
6mxowpiZ0u53XblY6OdNdG33VtN5hG7KbENRtVzv/tzQFwbxzB7mu8lDjIVWVG2HZM8ZrQaEOHzc
XOx71im7IcziqASV08eNTFCqXfMqFcf76I8fs2OUZRrU4Td9k/F2w7eJA+L8HGBnp7XTQkvhcEOJ
YX1+IkM5LkzkyQnVwz2NYYAqA/0LM+ywuqI4O0Q1BS/Vr3T3Mpfo92nwsYLQbvUo6WPmGG2zAUT8
mTahEryWvwhVW/g/SOr52HiQpFG4aA8jCtMEV7y+2hMS1KUbS48ZxYGI0mSdTUM2ONM8sdjFls/k
GyyflmEkPaJ92K/LBYBaPolfbiN3h0tuUMoStcAsxEJz1982vS8jxZRWLoHEqTwYWuUtLWjHv3sO
uaR48uzGZA3CxCtfDMKFlYCUyqNlzEiStbNjdayqLWfubZ9pFhsGUTE/4wXxMgQP+ZOCbLN8o1JW
ZVX6WKOhc9NLwRn07PR7bfPepD1YBeAqQUOv2BgcsxSxKpH9d4Z2MFEQp/md11vP6Ah4ZGRDA53I
81gF3cgs5VeyapgJLqAAL6VOyPYIljjIMGlw1lVTQ9eyE9Tgkv4WzDWuQuLpkkks9qJqEQrHWJoY
dZ/24XIcLbaHUcR+NWSkCA80aZnaYEKueEewJSCydIDrOy9+PHTalfw1uhCHSsKySJHlc/pp+trr
mwOm2rP+rkVqSBHCViDhre3KQ1LPDlz6lM3OOf0vQjgs4teoCWxGfjHunYJaWGn6XlQzvB/WaRYg
8Vzr0a+AIwdYm09CfbxWBVHjhjyydQik8gXPN0uSwXg9Ra2CZlmntDu+ETqWYBcBXAefdaV1ZhUT
3FoX77WdGslxBPeSJU2h/LTLA0AJFLtHSqL/zZTq+qOWPLTbWEPZUst1o7ApDltkxXCH5wxxmDNc
5Aj33wqepKa1BSeg099eUr9lIwzNoCkvnh6ERTyMuRNR0wxOrJVhsQ8qwKl5nAbB2jsHA18rgD3m
D/ffgQGI8IBQFa7FGCWsItRhUHtuWsHvwtD6fjLDcOGHMwQwUmkYTWnhsK/TTUN2njqWERSu5Q+U
/hqMwgg4RdRYVZ2gIGExTbD1/m/GNz8vRQTam+/XLAJLjrNnP5/oGxbt4VAaK9c901y+0r3GtVDr
U8Pjxv2wJDN6ohXywGLRc1if9pSQL8BjenLeeRG9m89LCakG8ZTiekYo/BkT5cnWhM9woKUlyOgK
d3/T30UkA4Lfc5pSDMiE7BKaRL3Pnfadp6jS5mb8aTLA2Zpq57Dwv90dotjyxtkXG+5GXshEbYri
HwrmuC1GEN4RALNh6hrvfJrFC4KmVmS1VNN+Q/Fi8mfPh19Y1aK7qmQqqa9HVZk7pwyOyOM8KAPw
ED9Abqzj2PFx6oKLLR5yW6sryT+F9/Wekro/60rLrXM45Ls+0vUP9WsabGgqfAYSOETXIY1cCl8w
sbGwPlyCbcK0BdXDGvdhthKOkzhEsqk1Nn1LH1RZkbzFgKTIsq316xGCIZMFycZq0hEwyNKUm8N/
H/Zmrlmqrjfzr9UifmFsntd9wV6ZmnI+o1+pUCvfFLU92NGD+DiRunZIRGMRTXYODF1nkKZD22DM
F50EeAoybJzRAPMVc2a7IBNEVFQqZ9JWXZPB9pVrrATI3cA0xDL35B5p1HniK+sUACeMkuiy4E2i
C+rT7kZQza/lgdxEFrAYcL37FfBEVDc1cIG55z8RhHAJMbVT40jNp4OYVUF4SP4KtLl/kq1wbPB9
aiBNvg+kSPllpyB/8svvanzqpybGE528zmwvC+zKuoimyS1A6ISm/QqPD9z1NdQDrJ62Un5v841v
hatqIw+tLspTnP6CgqNwBIxqIuOEVk9G6pCF7rK8ccgqWfvpToOqPf7JydVaJ61b+Tw91BMcQwhr
d3t2YvyoxeWlPaFC61yNQ9fVeVQ4dZ44Ukm2BYUoY+FK7Fs4XqY/VGXCVWqajZnWWeqaJFg6Cu1j
RCNnhCtExuQnc2I2xGyqqqfQsv8qKXhwupwi8nIYrexCSemeonUSBnWQ8VQ9/znJMLl7f6JQUw8d
NG2BiyLdYYUQudKGOUabG1WGxafwX/TeGkZsRNyepKQ2bd4d3C2d/CYPkvrmccse8kl0dV+6d181
2n/dzKuiQbqep3u8fy9UujkhhNWiK0Bj1RwdN1+WzTv0+cZTWMbhXNEgPGum/yd7r6VjY/pqTBUy
nRw2Gs0i/Yu97bTGmMcaOHw1U8VpJoXZ0lVWeTgnf5gAhwkWAbVo2XAFvgGLnLLny6S/O61Cnmmg
+nr49V3AFTDb7Rx66fs6cOI167sOqTkmKfagQaaCbVQLyWzIrkvanj7B310EyPiu8acXYSJDwRAo
wA6c3dTwoSFs69y40hxKGqaqoaAib0aHfJTjAkEbEs1HnmXhzuaj3uF8aKbhQyHAo5hcQiL/oiht
GDFFv6tBguTbJwwiCmZ3/KJvMVXhOtOeB4Em0mgVG5al8W9HQhDO/zLjiqC1HeWAES1ctgTJTfSv
1Aa5mY1yws22EXB+sayjHn7nfWn8mKzr/3HpXFyRktG+orM3ga9Ckf4o9QmdzlBqrLW1YlXkkLl2
9xehcSWs2a3qS/rhuSn7iRqVf4ZWRaKkqdfS0/fZxNNm/J6j+xg3kJE7a4F10HzE7x4dS13BTyqo
642Wlu53HI6vw0iFZg/lV6R8S5rQvykj9kvPPxqcKRAnjaK+IXN8lv87mwpwGRBVhjZD2nBxiKuP
+UV/4QQo8POhUyYPSh5G1kmrCyZ6xJ6cDZuxruPI4v6FTr4N3UA3TuEBlL3k0zZs10USiPxP9CAB
hKH3FqCb4oSIEd7WQVRlqUf3x8taUvo26S0yPDKacTsnsA+3m6Ga/YwdrmRgOvoZz368xiRWSWID
+wjiEVlQk7N8Pc0cFDZzd/miy2b4c6HHHi/XxI+S84sZr5qK/Xs2yO7O6md1tne5oEQnLxVizXaF
gbbwNrR/PmlwJH/YHPnr67ZNy5ZRwRPgx8ObCjJICClLLwhyb6GvtU71aExtACqltXy/VtEt0N0s
w4AN1+EFlDEvcpjL7/nx27W+1wACgQGHDbkBSBVa5Tg5UPY0RiKqlrALsBg1DsRVovwxWM4aeDIU
yXyRTYwfzLAwclPh2Z13+9rEAbC94dM+w2M0ZIgX/rup6Ncq9psO1azz8WVk7TLD1uVy3Jzv0lCv
yPcXEvA5sqKW1PGXWpyUPp/0O0qXenAQMZPHMMTxtZ1G3QAUzRnxUSvPPcV/N4UYzN0BEBpDkrcm
z0B9MRhBVUPXJ2VhuiLvE9RBouTBFdJtpETWZeDjik7SKQdbSjG6hO4Jm7IYqmT68GyIj1CVvTjS
mdwAwCtZiQV6/7zUB+fOnI2fZqBVGyjePWXK2oSRZCo4dz2sr9pfUE/2hl5P7dKD9sn+gW+RFBc8
P/W8EtsOUaksfkgtk4QEnJDL73kmP0RnllxIoI4E0wFhejIh0u7a5ZrKehcCjz6scs/2ABZ/UTsC
ZCWfNV7tPBuOMC7ALyuyjZaMNBsVN7MJbrRyeXjeWYhyYVcpw9IBkH+vRmfBK4a971OIhBRjaQkr
L2Q9Hb58uUWCjb6ai6e6gUm8/RZjij4op5kZkR+kAUobHsv2Th6K3a5qkwzXALlF/nsTlam+Fl1r
qlysJs+Hmj+/AiR8nDDf5XX9x81X5ac5/vxE/mU3gEXZYjyUljHbG0Hgnms/KC8OapsZ1PX2mfJP
tYiniK86evhyTPFkhukBlXpgePO489Ix2JC/SvAHUqKtEZ8Wxo1ZXRr3HXYfld8e7Aar48396t7C
t3UMDa/ZWuAPopj/bLaGqFTF47wbtT2C+92gYAI03vqpap7tU6+IcjhovVAHnuF7E+PDQnKzGT2+
TFnSvYLZ1WQYlo0dbKazDg9YeXnj5EXkqGiq52VAukABZA6sW8P8Twwov4K/gos7usvrTjaoohq5
1odKQtN4IFOCSenl23aWehCnPMbFW45BI/9XhTsnr7VKdWSAxAy1aNPDrZUQqVF2+4cXV2RZAJg5
Vtryed1ZMw76hkN4ZBH99uu2rcbiMScrukXf5oBsWAm1UzWnVuEsKbWnKp05OQFGMj92UY4sTT9G
+TSbv9zCkKEuzkgeiLT3dgc9O2spJhDcDPJoodzaDCPcTyLv0xslirtWTwjppRh6pZ6004poaWW8
gJyeNuiKkm/acUpCrzTzZSELG+HNIVUkEjoJdXqeEcgb+nt5u9OZWnJa3XVFc2D0p+MEEzHOGfyF
to2x3yRz0vtKMVXSLD/G25n0z+omA9KyBY7bBy36/lHoo02orlR8dDSp/fC18IdSyIbcgu0S60ae
yhPNGFZ4Wy2z4RA6d83ll+NA9tKwnHYQSQt8d0VUslhwG6CMl1SARHXrq7aAfil6mYG8gS2oPZi7
CU7W3bLiVm+ynbfMnM5xD55MuenDiE06VoZbuz5nI9j1vJhunRgHpnxRL5lQjyRISUkJ6zufi1QV
CGJC0A8vTICEeTJNw9ATp4yatABKyfpNbrD2UDedP4x/G2fsll6MMbSoQ6lFnMKCWVdXYD7fswsa
dmcjmVynXvByGgDWcBT4qMiXsD1hcZuhO1Y/S1J4JT/MjgumtBij0I45JlWf6M3jCLXkDclRLbqf
rT47mHSFsvKJ5eXV73RoZeyG+N/J4MXsXI0TTKKdq9rBW8rPjkODT1FM+aAwPxH55/uJwsyGv1JD
/cL9BI3RyY7t0PX+h/HfxHpXhIN0FHEHGgvW3fXM/3V/r+GdBDKbSnLRjnHBTfj/LS6+Yun7EsNQ
MDBrZQazjf75H0QmZWXDQVJZT9vPlfivSs4i4zFP3kGCgBs3wO1Fnul13YVwvZJKYkFIpXodBT46
afdWE+lBM+0luMulYqz+hU98kyj3WL9rZcRAMXmGHO4Ny5eEPuAAyS8XgoZi/Sk2+8m7A+bta/FV
xkZpl9fNkiDCTmhDwZralzlh/yYD4DeLO6PmPK9YHDAhJPrxU4dZK28UbyVFaRSN3xjBsqsMq2WJ
B90AZBL9psN3W+dlfb/ZrmF6RsaNWpQTSQSM5E/dELwDqgPy2b0e/Q8wqR8eKbpbOh6XKlGWiWfe
MPlaXy6Zx9pG7os9Q0wpEYQWT5CmyXYM5biU6eE3+Rp7Cl2YZFRAItALRzRaBQOxIYPU/7V3SOdZ
KPb+t+3IcpJKLles4eKUjHYBbB/4ABMmbWzwfJeoPQYN3sKrmecahEb5JdnWMCTpCOZWN8EBchBk
siTknSHaba+VKm+Avho9d6oI8GVrvqBkI/caQyKOYAWLC03GJZJCbEp/tlrVDH5QPUm9zA37XlLg
y4I+8ElXDhgfGkr36esL5c3U++33HbaZkqyjUyQ7J70SnQtvNpPG3OvEVp/othhPtSwSz4VgNid5
FmH5U8diJvb/18e2MX+qV7dVR/eEtzDffWn4OjtosdeOPC7+QwE5JdWPUZTT4mv4WLAeY1T/XclS
kDd5b8X2EhgsZhJPN0HVLSV2/Uyen2UyKeNcYUj4AAKs+Lo0zjzOq9kC+NrBtK4kjtliUuszqFJ8
FN8En15kSikfpRpuFsZVlGlRTQoxJzt5RfjoDVHu87oKa2OrORQZ/RXChL2LoiY1Esk4Xch7euZP
WDrF/VvbDR123AZ4bNCjjvqOsxu/ExZx04DZrc4dogQRML7pLkGl46Wwpx6XoAMotcx4bpdT//T+
3ILtSOKOYKbmJD+XEfsh248eVKYXVEfhB2DUWUFFKeneRJmSlFMuEy6nkxVafmi1K4sTqxaEuhdR
jgvNOhjHMcKT+CFWfTDkEYC/gEnMpflb1s1SuhLzMJJghxAOmmfTS3YsKEtGkHWAyaGL9TnkZwFy
JH7e13oTrwjDn/Z7sheGpMhUVhdL9Hw1YQAG0XzGy2dt8YVB4gj4F/nDagRsUY2xt45wU0EKohZJ
fQyCJTUA59CCi/JZJC9vcwLD38FUIJC2b3X+i/SOoyk09LAcoext8s4FLlXu5ogjdD0fcHdmtsYv
tExqFXC5RA34oCWcQ41mSXMmnz/0r1dGIAd11waInkk9ScaAneQPSd5q3HmFD7K/2DVr9ntO2Vpe
r01qStLwwqy/uI9X6lwZ0QF7izZhKhvIl5CtklwDyrERcSS5gpn9cDUKOmrKGe/zYDNEGdKphzBO
Vbq7Iba+7CS3FpVpoGd14zK47AsZVzBZLsHaSiPluUNHAvDEzcJcpRUtqbGyFqZrBHP+fNQigKl7
02zPJR7iwXOP8L7mtfF2FqKyAj6MtAYiUyV7JQ3QxdlgWSUFH+nUZwItWOZIbTazKaiJrIyIf4qL
K4VqhueEVJAKmWTGmaqgPgJl6s3YWThlO6UYKSp1kzEmWzswcH4afjjmAxyCuu7HwOuwu8crmSyP
fY+WbLrvX9RzXzgdEbmyT3yHv9c47BEdct0emU2a7Ypf1Ew0ACXfSk0V5RUSvEoPrT4sGMr05UN9
6V9NM+XSmnZ/OyFufi0qAI5rcKjooaK08Xj6ZuHCLD57oKKXgkmqyPA8ey9kL/lErkpcdp/pVWGP
Re5iRh9YSBObzkDctVqO4H2RZ5DLsEwYpQshfeKY+FTzAmhVNji4/6aSWdUGIA7YdEx5wO8raqic
QMwENJG48j/B9ejnYdyXae2gFsfwg6jbGFwFb11TODarJTBgkv1SuaKj6Nz2d8dJBDd0ZD534oHX
dNmzzUI+SY0dy5n7YAq6Nu4nHTUZepfyw27pURrOC+Vf8H6TiFglp5V+MGc1eo6Uq3C9T/pc6d6r
d/o3lxsR4kot3MQNOZTzwqVN3UWIZT/qJu6nYdKwPCwOUzeebETR2iM56D2rhmawZzSWYCdkFsmj
LRVmy4aPUt7zuvaiKxJiEDHrKBV36AnGGnzrfcjpxfJ5rhGzsZMzDe95+WpImKKX1txjW2MvRSWB
Ezv9iFMn/QYy+OlfiG3AwFfQKJM+NVqXFzw3Q78/IX55WEfhJXYghr6WQjZjVzKtIRJaj0jn8Lq7
K2iu7HVTGRUmPTsmCgvGjBfoakXeCKF573kDLIJ7OvjqYXn1JEGqfqeSHbWzFnsuuX/RGpZpMumu
qgd/enAncosWsMU/r4DuLknFUBbKttl/m8GKPe+vZuU23XK5LLQY30crO2yRkUdpuClKDm5oWTVA
92z4+993G+MTtC5ZzgPz8FCfjBW1tkYlpUHDHS/QLeY0OQavHayvexehmJtiHf40zvGtgLjKtT2J
uJk4IAoGic84+p44lBxx0IqyvVjPJm3YIxRlJyV9xtr2JUuqBFWIkjlKv9BA7PTNi0HQ0T+P+sxx
3AznABdBxTUI0kC6dsVjirr7zvgCoicbnEdy7vTOu5WL7re+uqP4M5ToD1AcKwW2/uN4BYA1/rLa
1GU+rpafSlWcdaCEmKcGYglWQYheFo9EWvJgjYxD4rYrpHZQ4HqBh/SIVraI7f2UqLHWUfzmfq9M
lMlgehHf7TQGPnpAVDnG9Zqp3qPqHEninq204ta4+Hfagt45kOYs5pZaksh7Y0tA8KsoVhOj8YTr
IP7N+mru77kum+R8prW8rSJr/AJoameciHs8+8ZpFTG4aN6NmzQl+fu3G9A4vNa2MeZpO3PlSQmJ
hWzciUWgCJu3a4h1vYSA4dtUhjdt7wjJ7bT+5YkczbUKr5oze1lJOmoStLMpguQU4rIiwqfy92bw
1d7CmOfwZoX+M6Hs56BIf8pGS68VGWGO/6Hcl2DD5COjjy9tgjoEb1sYB864H0Zb9BczbiwrdSep
AEbOHnSs/gIvwaxLJzypkoV3NAF8ezAyUiEInNYuDBk33qwrKGU0MPtZjclxx+Ebr4dkSx9+tOaZ
uAtT8s+HkcVohd5MqbhUWAtULVGMfmgTFqdDql7AjryGx/35gKEwkIGLuoB73EbW0pmJ2VAyF9nd
Lh73zJLJ60HaC3UKmp8BTAxckZfv3KWXyeDsd0l33PR7cDUYTUl7WkXQyWJjIWT8U7lw4t+Qd7bg
qOLM1FBiFE8dzD7l7T7c4mko/fg8aInaltgGfOQwFqCktVnnMafcKhVlcfoIS0GHazTROhQsTpKn
Jrk6hg1Ewlhjd35efLk0ACJHfWIoDfZPtNXb1vyL1D/cLh/MXNx+svFapgiUGO+L2qHHdJ6f93dh
a1AuRTwxbCqADkStPYWAaQWQMMLkWVeoB+XBZXOab4pYz2BYtgi/HfUz7M1cOcTlor02SPaaOXvz
/is8mZcUjAjt6i64BSFsO+sX0MJxQrr8l0w6hqZrPxbSinbs9IkMGyLVQxI/i5NBC+uJijb9XgoD
ggZFicBVhTlOBd2h7/gIaODz32vcgEtNx0Wc50M71xT2VaJ7zEpL0LyAI7+GsbJmTEQfkU6f5UmF
+p6BDwPyn5lCWP+a2mzc1oBVK6ITuCJd93SxOMigvNz9XByIShbU0OOEY2aQVMNAODKVuaRzWfsY
AdykOZ1lTC2lJUjvZwJBBHUq84bZVe/WRZ4V1gOyTLFbZoF6wLxPcR2nW62KvGtdQfnPhYVBVI4h
Ww9ljzOmUlLDE7yfKbD45dyUetK1Ntz7ORJUU8aadHOn3D+HiJWSd7eXql3LG4zTiMfLqOBgUwrQ
8TEGkoqg+KIj96B+zRERXWSu1Xm3dlju8fVcsRjoM9khrhpf6r0sgALBDUayMa/tP3n7ZoPoP2R4
iH52LFIjcJrPMasjYdtuPfKxS2MuSr9Mr1ZiYLix7kED8qapDuo7PEmSAbXl+KV2tC8iSTAokLd1
2g8C1mFpg4X8J1sCYvGH0MChM63wN+V7CXXU+/mP1FnaNZDKjl6vqN2riZfXc1T0bvOtV+9RxYWd
VthKJZ3cFWdpyYq3T+GJR9d6nfBQ2CqjdcklbiaquA+y1vtbOHQb4Ez02UTWCxDSfRs0VyO7jWLt
q7gkl3iaxWFHYH3qcbxLMNMHGPSEYEQfQ9JI4QnaxsSMRq5R1pozeUWq2GFVcLjxPP3ZG6qV6uJ0
C5SZ8+BYqmmZMFmTxqSAD1XY795vRd4Z9MAjezgd+Qq4Vh5JRgLLOWyH3iwcACOezno+B3XHyuuk
B2hg11YPtBovK6k6XbMQaG60duFF6BuAKKHBLGFEmiOad+xK7FEPp/uH1H7w89E0cNvGnZWCueau
Ev0VV+SgZuTcw/X1LL22cPMTX+d90yiOZIKR4Rn2gg5WbPgYFslHSaxavg6sVrAF5yOu9VKIeL3C
dp0ZvjdqY+Wy589uloJEMtuSOCkC0Js57ncWJcWtXzTx/5uongsJA37KOvZhLqQHBg0PAYjX4mO4
GuMQ/46f7EBBFzUtxDWoy8V35eFjRW+CKdgKE8wqZs5hgA94/Ny64t10ksohKkY/l6wZ+R0Ubv6c
X8asEM99QSODgp6vYYZpaVM9uNepZI43fEWL3RwETbJvgp7pYt8nHahk1Q550rtH2nzSDHbvBqJk
cT5+p+ypq3Gc8Gxsyaeb0eHBqQGG6skZDb76qaIX8jWlhQaCTefFZ/9IbAdhUz1jiaGaK4Vqv28h
oNF3/LBv9VzJ9D75pwtrlz7gjFRkMpbbqWwaBUN3fznvwZEgOZuFt5hzS7YQ6TmVyh3K7iityN+p
/K7xhIrCDbxEOUbMvy7ZUceLso3JvSdslO5aIRRC+YiHJiSaVWGZPbZZeYWr83plJv9dB2mAX3YG
B588IEBPQrw5nGZNoh1M/8u60xsCJgxCVMw0XgzbhjhNQpwaBIyLgcn/I4BtCm0p/+WtnSBOcvQl
6sF3CuJJwHuJz5Y/QS6/X21W39P6XTy75eipAmemkpRgQpmOMzX3j/poHvAAo5daCYxfvGWDY2sd
zVRrx/aNNvNC8H//ziJvw7b8Zyu1GK4Tu42ZJrPIxj41eHq5GUigarGG3CRoS0FxQC8mqkzedai0
GcEpS/9oMEiyIsGj6Rc8bKsNlSU9wxt1C6n4NH7KmfGIisUp3p/UN3BLfcTeh9rs+wLrajBiubZy
CH0MPE2KF5So8vW0isrfhE3+MiAKz8tzGC5GVEGpGS3t/ag2dlUEkDKY62UjynO+OTI43dXQqaFW
CdC1DjJ+XFMgyMV8S1AJJMIp7f75to/vm9NDZ1sMNO9ClB3RjhKNJ3s/41W6a+kt2wPTAANc+zfq
R4A8XXEVBTRhT8yCKncxzmV2P1+MNAeQMFRG6vZtKggj3h2Hm3PNfCcA7qD1LOnuhdsGhE6d6+59
Du4kGLo6nA7GvAjuD2Jy+ZfI85R3A/CxTe8j0ZIoSUAFuOQNZiIl83vqiowAOcFojtc0uO0tQzZX
VgpnRwp3L9ScOPQvpRY8Uw6xOY7mq2ffNmqZPQhQcRDXYkK6dYYCmT0SB4KaHTM0/z7ZAM2N/AXi
rsDmm9t8ei7nx77SA3V0lBEuxiNMKgiU7Xiw79FHr2frFdIFR/s9J6gkNfVl0Dky900OQdQnOnMC
uPRxUWBwuTs+C7YyOWHx9Blp8zjhq7R30K2cKMuMBmpDzUBLOlzSQTi+/H8ktTbVARV/n4EuUO3l
1MIrIf86TBHZzfFJ2LbISmShSAwchJ5wY0pZLtHdu9+MqNYyvFhCBL1T/ykQbj3T58GDtUfUzYCv
s4f+6RvcJJPNmfw1BMbVVkwHfebVRL5XDwAcegtGoLo4C+ZmK9xMqIi6Opg6GwAP/IOHQLnWcTW+
y6ypSzRS7ajdTotd63lypdVchWuTxuebjb0ics8e+nSJcYip3IApg3b3zi9on1wuqSjzBLfKs9ts
B50HEUqqPcw6GwNAYXxb7WthwSnJeQ17rHT3NYraht5sczbMv7XORqq+huxhhsJyAYmoJirbEm0k
1zlzxDLwDoEHNxsI1hdWGI8eYEfucs/EbiRu/yo1wTmTd8zX9nouqXBhZ6KIYu+Cgdc6xplyaOa9
95PZSBV6jC2Yz1lMtaWfUN+ypUMbBVnu9byr4stO4+adHY+Zuw1J0mh5wHJ2zSBQ6/XhHUrULwKT
PCWhbwpOx6YH/+vWXa8BTKQW9c6k2FgRizeaRwOU50e1nRmNyLNdxSm23oUJRADZpKFRWoA9vHIz
4392yX+Y82E//h78ndtw7oi32ldqfKDqXuc5krQ88+Ruvno8oWUvkC2EPalKxUAhYWfLuRW/mT2b
MgTP3JpXxky5kil9DY7XmFHlgtuL8J54RmoUi/cGMMbgdPU6PPPrXHE0SOVcQGWCJTGp/5NI+5Cr
Z3ESOINtVKqFv1ghQHlUWFstYqAfLcDg0C45oun2W3d083VxZwrzjcqZ3dmoYau4BQucSnr+qHIs
yXei3wm4ZKbvJue3bHMyewgF4FGLF36CXU74uV79ssHmhxYoVgZvjKH1clmc04KbqRP38GHWkhDV
UquM/fosQn5f0TZL0a1RwfgT8UEAP0TaAQ92K4gEXZWH6+qzngb1/zmwyzn1HJW3ul2WFRVONI/0
zXBFSe8+d9PNXK41aZHKdsIXg6RyUcLh5QvHp75GkwU7EUf2pOWrw+JWfMkiu5TmCDFJcleXCY+5
t7rS3j5l0y1uli7qmt9M7TvUMwx1w4b8lYznqbaHq6zb+NSPjGtaHo7F0FJzSy/dM1PX5dX7nCEK
JZQ9UAoq5k5o8q9lN2zNUETv3ux/QPB6E52S4Yxt0JOEyU5xKNn9L0gwBnTlSUoUWhun43FPs7+m
9f0wcYDUprpDpvUy3IUQ8VhE8OpIktsuO2xqHyrorRB3qUitqgNzpU434POBth5Zwrzbh56s64rf
pghIeYLXJGf3W4oMhM2KsR9jZXsp2jAH3Y4w4Spkec2lPLeyFFL8jSnBfn9nFoi16P+BnGa9J7Z9
qDRuQPSUEYk1xgLMHPsI3TqG6dDlGIMyJ1lACwiMa/ILuAZ2LH1Os0N87H9yk2OkWXW+RSRRmuKJ
Bk2BpKbS3P/aAmYadDkqzkSf9I4096tbb6W923i3gz0J84Zd+XIuuBVpvuKB9764vJzWJOhGc3pu
Jw7IxFQdvTnB1+gHbpYmARcfQQXjIxGHmn3cMyCoHh2P2m5OQbRLsP/lkoPFXOngstcYhcZ166f4
wx1iisrvjK1Rxa3gT5U0xDHqiD6Cl1Ixmx98pI4pWyIZ3OnU9IZHZdcCkrYjJlyA8itHrb/71LBS
yMzJsa1OVzOA0kaa28KjC1pkfLTptR5OxLP1DSaRf5IqPVcctllZQ2eTjNcLdOd14LvWAKFO2T2M
X5v546vXiGTA6HXe0O+99XdjgAdp3ioVkGI4nVW5o1KEikTjXcIADnXt4Fx2OZ0P0MMeT8WA/Zsp
1ZEaVN/Ee2PpZCZdAVnrWmwMWrvD818aLiSN1xGQsew5tyOD9xLRA4ioaJT2Nq43wPwokvGYJdwk
16Xl8YpgZPOaC//y7kolqXCvzdJI+OYsqoQJ6m3klb+LzdibL+hZX+69nA5q0EFZUIjRZdw3CJVI
ejbdd+Su93Brt6ele4LGGhObNo0ywfhbqh8pg7Ox+hvnzQEFB+ylVBdR5H15djCYmDNuSWrOMFtW
EZwiFRweiLemk9YnOgiGIXpkF/1WyvCizpz+Z2BaSlxBi0zd4J1kEllRtCMsYBmI6fm4zHWz+nXb
jbn5ookCcGqFgHY0P+xfBZwscED9b1G6Mo3eUspTygpJssNyGARLm5yNv01gl6o81hPXsCNHqmx8
0kinWgQR0md/cO0SECXJdxzgVSCPbq5TvKZidS9C8JQD2tVS2SzhPPWdU1B0KhjzI9vemMFo+mJ9
uYW505T4C+V309+emyTpJPvbIaPapHnRQ361UghaOZHUmb0IxjdvaBp5+o6CVacwFKVt/egN06zy
/ZrvPyxHijASc69aGBitlCxKfEXwUpP8TxWf292qjoAo8OZeevYyO32RWIuTIA5pfmcPnX8nTQxi
9VLLN9GzrmeP8quRFtG/w+uqhYSO9Jxa/BNEmpGsrD5dBfQBDbJTZXa7Sfsh+JRDe3zonZVbAWHc
8Z/6dtdETYjLUEIx19qn79rFpmL/4yqkEWPXtayLhygo6kTmdPmqdT3RQe7pHXVBRgAvU3eHZ2UG
2ZLUQpdGuI6+rJCui8+DXzMHT6oU68pUPw+wYzf/o0Imt78J4yvT+iA+PCOtJTp+nlH5Lnrnlar8
FEPdYGpcg81AlGSSavMrRsRSl0OF3a61223s5BAKBlQkaMbjBc7iKUbFBji6Kij68S1E0Wvuj3zC
r8VEx55c8jmK76HLZQyaDg5/utAhV1TuRxSnmdAKhA6PAyloB++12J/NHZ1nzzek1m0jqUTns9a+
VR67TyHGAqCxgTKeGSgoA/4NMD594iu43b1axbmm2ESUUdVvLZO0M+hSXUQLO3A6JinL7KUJC0Yi
rPuHFkurvT/WXK50vtJt2gqI/q2KgNgqxw23oLvKzvmi+5xk+4GPNLQdDhvTvLII7QOI55UaNA7O
/gg341dEs7S9Xb8J+mlkh3c5H6FRZsnCHMXvTnDmbAGzdkTbhgaFSuwPBVfGCdg+4E/84E1u1t4W
C5SdLAvGqtT+fYSJNVB6z8RDqfjKTK7P/8O25kPT2CGC0IS231xn5HipL4pJYfD9fO9iU9A0Ur0O
y3y7jykPzxgiR/FN+etUzgT36to6Ws1AxnxYSgZATRHKc60NSneo+FeqLtS8DDhs0Cg+vFMqVdhv
r0JtIU7zuatsDOlQoleEEBskHNW5LOiBrK6ohKEsmulHCRoaE5rqZqmWrMp28qzPcLhlYiVM5OTQ
4RlojWW8Sxb0PxYlCObvc5+3RGQO/mWc4ocHziomeNVO4d1x0PTCFFoXYGwKNDNc0m17j1GdBUIr
nuLFUkS1yMY/sk53JMWmWXkBUVntPy2MWZQXU/QAUeoFHldQ6gehMH+r6w0Ls4fMO1X0KO68PLM3
fYKBGtlPLgI3+bGZJHXFjnq/Q0crXDsZ9j/yNtAztD9XbmYcQBCbuV3xQoWTCml7Ff9oJdsDg5Gt
g0dIJVyA1QlAi2eoFAZZYmFQ70HxY+wWo0wws6kbLG1y5HFNR2O/pbeF1OfzyFUlUuQDN611mo/j
zAumuBxHgdZRn75cF2Tv5F808XKb9OJsGrjyOAU5v02ffoM6+9z1teIsOqQ2NvgpxkKp5O1iupAP
Tgjv/Hmvn0wG6J+Wh2J0dwLeAKirynrSAyIt87BqR/uyMjeNLVieBx0YBfQA1bP8VBU+hRv4+0vT
PSeHCDhQjH54kSC8WHcbCTQJce7yX3X0nIJGFv7ZyfCndWoyv6NtNNqXQ+DuwhwNFLH+t+2dAl0h
ZJHuG/H0kpa9nekVzYZq43ckRcfNWdEd4NDBd5WdLEjXMO4Jpw6aweXnjNSxS+uxp0iBigMNO+Ud
qHvWV329Ka3SkRswGYmUC+DC3l/739g0VyWXDIjL2iUruDNFKtSBbiM9pJP4Tmd9ltlgoA58SLUQ
Dy5nzACzNlR77Irhm/q7izUyGpKCObU+bytiPWrQFMVBAhqK6UlQtiBXT8OKA28rLONHyhJ0fToW
vruTPcoe8MAESKS0HfD4FFUQbfGr1DM+4ULuM/fR3STnCdyckxfTeE0XuQpX/Fnmqlsq+gxRAqhz
eWnisWlL8zXv7ttu2GdWCl0dIT6yC4QLVLgf6SDFu0RPTP2ZuN130/b7G9BdApWvlh8Nef4uP0PK
PrECKJxMSraT5Z9gAMd9HMWjy5fyuYHHIUf1gmTvFs/OuJzSBw4Gka1PENsXk7F0ZJGy6TwwrDXZ
04zpwFg9A4tUNZYSGdQner9/sB2R7mBndTP/HjCYN4ImXVzBWWFw2kRIg/fYvi4cQuqkECAlKelG
Zve6Dd7A87/QTrjIj413nvXIWN2RhgVCqFK/sruUWBff1NWVQ16DmbrQzvJEAmuo7sp0vOym0Nwb
v0isx0HnVJQcaRMU4FtPW3fmmmslnAMkbVgCCGueUSHgFr2tj4sgtbSvDsA/kQp4Dr914nyRiBBU
gxem8r2sJfWC+2sOQxxmrvg7gsxNWcVToUy6y0+5uqJYtZmRffli4MDBMSolewEw4QWSVVZ0yNiO
VgtzaqV22aySAR0M3xxUGwEOq61vzBDOvtLXdApK4D+Xh2cTuUEJ2pMRPSi1eMX5e6QnE/6kO5xs
pExvUFsgJDlLpYUKt0Tq21yOL8M1GySiFZF4EeYI/bhUj44uYUJfDMM6/uD8/DqqxxZ++P11kER0
mtThM40aOM5xtdGXdPllilvQjOlEBfAtQTCIrt5wH6V7flqEVHDiG0R8qIWZsHrU27CLidFHOjER
GE4Iu3S06MXjYWnCcQ5ie9e7ddE5/wW3f6+llq+S5n4edPRBrDG0Z6o2jsUI8TOkPpLoGjw4r/lw
cqk1cM9k08Fsx9berAULVRcfVBoeXMIPrhcQHhhrS0MLbfBg2jsq38vaF4u8w72x40ys4pp9bQDV
Yc1HpMfN22ClpplCKDbvQeh6Csj6w02zseAX70Lix1//u6CZRm+ZenHYG1BuqG8glAJ2j452GRI0
NdgifM0Z4EaQmZXqOu2hBp+z4kC0PmVmaYKiWUFh91ICRuQ8qNtLsk3LBFTpANPS2jABkSmxwpCx
qcxNqcuHWV4fTgz0Z5W0UKJOpcJFCon58DRxqjqmmMf5QthTQFiTvP139D7F42JRV/rQn7ZlFgAf
VSn0KNrdf2yuNzBdxebYTYM+1gv4psUOFZG9xzWusgshaDLTCZm8tPbtmk/SlurpNJaCBdfN+rIH
pt9h4BK3iV77Z5dj1NAk2cY68+4JqyKKvM981Z7CqINUrc3R+RUZE1EWU/PL2w4+L32SOnZPF2Ku
9S45w+GHXyk+YxXAzQBIxEWMSaugi2b3mwQoUr5CGrceqsrl9p6mh4bazx+GZDR4Wt3QX2YRXbcZ
PKqnz1dtlC3mVoo7sAKc7q3/O7aKCmge/E/8lwS+xE6JLP2TEianOxrs4aVLI1XVIxSb0ngbaB+2
zEa4k+kVUbaRwNs83VGV3hmFw0SC5YvWR3/HFvxXI1U1ZzYEgpjTB6tIJTuRbVUokbqqbmU2at7/
6z/W8KXv4LzLAV7yaYMl1lt3WtWLTNSOrBfl8Xf9S0pO79z46WGBLB0rFh4qC3Qr6PzbG/IwVKha
Wz+3RUoDlnvYyyJqCFqHPUNpuOyUf6rKLIdgjH78/IF8sbOjlkr3vMMFndlE6+OG3WvWnkfIwvZ9
RqnH3v08KMmgeYcu/+RL2Q6Ijd5Qsg8R1/I233pVq8B2N9k/e6dRIE7nc9K6l+uNqMpr3y3BCsyE
0v3RJa7FfZhzRhJWo+IjzyRQfjV+2TS+oGlZU3OFDa5WQDAsea2n+GUEd+nqiUEpUJL8/gm3Cnef
MJKkBdykGw8KOxr3yiXu2ponMA9v75lsTIlE4LX4eSwinsl1dm1+yfGKdBfMvrLgaJakPAcBDcb0
840qOqhizYlB+pqemUAKHAyyZJZooYzzDEXsjfAaMOP/Y7YF1NeKMoA+Co9XLHJ3OYqgFkQI7Atc
uKX73wBJum0VCNNZjS6+oUCCeMejrMDMZlzjlFLnNnwLjHzwRm7vwv0TMqDTO9ziOM7hJ74OAsZh
fmvv7m0HrvIra//n6y3/7uYoYbIMMXyBI6fDezSwWambDffycafVZtiAxY6/KYJ9Mh2GYACHP8OO
esh2lkooaIJ1HxyczrVZY5IFLCXEyWTrXAV/ffpAQn5xqmjtxaVtKTu7vzjAsoFGMeigOZ0R63+Q
upsGYCbragS9hNU6nDBBicv98PVgovabuyXFymaEQqdcGuTPR4YNjoTO7qK9W76TWDJQi1K2d08t
dpLYKsoxenEr0br5uyeCRS+HavOutegNLeo8XTzgqM7g7rFHwvV93RUcCDhfDAVaaTQH0W9gzx6F
WYk+qcTZ+EVQE1hYnkz0dxhvG6oTPzYEAI2bLMqso0RINsPxS3oHxPfGK7QtLVl1Qt6a1uzKVRQZ
6SLu329V/PPGnFGqFyaWgKLeIMWqZ1PROznj/MLD2IPFIf5qAqDyKGKFq7A0s+5FlO3m+F2n2873
TlLZPRC5P7wW40K3m/zr6JGLWTU2LmRumZSO9wZVDU6dhJHD14UePYVPTfUdNNisgYBzvaSsRZ7D
DxcjN1O4ElYx4hlGgSqodmi3f/6STcAjuxktIaaME2ziGyukG1uXIc41T64pMW5tKLCtzQOgtbOi
+snNsBzlYJTlLquOC3majeSmAToLNEFdyfpoy0Z3rKvqKNXFmWlw8Po/k6V5PYoYBUTeLkB89C5p
ouBYA/6hh+72tD1EErXw6HdQBqqSk+i7r2hi8BRGDzplF/ainZMZDu6LEYn6NSnclcN3vQ9lIk1E
HLW0XRaswIdavEPnyAJ4E4YxkxxFtevuzsY4rFONBec8p2FAzvM+K6FT7igJhCBJf1HNHIVh0oBW
LrL+TwuFPIDAGO4UWL2YuhpnhcduwA5WjTKoQf8v1lAcylqlsoRmv6crMdRo9ZfEmfzQho8u5WHS
k6XCJhrjDngN6edlU+/wmOJL6lcwl4PgfYDhfRU+QAWftm3AxsKY2+viSF1D0i7Yqh+MnmYEUWMZ
aXUUpm8+fLltxozJqzoYPjp3yPp6SdhcDWbm7QgxZP1ekcEGpnfnSWjT8MvWBQrja7eqXDIFKOGJ
rtFrBh7NfCEi1ouyM9mLRaJrHwQ2qRwuVUijqYA+7/N+6ZR9ZSsOK0mH5ZO3L+OR6YMX/qTGaWMD
Jyiu5slANMofJiIlCu2IBBovBMIhrG2zMt82bMngd9xDfXt/+E5AXyrDa52lzc3ec2o7AKbytwZY
VhrSin8TkOKGpY+Aixct1oOV167ECewrwE9In/8WM2Tm6ngt5FhZInFyiiOeGyeDi7dCQIHcLOVu
8u4KM96Y9lVFj3z5M4FLpocndj4wM5lp2J3PhXpm2KTjErlxMC9LQ3F4FyxJTPXAkzVGSKkGZK49
+xMYpJ4J5/sT2jz6eg7XSTb1yhs71rXB+JYERd1SgO4Y8XQcdDT6ED6N7kH1+CNRN2iaJOiUgDWN
ISZnPBOtrKbBQ0I670PMuyDh3kAum/uCqWsVNWFGcr70UV4ra+WWtVQbI9/6u8gbFa058ovqfYXE
cihNV1Uv7ucWqnC0pTXE3QUjx83Q/gl6XtC22SsE7DCiyyAy8DED7aKaCQGyy8aNiSYNJRjhYrbi
05juftIuMy6tnxzz6lRr0GXO20N04se7lbCV/1Qqz8MC/V+ZEoYs0nsWANlw4FtTParXgg7S71Ox
nSqgHlPlcailFLNZ9DY08QqKUhZJDPcIToeHMRnvNqRMRm9g7AoQVaooS8TJYfRYGvfkWzRyuYpZ
JHlxP0Jb54EKKiBxvZtloI0C+pK7mqwzsHnG1ZLyFikpEx2uC8apamUmD9kEzYjPrlFjN7SruYiJ
QO6Y+wRUZMe75SKSF3Q8huwe8wpymfPQXHhoKuChdbpsw3NTTO3v3TEexK335opGtwCI5gvl9uki
Al4zziYdfW7Ao9X096Q/jsQun2i6bTDff9/VvaKHrlXwbqBEzz1M0hFR7OXtKjy80OT8KQcIrZ40
X2jAfKohdrvT88T80Bbsvvb4f8eaTK2O4/VxYMC/pIJe0lBri5rvs78cgT9SuuV3YkTw88/FvCgJ
HXo+cetnQCWSeIOqAYn8gB6uEukEzD1Ac2GEWK0n2F3zB2/lo40fCHnxNw1cOR6UJ46QpUtLdDxZ
1Eetj209iGUmXpT+BTGLnQlMhaXhNUljKoy5FI/adVu8lMUhKIO1BnGh87GuaRWhr/afRx7h4dZN
Bm5WWrdnqBvuxTRgL6hqSqwNbgiEXbBuovJmtqup71SmNYL7YUIygnA9oszq+gp20LKSIl5BpI/p
+CS4T3Fuu7n4dU1+bsCNbwJFXjFBkzTqEyaYhfT0POHUekBUIlnzAtWkMUcGdKwHksigq0DRJ5YO
XbcaXU8Bx3rD8qJojZcA7XY3Yip9QNnP2EyCI24lCa+dRnguWeoE1ie2UqsgO0X43NvMBVqNwXob
GWBKhje3w1VobhP5lCgSi+rs3wJSS+uJvn89v3bwIr5axP4cTnysppxoQq+Ju4nzX03Iplo+wrJi
+mY7NwRkHDVlXjn3IMcrIFN11YJ0fgkWt4PlfDc/Qy/2JdNC9lfRfw9lLdeF5UTh2rXlWwDbGV36
2MHYV8VoEUI3u7tPN80+W/ku+WSxqSfbKTLl4QvKKEdt4QcGUiEhRPObVa+JitvzhdAjrs5E7a5r
WVAhX4p4e/2yBBFDFcyat88M7VRtzyVzLBJFoaWFMJEr4hPtWujjvYA8fPKTTkZeWAt7Bq0tPWGI
ydN0A1J6EeKyINwTAiO6rbjGJs31uCAAyROxh3+nd87IDjatMhTr69pmjcp0JAvy5Ipt0tKEhfpa
lkpuGD8jrpYZ0KeezzLa4RDqBcvDlbdAh9w4zTusFmzSOzYwd8pmnBKbrn9tTXThxVQMrjh11Wgz
BVcKU9yVWW8Q9Vz9jvTci/3Yx2JHAso9dp6bi7oqLEdvynrTvaDyinmgOxOCXU4enNP7FePP0pmV
1kulL4C6TRtpT0UOiRU+mNOioN7Wxi+M7h21WA1JAwWDOOTKYhgd9h2EpKAolDwFeKljvYnnCPZ8
buEbshNGqI9SfV9M6qv2o5uf044ApT3dQCADhpbmbRaNmvlmiv/2kWlpv0Msr17bQrbCsrqnQCDl
I78ueX/Zl9mFOoG48veMKmPUNTI1GG9kzZeFdX3Y+B2jKC9rD4AfnRiWys8Qq6nnxAjiU9KnlZdk
7zaF7J8oj7iW8jJUDPzjWELr6yeQ18xbE9a2xUy9cLRE190uPNu/VP+nZNeRgUpJHz0bL1Jg+zpl
z9ohfj28eNULAfWFXovFEylfPfDLwas+S7rrSZesjTbjAHaMNazAmd0WldFCr9P4Wh9uAxAFWYxc
Zo3qRxIoBvdwid92ZguBicC8wlR0w98QJRvSn0xm+UDvfmXvOau0PqS5lxjSf4duQoYneLmLAchk
MLWzwnmItHCvSs3GKqpQVBmFvADEkV/T7QNkLoVOJLIsWOodu5nNYq5t3HMcfNQcymdOiefg71O8
GUyMTbWPhYVyZldY8jCGNXk8WWp6KTQGqOIRg9/tsXIURRMTlYhnK0BbhzHf4dJC3GvESGXi0PAx
kC6GuM7v7NwTUEPC16iVIawrQ7r4Fdjx2UwFlMVLx2I25M0FTfBCKwsMfEDipKo6dREMsYJ6oA3T
gx3S8wRKhJSfH+Y0I+YGh+gp+6qADsUnC79XC8tVbwqGWGK+ryfP4BNmbyWkzk/rnBIK1+9z7xDT
T6IZl81EomPBdcLZE7fEamT20e8aRAu94JzVpHpSpwtfosMVkKDJgrePRwwotO+RaXSxXURutt2y
D9+S052EpfAxJ4UUExvwxXtFYrmRzgdU5Lit+FIfJrHwknF9eM+lQ0M8hkbhAQWmnOv+DZdSfpJq
uzP//GlBmbnP6dRdpMYtEtDgOXbckNzUx5jJepChEtFtJHpHj5ZOUCMFO8VLxk/2ubfu5EyeHlDm
Cgfh6AYPj7nl0++/twt6/pUYoLIeDa1lXhNiV8fYSy4gbJl3GvadZplb73q1z/sxuuC4fmPZmoNJ
i33KVyak9iq4Q3vRRL67cybbBsZiVMuHUILjioTf7lfbEIMgoMBxj2IkOCF3b3Yr/sHtUS3lR5Xj
nUlKLwNPEdGQeTto+Pdq29sqTYD/FZ3E59gJ4WTij9zHA1/tI+/ger8ncJh9l3SUAdC0M16znjYj
u9cPx3swxtMN1LDB9KLB2Aq6vcZQV+B3iNUwXs/TuO8p2COr7yoHlL31KSklTYyiowulJYcP+PwV
8YZGgow3qXguhV4o3EwpyRDaKsONIwt8dKTu6RjJUEb20Ohi5M0OKfoQ0ewwdkNKwpa+lAMPKei6
MHePN6MVSfPEYvAdIW6qWukA1xyTPZ8WpVFKECfti20QmcUufUydfgLU7n7NN7klDnxN8cK6wvUH
RQa3/9uxy9Kl8o6WreKl33y06YfUAUTo8CrcnbpSuJqUPe/ypP5a/YpudVRBtU8jLqjanRV/wk4N
uUW1BNyiZ8LH6xVtybKnLEMCWN0Ff5KXN8zxuezilfRtWTv+m6ZX2zqjtSWvU9/eN7if4NOIB84l
PLGrzwMje/bXZ2XrH4PYbj3INhYPnbERUF9914PyVaIFBEMd2GgLNdwzIQtaEGjEgl6hW4wOdczA
4Mi+tuEZn9Exg0Xfznov/G7RnWdPJ9xsVFZSfgGWvNBtMJ5SlYrLElg0TdKsFLwLkAK9QzigC+l9
zR5zh01iVNutNkiTTX5QyHtdjmZ/MV/czNlgRpi+CZJUkc3rsCbpR36f0kcQ/HQelMlG1dtrGj0P
0IcU/ZDDa7FQH03oGOFnf4SfNlVZWwY0R6+SaA5aWxZbtrWMFyNracjlmnk5cLvy7Ofp9qW9juhr
/B7/Nz0S27F2KyGLDf+TUo0saJDZvSP7X0JB5mtmBlXqeFZVEbuvpfDIgKtFW+/fV+GAG76DmOMp
awV+EWprzpGrzI36xP/B4kc4PVccZkM20bHQs0pPLmaUXLqdiXwVwcEUzZOUvendiFypx818JCOo
rRk4n1RhH7hpg3jipp8N0MXCHe0SUJF5jBSPIUy8PRQmL6sIwouo71JNV3z4z40AN2gMvJrtPTs0
Yo47YkXpeEtOpABQX7eDR95hxR+bChXbcifXu4RflJWbIT0olJl3ShBEdwTOPhM8L8OBBDFGWb8n
XZpXFc/F5u6tS8XRYzTqdO11fDAjIXAZlGBFPrjH04uyay8eKXx5k5qXDLR9AfYAQodbaPkO3Vb/
KlTEp/TFkLQPK+BEkG0/GM/f9I0gXZ0DmAAbFo4uvqdMmiEYQAQjUUQnHchkIrfYnLNyXlR2jKMq
ESnJm2He9rA2ARllZWs5Qg87FLh+CbqSCKvCYCno4DO2z96tEcy2urlVgSA25btfUfU0PSUiTcYK
o/hhC6nH1q34GA0rjpxVi3DOpu4BmgoLb5ejVa6uWspjILB4RdWGoyN9hxNhdGGIOCLvgsUha8V7
5iEmynuY0GWThDIRv5EzlhuTG0zvxFG03c2WNWbvBCq9FETtlLRyKxwdYOrEmjy2j1gQoLjCyt1H
SWFf2FQUMJG1cjhW5K81qYCwagc6wUC6G6TZHVAcg3reF3MWCz+74Xf4yesm780NKqvGibPrXr8w
zZMT/ZjJEZFVVrzvBsdDlHf6HtGvlj15XDiheFxMWt6xzGJhtXFg3aaEP+YqqcG+YMH7S7UoL/fy
MB6hDo1y/3Qwj3Nq5PKjk55tpsItXJiPyVWGs75UWC73Ji2kmh4W2k2rco9e0q5kdiuk4KbEUw8a
Mp5II68tJg4hLWh2EbgB6V/AJc7sVnDfjHtuhcFBuNGj+q/Si5BiXFrrORwI7RyS/JYRiFqd04Wj
YluGLBl9soXYtsPX+LyzWKWUP9QZqt2nQJEEUuocutXORhWk+sJ5seu2rgNyubVfSOtj6Od/viRA
oaxXMZ/4IwtM32hJmbqqx7g5dk54DfxpHNSqhI2X7of+nQDDLbbf0l/R0dx+tmqVcqJji+AoOxvM
trGkwo8CWwHKXS0NVnBtavlpDYpYqpnO+5sYvCuC3zVLIXJZ8Z4CXAD+zY1fJxi+bb0IPfXBacEF
x5APOQNCZPVdEXgN+k5d4Ujti+dPhTEH7Pvq8TKu82OwNw+p5NU5P4+sJPARU05VmN3Q0fBOwwoz
tvvf6nLnQHoRs0K7kJR13c7VdiJJ55jWABdCXDOETfVYAiip4FPG07bO7/TtIk1jZ2JN0tusjjf6
5R6xlBE5dJXlOYfIfgABoQszDu5ag3Y83LObaeOpQ4SgI6b/tlvqbBKg6hXhu8n/3R9QGsnqsSW8
9c9oiYWAj4F5WLYHJLyivt1blinSoTQ51oG4GevqQ/a9PibV9MBHiqkMzvIZ4KSDGnj5qbamCCws
t2sNwd7FOE08q1l8MsEHg5d1V5GTcqAbPr2JFK9Gxwoa/weDGKXoe8/QjQ1KS2TYCCu8qkodnHA1
UKmiFutK6fnsWJkXQ2GKd7560oRCWbbJcRxb2E/4xXJUqczDrTJKdlyYV32KD5J6ccJJps6z7dlK
yVAUVmi5SHaAUshv0sqc1OkYnczHh+7d4gztuiGn+Gn5H9E8PRIcCY7albdCpK7kiwL/bKvkXGCg
oMLe+ZH5KarwpPVkNU3pVbtyKsnsWTHPjDkDD38y6v1w5ba+PjymXEVsp0M3DV7XseJgFBUaLdhr
kGpoUqAktzZ2B3BDjGr+8ZyB4xptD4VpPrc4P09tcu5jl51+/QXanyI7xhsUsyB3F65f1D/OO+PA
0jBlOYmbMK7ZQ3/1JIDgRwJKDYo/mW3YVQuba5osNrMJjMp89BYs6kq97kjs8OpOGhNZmmwlgM6/
jXQnAzVuKzQG93Blw6wxlqmYX61YJyOlzGb3E+Cnjy11kAUFsBhuYhZJ4YBhvYk/YOxsN8dkEMzC
Xle32y5Exj58Uj5P9jt/UuNfdu9UE9YD0JSYBr00pH9YAQakCzPFVwYGfr+jmtvSdjlzCC+NTchT
i9r/XYusGdCVOtsXwR9URpDdZHpFsyXGSP4Qk8GVpp9t+SMQwXPTDscQI9YIis0FRl18SAa4AHZn
APb19Sm6+OUZvf4TSeHohLVQMmfTnkhlqTLejPEddLr43NW3ktg4AyaiWi9rk+BTn1RC2IpEtgN5
iyFkvGKYSNospsTFG+hZmnuWK9xIIJ/iN6PhuxuzzNWVUp4RNg80t02O5Tm8ao3WT4M19E7MuRiu
KaHZ9bSbsZceXhUJgAAr1fLBQpUR2emFnCwB1AEduLCZrlWo6+jmAD0RAJLEskBo4IS8AodKHDx8
uXolTh5cm8lvDw2THuoCEjnRDCf1AdgoikTqVyJoagAdaJQvOO/4m4Gbq0LEfSBTNaVEVj8WTjcC
5/TQEGSXKt/0OfmAdayjvxJyyCXcyrqRNvuwgLS5J40r6R9ej9vmKyCgHH1Yst8qVcTYhqCH/Kb5
zApt1OMCgeilBU+dGM8PBzVCWRFqzklhJkGsbRMQHLIbudbdwQyGRK+tmMdncFOSRLF2fHiwthRA
ALs2iR+k1sqILr1dLnEMasYMam2WxoaBCz2lIRdp5vuScQt1KNCOKuNcF+vSwZX3MIcob0lXgrB1
gHNvqFJrxwPIxoqYFWrX4WcFEUSB0i34YZ5Lm5urzJELB+RBkEUKot5+jg5XI2Z/v0QYOidd1noO
L0BbyZPDtg2h7ok1YS/a9suNWKJtCptX3vZMfucYnSENT9Q9JaX/jR/Hlr+tYj2fpaqEB1GbvkVo
MZw6Oarfb0x3L9Wf5jV/RxN6BinPVAChDAHit6KQWG2A2H0HPtEyZJ+7RH15n3AjycO2RIJ0lD9u
M/kqJtWLSB1b3FID2CUR0g1M6dXHTcSUCsW8YD33bCjVsOxSGtIGhb9UgyVjumb6pCJegBDXjt10
3w0QkSfNt83Ib7lJzxSxQYcqg7XnyNL01bUFWkQhvGsUiM5lwsCQMS9DqAgc5Xu08KnIXGL2H0S2
CXCNpSlEKjqSKLAOTI2J36SOtnh7mo+HU47XHPbly2vCxiU6YnvFUgiU6SoVUjJHCpKaxj1SleVO
FyH99iFaCwoPwK2DHetFfFilH60lRlcN8XW4/NBjmvh0w9koE+ndb3qC5Dx6PM/q1NgmlS8lBPvJ
w2CjA3x+cQFCN1+CKl/SYdUunL+Iur6S2JcJUR9hoCKL+2ik2oPyrk3/xkiFQaf1LS5tD5kgTKpe
LS2ZIIuN2i2E4a5vJ58pmmWaLtg3w9q0KPh5JeXKdMNiIjP4Nj+X8wTSqcfE7ITuTx4p+OO38XIL
nviKXp5HETiY0B3+/29o6YREimEML3CN6qrAIkUQ49kY5fW3tgKBCibtuy+7XVJVPR8ysL/SdCrP
moXNf6FjT2z78cDmz7gMbq2AJhOKxAQJqKtigA2I+R0kKz0sL65zNHPTFfSwOZJ4JFPoJlJQNBM8
hxhzwJ1sPIrbNd/KgklGJHior+uck6OQLM0bCLsnPl4XJDELlqlVzra/QIcp16GdBWXPFlO7aMIM
nPm4rdru/qZuPrQoxLxIeu/j4WCCI51qaAP6+CHAGW97OIMFHxlRC39XdZu8Ah5qdhU2uc0gO6da
eTtKDFCUqQfaNckH/S4dgXgIYBItL8hX3VEyo/riEjBmJ5HBdyZ94oBn555HURpvhwOZdEe7kOar
prqRsDfC1E+NmDYPdPTCqO0K+dABmwX5BxFiWOdiIXmw3CfqA3xEwVucKtTiGwQ+KocVkaJYKGyj
qZot/5kIb4/28CS5jfHxcgrlAe65ghD0Zkowm+n5eBf85zPJD2IjCQur7sek1OQKK0GiOmcSuevr
U2DmGoElFI8lah/EQdOlpS+3dLleCCbZdmtN9wFHYhxV3rNnn93/bOF8A530zywCizzfEdmL/KsW
ob9JuZo5iKMl1SRfMlCEaq01YJx04eYIQqiFhGwrUQqBOpgJG7j/eYMogus3GRkjmGeCEMqvbBpq
UtwpN9GPwcZIIxxYdOmXzDxS8DD0SeGJikVO9hJrD5kH2zFYJaz5OS9/i5XQ1LZ+j72PoUs24QpS
c96Y0c/gWXdb0DYHde2cIEXLgxCGti1IkSMaTBRjx1f0lGoQviMZ8WnT10tPLNxLAKnwyptzOTqE
JoZu6ok29PiF7blu+ThqeJ37wQEk15e6LolMPgR+wmbJzBFun1tODptb6gaEXrUx+yZsKIWUZjYd
w8q5tN4vcL/sb+wDzAm+EXq+fUyn9f/r6i1LS1nel5nQU2shkUXexg2CnmKTzhKL4IJAXhDEPsw0
4vvelkfiiWXUqp0SAiKO5thFghOr2X46kxMzG6hpC3LJ/QVjCk/JjeDTwQMLXX2oaBvYzqt4ZaIG
AKeNV/DL3OJ2bPJh01WrJy2l7qh1mcVV9HWwRJchPebC85AbeviAzw0KYyO2obJBItJAvWhszZm0
hg7WAXFMkNiCCd9aw7u2zGVVqH2Ght2sWmUtisTe7+7DHZdnDbvdsSOTt8gt51GW+EgGQIKd/X5F
WRARXDvmYHhU43u3GcQKyu8Xtxpz/jC+uwwS1kN+4HFisfsPt3Ixw8dDwFEdlZpMLFFXhZgZk9de
j7nhksutHSdhysBo9ORKio0AXuhHW1nj4g7ww8+/x7WSTLfqoxq2JgOkS6Yy6fQXnljkxzurU4Pz
g2swySOBvu5FGSJyPo9Ecj26ygIi+hglQHGFjrujGShVL+EZLA/Pp3wgznzPfhKKgp24442HrFUQ
FoEZmIrtCg2XZWa6+PiooZivf2YkvtgaDuBLVoSyZ9cc0WegiqPe3/RdLKLwBXDxasFPKCdUqzpc
/KhtBjteyM9rY0FGAy7XYHFl1azkITWZ3r427DW1Qukko949z1th+wtTfwFxBsuWMNz3LtD884pk
LS184Tj4Fb+qQxo3LKB9ewe9LuZ7yS5EqMKk88ETYuVZ5t/rwldqkkh7daDE99i3+h66zF/Me/9a
Ciw8HshSBNBmvl3cFSLtoRhRA5hS1q43ZjlHVjcdUWx1ixjU+nFAnINvEP3KaYstDudTmZ3TV4sH
lLDey/15Gwsv6iWOuLZVy7ovUxDcaF9csa4XCZVgjVRaWMR9vTb6tDaDl5mjujtJsniOGKIkTcFn
OlHeK4jLqVnvP2adCJt6Q5sTGMilzlSlGtHR0mRKJan/NMv82yf/2JvTw/og5KEiQeEckkkzWfNv
m+/SZUutaBm23wypItIaFfm7TSmGVk+w/kA0UXIz4il+IkaHq3TqtvuBN2QsSp8WxOhddAedmaXS
h5/mNQlYlWy1Ah9r1W23OKKjsjoIrs6svZPsFloM5V6m8GFPzRGmH61LOZh2VQL8KTyn5iu+pveh
IW/hfvxP87WKHrZuywvazAjFSsQJr3+VRHBwK2RLOql+xpqExPGpN2iwAsEr11gBc/ygQenlSJ0P
eVsFo4FdlNvp2XrVa3Kr1qjTWMuVXtckOFElR8QViCgCtTg/4/XdVKKLYTrwDlDyRFduCxtMuXmP
2O4A6qbPIT6hz+kU8MDPUqUi8HCgpZL3UT6FOntEWI1p1NBS7GWsP0XqMy6FNiNF6fcYiXD17ggs
R4N3N7J7NpKhbIUfru8bXHYmu96D5aw99I8HXM+QAE8Te9rdnKt7kUMy+tDJ8+hV86NYeQ/K+2oy
O8DvX4LpiINuEqFCdJedVV0thwzIeULrlDPB73Ke2hR9911fSqASi7zus2FAi5vjUcksSuuLCpVY
MC0gTSRtJ1JAQVMjfsjWlQg0K2MXp3cPs4XboJqt2pT0gBwxmc1PnHHo5ZGOGKAKJI6ue5wN38C2
PW6o0h2FLlz1fnlwevI28PRykEqHkSr1HHcZn/2il3wWWC0Z3ogg5gDWPjRAmjgzl8rbAflccIc1
jOL6JzVN2agGBN/Eej4sp3hDCaKhYjtmjTI7Hcnx6FxSpR+QyR6xYdIH2a6lFnDkXoY7ORmUwgAo
eT7tNpXIQzi1J9a4TU4V4er6TyLiVvt6wuFcBVVeQhJSbv4y1MdMM9V44AWX9hjClLK4a7EIt1Ae
9lEq77pNFhUtEZWOing0yXKmkqMjdXZtPZ2TFHNMYIJt+gjCNafsxpq/zxaYDHHXuXwG6kMjMCpg
oJsu07eg1wHSlgtQGuNjKD9ct3ASJCTYWpjGg3CyY+rGKj/CPDpVVa6zOgxb/butaXmA0uhTemSY
jNYFEUp+t5U22BRaRUTfBvqIzbfiT10rYkWXCk9AJqQ6sChlN2tWwqEhEvCO82P80v78m08bDkQ5
h3HEF4Yg3ZLZO83lt1dVgYewij6W8bqMx01Ou671u29g2gN6QSxyUy6hyq+v6b/hff+c2mIDFX/a
l6aKo4jpQt8XrFEz9G+nKbbNk949E/xsI74BLZZGsMJJDMLOhbZq2xLoCAzm8PzJZnRUDSXsiIKa
D0xCYXlvyk9fE7pjdP0JBExFFNhVEqRqJDUilF+TSE4tdMBowz9+fRTWC6TaNBTyQsrX/57vO0Mo
OWOoyRKJZZ8VTakxjS1Rk+psC9xrfNTaRdmVFHI6hROHfCUf5CdTqL8oajwpwi9h6lT2+PkMpLXn
HNE8LiciGdUGvaMRj3+/8uivNww4OTWulEfMOnXjUZXgQLfgBJliapA6Q88xsHJnk8pCAMoCVuus
68QyIzhY6RI4dMPi6/b0Fsh5SfjqCiZ+NjKWNt60H3SPAkNs2XGeWQU5ddbyyF53c5kESMYdApdr
eFe/Mw8jaGpqGFEklW6IihZvk3lktCR+jZodLHbwBY1hzCXL8kGbxZkG0YGxJkG69TgoGxw04g/m
S8KGbbxjceIMgOFd7H1RFFXGRB8AS6oewW1xOs/6RNFIuQz3X/JpWoG1bAQ8nDkMLHlXnjykRxay
zKRySfphjheg3+79aSiET0rMk3SiT1OnImZ6UMAKTlatZkzNNTPbPu2C+1Cb4hHf3GPFGBsR0UjH
jeElp2qxj2/wNg9tSE0zRSQHHg4U42gR3wSFMh9F7fCiwr2qv9e/5XKwp9Mb5pSqQA7Nr8ugra23
5wywIlEVhV82xlt5VcUbBFxLTDdICI95ZWrKUxGj0IuoFDH8hPx76Kv5jLDbPzHxyNwKpOJ84rvc
I9Y1bk00KWo7p+4PZI0xmKJ9+NY2PV7eMuVISb8F+dygl0p+7QK1MQYETlx2qb5a67ajSpMyeB3d
Q/CPpT0jKhVKfcEmZSMvlyCw9u40d/uDLRWW5F2jRbZP2gI4/936gs9rp1wMmgIKbq/zoBAzaV3r
6NqPjAwWazewuBZsw7AcG/NUz2A8Cwx9T4MQ6+D/1F0MukWrFYuPvoE44qFA3sRclRa647+cvu+c
Hnh+YAHuvY/cXmEZN/7hTOYCF6JLEo9Qma6bJE4Kwv1anby6cLAeFs0GNO7beycAcbDabB0vQPpB
D/69kDq+cDTX3UfjJxr2PsBJsueAc+3fu0+Up8EzXmQQwoPKlPyrSF9OGeMmi3v4PFLXC3sLWlk5
KHrl0ywa29IjxRMsbR/yzWijbZAO5tCYHGilUuXuy0nbr4GEjHbpVrWPtE3NtxTIEqySm5a76vut
euaHYtJQSTOUSYxYhr5ILRosB7EPgVHiFkxWpMSgxyMJnQIpUYDSpeoCSAePRneKOLiPRLMYpuIT
Ibaejmy6gLZvs+0vQ/rcDXCo/BeBbaQvF8qLQUrAVlcFEYfkIqL9MoHO4ZJZTjqkv17eLXXKUELz
ESfd++bAFhE3JURV8NrHq3j8+cA4HcravC54rcNl36cgtTqFSCjR2+Pi694LxjZG36IqXDmQOZ3K
TTdf+27rdiCLuV8vweg18M6BxiLiK2wtQ1i4VmP1yDmkHTU1ll+iYekACS0yWp9TgoNsI80HNSCW
8lxMATCXfF53S7gl8Wsb0QAtdlBUl0Gux3Hr9EoEJctSmrlVms47JiPTNQSm6KVWWiL1akbgimJ8
nHG/khuuJutqB3MGsFHV2mqqNeV73J4d8nRPmyzJ+o43Kx7jt62z5CgEkQ3lkR4eCG191xi6AP2c
T02+nLBZnpa2sCqlhof0ic2PaakBPD14RgZCsaONI1Vi+8wWcxhZOd/zkfcH15lLoFmuRdt6wAhf
4hjr8Pl56r98e2LVD0VHA7ZJzsRZ+Y5kMuUoR8+72XdDLlA3q4vWsfs4V6MJGLhdIRSHurqc9Ky5
ICb4D3UgxpYj69MKfw3q2Cv6ntPavHZrrXv31UEeuT43kADQKVm0SRWNrdYHETx5QwZv/uTVIx9l
A5ApT0HqKIN+YibQTqMF4JfqOwwFjh8RnkeIAc7aQ7rw7r7+uIYgsOoDTWIP9RZMKiJZTkDwBqrQ
UAkn9Ze7c2XUn3P6ZRdLEQKGW52k3sKP8Sza6B1tcDhU8qpPxymtjS+U0eG7LrSyiLgUmA2+j90e
ZNQd7dTIf7TgjQPhP6eXG0paLbBvXxTCsdQkysSQPzm5WQYlEj+LXpuJ4kGbXFAoK0/erFsEESW8
iLJK8+xLzDMyAi+Yg4YVRjmzY4iiYxUwkJFpy8CW1+ZIeqrm28OnwTp7x6cIdKJktYu9Kj2njXms
e+ImHHLVUp1dmt0TEZuvt+KfkW8uL1xEELQLm7sQ5ttDUD94VFydZZLBgL56cBrAb04M1lsSFXKx
ERPw9Q4fpxXKwxorSf4gNM77zOLnIk0biln7rd0pqKuZcD+so37Jeui6SOTPNaLMTgvd8ddYUWHG
6u5d9O4F3G0n1aD6AwWzuX/X1Sad8elsaSEOMabSXAAIBqSifcl3P7eyCkI0X17Anx3jSDDN52Ui
Cl7fzji64p+rnzT4oJuL1Gdc1b4wJT53MgMxNPtSWQMkOP7scpIp43dSlVc9ZUGHLe1rQrCxwgvH
v/5VpDzNpiiTk3ul4iFR0hpRDvG9p4brsd5DkSHmOjbytWXYWzAyluEA8D6FDD5rotuaAuQRCzXa
U2XlvH+fdT2+4keCqpUiZnw3n2ducqGJKUhv0i0yd77h74WI6rlygSMih5Q+FZqapn9yKwZkSnp8
tafBTshbHazdBMKFK9OpIU40wxuAYnPF4RiudAJOsYVgywXNlatFm0fl3B9RWm85iTEEXLuJin/P
GM2HRTaJzo6sCgxeEtZ/ikxj+oqV2Ej1B1EZ0FYnYe6fndv4gMYRTz+GRDg4ODPlKcfA6GQvserH
ke2CR55t0fnD/CjzkbAscJjMbngJFZGQ+EKB/yFB5mSu9PKVaql5pO0FUI7GewJUGvyrZcxdJzdH
3uEcjACXJ95ZHrPsvWjG4Gc8ibjX96aXXNNpOzH6S4PO7uG6dQa7pmWM3yEyjWpTt8yNbyN4K2jI
Pr/CdI4gRnAv7Nrvp7/Afi/cSZ19HKzC2fHg26KxJ5lgpbQhktEbI/mR4uceiYiz1O2hRuTGlV0O
apk1P5EkoLPFcJrMqAXEGfZ92IGaP24OLGmWOjlvjd0eKIHQEms7L4Pgl35ZnLMmlBGsDKSxd4v2
9XOI3s9meoRzDuO/Uu2K91dlH2zDywAQ7exztHltphlxk0kEBzOugQ1CfkW20AYTbIZpSrYb2HLp
kEG/1DeY5Hw+n8nEzlIuWTfKvLU5jUc3h94ezusLALy60ll7q9un/5CkUv3edqV8xlx+84OwUhkg
EyGyAkk60385zEsS0cPOdVTeKgGS+XtxcNeYNmbDnbJkI10l+vcGlTWrrdu2m7eF4V4ATWeZQJPM
N/G4X8w9Ev9ieAkhI3qtN25/0rGqJOHgAN5hcPtICTP9h4RBtwFCLTrGGmWodd4rRaFIizgZPfih
G4HNlYBFSjeGcrao61CbxzIFCfcb17mvMwkmUBDLjn8DUb5pKyt2mg6XHgkxKPGuN7uA/UyHnJm4
mqwJym+J7fP2GXRfcSx7QB+OBA0eULlvqKB/UvkihbLtW1J5Z/vHBMLubwUmSFAPO56K7s9yNaUx
IASJCz8r4G14H6mw1wueKreEfDCfYK0igCrKLMYg1aZ6W59YaLDfrGKOxXw73punVIpQgXsJ7pnC
y0bwQskBNusgE/6PmLBiMzIDrvAoUv6D4siUvs6A2IqnUoBapHO1bLvYF0kSkRrPypfEuwFK52eA
rf34R864QRn8+BS8KyqdaDWnWyVcUlnz3JtsdhpxQN5uA4QbQy8lg3XkseSjMyGtd9cLW4gi0Yy1
1vrL96CEl6WZFuMG/xzmIodkpZDhRSuujbpXNlCQEm22n4EnkxXWxYFlZol6ppllZRF2907Lc0k3
bwQQJCwCMDiHaPhM49/ZyZ7EHRHhpb3j1lxirZY3iv4xfafluXATB2Cz4f/tJAuv49C8FeiuPYIM
XyXdq7yngNyrSuWYXNpvwmmt3jfDZQAqujdJIqSKkxD5zQFPLYp5wn8Cs9iP13LDDfg3b9ikOPo2
gB1MZZykKUCNjQV3ycyGK3QHmhpdSutn95eOM6onjMuGDUJr0Ahlf77qaV9N4oP2x8m2q3WHYp7+
P3MM4OhQuJkGjmWPAxOmmgIuT521+PYs/4C0b2mULjkERAOMEVHWVNe9gy+0VQpE22WmRtoRfk0g
g6tBzNoER2AECVD9olX8rdBTnELDWS5/M30/8m9AvkZY4R2ViPIxlT0W6V32vgrF2kPouuSvXrnz
C7PjYBH0DOL0ud0AfeMSl+fm0zHTj3DbkRXUmXilyRRoaW/Ewu64gfjrTzbO/5cn3yYm9TQArNkW
vb+QOHsQVLWJvo1+FT4azvNTad5kMr4X99vQucz3LECzPbgYmVjJAWZXFnm8G+ZQo8rFT5m8y9q8
rJaHmlYw5+x/SteC1M2qwqG6UNNOpY1/jsyZ3llqVEG9BWvSMRQWAr//9pLVaIWMz+h51BNYMsq2
o6plMD0rxJwLeLS4ewn/UYicHYui9k/wd8pNkfWvo65Qs3HVBa6AV1V01Pk4I2gY3jTowOVug4Nn
qKoalBksETqrx0+UNCbdAqPUC/jKK1MdTCTesJga5p94y/JlRf7Pj71LZVxZtdZQSxdBCcn+/vzd
JlWUK7hn2A2yC4nkCK67GdYR2yekt5xC8S5P0julmatRHhx3pFJwIMbA/B8CG1AMtDF1PUZbokA+
Do7Q7h4jJwb9J9G4aDJzDxU9yLhIbUcdj6jNneuW9YHLoGt3tipaS5cO19RZT5ixBfffIERoQRlh
zN0N5LqSchoLg9U5an0Z3FDzkJqCk2BzUotpIgBkT/dbI3rftojk/jISmaFrYQViWoHWgoTJTPGn
kYpWlHwdUkTUKB5bYm+bn8cm9Vzvhf+qPjW5ZWMxcsJ90Bfj1KbsN6t2BQ4C1TS9ssRU9/KJllE1
i4KuumSaAtMg83ek2JB5Rh9x1UA46vD/RFCxGoMPX/vhGFOSefuGemYaBScw5gfWAPM08wZxG6Z9
dCNcxMdlMNtUIUaU99k8sEmDc+tUQ9PbcXL4vLaCOxJNxWruPG1rheVgrakVlL9C4/dcELSG4+x9
KmlyMNMxaxcyuR5QpZokDtcQluG1Bh0YUFjZoKWkSD8BUeFQNDSGGxcL3AoJhNPsTFEG/cby2zpt
Z10NgynRb8lUq2f/CPvWhEwtOPA/UUBYqSsQZCD02+fTH2LJ0VhhSCopmN+8C4Evv/fCzGTr82y4
CO5HDr8XvbRBsY+4aiX1vudk5DyMIpFNDmuEja3fvBmYK1doPQKj4cGuHn3m+5Nh6q56/X9/ZSCq
xA3BQmN0vBdeTYNCtLlCuETgs1UUzRs5bmO5lqU+CgENCAS4sLVHq4E+1MVc7U8hLzcrLP4CYNBZ
16KX7z6sKF0S0qq3YjooFe8OJ5cQW63IUqvAf8ri4U0f+zgfSNiyXLsivE0t3JDHzRFvJNkWbWRF
73cFKugzhszAS7IN8hV99JTNwXpvmjqDIuZ/14Y+X5IaiqdlSuezdTSiWTtd7cBlzkjLipw0sgkN
ERvWrPt5FATvzcfshPPMPbGwLXTBM6YQQWT73cyqRhXREWoUHiadvMKncbXjTW9Xh8FO0E34wfa1
x6BPM6EVlv4YWv8szjPKaDGKzR+rJJbuXXuyDn6Yf3kfEeZirjdjH+xFcBvNVc7Wja0eWazTneap
btjNUrkTZ3cFs5bHfv0O2TaY3tYbTpRO/cLS/7Rbc09cwAYhgeG58nm6kKSnfIYh6+5MWkuhCr13
PVGx4k+8aK84nw/aWytRYAr/+8xwTIXJnTrrq6VtfvK1C5C3gK81zk1aJMMHffd975qiA4tSbVwP
nSMEBmuvVN7tknhgHTx/V2ZDv0pkHAn2gH2jQ2SZ6IpSg8IDaJd2TV9mSs5qsmgh72KZy5e7CH2C
VTnIOoGW5MQZlDZNUSuICc/K3HkU6fjoBFOEAps3LfwdaoPLXnDwp7Coz6U80niVpM02GeFtsIkC
wWnZI6dGlB0zWHWWUKx0hNcEcd99L+VLy64pbPFac7BVzqVmrAtOWiD98UPm0gV0jridPc9Jjtuk
V/KDiF8LNAz24nYMYQwMnbVRsgXZuaWGvC+XQ7918HCqCVL79RULCPgear3xergFvj1BYBFYoGC4
AyjxLPzZLtOLf4ewZ9iEpHVGBRd3NbZjNWiC032Sun7bp/6iqDh0IlvQeX15SzsaFtA22FrkkZ60
N+CVdIvVYBkrtFJ8CMKydp0wXChlNTKN6vnd2arWXLqJJlxnUnJjwmeeX3p5DJd9To17ZZoIrozT
Iq3atEEw67bNl+QViwXXGIgkyzJfjqw93K/C4boHNKe9dIFMKBhBZ4KRs949o2guGE38dw+hSx9K
Q6EMvV9igHL0v2Sl0yA6sy+md01KWXQm7ghrG/VL5Ij3IzSQJaiFNqgH7l0j9ccQvM2ifh0POW15
fx5qWnisZG1ZXvzgMKNhm+rPyA532+SdRbK2f7DUrn19kTIrfysrrTVOk9t6xrjmAu0VkGdfhWuN
0OFuzBIOGXS9mpsE7WqkWhy5U15+VzC6H/yTrtxstNwvsiomxJ2D6YDtbjuahPGLnIZ0xC7uJL+7
qwYf2cPMBfu3/NdBwWTIFFLYAgdMsMlCMXpHutpmp/HNAWtoNd2s8/SI6RtzBZSv/twP/NVSIKT3
GVMDovx9jVEnH+DZxCEb7Pd9YqVswWFE56GXmfpJtDFw5i6cU5Ir8NptJh3OZAv7A+wh3EkXBpks
PJ+fLyVm20pgPaCQsgPenIAgjS95SBzYqMYx6ZlnyC8rN3o+Nmvb5KWHYHDUrpGnWrW8kcPLvWnB
UXGeWo5Ui5+NlLem4heKJBeWrhe3MhcnWU2aSKtd4e/Dl8SRrihAFp7DDuNmCEUbhGkrc0Ky1CAl
OZ8CbHLM1xPRoB7N3QnK+z3iezj3xvFes5BgAEmSMHREDlWob7PY+3dY1E5xP1WEfnsGg2Y+t0mg
CQnaMOlTXUdvwzpAJb8EkoKSTFKusOQMNSMwJkjDTqjt/qGve0p7Ir/mGmsrLO5kxbzus1/tIcrj
e0dtHlxAFem6xWJ44JCqYpJJ8P/gnWJBJUKuoOVB2X9fc3wLSJJecFAK/yZmZHJmWUGRvQ8fdHzW
1Q4C3xUiXfNRiLQJaYV18lSt43tMF9GJWJCO0Ie978NCFPr4nWlIHfGuE5CwyDNcXAPOmMefsgMu
m1IDIpleYSC+U+rIkkI4hyP0yWtX/EQyoO+NkrXJYax7lnCoz0g3imLZPf45ckuWfCKijcMW6Bil
aZVhlcBIEGigIayOlVXTKvbNudn73z9bFBdXMs+liI9pUvzI2J0CS6+aK+tL0RmlI05/EiVtIayB
9qqncg0LTFNAl2rkpPG7jZTsRPZZttz+J1H1eEScFjef9nN9babfs0B4a2dHQhwEhq6cDhLj/Wsf
ITXMvVkFSVHQMDP86GPskBBzY3wmJpKTFuUM4LPtELrr91fJJn8H7Xp2Enz8NpZddtBP5oQFo3Oq
TDNCVusFhqszNN+ZhtTNl22nccuIrFv1muFAApCebJTBxCG4upIGzCpZu5Y66rcKFInUDrbJSU7X
S+3/GGhA8MYMdHA4BlEbMudCGYy4+fg3y7Y/iG76TL6cOHQhJs1fAJn9BPldJ9mDLMdnhTUadRX8
BKcdmOJZdKC2XtElSv7JgpyywOAOH02bs8i/MYHqCYkiHkJswfphizaPs+OJDrQhduTqPICxxzk8
Vq2LNzQyLGcDQlSr9vs34y3lj53eOEyrdg7A2+p0VvUejwYCWXw/lJxvr3klfVT4KMi+lrUbyae1
iq8Cbtafco26LyzKDARORCHTlqknn04k534D3k8Igs4oLULkR9XfIS6s51/x8ajOiQen8iLQDQR3
1NmE5mHJpu2MzvA5eVZNVlYlvmZqiPmR/j+qPe6M1KOEj7XSznOAF3DzWyAIg8Cb4tAzAG7jOlKA
wnOQw9cf3J6midl2CmHazyysAiTZR3+mGin4GF2+QvpNf/Z5L4hYQc89DahFb9bLhFqBrJxX14zq
H1zilpmn0jLRLj8acisKDxDiO1jd6zouZKwpQeWI5t7UAmg3Xx41kwSP4kJ84W8jTxS11Ntz5nqR
v4FTsMq+YFz0sEVcTWHSexv1mfF3D5/KRiYzYjf+DZaMjQJ+1DEYSN+vS4qi8aPr+lh8B+HUAmMB
+yBWC/7S0smBq4LWeFZ8nBC5QDv4K0ylgx/+W53/dmojEk4iXFiYFMRzJAAnKon2ydxKNPl0QCio
WxbwU3yITKQORzz30kO6PBuTdChjzuaGpyxjMdtyc32o3Z+9uiMeFzN9Muo2vXtBW4mykYMKS33O
tpmk6QSbRl9kRCjXOPXTxEK11EpElUtkh2RHHuemmSc7O3ruxtug4ygsVdR6oWgif/sn520o5e59
5SiwG+6Z1G3hJ0V4EAC4K1WfvQEYm5G73W9wGRc7NPIkk5RdXbmm7/HyKPtp7x5l8NFkNCEqLJmp
EB3ajEX6CDJVY6mTUbTGvSpT+9+jjYLGOcPdwaQp37m01hOinlq1EdCPmO1lVRbnmcJvpylSSOhz
/4BJarH1ojB0EwrRU0wnuhqoRmVNw8R7VzkRHam1O+Uy4ReRVCjvx1dx8RE2rf/FjQ+UOqodPWLA
kS86V2oU0eIZQr3yVFQAdTtbG4uuRko+qra0ShPypLH4lGQa152sejQIjX1nNItWGivO2Os3i8zt
8btrZ85a+rXY/vWJqZXoo7jPz0YgTcuISA49oVqhMLEXZrrzBlrQo9F4L5+cnxvg/lsLIa/v3OBa
al0yrLQGKmRNXHfKtf5RsS/UeuSpttwv2jbb6Ykojc1FrJeEp6JwNkVe8IVucwJJ6riRKf7e/lEh
AORhmFV+egEb8Ep2R0rNnBA4xeWvnqWImyxX8Z5aFIsQZOkU/W4PW6ntBmmjZMjWpn3yXlFXIljH
QGhDVu5bHepMrLPxZZp8HpgQeJfmgQcaaX9coB4FsjdHiuqDEtRP9J8XWLMaqF8z1QoAlCAazMMw
uf6e3vMcPcRaRXae45APevvPyXNmiNx1nHGjUQFrkZRLc6K4TQDMXYTHOxeGYh+wLB7ItjG6fd2s
J7XC3nmziaG02OZUcaDM+FwNs8AX+2F4hUtSAOOSqDJ6OiqxYaBs81GIFDR+nLpLAGBmMJj5wJuR
/BTzsnJ1DEL63tGh/fm4FOiA34aiwR5HCsTBewM1L8+UUDCd+yqzJ90MzADDvHudrDa4+y+exI+Z
2OGUd4esD5v8tEW74sU7YGPbKST1ZOQDGayBEDOP3yxxsMFBBaNR7m7ihTEozUPU9JoEICgkaQn7
wCp2XDey0byQmacWJZrkvnwQiLXS8JYoAI4qS0ChOJmr8qy4E9bU2LMoCaNfrIHIap3r0rofz5qd
kWTJ83HYXXrpni8xqqNqU7lSPg1lAOXxkI0sOld+biE2Ce/EDaa9heLiDxr/Kancgda9AnEu5DVS
FcphijKpUsX9OInLERqiQQkUb3/PgAFy/EChoieAgX1DAug1hEUZgcE+KAOrgMcOWJGclMOGwhQC
/KPLx50fKWRLyvRhvDRmwwwFWzcafj5XmVlBqTZZFXHAgNX1MHdKXOTVj9JzOSogE/QmQDr91isB
rWScH2O1zZqvR8KBgPj285J7YwbfhdGEsHSd1hBnrs4U2wS9xlFaeJgDqtccZb4SOtobrO25a6vp
MgSwxHLZs5W7ugoj293w8LH9siB4CPlXLZ3ABUwvlY+nKZzRdHchYyOi2z0rXlxBGKJlianZJOfW
3YhvSX1KRb9k8X28TJkmgJ2fUm25g+BVLuvJadn02c3WPEeiI7cSF3vuaEQrdo16tM4Qsw2d/flu
JWGZr6ukmKGkRaOKaJ3FCQ0G5wOWGeU0A9Pejhb/3uhzhSD+n5Pr7AUEsErpd660ooY3HRBXWlXC
9BJJAYhcvbTdnYmof1YDjOF9tlLhsMSyF4wSz0c8ln6LVfp+lNxkJt9kUHGQwsMulL2fSWjMf8b7
suQHuLNVJd3ZOstBNqgGGC7C9DdUy3gR9fYiBXHQbk4wEL/eNN1QBJTnjQECO01zQ5GfVGtm3ndh
GwvyfZ8Rd61by+odEK7y84lYGwwjSz8NOT1RCX+Sp9DjtzAYDJQcXkuCZkVqGBnwhHo7kb2DO0lW
gje2eD7/oOImeQjTyZu/zY23+X3npF7t7IiAuCdt9FMwPfiTM7LoEvra/4r1kA/9tCjkM82adeJG
gR/fcdMq7YiTrbStI0kGYHdnD62dhiBk0Pi922mLFe22vFEe8IDmIVeJ8xyOSSXMNmY4Rahu34v7
fXOo1CZT8AcZu1ABPgIFOWyCNnCLJ4pqubCuhYqsQlNeVmfYiC6vUQjRmwsuHW7RcSa/HSUj1yEE
fRBqv8sT3YlV7ZT0h4zTW7wk6ufHTqIgETLJwadYWC1NFJkanyCWJ5V3ym4CEe7kOkjn/MpFTSRq
b0z11p1nq3U25WaAz2OekNqBa+S1Hwwfcp5Ogsm1K2G+wuCqZ0e1yyaVlUEcamT/P1gT8RJW5SJr
GT1Ak+tZCT+cm1qDLupFadi3S6pOdcET/BCT2C2L8iSzUj0d/HFehHQEfMFWTx0fbc9kXN0slSy1
iNQSsMsyDBJHPdwAvTBjdVdjdMcJnzaVz+lcyWW9qdIsosxNtvtwtbwkqO8mABrYiOWJVJGZ0DEk
ISWHXKBYLysLZjUTbgfr1EtDBchm/vXEy1YqLlzvPvQaZimVn/lux64Nto9lvWMsttjtVXuoFfw2
r3VPD6oO7B8bllcUon5INIqXRXIvP21rkkIgV3kDVW9AZErGkojm/oXjHICZNRBfXVHTn2z/IgL1
HSF5dA05fqrC4OulBubBv4/JtzZ0osme31i2xDWHYwRBjxk5AN+FvoHgWHqUs2/X1LYdq0ctvb5+
NPiIsoeBif4Sa9sVe87Qe2r5ew0GIna7vasDTdKxIOC6npjZKBhlBuP1o4xiyytIegeHSpMnZnbo
JcTwIG/85WqSSoGUWnSQ57/6FKNx3tEJit977ZgUUYPcAIyYa5V1Dfs69g3MMRaj4ZbPZ+PrPA0O
c1WO55UWPoHqLbG67JxbR/P1MVUN549ucAhUSrkBEuKjLOBnaEti+4dm+RM0GUzLHVY/bN/ESBNj
QCLa657n4Nen0Vu6za0fPvbs/PPWUVHP8aRsRzuXbf8VuyBbAbMP5MtcELgS0jdj7VtqKRnJ8NwS
pfanPW9WJg4wCYNmPqt3FeukpTM19vYWbnFI/oVHv4W/s1/P4dQCljAEcqsKMQBBa9LjK7B1koD9
Jcp9G8Lt5a+oIKluWa/kQf5mOgy9iA283lVpEQiqgX8bKGpRA9N7f+qr+LdfiE6n9skutRWzdxJx
GEYZ1/qNJe4dULnA+uhrh41cGrIf/O+if99hyctXk8EgHjJSfeAnkri0LZ3BXUMbpplQ0ihxQTdC
4BVog9qS6tpnhg1O7XjtWBSlOgxtinT91O9DLzL5EjE3Wcg6wQ9dQpFTTtWecV3ERA39KkvzS4KP
1UrXCKPN/CvD8eCjrAQRZvM+mJYc9VK9skw96eGehSELWRsOog1m9oxqMWJxZ4muB4wg1wnq3+v7
q5+JhhOYYmaN9F2kZWKEJr4ML3/amXNBWbemTt9EHyt+n/rb63frEJfCqnya7IJI2olbpJlzI5Dt
cwr7+ZdNUoAx4jAqj3Hf9izld1MbNKyxNKqFOzMYi0yWLtYp0vHSmLlZ0NgXGzroxgVRClTlZZd2
LXGqcNfJTH8mD5zWJmGWlDMoY19bapMxfy1Zg/w4aJnh4OYM+r4FUPX2VgJ2CLh+5vdbEhz7D8+p
KKBovI4mcmNch5sSKsgoJOeprwWrE2yArij0ljZkiaWWWZhcfCP4AlvFldEXQRBQ6H80U/xO6a9A
h2nZJX3EARY6I4A2u3+GV2+cTGSxzgK8+0Pk01knYaJuABy4AkqcAZYr5jAxHdhPgxW6sFS3baUd
3HLq5lHziivTRwkaPaNNGYPCTurl5V2jCQ9jkwT5El6o/VcYdKOIg6Xt6e/98yhXaLra7cXC24St
23SqtsnhhWdrqd1R6mGfu/0mMQHRwCoOY7SHiUfHqutC3YfZdirrW5QBcCRtw15nO4zAOvbokLqV
/1ukovkpE+z/MkOexp75FjRoTsgfGFMR0a7NxtDkPOy3Z3NPoU0R9sIVTMj0zo/smXXFexHKCcrB
nx573Rp16rCrJSFfsBgK8vkOV1Sq4b8WkeqhmMxjLscquDObtP8sWPMtipAiPcNJWwY00oeCXrEJ
4WvxonHZVtEjOVer11TyGosmA2A848bK0JbybcYUpSCA38b1ik65aNBhaQjrWe2k77W8o7eKubi+
haGqLKSK6sd8vuDjiQV44lAjSHNQIvlVFWL9qGWbvlROReW9DUIwx2loMYdb2JcY45wpcoxnzGOd
HM7wnb7MVNREh60wNxPtHOPSXzsB5x8+YnmKPCCzPJRh1KFvgkzO1VUrO5xI8H59WDULvvSzOSYD
MPymXcEtuKvZeLDSX0LFaS1QFkVPtObrQwoVckGmpPF9ioBkGSQb3IUu7GYxTaCmBt4vpdQP81qx
wNXRBgR5hTE4DOMWH6WW2ZEL2gmYZHkzQmRDGKkIaTaNdh2prDxKD2DRwblXCe/FdQhtQQt4+7bi
LYBKE+3s+oAlL13lkqjRG9SSyqSht1XYc4HPHXbrL7aLBvkeZ+VDCAi6y1wbxmTBF+3FN271mYL2
VHd3KHZ68PMw05/kNWV1Fz6iQFtDIuf1WBIdN24Nf5pXDQpfabfpNzJiAd/d7xUuGI5hpK6JV/ok
VrUdOKh2sRT+ZQeS0ZVt3/i+umW+kZ+uh4T6NPUAVNC9LAdaJQ5XUUVQtFZeMwV35SY1BNS9kbGh
DfjS9Z/uqtob8NjAYUbS4FNSxkhSc9z/V+oL77xIi14co0CmBGJSB8LHhrD8ZFH1f+3xs6NRlrtV
md8yFUrV5b1vtXaD/cxhYA7uCDZr30cl4nK2KOdyXxyTK+MEJCWSEWRl6zZIdJ3i5iNH/Aj87lBe
DK/33+XZTspzjGNnOBB71qmY5BJ8sKIJWYbNqsBrVsngJRN7FB0uq+6FrxSPKAsPZ961cRF1OxmI
vXjwn4h6RfYAWsasVXcJHZX02zPB9Wg/VTdk6qfnbO+282TRbCu6X4AgppsymFy2q9ffYB0pF6Kg
by7wThqsYw1p4To+RhIPwHJBfVg/JI4yefPBB8SrFeQ+E1ZOotV3bWVG4fpQfFmrhDGSLsCM+JRK
7qaKDrTEFbgR8hpytQKiw2Dws2Y11ZsbjI5vjZmcrSjdm3VXvtW7d0H102qyoayreOe3M86viRvN
zJcDISEIB1utWUGJRaDT7TkRy9ipSb8Uq+tUd3f64Itj8K1ojA3LvddQ1a13k+UMsxaDXNyheeMj
27+zvig/lt9Wr0uTrrg9POC9w55zLS8HZ71RrJnfVFU8/YjqKDJuHxeeyhPgU3aBG7ImYDsR8606
qpJzZsSCD33PqouBPVej/yF4tPhpxwxLPX7KDZ+kM1TCyB7KPexeQSGtFQCuKC6XMKFTDnEigToB
4AMODX9o66FuSVCOu7J8QKrqpKyRGAy3sTCTE5GLmP1U0B+Ho0UnxqlG/UNOohuzgoovKHy+xdUh
WycPltRyZuo6HuoSL5tPpEEoCgjR9mjdpMJ9WLuYu/F1JokGM/Q3RkY+axQYwDWIARSHAf94/N22
idsQfYhlzRIy0dvfy5ULluSsTYrdl4iQkdyUKncDVgoUuJ1A5u7zRWmdh0UgWkHpw2f4RLxPHVy9
yaJaqlevHVsDovRh3wg40nEooJ4z3M1oNX+ZG04E0OJ42UB8XnrJewFo0tTWfFkHiKk3E+0Dsxbn
dE4qhsxvBb/6xg3/xgtefDfvzydL/8Tsqm4NMmUcntbqEjHRB3w/rqSIx+IaQTJML4WOi1JNZNTX
yuzkr2p2M9WEufb8w20dWsXkyQ3FSuWijxn3cmKpzJ5nZ0YQpTZj33PwFeaxdY84Py3TboWTQsLa
1OkV2BxDa0MzpfM8V+v3TFCyXf0rfdGW7sGig0ccTUjmlXNcTOVymHc4N5fN0VpjuBcZYmJ7euT5
r5pTG3kapxnUFshPv8WW9GHS1IqeXoX7gcE2ujTxOOQy27VA121dByGg5pTwtcbmqVffayIGeGgB
PSupLzDc8++IxV+4hVvBIcfi2v3BGPPd4NmipKolsaNRBZe2eoH8lkHRxsrhI8b7V6vAvTnT137u
Z1AJcqp2OmirhyB+qSYCW3Pm+1jLv07shIyaZL8HwrtgEzeKFplEEjh1UoYwo8vTP0LgqmnAQouf
M1m5Nmq/1gcNS+fHXUQRV5F57pJJIQXcs323qnRFt4km2jNYkLH4OPjvBg89faqj4WAc/OnfU9RO
CTuuPWtYm+Ra1yZ3RAiLmePTZqFD9GA1Q9QcUuZVPnHH8Kh0J2KI8nkzLmwsmNg+FjLl84jkSsam
lvTmwZwXUJTe7D4EWQi9cL6oGZl5IHcY35eVhW5LlujG3+suArPcHb4nBDSTBBgH+Zbco6rD5ozT
tAAYqFW/TTk0TTSXaNqLpbRNhKYGeYrGIg0GN7RNzIrPWrNPQa7jIZPH+0flhLmxYz03tJEV/bT3
byhd6453MXzEE7pXa/ktRyaG0BhBa87dWac4AOkhEc0u6fVD5TBPa7C8mdEZkaFOmRcWFbCQMQ53
o4oVMuAyP83VdO0y/fD+brMfNkNES+M87KYTDUtwxL7Q2rHUpBk0jrEFJ2DAz3Y9tIEBkTco+m8R
iLulIEYoTYZ8Xd6R8IjuxYUfMFWQVwhzZ1+TXYL/oBWIovDwjv6s6rqT7KqPlX3KsDAf6yD7FMFQ
fcdjtnTnx5U+Ixn8tBAdhkVQhhp7BQGHuPsE+02BqZxKnQAjILcR7pRBPMvlIRZeXHYnr4uzPd5w
I/1No4qM/Ur4QMChqEmfK0EGLHK6UI7//Lx2kmevuCNrbdXDIFiFO2UXf6ELDezCyEcb7vHWphyu
dy2iysEgoSe08ybkspF1r77jOFKfPb88J3vXI09ntvI0eU1GLHRNc/Gm5v4yxisLkZaQm/PHE3yS
yMYSsin4AXuRYSqGYey/DeZKXcxEbSgh4O9Ex3hRc0qHUPe2GSrDVVyzjd+VreoisCofYNStg9h9
JbXDKBA3r8bF+fBR6iUpVjgu7XYbbFTkerI7S/PlGAxuKR6+hMHUAzeeOcytL0pPWRoGk5TV5X2z
hPpF8Z2kzwUXSIS5s+dPN7XB9h8B+ZcdJ0TY+IDt5xEaEauEyAIgYHN/7USas7m8GtFWfcgYJzCz
tBlWHgfmCfeEVodxfzahYLbkTOH+EuO/vzF8U9zt6DjtWwZPYQbGr6bSqA00NUvIhFYPWwnug2jL
TpA1NNulkf65LB7TKKqhrsPfksXacdFx0ZFAhVU2+PEhxyLuMgv2oX5wJRNXoLYFPnlJvLUrynxP
o25l0Un7+rIaoMXT9rF751tJ3sNeAg3xCkNbSgmwYmGEr+isAefZoGTWzAecI0exzxSArteAJOq+
g0mss/ehHugEQt5+AKAQMh2NSfMIfgXWEPiCc9J0hYdQnfjZiMdriwBp0njZNg0znWo7KEiTFasV
Qg1XrPVlgxF0lszOsDOttbGbCyX7k0aDwXRBV5NpMyQ6fJsl340cF3VR/wcFHwyyss00JR9fVqc0
hXtdA2ZBgNiw7ky6Gy4ZDLKDbt7M9r5J28J89wiR2lkQ2ilStLKCmOP0nhfqUMtCjbq66AySiR0I
Wm73Frs/Eq4WT2P3kWmb/xuc1qAkHWWBPybCvzqXasFWiBH4bbFyC3ceNuu5QfQ/QfX2zsecErzg
N9XQygvAk3HPbLjA02TE9I+J7Zpcp8xP4Kan/4fYN/U3TEEBiL4ia8fOp9aaWpGLPeYtV787bZX2
KBu6OrX9/zEXw1jjdKHsKknlaot7MUvEl/CT4DKf38AWbYV8a+Q2e+e/krxOfFG4OQ3iFb15ayBp
BBXEcv9WPZDvnPc6egOgWJpEW21K2wlbxbi9k9LCv5JPO7pL0SvWBRBqsWGgeOmgJVJ2IlesVNVa
SzGdCdyyQi3zKUe7T9FS7mk9zgllGNuLErMrifa6wWCSyjBhpC99iTe3zHE5k6oEK4r6d4W/3TYb
hx75gPVW2cPsaEdi4/7lvSYT6Icy9iHVjjYGF9hnUQCOAK1hh3O4i+KGyl5MmrTyREquAcCRcXw/
D+crouz40YcY1oeSgTqFMVrriLqLskeXI3ujbYaY/XwNvZIVWRUj0vELhMtWvq5yoNGULr0GFMpy
w55pclh8Rn72DAzct5DAm5/jHBJp4eQQTuFcMu3NI83EJq1hZgBBMncXGe45SFefRqhDl/I4XbUD
s+TJ5zIbxBNuAkjvAMuxgGBpmuZfVsunfqzvMXC5sdr//MBFbyN5sZlIqZEPPlUoKKJU1Nbkf2tk
XHagxVbILv8j1XMAUOCHOqI0g/yb9gzN0nkUU4jxNUhfpwQ3tVvLUlxbIZsZyR7LqL7ddfYiOniY
ENxwOV+wCkiWNq4Z0QZHq1ZCxvWMEa96cdCeJUUq7JvxMc6KOoXvjxLUzzvbPBZrxkH/mmFbWJxl
tiisfB05iQoZJS8/QIWJt/MTzlZS0me0U+H91x5HoYb9nHAl7TP6aCOdhC3Wqq4wTSvpC5uPBS/j
0EfyAP411bBKGM8yophYU9zK38Y/xg+nScVaAEdXQfwaSq/rg38kayT1IkHOC2Wq1QQjcOXQBLhy
tjXdy45LWKewETfWom7lbAvdsebvSph3R5PzJDCQAEGKaCdX2I2YeGMCaAHgDTdSk+uT+gEVTAvg
Dw9VzoDgGr05bDge3W+Gxpk9abGdwL1NzqK4aZqYDbhBjidSoqkbmkRr7nVtt5Aub/OcRpVbm1Yg
zJlto/OZa2rUpW/nEMDguRsvHEOTn0id+SCiODOUufveMkVy2BRPGij2qmpjWIJOKhQkv+kpQikg
qOAjLkwTPJ5ltEVf0V8bS611SHMI6JoHjW1Vrr1ob1eyLjga7dpDTYN7mcRasOrNsH2vz3Eeslik
swJy6o3H9iDE78zhG1EHCt4tTnbzRZTbtdw0ZlRCnK/VgfZNdtLgGVOWDjB4ANVEXb2geYSkEHZI
hRjiLpX7z7q9B+xce8a0/EtfUBCRTU4kt9D46Ssa853tEk7H+ukzQh0Fjpt3KC9Y7ss4bI+Rb7BD
CGaxJ+QNCA1iIKKlzTU+ePw/Zv7HphOrev4GSTSjpu9xoyJxoMZVg990WrXT8htoP/kigljeO+Nv
S8pCy5aAo28Qw8P6AFiNvv2Py6BtF4bMOAEaVxJS4XzC4i/1etyUzcr/Zsn+3ecD9c6LEuXJXgMW
A0Qs7J2OgNQV4iLvHR1TbdLvh8H9ZhffGmsxgl+H+sGbjiTkJ8DjvpyAmTd8l5oeDJdW8j407Xxf
/Nuxr7VR8I3JfbTIGeNrMViZd+EjFVwqy0BpFV52qVqgLh/RmcPxiRPi3YvhNffVZVVslOBzN4Lt
HTEnca2zEVCzHPcvN8wHpIp8sJUkgW7egowNnYlL/N3ci+Q+9KbZvUj6onQEh4G6+1dyX9qKOau8
PX4NpsnZPuHr5R8W01SuzQXm+L3+A9LAgy2PkudZiJulbXs7Ut+fcVxXtow7XcBDR7lVZCnGdYMB
dg7vY21YaEJ92ToMLG/6wPbHInuKN2N2YMzdI28KH4zerc9IDIRE4zf9rcGq8bKdxSC1eai5vgAc
LISTm/X7iF0zhdKXLFNcJhYyUu0IxbmZoDJUAhIMJ5IRlGRv7S4dYhCuGEj9fCUq2Mga1xoL0egT
AZzGF33fKtdAZEMk5maxN+RwB1F39Ch2kKW+CY0Ub5sQgDXuxGXo4rVeCoth11J3zNUTWW/Bu5w1
607Xw2egxWZZMGwrui9mEKq2CA4zMh1+f1LHZjOze4KHFjDo7tjOT1RpBd+cxjzDLwkCBSvjZS+W
HWy7lbH/1M6UFtkh6CQJMQlULjn3j+6XJ1b5Rq95Ac0oSALnKKhqumr5o6djQgPMiOieT5OCf0Th
NclPVZyaD8RSLpCSISASNRxlj14b1GMYZHj+HwgMSV50a1Eul2SXT28TzC0aT5DJOQXG98/Yi/6K
JUstr6PeiLrYS6OcZQZ10NScreX5z37bygBnzhLiNCl8OuMxOHZCo/IeOT1hgM5fEIM4Wezjju2y
M7ywo617cqD5tD2v8JmRPWXksilaAw0j35fCAndcvEwGQQX+o3fWenS1zTyjsqQS7HhE59oqXyKu
4CTOjfQUfgnQKkPxGZ/TlP0YfGg7VDXlF5AXrgulxOfHFObm+JqVRmcVfOt1lZvOVHoeifyFIa4b
61srI94A9aovBUg7H0AiFAGt3TPlBmo8doNGGnaLu4CBvqlCwnemdzF+M+mKkMx7ZbOU+94erdkb
xBX45UzJFlJPju1psWxopXX1sw4W3o3B3GgS259UZmDbepGysfMrj/O+4gKhwRcCdv4z13LhHLk1
g3B41v7228tkPjtB/s5fPYHw0AMleE9FzAe9SGNYfKvAXImwTBrB9XGMcZwHLBi0fZBmX4xQE2d1
r3OXp9+uumhTxKd9JWcP5fpt7pMuDjAvA9etVboJYQMAj2cpM5iJMlpeOdVkvDMDgc+Fu1VgBZKw
EXVWQDCnMqndUMKf2Kmrw5tT4tyhQ5VwPfc3fQhNo74iE+fwwdeVqhZG+q2Yj/m7S+2Pg733GmBQ
+f8L756KwATiRxTz6mymuSr9VmWFvaEx5nmn0Nr0DixZFB/TrmNBCCejZ8ozcfCxkww2NS2EC8Zf
hWbwIl3PdEfeo87pDn2dp6p2L/UVxyjL97aqFxRfSOGR2YhQneJF3tMGg6ZtS24Qy8mJ7s5iDkjo
Ukjd5VrT8M60o+xFton50VKpGTO91XbLgQRFxJTXlnnexGj8D66vm50sFmjGEx6XcCSSyXg/vZKm
7dZDhEeClZUqNX0m/KJHiP0arUTZe/WMJ8wf09A8/vgWW06LfyIGnry98QcucB3N4vuWQ58k3pUA
LZQG/0dDK9fSZYB9YMeVp4Vd2Zlr67+dURE9AAfOl+xXJAcC711MjjO+ADud1pHWJAY6zxWJ8q22
WLOBtnFoIjIiJbmr9DbdQwPv2aI9MLUOClBz6xePwtjXiqqYoIEjH1SvaR3uHoTcwOfrGtEI33QM
OtwtP9C55qbndVz9iC8IprrC/ksEGrEeEkx5DCS6dyesEb/ZUP0Q/IHOecwQYrpAb77EXtZzQiSB
JLLmoZyKuARPiTvVV/3ro+fOyvnsmirkicxYgj8uRzxawqrNzGwwNhr0xjgkkjXdyZQwko94Cmvn
uT5QJ7Siornc21eRt0NbRi/58C6AF848Dyr8hZ1ck8nnOJtTWcE4mF+gG5WxPQZ+NkV8enlGuazY
uy+azF2l0Wxooq4t4HSY9o16rJan1JMC8Ym7vKh3JrMFne73oQZGXPN29BwhVYuyPTz3FoBfhbE0
En22zvBvLleeaMRkMCZFYWgYfsO34HVKtuHRn4A3GlM7CfKEStGhC6d/Uk3qkhluNMI/C3qV25m0
5usJSnw0WAl4Jp/Pyhcj7RGIY+mgzCw2hW6zZiOG+4YoUs5UsZTneXOTUGkkj/ihn0/IWGI6Fc0s
Ew5YcXAj6mp42pFkGA3i6Sa6wsW5p5qPfojizK6NbZ6z9BgNqFCB9FHowQdS6ewaguc/rbXm2Egm
arHBogbLpPaSZRD2enNkuMbCGAts8odJkyY+ShxdJQDdKLfvCwDaeJYbp18rGvtHkpJCisiEfWHF
+9Bx9J6D5WNiciT411INhgOH9Vi9k6AdHD1RIOE6sIJh3MyRCQJrHryjyofaGVcFRAglz+D4Z8Cf
x2aAuk1ph7dqxXqlI82rc7FXIR4t+2XQ8uBvP/7ONei2IumZGs5QBOzp3MCtJD9V2oM0p/QVHBxL
EBwSXC0wSjnPkIzDNqTNXUU9TPhCkMCARuMdUkzMu4pBw4eranZ+KMMTNe7ak20yuRmEREyxN/8v
AP8isPxsFn1t7nxs6fn2VofzpTH53w1nHIUIFE1oj1tCIFcaE3lDMci+Nj0p8Sn2qg+A4QH/ym9c
W9xDHahzQrcFqP9e6Lwv9MKFtRVyDZzVTn+r8gVaXdlv1kYCQf2pKEm02PZ9HtVX2W2W3E71FAG1
N4fk/AXeDCnndkpAkOuRwx8aWaOiyUoBUFPgjFfQHRQpZ4+TBhz3tnPIJprPCI+p8m+BIBHv+MTc
p/7cWOpsYs937w4B0VYbwJOeJ965o9GPaCXJ6+Vj13eN6eLhdz5QNbLxYR5JkJFSfE3sA5rSkqzI
3lAc9sN9fvJO4mivTTaDX2DR4d70LmzbJ/bA5owPBXLh4XRuksF2puwOivzcMKHoRx9BIrhJgTE8
XE8ViLYqaAl4FMzQMr+fCJGzvzpoiAnzxy/Z/bnIcwa/CxbykDnw2CjXMqBdoB6Bn1Y6/I6q3I2S
d0o8Q6pibcamtsD0570HlmTK6/OuOGx4NG97AiJB+O44pGmPTWWYog3dNlddMZug9nFDIHDZkKAT
iVm33yETcDh7QHL3ezGxBdtzTCvcirwE+QsBCaUEc1o4x2cOF1/gnpAWsA/4LVohOKT0eW/nRiQ6
vzyo/HjRd/hsUKbS6RMU77eLNbFEnYbbLFseQCP8pN1pWJYArED9oVnD1BJvsTlZi0cv9UfieGwr
UwWbVho60Xqi/kimEXwDdaE0vUdsZBvkZj+KV3pL0ROADgPQj6HUNXvZWrJuz717tPd9g2DFyC9Y
uR5S8fLW03os/PkWOveHf0ow4cMc8W5juuuKm68oAZn0y70/6447vfZ41s2c69IffwtEL62UE57V
Mw21d633f28VzGfxyIXTn4bxHQ5iz986KwFgtF8uT5GF6zrvkHv4A5CPRNkcbIdBtF2pX45m27ps
/SquFnqfZ9YKX1RsvxBdVexNAktvVA0yVH9IteAn9ffLHdVk6iFVksvhYY7TRJBmsORwiQgBOMfD
uG13qHx/EQysegUstk/tx3gEmomzNen3PHgHvJ/ygU0CSgAm75zOeOAKfapgm4ATIX8q6n1KmYFg
zjVS5LS4fkXhXA5zpXFxhGWJi91s2kMwK1O1RGB6UeqNOBwX+htlEb4Kgm3ngxtmLJ4hEAKfs9sh
VpgtaUK8HXwq4gSl3JMAH687nmNcf5+Lk4OWPU+C/21lVX1bpColBobcomZTj71IUFIACiaHCFoB
s74vZFOh5wyW4XzbSZXKtZJoP8sFL1QAkp0U4Jp4XuLbospEEL8uyDvSr/HBRPhEcKdxGdvekokR
5dePFa26WbXHDNztgV986d5b+hMNjiKDeb4iJUV0puqLh9hibnVW/8IYC4VHVnpkK2BJBsos74f2
mXCbgJy7Vklsi5Oxbr1Df9BUQAMTDcoEV8G8fskeXajjPTcA3KbnoVmcEFUMIEPv4bx7M/PCm7CM
KWIXGt6PZugQSQRhnn23gz9d1lxLyyUz765h/a35hmM3rG8PKGm0k4LER6CYTj78B3uaT5jduYyl
zAqrYbJHpvajvmYufMKdbKPUlZwb9K+RPlNMFT2BGeou0DRiRVJbkM4syaawvd2yDW5lhoXF3Dd7
Dv8mKPS5Bf8Ft9+rNo4ERvLHuKEPcHAqKtXP5pNWeBA15JrJOixgLdV61RyQI2E64+Opbj4X5IKP
DUFXa+ynyWp/0VgiGwyegcwD6onNn3setW+L2Wot199vDfOp4eg31x0TyMVS+VQBBSU6m2tYcjXG
hSCyK5nP+NCOWvN6TFTHIFIUGaiHm7sKuelkn/cFHGN/fPEF63QM1qiDFjA0JLwvR6GcSnprLtyX
VDXcO4T+MpfATpH4CI+Y4zXWhJcwe/14ChhvBGrxcAOiU+yH/HKauXa0FHpyMf3haaofPo1BEY4i
RHJylIIj7TRAqyCLQRWtrU/KEwmCXxCkj/djTuEcoBN2/a+GwfLoQ+cDMgbiQIRSEUGHOVDCwNMo
9q9ooFjj+jcp6gIMij2bbH97I7nJYi3WWTwH5tBl+W9WDj4wwgmMLFs3iCNUoDMlCfteZNqMRBVf
9DALesAu63JeCpYxM3WsACsLMBi3IGXHn4fM+q53yVFWloFj6K25Dd/L6UEgLql0xRymXlv1kVg3
6cTXRBDiEZAOav1j6kHfynUnVGZtgn9PX//lwKAs0cguXkc6P4SMKkrL3a74Gc8wVb0GbQ34UgI0
xAsMb43NtbnyzSfNQxjC9/4WdpgswFfqybfpP8mOsBK9ia4QVoOHtmx9dIy97fGjKIhJyzlN5SII
CVG9COdEWwEjc49DpIn2429qhGNnLIJd3GbSJpWIorIUekzRCi1enlbcSybr49+aC0SK0c0nkMc4
VhqGG7uE6On/YPPAX+3Q8kiq32VnU2wRWJXczdx6ZeWJaI4hbivBkcUFED7w/3pR14P/s7PlMjz9
NwIDLs/hGYkUho0urZN3PI81oHz1EQC7avAZuaQ0i0DqerJW2k7Vz5Qr20+ISatTOVi33JwNbPME
vgP/3KjZuNOLO26HjAg7CzG//u0I4RjoAkH2iujkDKTigKDsHsEckN4T8G50xTj9dJb547uYWphU
e7UfWpTGtmvsnAmpj3ZwqpM3KhRdq9v28m9Y8KPMpK2h0f2hS0VIumBGXu+k6L+qNVc29EJ/wZ5m
luNWJh1I6vritwEyMCxS2EEmppMDb+meGYFAIufEunxlIUK/at/StoMag462yeQ07zdnS1/wNVS+
NAUSe69yE54k+PL6n1C8qSL1RBMUNSFg5FetTDqcQ5aOycjlTGHtShyxRFYX3V8Kz5CNUikFqWw0
EPNe3c0D9uqLsbZEiT6Gi9nMJuRHDHh/x0kxZCi04WrAmLpcB415SqTnmUNwOYFX7DfRDPEFZSK/
uYp4PsjqcJdoR4C2IuxQ7VaT5WYiNtCGl18babk+bR0tAgCd4Z0OpvkmCPIo2Q/t+c/RS5shj1Yx
rQHUELhjU+zQcbfqXU8n4JY1kZPFZ7sLNgKrihV1K6/PGK5uDcFC19PujW/1N8zaUehTaBkza/Nb
D2N+AyvAdq/VLCcYu4AwMAj2GlKpOeFABX8Nq/q0/jsEf/fFApTjhALikSjx+sGvUzNoSIIKE3ma
zwbXvjuFnIay65Z79T5spnF7YEfUZLR24FCF+sUo88ojcbzD30QhAYuReFDad/AngTlw5fqIYL+9
ZMMrkbq1aT4TjDDrUjxW1Q8QeZ7uifaLevRysh0jooCaSHfHdev52tb1K4QvotZceaZ8KielfMN8
rX6zr7r/elk31qqVTecOfR7w+I/R6opi+O2RztjserpnvX1jYy0YjSs9PAPa8syZsl1kw/yylh4Y
NXoo0pbPgjZCiuxS6hNspz95lrGkytCWUWMUnj23dX46o7j9R+gH78plRaTz347tUy+8Miv0Wxao
TaKgwd0cVvMf7ROXMfnj/CjRT0c4D2+fKQdo2ZEobhShye5Xqo1L0t34HMFsBFboJnNnK439D8xz
/LOAmOMdD11bXFtEd98ywxIoknc6+5LkN08oQRQY5/MBkhG9Hv6dziNYsmwtJlfYK0EjJvChjyAn
aQHgoJTfVPJRl7LeNCMRxzGCqnxp1DqlrBPdKt12FqIrbxNGgxlfmADSMH/D/UQRvOSpkJifXkuO
2D+m52KmPou9WLDSQ634ccL/EAPvjGcKBdhUeKCRnbONIrnNjEC38x1FanaHSF/7l0l9OKNm2keU
zQxTvayyRgf+bJjkvtaKutilbXQfUbbpHEL/y5/T7AF24A7xvYXprQ4NlyZyzZc0rMi4HlYhDM4l
tZpuR/zFW7DWR846c3pXfzDeLuxcfmK0SW5F8CihcMKkg7/Z8QKUopNRAuvKo1tT7do0A6bAF+L4
suFRxx9jzdvfTCSIZx8C5SynXbFN/XZe17CudMf6tO/0f8AIs5Kx+X2vQakTUBIZUzcVSlNyvbe7
Icp0KaOrBHzowwVo3FJobDRg0h0SJ+vwbKcjisJOAaU+2RClHYB6q1ndH/eOvIxyT2dNqQBBqg26
30EVsKXDNW82bHrdLJl4QeRc7+tSZedeiocNIHK+zauRN6SwhUl/AnutmO5inp1pK99Rr+VU1yyG
4eRbfmfz3mxUtz2VaLa6S5A94XTfGQpQXKyvFlXBp+dVvh9ffc6MvQww1ogYJLxW0yAj0v0vv+QT
DNTMhq6Gvgd1kj42XJvo3gH0fcy8Pz/AZZpygnx4GL7RuEfAxl1FLzitrH2jtbK5J0+G8+Y0O5LA
oyudyC+KY8bFrzezfgBs3VNrEgPbABmQ9lIjAGQ3ztkJp7mZR4TUcfthq/mRNhfWuf1eqELLAhtk
+AYAdWz6n4ax9GtaJRstVEeHejJqQ1GeihQS134TYIUFHEiIbJO8CPTldtrCPcz0YTBeCVdJp6PM
tiekof/Q6U0+HNUrgvMEvdMiNR6FCa9r+UJm7qhTqLxelFNnPeDgehxJdlyykWnepOqR3b/JG6gK
5VmXw6P0nYc29VVa/z70fKD2TXX3q+f9PyRgnY+jBT6SrdRC69RR9GkOOcNXR2wU21WJkzpT07OD
sauwEeLa3jGj3OsuNYe2F8w8Zgo8GftPtfHaHu7jpm5VMBRDr7lpOmNpCr+YS2XwN0OYdvEu+t8o
xD+HgUBA02GL1kNJ6jO7NyTFWCXHfgD+DdR5JqNL2iUoXSRW/qDyTtzFmTGY3H74m+L04PDSmkN0
oo1FWStzmE2qjYBBPKCvj884H/qegRt/Epjqs3gTj6gww4jbsA6UQFdGNbwxrnn+k3m/XTOjk5KM
xj2DCyW5uyYVyNrSols91bU+FyvN/utXeecFo9nDZAyXBqxR9HgX+sXUJTRynZTDxngaFy5OUiR4
0CdiLu3QJIdfpWeQLXvIZfuaFuww97KY3jmWl8DMoaitFmCeB4mbNhvFMw7f+j9Ny38kZ3ITFabC
88fDH5osygIgJFzyS18jBNFG7j+zVtBkdpmDxKwkORGPJrzUxbYI82YE3zHKDkV6iJHVX6X5LRk3
kTFNA72XkBvHEJtPlIQyPsD0Z6E/5cJdwfGmuHZbfHXtnENUOeI0ROSHdk3OZhG+aImlwYIugl0n
fFGyU67a2zmCCNL0Edu/9GZHUw/V3A+DUV1tlhAuuUEUh+4E+qCKhBIzMt1MM3guUHqvvrPWNI70
Dq2eusabCtMVEue84rZrXhZcMYPBMpiUzFBoH+tgTrFbMQcEKNsfThVIigwBz9VYMHLiRSNVgeLG
kjANGkEFE1GR2ueO/61O4BNKJ3STr9b/0oPBuPiQINxY41UYXG6oP6IeXHJXPp7Z+8+Km/6naq7A
97wQtwdVd2L5hvzavbSmrN60kK+IH8LgANkRPN2T8mIBdaDo1O/6pRNeLqVrIkxFnyGryNu8SSWq
WZPQNIxH/dzkb52ZhBUczJoqF7vA/l2tQNpTty6t6dcP2AnoxycFwEI4E4isj9Ym4JJqKY3Vl53G
c3Zmp7qIgOyW5JDmER1BbXlIUWAIU1Grxa0b3nHFxSW+HnTHJnxFo5aNUx1EKTZ42fpm4Y5VTibj
lKaduaqB7YxH3X6ol2tFqE3RjxSYNvr+c2j2H3gNORay3jMdOTHsS9ltb0I0EtVzeFtEGGOKeutJ
HPSXcVSdpJoMop5dnj4TyDcZ+LqgwOqgT9HaA1ntvF9v6HlZkQ6f0fvsJTHTgWm96qVNAc0wF+dH
sbxaGbxg+JGrzTOFbVltrNtztAVBdRqCdOri2uUVtZXx0oKwt3OPeP5TUiLqGA7aIr2SkRfzeIYi
+NZDM5+HMYg+asvfxYny9dbfVBFSlPMEQnH7D+EPrFz4O8rtV3/0AkbQnA1mwhoW7NtZotNFWR1Q
BItsTY/AUcPgNWAN+JnsRa4eIr57eAUxJ1plOog1DIu3YlGmvFejNmfNYR4SA+Chb1WxiLU6lAz7
q3hzxaaaYm3iVcLAcPA7uSWzytPyB2JvkpS/rSAuR70ox25mB+BYDf1I9GlK2aQyX1l8DDa42VyW
daGkKZjTgKy1PCjyJdLysCFauTG7EdwZLw71Ni0W8NWNY3R9GgXWD9uOuqkLIXErOJYlZ/tu7iPk
UD2CazOlfU90655EQiTO1H+MIsNNS4FtoAO0WWnXFVk//SHmk15pA07NljVBy0SsmxlVuZFh1Bl2
D9NZMjux6eeWrKLwacz0nEQ7daJo47apuPSqxqsI5gZ9GVMQ28CjHqg9K0zL0Jrb9h6ZaGkyj2BQ
nUqlNrk/tSanVXyvIFMP9kh8ANI7RUuUsEWrt7WokTad7tNSf/wyPsl0vOgg54kqRMyioFsh/Eo0
rytUqzVEIlJXa9eCPBlu37Nhmdhs9MM+zMSaVh3ZqX2D0M5SsIocOiOW2sL+MTGda7tJNUkVpTe2
P7fGCdN6uK9zSl4A4zY8ghaUDvhEiMrjl37rcI4Nb8XS/+yDL8AK4Tx6PpDMWQMQDvPrqOoK7ICL
mVzG8xWvPt4hYKlAg1FB2Dld3NTlcWqKNk9NoKD58jwacDznfXkUsz8t0Ns1vp6o+RSQb9+oDR4s
UBApSd1P68b+3rDdfa7x9I+oWYJB0urg67QsGCuNLI2AcoQ78RmWme+tZ/CwNcptl94QxcASzZJz
Py3IvWC5BxMyMOtByDlHwJ13iHBI0EC6X7MZmItkUe4R4bOSgIssgjHZgm3XTdvoIoQQvgLuutiY
ewFCEOBdPOZq4vqT/TTS//Zka+fXir9QdIsdOxyCwpEdQMn7PxAkXLNmeyw4jgqGd0NYtsnAAtrJ
nmtsrtx9gOZd2BuvvPsGpUmNPOUKYx+OTVMydDwKjMYSbyD1BdVBKsFTfztM4HGnCXYlxPI9QQiE
NfrbEwrtElFhHnk9E9VhF43jg+1QahZXLhX+o7Lb8n7aYBnDe816dshNdc9ttHjbKNrBRBFQhkGx
JqqiS3xtDht7c8wDjGMzrGy+VfkU2dJD+EFCs4292Ry5U5085zvKYWt88Xi5/aUvxZWTe/YUFtwa
sypkkzygw5YS5Yc6KnvSeI5O6OrXaukaaF7GG34TdByFuVz/YnN0P+r15+s3Z5BVAeWoW5poMVK7
m0LZ5aUV6Jd8MNQtlTQTSO11AvIMFQoxoVVadRoCNtLVBj05br+mRCdrwn42nocTps4dWshhQTdS
pG1BEjzAnI3zHXQQK+j0jyJE7J7VmpO2D9M5XlXlI8C+0G5GgYkA8Y6Q582cILCHdXMC/QqEARN3
YqPTx9iHINFST4njndEiG7+ZdjTjdIyW7Aa+cyaR5VhfRHeevAsYK1g12vLEzCRLf/F1waL1bFTt
J8ZkotrL/pSV52W9gX6Qcv6ru2zE0hr3JY/H2M6sEzCV/Z4HYE2AtCmKwD+kB3Rw/TSTUb0Jm78X
s8jG2J6yyNBjltk0/e2hqNd53SQu1Kt0Ls/BFfAX4JKQbiIOe4hpuElFln71rp/ESiqkCz3uZYvC
cGVsiRvxIg1I3FJWAcjmaw1AS6B1sIoLx4j5AX4fFVoLYcIhp02Je8z4ick3XU54iKCkf720788U
3blIdl7Mp7AvnaLNzlZMa0W/tY68TiT9POjc82YlMsNB73s0q0ChS9L7Lpy42zbYHrNC+rHsrDT3
7e6RfdFWuGhEwusTdFHhv7H84KFj1XMykw6ifUzj4DYKaQBg6BaLgdwgjZyCU/vwQfVAYTjWJj4+
TgI0XqwqDDJtG/+zJczjNpq72AUjkpitzjnqAITdJdXl9GiCzP8XVwL2RGKDatQVl+E9Cvg1MBCB
Jz9xZNwNd1YH+j3EQwPXkpA4ujDzu4i+gRGmnFHHzw1XIHrc8/W65kT1/hLmaof8NAnvUWhdHmIM
icHMnwpMpSEsFFn0/Jl2xkakaOv5hH2flraHUKyCWV9mwzOJ+ibspSgKdz2ZFhmlseGAuNdHGQlf
Mo7uMtszzyOGMLBzwqfa+wYbA3hR2/6rklTpcjOjYIAwOlwbTT1su8QYGyzPZ+16Tv28QBx7j2+e
F7WXY7EIlUIf9XmXJc/njMohDp7moTH431ZVi3TFmid5Ax5aS3wIUABBgC184n/b4jFodoeSaAmW
z9nG03Z0DPnvIgaigDMP+ZRnfOJHiNu43lOX2AfQnySlG9oFppMZlCeCqzB79zi7AMsLoBx2V+sL
F8GHqbUtrM7Hjoe+AzkZHIJUQfcp/CY4XJFWgvLUB/eGVF68UH0GZ2l13vWhMJvd9MgUfFft6zoi
X+lCdxG20IIRXQVYp2Nco4U/ofWc7hh8bNCoyYq9tvYPf0/yPWuqeGljXTqyvwjYM7jDO1uea9RF
KXfCU+F3WkFLhJUtazfK++DwP0XKPiL3C1CzCzjnK5n1CQnkiwQORO0E3gjVPp2EhY3tq/kAJTaY
zL/tH7LZRXmZimK6kPPU1bHgE5x0QqWollCLceKmndZ8+zOwzOaOPJXi4dbfAr2qmQ7Ddf1VUKHy
05yMG8jiKx/TmfBTbkcpfkccOgUnsEw4gt0zAPI22o8RzVpuNjvZ1MMCY/FcDiIdGqH0mX/9E/Jv
/Qu3fyvKONcSvwrPJbNvzR1ZZgtNexc6Q8kszbSYtXLCTFJvUgZx4u0uLzvcmrbArWX4FAR3wIpI
GhWjuSzWFXctkVZ4pkmeAWn5vdqyX1OjgxYkegLuRQjgVis6yol/K8e7bLU2YeoDzNj9ALeh07nv
CdWog1dJSulxaEshqqzxLjB4IYJRVVTkGJJykwRabInx14Zfbdk6BTHaNr3//hqb16GA+fSJHmJW
I4FErB6ve5Y+xo6dl2fQPtQlixEWQXkoQN6A9wHwoYrV5kr35OT9/Mnj68Kmfv9LYbQPP3RGWWO4
+Rr/+yzVn3j0HigCzX5gpnnPI9Oh+4no4URZToUAtqHUoFOarpb/m6NMYLXtt5/oClCmpvRbxam7
7SejE+/l3qSm/+S2TNNEtwro8/kudONNNqKnIxCwgkih+CJdqLGHtyJCtliiQfS/mPTwT7pY/DU1
ayiCWG80Pv4eoizAp4b9BlgZbycLbqChqe5kNrCD4GqtDCHAieJH0rx38+lmkvGQFMXMl6z25VD4
LE2Ug+ry9f/q9gCvfXucP29PdD7M3H2p2fRJUJewdZi2VyCfgThz3DgxW8TShVAvWfVbLWlhYycK
8zxbPCZYH64Rye4j7Y3Jj9Tw01VdPU7DmDqwTVtcM1FBBwsd2woDAmct6RQg4Uf6yVcgEA2JSyYx
Fgtyf2fkIDmmWLQbKIN5cqS4inxCH1yS9qXxGCvEb/qYsCx+4jXod+vVjdlYoUKRHOV7q5OgMy+N
/7HwoKhDsKaGyHiouOqzjF3/mMqqRrWKiyhkVZqAdaS8pFJfXZ3k1nIw6nyiOD0AGrJ06DDvS8Sb
q0N5swI/prXm4ChDsa7k7T1ceoGMOM4qoKTfgnGgR+te4dZiEr9TUryyvicEUuVrOwd79VXh8psN
i8fza2irtdd7+aM3hQzphsufGfAr5OfuRA9QVajzz435LZR00PBx/dTjakvDq3/mybCnE+wkhwdU
v386h0pBB59waUYe/mdX0Ia2rMaLS0wzH8U5WrTqoiXmF2gtnoeU2Af+Isf7LgJ0NoKXmrVk0AzL
4kbPoNDM/ZsCnQfqrB1Z0jghdyJu6xRT3Nk4LqCITuP3Ea8c/w5zBRmemZpo6bedQixlezzHEe+l
A4/dEU5grfl8nyxup30ZS1Drm9+hxbCMR+znLvWuPsmh+3cc1650TbDJsw4IBfcAQMvIyeqWBxuO
wLmjdC2Nq5+68A0Hqh7kgLNTdajQ37XbxlPHCFRhP4+L/2wTKe6BTlPnBONwRu0c18pylStJgBgU
T3nMyMg2AMbuBsueMkiupMvWlKsvJAQOIgB8bsoL56tzjqxLo4EN5hiFl57OgOyqI96mxlH1k2B2
2456Oi2vQO4ps/OmEPwIXb5rt/2/4m34WCyUyKwudqb96aTn22IsLcwAtFuFWjaQiXb3eLMp19mn
gwWgSSp2DouzO+D6xks7OY2zHV18mtX0pkoIONm3N70E2Hxi8aRfFplKiVzfASePJ47HPNqZv25P
W4Og1ZvyMcyYp0YCu1/YNoekWwcqTkb3mwk+x4Ljr6VeNPIbhK+A/WORX9ToXQPUjqifjQosKOQ+
lof9K9i+tYK/5AwJYEJ9xGmTnk7taVbHu1P2Vs5rVLFxii/94aLOD5tdW/YY7j7Q82a4oha4eI8U
J6DLAdlu5uJQ4QQrMi1BVtjwqP9R9peBlh92XLhsRtQMbTUrg4gAZWATBKy5rzBJ8lnWeAMEpBQG
4z1v6pJx9WiS+5LcV0NSnbq4rfdpiToTzHf+RLnlSirGBi+UF30kFCU3AiJI3mf6/5z+4PfNWrVS
NhbHhTQYjyRxLjJVG//bHRApwScPoWIkV1cvvPvL26WLdkoP9kwna47e8gK5fqVlc470rj97PPjp
oT0in+4SinpujbusCJXgI5ypjjsmA2cb3i7llesZAnAHzwYcTLoEjVarKWRo+fZstd4A0uxypj2r
EYAwn8AWka/L35f/It+UQJ5+EbBLH6HKPo6aiq+lt0JtF+QsYxWowQXBeFJzGpTVrsrsd/fLz2v+
YTtJfL5H3Mb5kvO4PBFUyDLh5ecix3jC7MFok5F48mGhZQneaVWDC+NUVs+W80DxHINxtRiIp5Vy
0UlvJkABgrSb2dN5A77JjbjuC76vbpYLdKiIMKImkXwr2u8QMTEqSFugRom+djynPGD1vdC2WPX3
baHt/+zEYHCTWbw4uD9RfjT8CS7ELVb9vekbB0ZjHBAXYBuf5gaiJNutUvIlQl+7ndqVfFxTZfha
3AbYi2uYZKQ8V+N1OVljiVCe4UVGoa4d3kqyw4evcgZgp9KtIH6FUR9Igpl8/D3ISeVVXuQd+v2f
oysaCpIFPkPxQs5tOHomgakMJWQ8mGZb+fFdHk3fL7HHkNpjXl8MvbIpGC8bvVchsMn0QGqlTqbO
JRfrA/b9Hu5GOCHnaSlD1XrWRhuyK7JLjW30nDNmnexLsCRfA7r02U4BEjdQeN6ucMnJF+TcDGEF
0ZFzePOhdq2zBtLJrjuzdjQK5Z8tVPKzkdexqRTVdVmZ0yY9P856uv4qsto3fr3wA5L3eFvtl9ER
8UDSaWzmRUzZunesFowpV2RPvWPkuCqmg88QaPqTkTVLhu6LWZ3iGh3YS4YpMW3OMKNf7PmKv0KP
3yUJULOnxBs+r8b8oEUMlfP2MHDyzP2zldO3ebrojYd2YaEYz5hvedGgzbG1pj0A5s0wy1YxlZRn
O4fpIMswUwpkm25+C87sv5WoXYg0b9n3dAhu/Hbj+Ea9pBTDXwB51d/n3Xz00xK4M7+hUQgcOXK1
i965pKNtu+xG+I4Pt1TLsNN4FBjWPB7htpAYEE9uUV0lrdG/px+a8XS84PVp8sCCtL0ifp2Xw2mA
kZA04wNrCY4ALcUyuwrMOsC4MmUAN85Y4h9E4d9JNAXLnEUEASi6cWxIgu8deE7xG/ByhhV+HjnR
iocF5uBQzgK0e5/zPPPE9qsD8bI2I7V10oFIXDB7nXtd+mfNz4UXnx+ixKP1yapC5pGaYgy0056p
Heen5CH1Td76QWyuWc2dRxTI5HccNneadaSEmAQWJwUsbNoezLWGDfSspfMO3WFjljc4xaxYU2yJ
AuoCP1Tlelx3NpfLXQ35dEkTrvn+SU/yh+J6tSnlFLru3Q7TFGGG7lkGV4QaqK9AeVKEhGNORkMr
VXqTUoTT2WbE2LRK2oK3a3ESC9ZtDqF1j9aSpfKMhHOuL7sqFBuQAmubIG2CNiTcQ9YIAO1UdkyV
gSvYQufYLUUvVEWlKjezQP6mOd3yiNs1ccG5KI/4Tzq3OCq/g85iSQZE+bB+GbjFVxSHPoonMcvX
Dq0yD/4Q84irAsvM7Hs870FW02TOHV2yCPlVP/qMDrHGtTjV6J++DKFmPk32TNBvxbCOORGpOKeq
aAosndYFn4px5DLYfJAH12VM5y274Xouc2VFPZ6De0vOh04EczSNrUTghXqMtHRVKCNtmlhRRY/J
cSjns6dw8yPiW73ZJotn+3+4BuuTSEZkUam/CcF08+WicQgJ0V2UuPhOmHVlbUDZC10dSB1E3W5h
/u709ZqcybNPttl+fJguvsBe0QQyNdFLo+SCMjFSD5Uxwz//lOYdm4t5OWBbHP8DwiUIdbI41clO
HtycZW6ZOEhuDDIgv93x7l3192DYFAPPSqh91be0Ub9R8wk6joVtXo4ddQAfISWZrgSAwkHotSBE
SSLSxv7x0Bm7ReC+dEL5L8kHD7+pkH7DJUGzz2uon4ZSAJk2oW+HSlZowEF+yZIH2it3UCgREsCc
8wXKKU1CWpuSspesJKcS5M8qMsI9Qd60mixgX0INmkQYi/lh2+HUtM04EuVF4qHGs5m52Q4WP/xb
RVqrQP+z82UkYZxvOIxQ3nF8ZVJUYHAxCo1TqHoqLwOPqmyQeu1El4IJ2sqelxuFFT9IyzSjPkxj
nZg/s8ZfLMSnk/O/aUwROMSmnW/gwVH40vMXidoQn0FYb/TV9DhmNlW02MZXhGy7hGu6/CM3Uo3I
+Jn9yz9Wm6QIUSvGrVYuKEYlOU7ZjMNy1GHObQ8ZCU9KqyKg40N7HGDKea4jonhzAcexzhOi/MmJ
j2FApr7JTVQ3K4LQwOs7MT9h5bYZHzwA5PYO/cEFlKKZ62a2sYlGuqguLCpoXFZG/OerigwfxSIr
cs+vFXakhRhtH11GXr/tOPS+K82eD2NKpmu1tOSkkRdYjIzTzE+xyLq9/ZjT26cByVTviAGagd0d
F2P4F4idR/T48THuSQhVEtmvw8EGQiJ0qbRxXqPcDzpZbuvjfXuoFavkAQRUn+hHON9Ld5CU4erM
SAbFkgK0T5ds59+AL2U8ZAEc/SgYTHix3z+a5R7527uOHqzChmmLBGFqWxC0dFGueecePwbnLA3b
2aKFiKpyjjhaatgaR8kv3dypngZVoetxq/eRsHE6HVDUa4mI0sqiHQe3fwR928w/PzSw11Azuwh0
dAnROkwpNdQMLMQps8Moo7eVyvaJU4ofzograqT2bjqpTPlMmAAzu3f36ot5G5d2qky8ZPyHZf/S
CalZZ0EdwpmxFAQBSDo5a5a0ZK97HAc6ufzqtIIi6oRv8mSMV9YA722plY+8L5v1RfEfR8rz2EH0
8VfJFcVn4oM94qW7TxdVg0ze1G2D3SNvHc8Q38M5pBHamDH2QAkIcU9CVdAZSI6kBUqGGrIy5S49
PLnyIvxpIBRy9S9HRxSDYJWnyL3GiECbaNCtYwoZ04dwS8e5+JLLw2bIcdbOiPf7l2x9iyMmol/V
4QzYTD9WosjDWzNmDjK1qodF/zX5h9Xn9bIIK/uZ0br5koYeIgV8M8B97nVg1E11gPqkD7eXwy1y
znY+i9zpsLxwdTpnDVQwhTv+JLe1QlWhqR7XthB1xWr1vou0dSizRx8UI0bU+wYh4PTPbdMBwPld
rxftJiqTAq6KiabJCIYZBl8MgrQrCRCHDTegplKzg8+mcjwCCTUjTjB189UOYlA0VDqOfUKipVxz
ciZdfBjDm2snJOChMim03GrI8BBYFPk2dXi/h7ScrGcQzvxkhBgcDdkV+KFnz+CSVNg6T0/yf5cO
6/zzy2hsKRg/bqqVJJ+LoYih9C6pmdgzI9myyqj6sTjO1oULJvehuHUiueqW7CCR9DgmHWbztUPU
fUwm/qDzJJCsCrV+8fmpJ8WKgZv96/NpLClDROKJANT/I1t2K7SYAElZoxl09rmOKn40lv2om3zy
HA+29l5AgH1PvQkbS7wQlRWaHapQznxZLGFoKDcknoWILdplW6Kt8prjcfupB79eDT/QXvhRh3Aw
nqxx7D08v5A/qs0sFoQ9qVtz44Snq/jcHrK4m0pXJf+NZKk3SaF4qvfnnFFGwWMJYjHOVjpFplmN
EYDTK1cSvemXweUJa3bmhM/U5T84FexZPazrifBEdGDPNHgIF9imoeySG+nKJtkla0T4B164Esnh
GUwqGNekrXbS2udr41ZNzZDOEDe2ZegvwZ4RafIGc+4X1ibAhQk/BvQ/DtNY6PMT2SE88CgMqxJy
mrkvifH85+aU6Mf3xJcAvrhyW6cc146NwMlPMApDvAB6YQDxOVUZRKOjnt7pL1s7LR9oZ+l3cEUK
CDTqY+jyf4hAxSex88Hj9jZ8eC930W02Traq2/wMdHmJfXxDxqe9ed8iAVkcL16eTadeN4iyEGfH
7ii6H7epU0Acp5jvyVbu0r9T+bbTW6mmZNoB4XhXZZw7mdeDYbqeR2WO2555zS16eY78uq4gWvnY
cvO463Ka0nwqOM5/KmcYOLwlA9SzXdZWnnqTNTXUhhagS7JsQTFgDFgH67LqeYg+9I/ba8j+uYl9
bA2OvRwy2Jnkyt2BKl+PJcqamL1uc1k/w2+wdpjnthAorjRYNraC09I4ShKj0DpPfjo2RrJeyP9H
G79NdEA/RecSv1prLPhpOaMMndPgE+TQOWTL0C7dwszEaA8XiqAvMaZh7e99j6TAGrC4mfKHxCXd
YjXo2zIyycCx3ag7EMxQM190fCmamQZuN6P16fqNhRR0L/Wm3H+gxiUH1S7yJtsI+8eUXYuK0P9/
z9iGBP9/u1Zhpis1vOJOZKkv5tO+cyvhlv5R8G3aYK0q0UkYuDCV3YvEfOZI/FEpGHY20OsoY8yX
LvkcandGtXWZ4e7qFR/8f1jweViBgA/iaYNa8BAsNujuZ6NlbdBVBUM3C6cAFxnA3vZ3WL/ZhyeN
DLBz1NhPLW5LfDOpIm8SqI6sBxXy/+6zed8eJ1a13SZ+6qbhVWvwNr0y2bsahS2YhyPiVjnDpNo7
qP0UxwdCCdpWZ4pfWf7Z1j7C0ngWg0YQDFwBwzcZAZpmpBk5fP+BBMZIjzeSE6MdYlG+y9VpdX7a
ptWxmMjj3wNlLjrFQ+G/YrN/sQgaQTSmpO/tF2vxIysFAmEuYsGw0FJaPt0eKY05fgO2pOsRjHgp
JAytEw/NJvSyvskjsV4Dnj5XiD8a9OFzPwhK1Gog8tP/nEBuy1myn/6AClSZYyqxM00ThdcVHkP/
714I6v6S5Kb/xNmYrQN4RELYmTg7EoljS1SeF7gn5AlXXIvx+r/Q3bhmXDQjdfdKatztqK3jJ7Lo
9wRmW3GDUBJXXOVNrBiF8h6qYPG7+3YLVuV15X0kDocwvc8pkqqcl3vIoBGweicS6F6JnhA7qETb
yUTxkX4lmiY74/4wUv/hTPgyLB/Daa75XI+cT8kWho+W0su3itC1LZh+bsVmUWPLJ0yTWCSXPr9g
dcaJR9x6qrD5w/t38hNAxJ+T0A2ocR7LzU9PzEBdNNQNci2kfs3VnW94cyKpfHBrxbhPDhp2EUsE
MhpwtA9343FGUcccxTmiaJ0h28AgEXGUhoxYq05RHnnA/Cs8wG2YGfeP7ekJihu7TVR4ZnSSoHHy
K9PVdd9dVb9F87ra29XHPUqOo0VrdmEJEfM/co5E4dVMoynHKeGJ3t10LFu+4/ufhwotuwGsL1of
8hw7Qauc4hz1xDkXKD+3gH/A2IwYMYMJhReulHIXDAA2Lu86pGDlA8SyQuK/THY9TaOFQqqgCwKt
IbauiFo62Vm+FFH4N2BUa5SHmr1F51Mk9rVTejbUAtP4e4BEfTRs8wnDyotbwi2CD+gQ7v04q6YL
It+nDzsz3vBB0EqB8AeeR409ty9dOKt350ELovoImomgoMTLcgbYMiJjaARfiGLS5t2tJPDALgDK
pm5ht9qkT0TNHKIitQk9Ljxpub5G1Ad4F5eHWZiVnbu9GW3eaUS3J+v+uTdCaWRtUFMcUxrqCx/j
uMq8oACdlUgQz8RrTLDtavGaGyR0E/xpmoBA82aqehsBGVOUx3Wp0Oapgi+hgoaJnAZzE+U9Y+pS
/XK5XTWfxx4wZ/JEAu0gDkqo8fn8lodYK3FBkGiLjVgIJ9dDyQDBFLbE659WDo4NIE5pNHiYdxGV
+XpudGcmrcvRGaTxP1XaKxyadZfdyNHQ/0lrDtB2bFrAypIfIxMlshDwFUbnLCv9y9lZwrxcTIsC
GJm1+j0X6xxG0pH+Cxnw/tz3DB/tccxdtS7s8dHjEg/RvQj3+6h4fhAiNWJpnEYZUrhSX263gz2r
kpTeVspzi2UpKUmc90i2bnpNfbYPqy+0wh9Pt9pKueaLfBYnztAL/3Cb/yCfk/N6HaY7Wx73QlrX
Zi5/qlv0FG+yjNw2jTu1azkkZn6jbsdAVqcLmqqzwVFXmbT0URQAxiwgNSGYAOhU1X4qD6mAoFnT
vjqQHEEKSii1Om7rIT5goQ06iBPJK1zxZlzijbodYcDbVlvMfcYfTvEVNmHMUN/NDqr43kDSx+Gs
fJnnW+O75y7s95cazmWX/viHC0u1d2rmRdUc1z9ySODU8a0u8ljIXkEA7djEed4Xe2DVkRkIx7Fb
+eJrP/SdXx0p/iQpRbytOEH8AZXmUvfyOQ+J4u41sXJYVlpl0Zf2RXshzMhuiKSyI7QInyaQiybO
HCdDJiHMnMQxMdYGtfijGEyZ+Laidd9RDeIEB84ULlM1yesJ7LpJS0GVnwOLoO5IpPtg3ASfUazN
boNk07jV8HFxV7phOPT//QpA9XOafQ8CRcCX8vl0NJv22NuPMBXC2lxI7cw/Clf1r0NbkNn0o/5G
/lqajdLp3+CX2Jv2Wr8y0UoreGM8hedbpdaU+L2IG6b7yvHwfm5xbigKN+veWimP5n+kX9xhy05O
VCuwXtMhqUOYQ55uxXfOD823WiVJb+yeLO6mctHryybz/FLX2X5O9grbjDcli7sPUbCgY8HWv6UM
Z5aQR+r9HODzYBHSUoQRxDe0s3YORjK8XEXVjLysqUFxZ21BoFkoponAeRrl+qbLsbN1deJ61Yrd
hGJ2hxlldd62l58hRC9qlIhXSkiRV8YYrcvGCih6gaav/GcGHbTT8PUfxrBIA7QDGVVJ1l9KXULg
QXrpYYchGggjjq1jAHXREHRIDYhnBDwkjiKTBceEb8JEYMPzBfF4bKcVxqHAyvelHkqqWvdlXZHK
4OiI46CeN/mcsUeIfpmWTpKkHlcf7eX9GHNCuCnmSMqgvgE5iGmBb8AxnkG76ZSTg1p0H34Pr/X+
xMq35yHUNCAkrIf1/m7YaudFnf4nlXAZ01t2eEFRzvaWH4J17CzWiixDXIEZsbGEiFSOquqiaatQ
lmDGWp+0mFp6aHDxD+4ai4Y/fWXzjHNY3d0uL7yFfgcJlV8l0U7QUO2NnleurWx7bufXxnVyn5jb
sTy1YvD95w8O6ITbKOtTohzvUDp52lbK3RNoqStdPdIpuvvg9LfQPP0rRIzNsHOsIgzxZ/qLPHFK
dJ8r/QAuO7cYClNEfY4FOWtjptqQd77qLXK5JxIyNPhlHKJOSKkEySSJ3arXdgMJnX3PCYFI/c+9
/M2lKummAsncABKFipOIiOKJUk7s3s9RnOhcbdaRZDLr1sZUXsbOgEG6EK4pAYfHCVrHfMhOtBHS
gwUJWwMTjkt5ohx6I6dWAYBgBhh25txUXc/OXa/whGYSXYiems4R6DLYVRkN3pQ89PgW8etjqJkf
gv9ACalqPkvVJGQxsKbwPSXnZLT6PdGEGqtDujE58e5ekUm2htVK4PzVEYedM7wbYuToz8RZecsh
TMnv+2GyeauApqAoXOi2BtABDWm++XNIRnTNtJT22ZzSE8fnkFYkvPt3usCfb1Ub58IXj9a8Szz8
dyfJMjTkluVFeTSGN5f5CBv1XmGuu4Nmzc6/7LT1Cn9MrtJLgTYf78ZmOJuP7MNjdm5wtWmPZkQg
lDZ4yu2+foE7EngS2ueM3jJkcpsvUd+VwG1fTapkOumrAWnLaphO0NlyyPumJHUssgkRajwe2tIP
pAJDzIK/i17JSpF/Rpj3b2xsdmpvEROC6JjiqvUTAX5N0KmOCHPKs83lsIxqd9i7k1atfFhTU9LK
c4tbB7cTmmxCxQO6euF8Ecw3kbC7WU0y977hx9K5yFisJWFAFsssGShkleK1EUtJUZNpoIaelHeu
PCtS0uzxKXrMwQ2rLT3DA2H1VHzRkMZ6ou9S2mYIzJUiOxc38/+tHPFVzSqKZ8jB3eSEjJjIR0Yt
YBmZ5AksbYsxzwIZ3a5Xhu2ErimRYIHl8CUlWz7Q08s5c5/wyGHEqCaiApfsFr4B29Qe4OEWe9Fq
IwELkasDdTrM1B04mL5BOGz00SJ6fNR8tZMVwMrj+K65dPzdDufC2GSfL23hs9iKHIe36OBj6NOx
jjml9mRXl3V/qPFKED3SpxZHLqytsz2B4yt3BGcPBuhc9ZG0blC1Nh/SpsrgSgS8nAuYX7NP/0+N
BKYf3biw+b7c8RYeoz4tO/qRwzNiWm1HHtkPVQt5Pc3GQlxXfxEJJhThmpy7XyBNJnXV1Ahb4qpc
S7h3O51yQb1qXoMAY4uGBg04zUJvJBViXvrBuipK2ws+XAIHz48AIeKrOTedfrV7GP3mlhMldc1G
+otw5HWfmUM/haKPoj9aomZk8MRTDFkWPzq+WhsiIlQwlKD0Wq04AP1CxV9t9fSO48go+rEvPu5/
DI8toYv+ZFMeaZHm5flaKlswooZ1tbHbbSJasNiXwl9vYYcHe4NZMYmAwuULtGNsXvsvE6xlfxeZ
BsaignfnHLL4F57B2GULBARWcpbL6QOgPh2XzYcW2BLCvN+d9weWJvqbIOlPgGFlB+m1miMgbNeX
ZB5/6EV9sZWbu5lOJMYQS33aRg5i9DNANyewRflV1thRFsGKvM6iK+QOdU/us29bYRsuf+r0+Y5E
3/KBbxrm8nAJ+mvQTfs7WyyAPeqcx0oWoyo9etlItkSXcYNeDw4c8qx7SVTKJUJlpFoBGKt88fkR
OpYHFuFaM+EIQsXQurscK7VmfTcn+BJx/JxENDntBrfUcFShoAEmrNphBkSj3W9nBOq1xUXCPJ72
m1XskCnKRmbrXRHX8v0GqFYRPi7YI5qUzKKBj7YbbXV0yGOWek/bkAuC5M6BxsBycudfXb8ghyyb
BZ3wO73KseFl3Rz7A2OaREZ8mESBzlbYJ6SmrPwdIbpvDsShio40db8TSQRMXPBAzogz98U2Ws9T
HhZlrfIG3g23/OpDOA9fuLfAMyWVO5voz9Jxi2v1jjdYfp5VDQs4wH/eRAOqt44Qr+N/8O61onZN
D3BKXaTD7v2YybEqOL1jksjfyPhPOMEph7Zqus7NWhPfqyBzB5SvM5J9qeq2oLgpbCVG4MavPRQh
3TFA9ENIIcLPLg1Y9hZLExmdGxG+JHw648iWl5FO04kB+bjkoEAV3NhaymUUF7cKR4DCWccw+41F
DOYdPphXwSy15Yxzd3YWmpksx9mNwFenlsEtemWzH9AP88Qw8J7OmslrxFoMVoa6upJk0tdA7C2C
942f8D2Or4vT4ih1wjCaoWAnKp2eJvR+rYYDnBtSoCJcnhvqam5daedLXT0IJnMl48MD0NShZSHR
nY6oagA9rM+sPFUl6KeQ1PrvodQimvIn0k1Bb4XUqOV/RwGEbCxOCD55d98yr5xdqGKgFI1ZzgnF
Vq14mkryoEgiGKBYRIwe+jrtNlV2ZR2AM+TLSSOwcVTlYXIQwC8UUpPivNc4pv9pEDEHIW50eHR+
pBn1578H6SDY2vp8rZV/GUVrwCtXjzC2A8s01tEm1MEe7EVDg7cjU1BOdeSpfq1x4S6+c394hDpS
YAXqdzY25A4Adr1Q7/IwO7BR58JdR2cGW91Tzh/ylVSAhSAl0dGK/fNUBIpQkzkq7lSe1p5KudOL
ko18VZJsB8rzAJOhaf7zOGaycfkgPMaD1586nuPVqjR6a9tOksMMm0S9pffmKG/KqiSlWvu28Yc2
nNUOjgQUObsFzKTy4iMBeXCuzxe3kozm3RjIcbInsnzrYCvJ4UzRRpvACMrwPGLUzOYhfYXxTeNn
qkCCtnGr1QKAfoh6lNvbIwSUeZiN18fcaSE1wGiANSSm+1P7ukkYmlg2VmjJUFg0wMIZSMLrCkLd
rVZFKkke/N2YBhuU99JhjdUq7TWEbg5d8xkMoB3EH0x6TMjQO9egueP9gLHkJ0NP42szyqHx/PQN
hMOL68G7fxigmW3ZtuS4/3OMH7SvyroUjIE0BMifnOxk5kXXCD2EfNGzAAXNFu6Yft2nPAt96ohd
A3vW/wr8egBEcLYHNOVbqI57auP0x+NKp3WKkdg37AQfo8DouXmySdSP99vwWQUswfik542nPpuE
8LFEAy/iGy96ZrrXF5+CHh5jqb29w9UdUhUux+ZCjQGgFbaJmEPdVDdvvaOhUoI03kncVT0KSVN+
St+PX/CKduAZaNNaMcZwe7fonAtLJA+Rrr3e0QyTfO52HDOBPn5MLtM5lYVsYM2Jgq7pmuSLatSf
NL4jCVCqeDQZ8Dc4vHOqxwncwL+mizYqiT1UR17uQP96XelwCb1Rf7raAGE+rfVoi8w9veGgrc+3
0w2MRGNUaJTJ2L854IZVTvoojh5x86ipnIson7orCMaKc4XPDewU8DDt9goSMGjflkVzRJZa9rpn
Bwyf2p3cejhswlBqWrgIz7APKkbsODi8IDKiIe9Ca93VCfrZ+Un+xrfpIvGj0SgfZJl/xfLusVXD
YenCM2Jwmkfz7jEc0kBgH1xoMvVswBvKAsozaDVFVO/aeMAHscvqM4QvyR9j/KuoJhHDBHAR7PAI
73fYJ1hoPTP37fPC7iEr6saaL0QDT9Xam3r7uMh/o8RAkVdNk46lKUnaj3me7rsiaaMBCv6jzOdG
aReXbCK8LziNF5v9yc3Yhr4LgxYIyWMDlJ1kjvzGldcPYa/YmeBAW4Q9ZQRiJOZHy7KkaTusqPul
EMwvKNeGOxx3ITmwszxbdF1LT0tJ4cX/myHGJ5q8QHiBWGanCMu/Fd/8pLdFqFAQTSJ3LfjUKCg/
TiFdMdw+s1BWz4NnOB8bwH58qbB3PYzgfS30dFd9Xf6X8YfpS3qd5N36Xq+Cy8EzhXukNyGHBhlZ
0X2X7LCJQHPuy68gkadbQR39ydasKPFdFVBiFda8YFh6swi+mGMyfi02Bc9IFAPa6BVjbq+2Fk5x
TvNZP0pjh3nRa7yKrWJhsx8KeP7ZaG/jiHM0kFK2tTykpUtgbgw6GHeUzB0354Ka2W/Izf0Zegyb
QMbb0jqGPaXvo3ojtfukrLXsCX90t2L5dGMp7xV8lRcxkxXwoG4l1HLjogB7+mFE5/326xEN7gc1
kzCHW+pCw3Gd2D1vRUI3oh/80eoG/qkOF0fxLKlSNZEFFuWsdY5iSQj2jnav81EyI6zC4alIRnZc
gtirdim2NrwXaFJvqi0Kw1mfO1X5zeggnwmF2Tl7awtNd6nCHJrAH833/YXC6EmsU30lKtfFsVtV
7VGeNM3zMLviudYuUlb24BQyWK45+62Ee1FupBePIU+TGAI16mcUvFMU2ArOZ/QJTlTbqhy1toc0
GhUyWOCRH/Ez7QAz3HAe+W+Qf/O8b2C+bGO2G1UzMibphAY/5AQKvmR1opVrgcV+z7RSOWCiNsOz
kbom0mdMXEwVHo9NaOL2cB84MaHV/toR58ys9CkDyVA3vexyYdxHgXOYBZRtUGZtpfLa6VPtYL2k
SlVOMl4rKMCxOXOij9NYb7ufe0S7j3EB+tOBqkxqDfLqVRR1pvQUxZaDUBYy7rlRU5W01NtnuMf6
sBOwYP8zffwfweNJ5hNjc2rn76FDacVB2O7NoEgMMjMpjpKqzsEOFKgmpG0f+kF5bihYT1EvlrF+
19WTit+5SRWyqXpKeHzgFK/cWSaZRs9tpDZ51hsHs7jd1jFhaKlWx2KxW3+TzCPm24B8S2Qhbtt2
Ru+ipbuWZ7BoNwlwRYQDTaMoIMbhH++6gVDLAWYduMMHldv4hJiQEfA2al4wzZkb08ixvc5UwTm8
/WRBBLRccmiL8kq5pVXLZbGOma6eSLLOrgrPS012g+WcoovvtlEmd5rnNWiqMURTKmDe/HE4sPWR
5eEddccSy2j9uYR7DWbirFele8RS3aQNfkUxXNS5ouO6NBIXjjXPX9iyXG/zc30xM+5A/2Dm/IK0
Tll6pN22ZM8brfI7vhK397iZsQRcgnOAnfVfcDPYk0HabX+laOc+zbebvN77kylWk7Ym2Fzzby1e
vXcJbcrr7TM+r2Kh6jMb9Q2IXo0OijFzBtRX+Ht+Q0Uvxaz3DbHtxrGdh/eZnKJ9CdV+VENBZddR
kWjpXNkkwF+GcWmUl9VznqmK/iU8xGgCBKMTG7EKoXAlmadTDjSYXq6z45nTNjBGqi8GC052x9Ub
CgabmqzG8tu+WWVyq0m06TMeF4kyOkuuXMvmm0TGmVnEh/lBRbON3ldWjmBB33bKDQhkrawb/4e2
JzyDrvLmsHnv8qXZXVywJkm5NCVnXY+VEzTGHIcvIKlYlW7QiURLBQCsk9WQVhpaxtq4thvnOS20
zg/RdsSvNM1mNBIBuVb9uuCXfKU6N3FWc3V1wcQE4D75W8fUPk3fUI9bJyzxyKvRtYBy3x/tQa7g
hATwZpmZ9LKGN+ljh+wjKOLt1kDd1zDhc5uc3QcaBzJzabz8DQUQ0iSaXdu88MD0IVZ2vcU6YjnO
91vGtX6N4KQF6YYw8kKDuc69NhPCBeIVfxNNiYgwyG2X3S1J9HuUASUDR9L62ZBPOkwk0ACCzDT9
YvlN/y53pZvscBRmkuRHIpQ6aqoYcmGdhKN7AFqAX0fXR/9FWbgVEgeSLxXWz6Pqrgi97k3Uvo92
/uVu1qxCzXLxNfR9gBShhzCWkDa+V5TNGkj64kF4gEhGD1nRShozNDGTNROl+M2IFJnDIawZe1em
JVtpRqoFyzsTp1Bzm6CuAh9k342xBlcTv+vZ2TSgijDvy0RXMY+y0BMUxD7S6hSFx7kusZqUCOhq
vw1kwi3zO8odWWN1gVDk6mHYCan2+5YUTj4TPxJ3lX8VDXRyB/fDt9MugnMVvGqm9ztHuY6cC9Mg
ePkCvXDMButQvXFwGxgq5bJtFXDoCM/C5t4tkGibwu0V4D1KCEBqx5sbfuUgV9kGQLh44sUYfvi6
eVnrhSl1PSztbiUlO7tlBXXY9ePVb5RM3ugKNlZZaLQ8bmvIrPhnCBebt4xw1oRePL49YORTeo6A
mf7WEeqxiCbdMlW7zjYgT/mk66+E4yNUsUXO3GD5ZWJBPlh2Mon4tgC/Njy9j1n847N9r1RFC7Kw
CfRhLf8T6cCgNFDqt4NnvgUErnw0+wAkN+5JP541RG9QFOyO7HJtl4Ex164qElBduyj7vbHKkMDt
jHVavjx6Xdq7AY11ERQ1hE8GgXDtI/6CVJEI+ZQV1hRzYCSHKQ7j20+wYOoGCjvSz4hEMBv8qsDv
KE24xI5cdI6Aa2khe7ZpMPX9zJZTUiAygxbZRSOFA4uiEctv18m4op9u8YZyCTTiWlRqEku+DCSA
Nelyznwrpuwyddf6p+P+EbAacM9J1R+1wwKb8r0KuU0e72MMaXI+pkQ5bQA9C7x04LIqTtaQ++ug
BdMw4YrIy4wt8qlCTuJk1HGwcCeQgHedqfjyP+jHrXbCt2GzYoyPUsrq0LR+E8MQdYA7aLCY/weI
ILDQYSkHlX++FbgqEdjKccDn3iQ/SjRXuV8Ce3yfgT7LDT3Vz5kIJaO5pKwy8ILXgcxC0piz/e8y
7TRAai8F1Z/Xk7JOcC98POASU+bvbx9da0mfNj+dcj5JvszjJ+dHevYunQVrvQxEdU+zx2v+vhv+
YwizruO0ZERbIykIBIRTU+bI5GdyytXD5XoZxnnCWT0wWoq3W/TDsHt0Es34LYFKzcEwY9IuTVF7
Mn9OgDb1cf7MD2zCtKkMVgNYmVkSffm+hsoZz3IegCX/MBsRgFUdjrJb411WsOnWVd/J869hr3E4
xVRkfUyzx+dSfnoJmMDyOayMR9+zaYY+ucyGCMVTjXrJvpRHe3JcJZSnKCLa/ly/igowhVyNaOgl
0yolE9I2GQ031HCT6F+e6Mw6oLXDQ1fQYiKhNOyfrHj3oFOUQbXiJ2J2CVrxw91JawPQwvdRevBk
04rygd7j63afJf8dNlYCM9TdgiyrEiAIj+II0IiXkQThZEPe9ZXdnB2x4nVNDs/E7cjsKmRcfrIx
/EtkLN64dT9vqrKA2sq6F2SaLJYpT0BXdi/8GWicJk6fw1T6L2IAHgQ3+MA/jThCtasodAilCwh1
5/Fw2kQKppy6ZAlCrSeLTIVqOecF5mDIe+paTMg66vOoYhp1DpkPdjuJwJJUvDLf9dxlX/PigphP
Ax3131+1OHPHu1yNZNMcN6gn7ZNOQV9r42ghdIJb4QeYqnf2NLMGnkqHYlkGofaK7uQQF0Efbqfy
qj1glAfxJGHYNfW9USQwhu++i2+b0koFzYTz+s4cmgyM3EzDIsUt6N8i3So0X7RMnPHw6nZdfxmW
sysrm4+TFAe6dsp0QmbvtPZ2u56LR2kicl16DiEF/MV9dn8wC+IhRvNPmBqiTBnMy9u02L2ESW65
D5iPB+6FoHtfUhZvuw1P7cwe0C62nlK+pnQvlJM8Ba0J6iDflPQkdcZfa3Q1CcV6gQg5SgSzf4P8
HWF4vWbemg1Zrk9P3ilmUiLBDZCExBXPTL4/LyUQO949YJ96tA321cX9OCHcTu577R2yD8OnuW25
VsyX04XVftFLaJ/opPIhXo8Y7esC2Pj/1bA6xScP+Gk7Me84QHNQCJbgOJkzzp8ATFPO/KNWp6RE
YtNZKD+Ac0SyJhSAQ0M5jCkp50Pw1sr5isXAueocVTZdoVu74kEP1OpWBR4LLzhvkUoMNpliMYXO
SZItRC036je3EC+jmAtwoC2hZZEf2ivUfVjUKZkTFYew53ab7asJHq10Fc9tCphfbF5POzgGQmz8
5DGl9ShNNNAx9q6rNZzU/Wlh1MtOM2GGkf3R8TsqiXVMeyQl2XyjChpqv4I0PZP6xTfI5vwz7X2x
1lVYhjDHZJhvKagzV5P4vUjU3ac9ivoofagWeCKqicXyIcvgi/pca+xLayvnkhYEl1hbjtaZvCqT
IuLUXiGrYI5aDBEqJ3c1vFXEyUdo0HU7F+2WMgnqtCWJTt8NUDtsq+IouPDPM1tg7zMuqAIEPL9o
IxX9+d8nfM7EVhr3m8S7fqBc5Lojggh1dgR5OAqO+6a76s7pwv6ij505neeZcCfsb9hQi6mmz8gh
/KI4KKO2+qhYwKhrg4S+dUu69WWGWPz/7Jr34AzJd530f1G0EGR4vWuVq2ZWaH0o4eTCBc8lSDnP
uzB4GRkreO+TNTy0gdGniEqjXSY3jVHiZioHnxiTC+cEplLtpF2x2lG8R2YbqhDroYSmVutt6q5z
3M6LLYkd1Wq9FrRVG57zFUUrRWwf0MPr8t54AUyiPoP2OWzbFHE+8U5uV+IH1knvVmd3uCfzK7sx
V23IF9qxP9VsKWXk3X3N9xkiF/OeO6vkOqxt5EpBjKywz/0QvAoLe0lDJtjlw9/0KmDD2rzVEc5K
o/E6bDljAaOPCalnyrzvjWcG6PnRmUf42/sEsGp7UfBDIiBLaVKTrNkcveVcLCWMwoh7ncxMbEF7
DfkMohHI9hHQlIVTBKtEGgdVrwwAmDvL7rxepKeavVehWmDpJawPZ5ZQ/TL6JnEvHTBXLiu+4C0c
7njiZwWW8zLU3SX3KmW8/st2qlRPG5Ou6eoMYsUd5hTDyA7yXfGUVMlzl35FSYhbLQ+BnpJ/gn+u
KwyttgmBb+FjHPZRtMljCfDTrhFVLasGmAB58lqWKqJUYiJX+BOt545VRx5k9zNJ95mmWWZbz8LB
pRpgBDBZWFXcR+cBClSL9+LE9GSLop8NBqPwG79N90PT4OPRu/m9Yc1VtY+JwLIoaDqmxJqC14GM
OLurS6DjrufC6GnWeKS1Q7W9wNt0vhvmrUhzmMCfoKoJzCB6LDMG/34Jdj5i4wRbfi9qtrX09jJ8
TiFXyf0o81luUcX8r6wyG3XuWr/AQcTLAPxiLO64h4X80fGtnImFXI/bFcWK7GOON2TQ8VsGOOq+
46lfF84qL065nUeKBu8WZr4xFYu40mG9e7dLFesOv4RhwRmCUrfzvfMSf1t4FKOMzcRxaj8PJMVb
67AnjXZHGTCP1ejh2BJpDk8+qSFCuz7SXft1A3vSOCNIx+z1dd4v2kOrCRdoVvFpHx8MSKpM7va2
VJURGl995ufcBFEldzD5C6rToNhOfKjFjV18IW5D80SwN4XvXxFGk0yffagF+yoprbWLvfGS7jYl
cwsBL2RLMvvOGjF2rHy2iXZf4aZEbJG76gzwahtf4o89b+0ypsz6zdSIG3Y79cmKe1PKMkrcjeTi
bCsRGgOirRhddTLY1qSyal2VoEOOg4uC5ZHDYWk5o2bzN05RVcmBrfWpfAaOqUK/hjgpCrgushMX
Gu163bszv0ncSAvcgGiFoXKGZzL1/7yYcK7C98iARXFBWJeVOdOJLBcbGNgHS0akx+hOWzmDTl8e
AGhRdRJq/P8q99+J5E9Jjer3qyUUUmKuQrX3R8yJM3LXiy031q9WANSzITO+s0HOnPVUxzeKGArG
TccLy8sEg4uK+YW2OGBXRHepcOdiQwxv7vlBUNEolcttHDLu2PW6EG7yun4pc2Aal5XtzD/ioOMn
fIJIiwBWJ/VsIWd233dMx/HkFIODfldv/qWQm3goxW/jYZYMLgBxsoapNo4NaMVoOKTRuMk9Gsa+
A+zi+6vzqtNsCCNmiIs46qxf8dBJ47GgDWpSblT7YFwpm8Egofz2JD29ZFrJfT27Qg4PzkM2ctyd
YsTSxrHzxHtWbELTGKblDq+61mAQlZrycsiynzg70Q5Iphew2C7mlJHq/0zHE9ayHY0kGpgwFuUz
6q+G/8z8JApHSh3HaymzBCsA3+eX1Jqo4zvJkl7OC3vMOdk5EXXw0ideC5D3wMATehfrRjkLGd6k
/O/xiRgH0+RZ85QIsUwkn8xJ/26gH7AIgN8NBguntGM5P1CE1TUTS4+kvhHMbAmUTHsnmaI7nkJ/
rwi7CJqZVPmLeAWWHfXn27vPztfjzBIWNsKZ1KMahbSoJpCHd8CsvJdoq51r6e7wLnHx3/Laz5Sm
hZYfjAqfk5jytJX6b93qFE+0HftTnuqxSxwRK0Z/5mUd/aK9Z2iNtgR7gm2NoLOEBZcpdmVTuZhA
6RXcFlAcJtq0KG+YW7VfS2VCmN1c0O8ZdQDtwGmcN/OGqBMFgHtldXG5O2bTEzpHVBQQVDTFjovb
dufD+Y/8Z+vsAh5AZ8kF4NJRnY7Hr71JFiad39RSfK3ua5fgDkK70B04JjPgRkL0+6pC0rkW3817
nUvTt52RCU9JALZ025WrBbyLgbQHd2svk+dS/Ce+nVJNAGXXXwEBYxXPK3/jiCvg5gSvAr7oN1ka
OPw4hDjl3mc3ueFqc3rzQOHr10qwSBo20FUpGtLgjHHzsJQOFMihtrdvjh33j0EUVh5JaS/Tq9t5
ZuTy27Vfzt32BWWDKZJxny76nQhUFyP4D2VH7RiYrOFZwpsXsBwW8S3G1GfEVTngJepa+TAFmn5a
l7o1bHKnZVdiOFUZRKPG/x55BuVfLUQEFbjcxkspOEMAyh0zSPhOVPDurVm4yowa0r6IvZJX4+yR
5Jyj7hWTuB44YpQ9x2hrwtIo501NsPptc7CEJIri15+1b9BXpP83ChAQC4vMJ280pCSoYkyuPWjV
V/fraVdiZ0jr3RAs/hlB+XMldl2TYgpJMwyOdoLafaipcVmOzvYA/wJf2gKFsNz0n1NC+3Cr72FV
noDz+p8E2oOoYflArHo7FwOAXqmxgWgHRJFxKtn0qjUyUnd1xubM3jkMeRN3Pd8jDrut8Ht1IBN9
W0m7t7a2yATFEea7plgrVh09AOLK6sFfpmnrMVgFL+iF8ubwUT+KBL53o2nbXdbAEK3cMxO0Na3e
9V+06ZnNSiSsbmqoHjItbM+DzIcPczsVu8T7+bGgDeCoiEGb2RzcdV8cswrj8AwSnqUpAizP69px
JQA3+KMrQ+rlMQrxoL8RSCMEEoUWjajuJNKixC+k3uR3i3IkXmG9rOLyDbvgVvfKRrmDduG3aX3R
x8Q27ah20PM5nAoO7KZqIt++LHQgrynwodakCcAcSYApCU8XmxpR0lWM+xN6JmGDSLE0LGoydmZP
wt4U1Oa3LS9vGYn1yUGVNhc7bc4wD1q1cvf8j7dtRZcz5v3Ixa7DIHpgHSRP8cQAc1NB0oUUSroc
So3gu6tOgDvwvsVv8JCHZNqG+mfmhjNQ5vwa68fP1Ndopska73+UhKcr0/Zi6qe8lzI0TD3DFHik
qtrBt2CyipQcdeyGc2qxCQzMl2FZTMxk3iLI4DgLdpyrX76RylJRpn/8gRQzOjiTKBck54aB39CN
B6lJdhlKtH2+jfOGR8MF60N19H01D8rkKZ47eezE/4ljlADMBuuAvx9Aw15/yYOm3iUpBErfZEOL
F1SLDLqukQmki26H4gH1c9MIrUUeCVlgTEq8KOsN+Ya8mCR79ybdy4ZiIbNS3IjyHc7zwLPkg1rE
mgGoClBpYQmEkAd4Vui2juZUXM2A4yb6y05j6xyhij0uDtA6dG9TCah5W0HDPD76iChCBk+mFPxR
AjxRhTgkGmNlyJKBUpCeZrw2N4feuf5zYyKyVm8zCJZr/dQrxeA6e823m6EHIEJVPhr4zinyA1e5
Hunjogs7T4B+7HKj8ukq5PfPJroqUr0W1WCz8mvLOSWAxHxyQFbUEwRO8A6CFR9njCSQ31Ifo+l3
b+03LZ1eo/IADRRAwNILKrPg2R2it221Hqi1xdXVqRoAAZ//JfcqHQ6CCr2IthnPHhPoM/8vQ4NL
pkeC7OSIqJKMZh1t0K2PbZacvDQuP6oTuLZINRT13L0JxgKfg7n7Kb9DZzMhk7n0R6dwjoL9BfqS
12KfGE1+5pp1TEj5256VxjZbs7g/m5oCWMrDkwyiMsFtzPplrbYlXu+xNSK2kosCUrmMtNMcTCRu
YLQn2q8vFlX5HUTutbpEZE+sAGETunFSCLsuUgaK1UCDhLYe2avMls2rxt7N7fhh4r37JxFwmqZH
mn6umtV0dmM0AW5Kzb7qvOQNoe8OHwYju9o4siKGk0Fl9xDx8woON3Y4O3Qp7TrwSw/lVf+MYO7v
62aWMPw4QcSfWiLmHu/oTtg0nwwfqqOhVHpirReW9fslU5l1v3mVQPcLYDA2O99Q4ZmA57Kvu29x
GJRlwUuT4ONbBrMC4VLuq23Z0bQHMLBSA48JTC6aFyLhw9OjLUk1RyU7v64i4GKiaFT6BFiFd3ky
fsCjT8DbQOXsCSwLJODZwdWoxNCzH2eZFW/JNj/Ye2cF1EL4pUYy/o5s+6C9ZscQkKvrWlzuPAkx
nn372Ohm8rx77cMhotVoDXdrqX3xHzPgB6ZIVqxIMn2NI0E5++vSuU2CjlGe+bFp18UnodhCHxxS
Z2C3jd6oWtmQxR5SGeyUF6xQvJAfL23Ga+ozgy7Lu4yNvcF9HS6Zqj8I+V4t99Q8cc2IagsguySR
juRRLamxwW3ZhybjPj3xuugNEyg1d8Ncy0asdQtk0yKLxM1+dLTpmdilyQVpi8wINBka7Anl7TzM
mePstza3tKTHlISg6hyXsvgac1/SYDR7gm1Ll9+QE/mTmDShzC01EqjDRGWsO81arUIDSzCOj0ZS
Wt7/UfEM1Lvu2Z0yDsnosZqnMjZsOVY8cheVynhZqAa3uy2Mvyebaxf4gHNOxlnBOfM5pehRVMGL
2BimAkB7NQEaZ0vkiohzJW1GhqCWKocvULUPKQHAabA8xb3nWWIQzR453C6s1hFSX9/E/ufqGfZv
SlDoqBAn9dZYNIegiJNWEZCGxpvNn4ZlhumHkKS6TgBX4CP/AMWCBeLtelRwMh5TojNQkgNsSoB5
Js39FIY5bVgOpeqWEI6Ui+Z2bID5ibr8ILdNtJ1jeTV+1XYbv2+mSUG87wkLAuEPsV4Z2xLxLiE3
3rgAzrGRZwkV1ZbG0LzKB8uhdiVI72YHsA/gVCywuXh7aTjGpvgNy4RwRcVQ0aB0brGrqtGxxPkS
4dwuQ0d39bKSWs521RbMOUD/35rp3NJFY0ggUJh8M+8LDNECLn3NL7odp0lrNkph3mR38ziP8Pnl
zeZijgeRQKta93BDqBh6KdQ5eMP9VVTX2GoFZ3oMgBR6qRcBoPMQ17XaqVOZbkj6uCH7UGWn4P5A
DpBQDJp1J/JwaCJ+DDLruNfNBdLY6HqnTPb6mCJXGTg3kV0ieUs0aDN1XtpXAlmPPNWJ3Q5OZSCQ
x2LzNRxQPmGO8PqEXcqQkImPMcyZbwBEDh/1huJ0F4fSi/h/VmJxcf7kkZSFVqdH5EpaLSXUUvhe
QR1mnFLuoMtrXQPWUjQBQ8PY7DfiZToTbY5WMw9o/MQVi1qNmibmDXu6u/JiXg+5b+I1mtdiU/V0
mpVDwOQR1jGnFwBDMs54Q4vWw334GENoyeYG/0I3GNrnOPI4mYI0yUuGem6GEnGsF56aMdnxQJU1
ctZc0wOrhOQ+2KS+QudyJrVQ/8rx0Qf3EWQ4x/UaKlx7EMzx5RLNUNjD+OJeTuOUdg3BY6RfPfn/
6u9yNQeze+KVY/XmSIe/RvCHag4Vi+iJkibbGc7+3J39+aUq2Kup3NlZtX51NYjc96Mde/ivL/4t
7I8cYRY/asdBahv4XIht/5QhPlYTnMiJo6SnYzb1VQVfZgXcCP3qkfh1ERaGZVBcxf+S636XmHGt
VfXR9SPuYmaQVE8ALNpPu0htPrqUGu6ovFp07WxIJdYmk4hwkGjhWv6PVgnKTw1KgoRqKT3bog6a
RtnAZGGwiytDy7ZISY8IiscAzdPtg4zzflrh3OEuQ4h9B9HEp6D6E+bc65OV4Vc7cz/s+kY4tkwN
XG7fOq5DFtcJq3d2DFyEIvavj+FjNH0ZECWOBMBJgIGQDD8bVOq8x1x2wOVVfekAZByvNC5igxuH
Rtd8p+DO7QzVNGfxNvNaFJVOeM9OxTP9kMdOZ318M0ImldD3tGG+ScXZNs8/QIXeeXYHBN5c6T86
q+4fRV3wu0u9JctOkZ3MiG4bSxk07X63edEXlDZWOLu91v6Y2l7/pOZPMegTMtdDVOtYy5hC5ABy
PL0aNkm69OttLBH/3ZhGgKX3n3ryy31iWcwHjtrc/nkmz6TgIV+sqew3omnq6WdtPiz9w6uDUGRv
GuA4YvFNWsC1VBUyMKyxa8G9EXLySBDH26MCAW8WXMcizBxlcAekdY9O6+XfapejNq8GYGtP7gof
4epXO5JAluTkGnZsTsYdLhLJfconSJAsCkI1ZRPXTi7IgcXmFAkRIDc59E9CI72EyGT9xA/JM+b8
rotwwrcB0M1KhTYRFsY9NlcJr0+ovElv/DgXd4nlDtlfNZhs8BiDjQsMlWy/J8b9/5ZreZ4pQs0X
TOjxXemodC1xr3cZQRVUtWnCZuDyGP9AIOCUwiIBC9bW4dDTkXuRldErJ3odH0J3iw95Udrn7qY6
VWY5qBVDUjHwhdmPwV3PpvcdXj3hB9ybFt6UlurIRNDvcNAkO1m1YCZtFiiWx1sJgFtzavNLHTco
f5twIvJP4mKCOHk5u6vTuQcZJbFY4ETHPuDsyp/6DwHagXhUSc2kdI2CTtYejQ/tVlLjI9vwCjuK
a/HxUIa0HosQ16xNPhiEhikdePTjK66E8O2VMTcN35kmBxttk1yBqtBOdFuAHPSlFG+IbZT9cNV9
UIp8pMfS8JakZKcMfhlMm31Zi5XYwXU2k3DYYcCJIPooen8RNO0VW838IkFMEv+ipu62sX2c7LzI
4SMrQoaougWIc3Efnf/a+7K1VvgqTMk24m5Pm+7qrED0pb4NvxfSUGANCshNBUkKO/OfUuB+Idlz
199x9inoQvtbDtIq4DDdQVunCNlX30CaaRtmvqE9wmwZ5SQ8DC42D1zelyjZ1UYnJq6qXNxHFBvy
HJaQk0AwaL9PCwQcxQKL5E1U7WP4bZRfPK1ptv5yVWdnfKBIwmWQZ+3Yi+8r2i8UBWe14LsWSqHS
gXfxBk53phCVfTNTKaRyYZO3QvNshThlTpicEJHWXCxWvK7p4r8wtSoSfWYUqzLhP9dZCrv0Bnbe
Qfo+OjhFjKP9fiQ7w+dlBwD28OD5Dcgf3hLL2tRX7NxWIYISwU4k2XJFJKvPQg8aBsbpKOXiq93v
uupvQtGP8IfUOrf+dXrGcV4nSirSXwuAxZaSDoUcMvx7VR03BJTlAeFTo8l52/zjQ+iUCobNy4GC
mCj2r2waFxeEfDIRlvwQH0FBx/qK5UyefXwxPMZMVfsI/Sn8KEshe5zxs1g+CZcgh+NX2iVVOKHd
x9HsPN3jD7v9eTG5NjKlEkxX7/k6f5eLvWC5NBLTwSM6pmjZIIK0scBnBSrRwhZHhvTQyNZ9c4GJ
nIGI0HdyoGKX0UrFHgMwtAb/lx4JW+gUPUHeolTHigOc7BGqMhWdGYg+KjD05M0wNx5gx248mARh
GRbE/vWdXoO5P9XFjO2IyANAxqd1BW4ODzQ8JOS/LYv41SqabE23AURQ6zreqnICLNSJ5x3BzDsl
0O3x0DEEa5WKCDAMimp5Vyv1N5Ybn99eKQDEeqP0s/dJiS2R4wC84YodBQAs6NGC8DLw8o5f6VDX
w9hKKZK6eWaWUH5DsnJhRs98aKiML3dkE2drntIp66jy2N1RlCeWpuWWJ6ANilyGDzOvwzNXcmUf
BCSupKjrbzUlwEo1kuU4XvQRceJA8E2YaiVfg3ZYbDUQNzydO1KDS8FTev7yyxkuU8X8zPTaIVsl
zYgFy5MURWk7JZCgw6cXmMK3btRMh8hNEbIEE5oCXnA9omNsOrv64QDmna2u+VYt4P/yjzGQh3Iz
k14pmNwar2Qa95xjM7G1058Rj58e9P8GCz+sVCEJns0k3eAy/cBpzovDo2bK8fZtMIt87g69kipM
4cgwRmy4+U3/ilgBqiRr0IgJIl0vLgfS53hu+BdLIrMRJ+sEyPz6nzqcLdFBqqhW14QWYACvrPHV
prX+bEh8hRhUHDeSHF17jsAm+3RhPb1akwwwDHCZnVMQ0wup8EtWlLx4OZk/W6TU82MFzqpsa5hC
xAdAVE5fpjHnnaFwLuYaS2JLDADlXRf7A5Gv/o9bguwzE37IyjdL1otZTipSEuOAOghcuVRosiwI
kZ6+MWqzyTu6Ms+ZtqXvB7yTTJQO41MhBnH3WEe7/QpejMDCwOutwE5qKN1HL9DRBdKpKStkeW4U
Thman+2fGrf4IJbUg0u+Tcwhu1JapoF3A6KmVKPwQUlUqAxfNAIbm2Cuv3KLSlw3e2OtwuPcVs7u
DKrm19+85V5DDB9DKvPP067vng3DltY/CSqwzlteBK2gcLWk+zeMinJQfK+Z2gImeMUjM416Gj68
9ofOeLYw20Yyech6sJFKHniFv8Xil9sBYK2O4Mp/KfAOV6Lu/TsXhym7H7PW5MpQN0ebAvrAJhSl
cYkmjXD++Dky6eyMP9RkV3t3zbM9cJs0NCAyipWX5EyLEPjp37O20abONlPgkjX4iAn8Ehqp68Sd
QMIgpc95VCnaXED16gdhMcvVs+8ma4bZ+imPtXjQQ6o9cujT2xN3GJIBHV/+1Ym4Wo4+XGYAO4/i
Aacm9vzeg/BqMG/Qu6/NY7faeRqGki751EVNsoR6DpWf36LD7oa7/FhpdnCkJYtRr0N1nzT48wY0
Fjz1SqM2tHLtx4z8SBlMKJfUdDQjXzIKq3kTHX7BRZkr+jgQH00N0vupIxusMuIlXLmSiIstRtYc
YDI4pI/ZXPO4nJ9lXOhtNAAtPpv0S/ig1ANXk32P/dGrF+lZJrHCzDAHZ5BRY3L+ys7ZchxQ8uQL
/QAgwIi/VsZ9gMZkldwR/ox8wHIc3CGxZwrwOYftz2syViC/oP7Nmexm4QeaEgCDfAjnt7u7wc+k
Nzp6S10QV17vu+mzQ8aFNdTMBT3TTSSvgBkQrWXOIfCktgbNdL38iX4pIBvOevAR4prII9tBNdEj
OXnk3gocRolWM9OJsh1XgQ7kaG2a4eytJebOCBlUZ8ehHqIklJ1KwW6r5uAUZMCM4VaFUbPRWp+Y
+6OTIKZ6EbHvXK35ePSngMKGNwbV5dVf3qjm9IeJJSzKjhRDacRff5CxQB4sh6LCvkouASfJ6rPz
Gh9UhWCGwXFrfGRJ3zX+Els5TEhZPSfyuA8cJG1Vd/qt6+HLmpUM7MeGjQGKX7AhnYBrR8D91COp
PO29xSA3Bh1ygWhs1NJUmHrC0bM/CcDaGa4ZQ4anB5X4i/HRv/wGOW6v+xSbaKfD7cvEnhm+hqB+
S/EyVKL8EsZkV+BI/nAH3CxysqsNCmHvW35OCduaHl0yQVU6WvPR3B1my4Q5J2IPoJAkUZgV+YGt
uCI79NKJKvuVDdwmvh9S1KRUzan93SSLSx56ANaHskcfntpMBdZxNfBp0TjKM/H0y9W4/oSLxgtc
Hgp/uvy/6yyQkmUvtShGOy4RPl9adcWOOPEHOi0tMpmoMmkmosIkP+qwaAbA+9+TE6mqnR/P4p1h
PDlkApYbPSdKKf10Tv+ss5B4nneAIQSZUCjqRLFRT/KkC+qGNV5Lxvjjvg7PLfphGptG+Wum0sCq
nNOIRbKl3mOJ38IAu1hJhwzrGzOAfLrLKVDZ3vhMnTJQrQd0xJM8I0Y5+3J45Yj/Pxcoeky1FZ5W
mdGp0PNpayZaOhblIwbfNnkxGpmOBWC/A/6uLM/1AgmoolteTnG0Dn7M+0exTkXGliF+wjZ8PBdD
Q5TvDeriF7+i95qpohsiFeUmyBGDQR51A8RTAvBQmcS+mWMrQ3iiieqbg3u1SqUkptMLdxQ48MG/
EYNGPd4JiXRLAQd41bAIYGYHMgZfJTUtjYbJaG3WBc3IC+rNHxIx9BV0zjdI7p/oaavVWHIwPODk
JFxE+w49e74aazDecqcjjWgvuqlBaMofigUFfPXfK2nS6ZO9yfXIIgrMdsdVuMlwiMvXwNzThl8q
7NPbKR2UnDcdkFK/Pbb79o/HFbdwF8dyWCvT8luZy+MfogUBnOIeWJvQfxHEFzpVLXbXQTN9+PHy
zzAVWiowXLoEf5L7Yzu5cAYj3cisNuYqz73Lfm0KAxoqNLy2PDNHlhVvbqVxI0rqXF9q916rvYNW
KkylQ9VRmmGP/xu0E0uthJdkLCPflWF4ZShmwndIO7Likrn2j+iLTDf4Jhr7JCVwzDDiN2laam4F
KGMj7aHTNkkHslbrgXwMCmC9fV9H3mweFjoNZtEUuDp3MUkH+8WrMgvoWxAIcZU/E1TOaWXYRC6p
IxOzwAVFRUgnLcol1Dr8ip5bahNLZPb1ANmUNQnnI6VzbcHpSvzpYgNGnsqLj9U4iieEBCZGtXPt
pqDT4n4Rb/W9SHgryDnICpOfEyLHPpNkqccv0OaNAHKb8dohyCghkPV80jMgxt7yR9BYk+eXiqEC
1ocFzHb3t8OHahZwOiiP4eWscpMxEIiuWQ7/COW8hzf8syHxRRJtEpEgfKAN4N0GTnkfvUqB+HfC
ENMcERC88Szrt3xYYybqcLd8DRH8RvHzKLGcoKf0qgJPt/PFBuZrgP0S0mhhxSZ2OiTXutSGgWUT
NtaS58HymlSYaOhY+s9G4oimwp6jH2EeJ3FWL/MULTT2pS+wlaHrpCnYS6tN97HHu46c7bbNShRL
XUNLAXCr/vMBPRQsjYOg53+ctrqgrTEzoES/NQVd+F8gzfPB5QLzJPSZB2EF4mr5yqv0Fn7aOA3G
78iOEkvWTB8TlyS66oGtiip0/zGoFwHt1wzLp4xs2JyZ2z7yQzloqyMeIylv+6dmKlNVe/wyoTnU
vf3INUD0h16R+i0DA9rOIyVKCEz5CfSfe+RVNVbHRSdKxmo2fWLtmk2wsfLuOXPPvxo0NMOhDJIS
91X5sddzbNtGmNKAnC6+OVFNgf7Sef6S0806Yt+ePfUdm7rvjwrfuMhwQiNPyGuTQszofmNiQffH
Yz+3Wgr9FlSgwWF50RpCsjLBX4SBQDMIevk5Ldyem2g7pfkiONQaHQCtfMh/KC6eHtz05qzqwHSL
Vy9+M7Egonwj0xH5gW+0j3dRNDxj9hS4xWhqcMwgRjYOr0067aU4skfCkabZ8dHTz05Xm0pccMNg
koPcHM3Mzx9chHOo7G7Mz/FKH2pwBEjg8yNxN76ETxo5JgewyOMxcleVur1OQN7AsuEEO8v8AZjm
Xc+NBZxGH3U5NhIfWp55HC2GW9NFML2/t4f+vikQi6dOsuGknv2XhQ2grDfbylao7n0K/GU4/W+G
DBhGQxgdXyVrBkpsoY/T10QZVsk4qnzZYG9DqrJbpkpsceEjsboMk73mg8rADqJEW/OKlS6EuQc4
jHteqZW+6uYwFWvao6Jxc6hk6wdji5tTW1qqiZy2OAFV9x0N/po5oIzqEHfhuDcvaoiRewCrKnxn
S1H/2SZwuJ780C+5PFJ/KwP+mBAClg1SkEWH7z44A/tIA9HdJUp76MsgEGzXEw/rRuv5RomPKP3K
aBO6AeRvSey0R2/2VhoUpBYWfyTud+FXHY8z5x0S6ULl0sWhCVQVhj8oIx8s0O1piMazH6ihqOeK
+pvjxb0itGmOlqibvA0jGsdoaRXhbKHahGKhUaroqBEUWBuOCcwRsHgILzHgw+weo7MJpn/rnRiw
hcGl8iLZE4d5+kZSAQLl4OPmikqYqnKt6QPhMcGJDgX/kPlQPAygU3fa3BzkDngs/HjnLIwztZQk
0aJSiF+7+TAkujpXehBDDGOIvDn5BXaNR5WlZZTRi4dS9pbSV7RVdpeiNAe6Q1YQe/wE0c5z8YJj
39IXOE98Gt85jB6l4R3wUfhbEqufgm3bUvi8nuvYoluENjt4FQR7w39bDp2KO141Y4B1XPrO7cQw
Xi/br85IbGj2V8SsRQgkIHvv8pTRcTQRys37+Z2M6yOQGuF04wvMYWVwZVsaq9NTYIpaZZgone8J
yaATMSS133BBrnQx8nBHr6PMP1IiiMkc/QuqdiGfasUTJFjz5LJ8+ko/XcIdWcW8Geo5fu+LiPVc
oPDEJtosSrw6rFZAFy9xoOZD/OSUT4sdCNdaCeARWkkC1VGTsz95wFaZInAyVtAXe2N684l9RPbQ
wgUOa1YcHsUMPGhc25SemZjtsGqUutbZSFBI6JuA3nthky1B1e+eB/SSdBYiR2Zm8o7qXsYsQXfw
TcdxjCgoiXa8pOHMGaJk9giwxODa51YSNsz8ZlksYL0LosbtIshIu3Yz+JikMfGliIWvPNX2vcGh
q0IBohMyO258LF5zJCw2z/UT069OD/5FPgQ0tBYUF16KQdxVCkJWVY6CRnpidg2U7zyaAkPvMUPS
nAuVl3TO6wed4FxcbmzNkQr/MO66+6hLFKQyHYUomrjH4jKSyeiaKCPeSKqBoWWT9bOwsOKvo0yB
9/wjhw9BocYMxc4PX7SO9vZgnwvt2t+8SbXHeWa5EvRbDyMEBNgMMfzjUhxUAu4UdzcC+KZ1Lk76
ZgS+KErl7Ybl2P732CgqnQRBzEJdyBHocLZKejhAB6FAZNXIaZfznDp71DFNty4d+TlWBxOYhOGt
IfY+J0scdOE41Pl5k40sVpqTVBiybAfFk/sXJLt62X273mkn8jA/iNTm2Q9AJO2u152ySev9qGGZ
7f69dbS/WIMSk3uf9od3etV2EjzlShWJPblVlRz6JdV08++vEAyO6S97I0srBmPGC00pSlCepiPW
/F6TR+9Dfjn+bm46AG8TRsHVUzFUfY29XOB2+btlfpOE7NnXup0Cv1o7dGq3mB69JP3CJMZJlKoS
PHN4HblTMzKc3B+qkWgCRbQj66o3ptZYN426uGKtSQWLxvkVstG1EkKyuPhZjxlOFF0W2poXB900
pGxsmMVEKKGTxSs/eruDgq/rOLP178gNRTmXDz6KmrfBLW9/VAJS2O4lADDICjcqtbNPeSUS3zlC
lqn/OBPN65eiSLgEFOf7GhLAcqNrtHgNVReZ8oYsSb7Szc3W/I4lK0Q2HQg5HWTOQ3IBeXJe4zru
rJ8wTiemH449dHKxvuGGhD13VRAtgwCY1fAVE00UaT4T4KjMbiVrBKFPaJLU1/YH0Unmllj+/uua
YXrkSyNl6UVbezD0luBnktvdhoL266kETGN38jZIuMyPLEEezFK79HWE08k0YHJHJG9qc5i9KDCm
TF5b+rBBq6r2qCZ8X92i3RPoLezs9axW34xjg6ki32Ir4skdof8RGB3c8fG9I9qcSf/cVK1RidKz
i5ycX1NlD0Gb+HFEN5stl4/U9hZv1kOkZqWKmFV/hpud7UYxdJ8a6OnezsoL4iim/22TS1dc4fA6
McLulhySyXdhBKSWBeOgFqy7TijArxNR8084CkknxWeOZg9W2PTMlGBzQDpSuHv1InkDHtbPQRf1
rFT+ViRg/7NbIPeaJabT/Bl7V9l64aEeGr7DiqpSj8qZL2rkn/o+PdRj1G4OjNf6Ei2Av15H8uMu
CIowPJ3fu1XQ4pSF0azuaa5fWUYrH8KP9+0Zdc2/IvEyeG63DKuQ79Rpe+UuMijlHdSWiskfm9wf
MuCcMBFb0O8SnGJFKRa7v8tcflIXuaxLxwJqMjNm0ca1dDxIXq88AzZv6rlTXztCEpHGLJJclXsb
pqf9/rR+fWlGH+LT9n2m92bQc5sN4CTqgupqySJd5B3XjjKUbv8FJKItDCiLEUqLahU2BC+ehSxH
u7eBSIjgU+jlLSmpQQSFbNVN7btsWLXD9z9aEKTF/cidw/CW3+M0XtmeNwZe5BnEGndoO5kKIg0m
51t+0NEOsU3aff2goMUL5S5ZYdUW2Wum2Y4HDt9kYvpZXkXiVvXfRekz8dFCzzAtANYyBEQxyIJO
8q4A0cbeINVgJyU+TFkNhNq2B+4idfJEat02+Kt9EXT8WMx09DNUVhaIzsoEBIVHRL3ixK2coRpO
VvY1LquE27SQJxUk5jVdprB6EzH0V1iwFpG4b/faLtSqvDEAfNGmi3+zgUpfeEgbbas7LYYDSDMn
4PpmtZnCv40i8fhae1K/sRpD5px80hutr9f5ZizF13BDKohI2dItFiAP/jqQTBDxRHCT8ketliJ5
Cy6uZnPGWwcYwKTFKuXxA+vcGGq/Cvbp4j5Zcg8nEdYdqlmxanOpbg7AsNm/jZ1PViU0Q6KVOa7v
RYIlfeKlVGugh+aa/oDaxmkfsa0M0De3RZAOQzIfnooonif6j52FN1TiZL0QyqGADZMTD7DgPXfj
WS30//8XSmNLMOYO23BMiQK0XJmsI+eq5ey190lt06LX/ytgjgvbXnVj4uPcWAr1bo0rG/WyZofr
025PJHi+D6NaJ13JNWppeqqS1hDonv7WWnQOYIeVTJnZJ1VOMr7kPJb+PeYuEPbshQp3ccICQ7JD
zIoQyJCGpJ9DWeOrHEBULL5VrrK21SVRzhXaci+fAGlnt/YnSkRwx8xIsiB59W76I3EYSXtWM7uJ
z6pbIYqsfyl6i3p8jisWmMfrzUsvWZxcdzIA40NW9NEPWZGgCcR2zriKF3eX84LonT18eDvtsoXK
pjraNdcjo+4Rwq4gFCJMenhYyVx7+tpcxncSi3BaHqoTJx8VFsytyhMuBx2gYFiGFvkY3mlYWhAX
rwmsS1qcqyePEYRuJtRPqR+1xUs2cDvUmqApmO3tjbFi/eZkgxbKu5Tv2dP0Qi4SObvoEO2WYEBd
y1WysWqK9VixFIYnG4s+kv/ms9GHjEQISv43izyvV6L/e6dS7rgF2vEpOpnP/YuxSdqSTHTsG+dj
S06MU3mko4TCkKlDDuVI+1Rp5tkqnJVTHU1qBRvJ7YVFSQTzP5Ai/J0wC5hYOq7QYbB2qYQPjZH/
eCkFWsb908U9mRMYb91HXsFQrHEqxulm2+uPDzrdEslCQu2qmgDjMgZMLJsVGhnPwsZKxvo5qRBM
ge9q0VQ9JmQHdi5BISaNJsjnSzuT83gofAXZwkAj6XM5EaAAsVB/4DJS/5YLLa4suR0sBJ0fFwjj
R/GsQT1e7WR3QhIUHGTaoYexhDnsJmEspGIJPESlotiRwq1O0hItSt1Unb4LxOYLluP/mQgu9WrS
LYzs5dktJQ982MqvTjtQdVEEtb/KyGZL61yiULh+FaRYxQ01GSJpmgjbKgA7dVz6n4AYnjr07sdl
RtPbVzDXf1t/xWCVPKlEUIVeOHkkOUWdogfiws4QigDklfVVFG8BczDQ5N1ikfxedtD6W27PAFLS
ubX4Bhfop1nn9O+pkCjX8N0K18Ty8BVpeXtjVyy/nV9gxzKruItuzeMXY1L56sbqe14GWYUy1u3d
Di5dJYREpmMmEJw4fUYOJYdBNPH2zbkbf089ZU5QoY4fx3vV/qM8z/C5zfIRG8VJnx7HcMZiJOrc
7pa3uD9jehYKcPmtsrY5wIazP+aucWeRmC2/m1Haji2bQbix1BmIv22ljRNKLE9sdZRb71wEqwUV
VQ+5E5Zfc7mMB/8PA16DfMlhZdGpML4OKu4493d329KYbcSM5QDMHhoZ3OrNyBAx9l87ztz0HjwZ
rHUk+cByN4HesIoBouR2AecuzKldofQJII+U0g2yZbICwE5AyigEcaUMCIXIUba/0IBlbqdjKmqR
OfhU6LEOePyi/gtDdBFQFcDNugKtsHvuoLwSnIPQEB6p71GFAwKU2kJbcLQgARoo1YUUL0mThSKV
6ADIzK08FX3Th/N96m9QgsTDeWliJefs0H1OZ5AaqNrmopUJlKGRsDd3EkRqB7ssXHbaMuz9osHO
2SDsT3lxpo/wU+7aSBl0cOlLwDlBBRqcL4w7NROLkP3Poeqa6QDBTnwR4UX7cMh1IRCy8yzoEO9G
lDjf4LwP+Cr55+ilveM1e4+5rsxA56ftKe7bDk1Q9a5a/nyiEMY54FsaNBKFCw9Tor51fUoCstMe
CpZaO2uN41D+M39/qcBi68tMdHjORbDTtNo9ScCydW3b6JER9owJIDTE0YV8+6wRnrjMfRdqDM42
pb16XE9H5eajprl4TDX/qrQ4OQSCFFjfOB2R0WYt1AKRpFgBmzI+/c9kR4PHQ2gL2jgjzEqhkton
JZ7mzoUVF9zLcwSMk7i09ZzsruXkEFDiDNyNwO43w2HVD51kcX1vupO0Wek2ckpau6r0M0iF7JPC
rowLJIp0U4fsWykTYRXmrCPl0nP2T8pHZRt5FAWVkPySpgP80yvmvx3wKieRBud5bcCiJhS+B06b
1se+KE50JbL8HHQEmBc5xg5Pklii0WUaPj8drVxsIH8ugdC9gE/1+a5FgFe3WnsexcXGn/nQYJ6U
kdzTjhD8UJmsVXpO8r47+UlOgjDgfW+p6IwMO3ZyZ3YMBclnSGHqO0V2l7cO2EJLdUAk0trlGj8R
7HAHamfb4XULJD3QsWd3zJBohY1kQ63pOF1vcBSa7WQ9WyM/nwknCu6SarBMJZZ4NtnJBa5H2ZTu
K/l7XjAKaXC2CtKxNBy6F3AMKGyW1HtMRmMdE4AiHKC8carIB1oz5vYhWhrhzZ/ZEtJ7jx1u8eTj
7Mv38k81ZpkyuMEfeM7w6KFC2YN9Basdwt/mA8HjEPk/YwvlgasVCyVTKAoPVysVBsXTR4Fw0MgM
e42FyJ9/MJNaIAAM6Y5FLnhXU6pBfRnoFZ2CTKnx8ZY771s0vUJcDHJDPgSvvj45m9HXpea4BgRU
GR/itqngBqfRq/QkmiSYyWqS3tPcpxG/JyZTlLtLvJ0YEiBs0iEfajebz11fwsrsz7gCUJE3Ow2f
G7u71WL0J5Pop6ieEi0y+Oc8q5pPA6uTAPPOqx1zUkSBdYUorOh0dOSm/dDxUiZM5Ni1YDCr6D19
NPWjNZ2QQWPjxUS3FL9vVF1HNo3U5TSNkb3p0oJsqqajusg6GnNHiu49CGyMGLt9nBlImDzWxDLt
zqJUD4Nlwoev2GT0P57MY9GN/eAiOrXtNjlAVr0IcnTcLB0ZH9P5jGPIWt55p2qve/zEI4iM2iSb
ZaMTvgB/zOoerdIyqspDMlXnzsJD/DtK/bYsR9jY7rpxXhxI8+3QTa1SsUUdD5bgIh18GaA+5KzS
xFTO9sImmOXl1gQM18SFYTnvvs3KHDyTdU5OnB0jeeGjcq24L3cvOPRh5sdPKA1ZpldiQdFgWIR1
UDM0Sk7a/ZShBFQcya5I8YVJKVQQA6Si3tCQcTkofxgXJspq1DLBxugFsSlDgg/bmJ2K5lIfsMtO
In18nZy/PN3MW5pSDH3XUT+Fj1dq9UbVZWwpSkVmdESQXFk1b3K5SQOL3DjQRDqdIPCbbDw63U66
dV0oNi4gXmcnxXGYRuQFACcjUCKzCzMrk+b6JoB/Mb/flQtA1sqTNuyvZK7yIPa1NrOgLvFleNK+
fegRIIDnqXIwC7Yq48fUV8LWujUnXmurMeH8p/U/TgN1bRJWuQXyg0KHjoMnBDM8JeifnM/3uEkb
1q+5clECyBo8O5tTqRZ6e8HD2qowM80/e0o8yEWGaRAJSNJ927NLCDuzOoy7UBH9I1zQmcDK7LQy
G76hzJf8Hzo0RTn4eoBxsUq0qgR/SHY6Sr5bFlJc5UfSQnadBKdXHkYaJoXwW60nEcsfekzpPEwO
hMeSJ3hISX11sxqjreikqLLUrKLwDjwT3QOZhFuPEU4SqvHD7rR1xmAlcq4ZSQu+SzPQhjkCQWkJ
hYImG61nGBxSZfzs0TcCXXe+2l0yFFmtzH2n6Z+OOGH5RI6A0u7BL8f+dUDD2xOoA5jLqspag88+
Irtc0CgrKgMZnWpKlQwAvilkDy+L/T0jMxCwTViYTy6zuAloHpStlCFUIVH1FqSZXwhTjmmITW/k
qTt21jXe9JnUgO8DWSOM7kgVM3CEO2YcYg6o2HZmWpfb+pPp+v3rdQVZlGKPCD0mtbzl4RADqtTa
REH4O2uaz5FnaBI5p9loKgpPAiYXb+9T1/pWICtLCDesxHs9oCfgDlIII9QetdaCoTdHdGXAoC3g
pOMBm2mN0npoMkjMaatDF4H+kKA0kVlaHVgGhyHkAJIEX80vdzU2HcYWVQ0+o3e2g5j4qVu+2WAN
BXG33VYR9XJxnNtS6C9Voj/ftuAKsuiHY2Y3swsbq6+cNB7qgKjNsGk6XNpjVHQ1DM4zJP7mzD0+
JpAzzy+BaGCndJYUu9jAIshJYT9Xf11KRT33Nb7l/MxIWKgpdix/pNqnlYx4u6kSiM40iwQydMc9
NrTsBx33THL59ICVboxVAqWSKt4mFSOhucIy8OXFWpL8AOP950ZeSyY6/khXHZA/CmnvPhxzQiSr
+Yoz5eKC79u78lnh5MHZySg1Ya/CJog8Rzzuv4y5PCTq+PUus4CDSCOJps+yv1MIQLur8hCsGH4J
HHXuklR6agqt9KPwaMR/B4WNA05Ojjp3S290Su/cyIsA9XkWLHoc9w8Tc7Ed6j/WyJfMDZCxubU2
3ncG8wI6RJNX/SpGR+y4/86JS68PM5Z7fUD0mW0ZymiY+MUk95JP9cYvfVqpAhwX/WbYzcrlrjKs
0qfry9qmEDf6oRzRCOtruSUFlq4r45PoqpfaKOH/MFfFieDYIpCOA04U9HOBRXtN0+K7kPDF4Gt8
1M2jvsj6l+7oInjbMO/syNs8wVlM0XCCEuq+b+1PggY62UNJJu3SSMepRN81R6v4Vo0lE1iuv4FE
vGg3pX1ZZiWWkfmroBJBKL/u5sN5sUTuQthQRggsE6NQkyFNSbrPXm3Ni3cUFiAuoSomQ7KRO3SH
SugPmqPYWW7Q1OADJEyM9LdcDUi9P5dQSBSOPlIh1cDJbaWw/2WZd2zlhRGr06NgOyVr9HKgxThX
fTX9HjfynfaEroFFkuGPUvueARZk8M3kjMtUCZ04EjLV4t0K6sJ6xd2O7M3yk9t3472g1XdtIe2S
YnK5B5g0l4ymjTuy8PiO34D5VV2w0STENchGS9ljfkKLqox0wDHVOjvJEPUf4lj7AuPTeuPWAeHr
IkhZxp2aAV1Yud5mTyRJNH5b0aJzOhDHaQtP+YEeAIrJNifGHpcB8ZJwDC1IKi/9+3uJruNrJDN7
c/nqOmvIIJsLKoJpdZq4l1M+qW0GZpWW0u581S69ix9tn5aqbJXzBCQQnnVoS8g8gnk+HRqjw1q1
5FFdbj41CPJJhAJQ9cyc8N9Fssxil3s6555Haj3gQO53cQY871q01qWJfAS1omy8bI/0ocHfOvZX
wEJtNIC5CzAflKKpgb0Ym8nZjCzrHt7wKJqsC/8H9tc5WHk0W19NAWyAuyruQ9+Ah0/dRs1Inb61
/7e1F9BX/VnNfwcXXqx1OMuitG6NjSC52zrRb60LhtNSxhjbTo4rmEvF93YQ21Gq9lSNgdWw2LSY
GNntqtOZKj0jfhIFqAZRC0h3fkP0jcjgO+wL1Qs+PXNXVsw3RXWaSHm6YSKbfAr4tptLpjl2m/MC
EGmhG1f7++xUmz1VlzFC456s08/glfMFnFbEh9Ynt1eCkYifA5Ge65W2znFYAYiumCkbyR4YaUq1
z+0ybm/F2nVKqzT4iWPNo/Lm+/IgCHI720VJRLcUTj5/46JW3cxWYZIr9XbsaT8CjqKoTm65Lm0r
2QOlze9ZTyZZmTVZCmy9jTitF+Fi8yoPBBT1yb2NC0ZoiAihcG8WS5CskZFQBwzk3HwUAAmixlE2
Zez7433it7TRe80eHIYqwVk5KdhCNUNoNDN4p3mJhfjfpw6CKUUdQDZoYrkBOJmtdPfXplrwF08i
Xd6B8vIY92ylSpvjMZHgmug9AqPAi/fmsrz2uD9+TXro7RcOS2fCd4AaXqoRp7L6E/9Gsch6Fm41
9Lc5ZlZJaD287KK18QoPBY44WYp/MIOpGzEvAhx52Klmf6piJ3A4JiR7BPxCxVDdKgFGedCfcghW
x/wCbFv7JCmdpuGwFTdj9yMwVlDHuQJyT6fRTpgXEYNuwiIZx/u2dZSQwQ8hpqeSXWIPsm4w5ajq
kvp7bzhu2kiadK8q5Zo4y6qavhbLwzwJnkjZoShT5IzXS8PzAevdnUuOhqzKOV381eYEteLfqaQD
nPHEzVfhWtphknbnJTUou2M53g91nWmNJoRW/0W1J1w7NrrLaQA32k5Tw3gCjuXqMk14ea7k8YWz
UqEqPh2J4ly8F8aTfBtUEsluTdklba/BCp22bFl9R+0CrQtPU4rh49Tq0NCgAQ4aGAw4InJiCeR7
FqI2YtLfTnYmtST2ZEOwMdGaiQJtcZuZqLCcNDb3aSw/BafR0HvKJZDpq2IcRii9v+6N4YjhAkNe
wmNLCU4FuYon11ZjP5d9EDf5okpIsYL46p+DpWA9ExYdF1PrcyXY/ubrkxk4ddijYS09wkC57d7e
ukTrnlYmDBdG0dsuTRtCLTmX1A6Q+hzXaMj/hZNHll4eWBCyieFNUjs8NH6YDK3qbc4clTJNP9Hp
E+bCT76PYJ4jqOF71IoWWpB1nUsokNRjZJnrcAVtUt44A48dHyIBJDUJ8t9WC9ZVd29CLO6YmVXE
qfaO7VtCFh8rRIYNgd7Bp7AvZlaXKqXdsms+GsdQi9Vi/E8G0UrbkFzvOeULX6G6fgOKUBApzbuS
z+y4AaqfI7iBzK+xLNrZOr8VOuHNmGPk5xDhaLHBe+GmOvp9wpxaUUzTfAtRzkyNYmSIciLBrCOH
MB1v5bpWuOZNm4BexIwUnXpf3zGaPdS/b/t5RN3289DJW3JliXOYBcdCy4US3M5rFyG3SjmHx6E6
XjHS2Ess/B7M4fQGTG1F19dOvYnTYwGxgr619xlvBh1O8ajQt9AiXh+YrhYkSvwqjhixJ5yFv8k/
3ogYH1+i3zLQYYxeTyOn1taQNcpky/yLGh412RInRFMslz2+N5zjRnzBdY9fvXHMgIWOmtugByVx
nMc0RqKFzhnG1gpPEvzQvWqQQ0U0O7Qxzq9CIbgZH3nTU8AOrCxEN6Ri4X7reBwyPUtlpfiitR4V
3nWsncflZskFqyyq7TdFR4kDcyE9f7uRuTOJIJrplpm7aFXyTSPoKBQcS/+S4BfX0umBRT64qy1D
mTh0IDABclCZbZTAhY8EsRimx4RFR5Sbe50q1ZZRj8L6qNhKzIFmJZA9ZLtejWBxwKXUcGMje89S
eaA4BLah103/36Wr/5+h4dhFZ8d/l7rNUvKlntGGhWyEuhxGdge0HroClosae7WEUdkvEc4Wsh26
sLWnzsjS6Jxc9CvLwcCEOvb2NQDZww0E4HmTAvix4tNpCsVlonGbV5AKigiKltqm7DSf0dVN6e0U
pI74fxX1RIv55yZ2QH+NtIyTSE+xfyTe6bzD89W+0VDfGwHLPHL7/TpMjj1ZNoE6c+ZNZlFUMJD6
P2qfN7mOpm++VaEFRpe0qICTHopooSudU5azAIoAz4gNOZESZZkrI68wGAhAHFIj/8ChRfUGvuiz
iyTQpcvWZZjfnyo9GxfVK683PYqDct9VCUFmt+F0OYjEajCTkVA/ClHx3gScglbGKHZ5aIIMpxUf
X+s7EFUNNm6v95Ez5Z/sY3w6Vl7uf7PWjhWeI/12SV6WgAU3ZveiNoJ4z2ka3ZAO6vZ4M/47qJ9p
LfXiOcBSpJaESfLjqq2ZlPNUF/qePwcisgK2+NUUkTCy0ElQY2tAWCL8mB8OctCH7vOg8xjR21k1
AwHde1TYCRhGYK9RiwTGiG6oNVAZtJeG3FIW64i1MdejIopsQ5cqcmJqNltkBxGoJajvsCbVV1IT
KSPNe/NxM3Lkt3VF8N/riMbEsb6xK7FFf8S3p1s4Ovfg4G08BFEWXEX+wZH3d4eIdqS8s+sEBeek
e17O/CSR0sOWPCTGYFCpMTJxlQ6wrFZKOqNsu/Il07hb43fASwNx0NPe8FUwz2u+ExNxuVg4nMAy
wFHCUY1TibCn2mQI3U8Xpzspn4XIuXdk0E/SjM9A7bFmOXjbiWV+jM9Fl1lNM/GWmay08CXFPLuA
tonzDfw/7EoK2q2c/uF+Ml/Pr99ii9SB2ZZ7gKusSSJwf0i4RMLPgn7+2xvg9qAQRGdUYV56Kkji
tsFQfPhYTWTMhElCtciCDjTi80aOeMbh6iicGtYcK7aoHivuVFatPiXAQFvFEGuWhfAtPWicP8VT
neGTqJnwQx1qncBv1dor9GpHrBp0PnxJ1SGPEW5t2SxSAXIWPDwdoYB4Z6pa1O/WU1SRnqYOVRka
W/9rz8WdEcLP4xpKu72cH6O1SRvzvf9ng0QtYLidqBwWfyzR4DyTuTyH7epP8xWDV6GLiQfhA+UK
28pCZIXpoLIm7srftbO7kU9zQikHaMwfQ1f1zXXxXbL6X5AuVfrlsdyFLU3pXKZb+4mJI41Lk1dQ
UT+9NgOJBGjvwx6o3KW1oH8OU/W5qNckOJ+ylnNMXKnyqaqvDOKtxjjqeXKPQRkaSe9XdECedhdQ
/ToH77fnqb48fEpUfrpIbQbMIyXcoTtOUovwLnJsIVyZDc2ueG8P5qaMaHhMew4oBDRBALx8opz6
+Hsrn4nCYTuREOLXQZPS8x23N1RKVuuYJbYXs5vjKrVbnB9RZ37i7eAx2v90C1izGLli5Mmuzf1s
gUcuDLU7ahbrjTvI6qrtFFbPbiNv7hfjbHNIig0QbzcJhiM+jJSEKknI06yTQ/OPl7jBI786o/Z0
L2XBrortoueu3sjhJSrTYCO28FL1kNDLbIB03GkwKojw3bygjT/Gslo5SEbNKHkhONxcLxo4nyqM
9US9pzOeKprZF+lVkDfvrLuZJWwM1CL2iCrnd/xVZvVPO2zXFFJvR9jKRC3Zfb/mdZKOg6kU2/iM
fI0x8ofkCrY+K+PV6FBctzkmYcqDKDd3AoiJXw+BRjDY0UGRsDxQZ8UHfNCjkz3ht7XBYTQrVR1z
OzSe2w4QqymgE+e9tifbyr1RaHYS3mlfU24gwMqHZ/lUqopddclQQcqxekcaZP2WlilwDb2C3gD/
IEqdAGqlvL2pzn/7Iu5MdEQEcXVE+BRMGwJCbcm0NAMs95wnIro758MdcJlBZPAx/MEVXD1yiscB
mc/pRs7NbG1wU6uQmrwDbk93cti2TE1itfDhdZRuwnTlrQhd/uvwlGM6DbPQBzG3ze1xNKPGX+b0
HorwnKZ++vV5VaDq3E0DLYlZG2HcfSYaYuzLDpRD+YonJHlVGjR14L7VHKiXmmYegBxPXYtgzccL
UafsLRbrjVsmf4GYNDsd23Py7PF0QIyw/jUNHhyGocB64QpQRaAwiKsVwG3Mtno9JKlcO2Fs1PZX
R9W9IQ/LCYuXG4R6QkMhgfsDN5B5z+sj9GrCVznEW9od+o6y5TSmAuRPfPW7mHb39zDZs7bjoegm
DlQJ6LmAUcpmsOfgOTif+z2T6VQfhduM37pxNlWiPis4RuZruyVnA73dNl5qiWcmcsm/e5d7+0/H
4xvFjmU3Zh2ybd84vJeqK+U7n3hB2y+Is4tkMpseAJZMnUI5EiEli9PO0yk22zdbSi0kPt7kyDND
QNhKV8CHN1LsN5C9mDG8KKtr73+rqp+rBo94tHcCIHTIGToRrS2i1pqbjeWvN6Dnu0KjcBYuO9Ki
+DNnbP7NTfW1sIgU8ilzaK3EyAMv39tbQy5EAyQNtn17lRJmqx/Tqt8rP3gtvEevp9E3vRMEE0dK
ZRui8P2Q1oMvpTvn9JnaHj/Hy5f/03QKLj0v7W3I2QoGXRLYE25YtBiHbshsfR8Nupu1CpZDDvFo
bHqNpsS9SvNjMKAhZODTNjFI6z5FvSMNUFV6ugGtqiNYtcYA3bWpEWPaGD4xLl1DQ/2Kf/ge1BoD
kKcGmTQWSOHvlvoC1/nSj0dc7pzBiZZaItp6EFSyjySfa2IO9oUZF4O2LLyZBjMgJ4A3l7oOh6AP
zv0FGoPb27TfubxOIME8VboF46bTtAqsEqPUlyRMbiriSi/ol7QG63eeBoRjrvNxTI3n7JAOilP2
RQJ5clFAdYu0IlAlssf1PJfQy126wZJDWzOQUNrRT6ly3HyWKFewWa9NPvMVyM5JbEtSxDlynuo4
n3zhk2oF0H3Nn7QcY/PlqfzKuSTUsxV/tNk74KOFjaSPRZkjIU9y/+oVIodqhG4Arw3InZTyQsPv
8/UwsTycMg4KLyAQgxTHq/wMgr1FZp1RQ46JiafsueDrblQL5DZfF2NIa2iXf1AmFQOB7TF8AzLd
QsTW/jmi3t4sPwaqvEZ6qC42xIpco/Tin1lUiupWe3VH27IqUVMH3u0aXlJLe3N9BLBQIVDaZ/EZ
nJEZ9mr4BA80jOa4W+uyMOpkAKtjXzDJWhl8TV+hI+5Ob75RlhkaTwb60TNbH7P6GxH5Ckq37LPY
R+0L8f3LwuXw1GVuuwpvEvKv9W4fam97tVkC7ghwNwpJFFb3aM89ZkGwCTe9wUMqSg+BJcN1a2/r
hTqf5AASNrOPtOideqmLeBcqml/a+fSCc3f9nQhdYD6AG/mC12hpFHnfSIco25licPIF4frme1lW
4DRtwiLHnprfYFnWpPA0r0XOW8HQiO/67cM349JJMkg5Uhg4sTJbmnNwbLTWarF2KTx3OnaAKQta
ykCbYi6EcHVqR1WxfvxIvaMtRQYtWD+VQpzgz0XY6tvc4/w5R/ABtl3OxuvBEvaQS5mgmrMMcy1m
WowjgMSSuHKMbj7XvkhJPvCZWoM8ckNSKLj8SzwIGQ05nkyMBnBNxjdOZMFa1NMNFJmg7djfazg+
jQ7rKHCDJV10ru7qBM7/qKOeiH5CblNhdGEAkBfYd/PIzhrZaA4jWKZZBLUYnRgsSIA/FbNB0qwS
3yjGBf/JDSQeBwi1pugSab7IV/q5biqEKyWsf2jO84n9Yk6dxSQGi4AuYPZMJLw1+OgF/GojpZq/
illQDCVUqjUrFFBsLYd27x9EuRwjTWMSTGIzvaVijktr++YAPjpEeMKluYPdQgSwdJwcpH7tAsqF
F1ZAnqLuDGRClpPT1FP6nlUvNC+/tqAogbafhAupobw0ODkr7y3j6GVVfB2VpP5fFNetzieUkBbY
V7jwXX8oRTyAsvVD8HFV3V65hQcJH2jhXWxq02R49GU2rxIcUfB26EX5S2frqDrYo294lG1y+quR
y8KRxrow63pdt95BjBkCANlFhpZouzLHuZOjqzjhsXPSjoE2wgrpE8sSsDrr56JebJOtpJpXoFx0
/OXLsbal9IGV6AcnceuFcKzDlLieOW8lpCVYorDKYKIRnXF3mDj8APxZYRzKRSSpAWQciRAC7/n/
TNnRuEhs3gN5/yZs419EXewtTCc+KHwp5HGUOjsDB6jqK6qxcqBrJsObGH6nK5v9II6YiiAPw4+A
giwZLF/WOBY4KfpdJLXROSaYEaKoepEPMU1OHo0SZ4Db7pgVaXreIew13N3lpqseQi9Hwy0Tm/cL
IlY9cl7/6cI9xGwl6z9dCphQxHarJByFnpOa7w1mGOGaCSIG/pbveIhLGb4rQz4sU9PVfNtStlEA
5+T11M21ntzxon/cyRhHLp8NaSRJ8/pzT1XjHlfjKvlUpxjDmMgTQJ0SAauyrHuHHVVHi8nM0V+7
iWlGbvNdnIkZN+bASp1nP1dnVwX2JvpRoRvDR0V3L94gWsL3VQCFwDvU49Yvs8V7oU3G+vhyoY1G
RjLKBz3TzhzVIcJdiagUOQdyoo0jXFEIyotv3MxIr4hEW+q16xTWVWH0QDos9w8nUSpyHHUNQzl6
3TQRhZhFC01Lg3otnEeq54r67/iEYmppqAKX0j4xrgpxOBIEtYAOXjd93LCAgA+P4TflBFc/XQT1
b7H6RvXCIFJDgA3FuCMWMnXjkLxlPCOPjVC0ZvBd+RZotgC5oaQ4rD0lDf6QuVDNdMb12VY449Cn
UMeGerX9mMTaaAtRZ7vfXk/sGc7KgDnO+w7F81ShxRM7BrR78pV/qqgj0vXHmwFPVYr6XaBOs/Tt
ilK3eF2sB6/9XQIdSk52nnItcEBfjP2dF7p1Ds3WAHLSo8SvkGmY7TwDZ8TwmMI66WjsaiduWn5n
cyr9fpQ57PpOlSFJAim6YSUMM0xy8ZQZblVSIC92SEcyzadUHwpqFwsc2ze6wQG5fe0SowIFLjMd
B4hUttHvhYhlZ6eSIDqDYc/ejseJvWEzWMYBRCoyuAs34QVA56spZdW85cuZ6sbkdCX2AohKxxei
IA7qeguQ2EvzZTMREgmOnZnoIWaaBHqmIuQn+0uLhZzDKczPvRYRTGOXpoRfpdlETeaBwz93hyFB
6TWCG0gVxRrG5jbJeP1Aw7CWBpzVG3uF6Y1N4z8L5xWMzwBUeYnAHt9GiU9perZPG7EyKEBCl3/Z
yZGYFGg95ysWXhJt9vV7cKyvZSwhy7wcW29AzOnih3c3YucYZQ7oPHjf2vStqF9Gpb+Oox1v38Wn
tK9Hmpbdz4GPakUVCPuLAufLb1SGvE+DwuZFSzGSm6Nndj9Lmupmg5xGmAxLAP28qIFBuG9JGodm
hNj733NUsUCibNJS63YrpHLgO5pUK6SkE3U1OFrHCzPtbUUMixqZYtH/1X1ylbzMper5/nA7vltd
Z2xApH5vlnAcgUq9LW+PeNnx6YannakaUbK/CeqLpPq78QDGVBpVAtgxsSDTGbvTlf9zflkGwP7L
5mIi9o/AhyVtI9EZy6mfQN7WA/44A0zw2ODsrvy3ulTfP8lNYKTur7W28ES4GrT5WBPGJ5WJiV+X
IpdqURbWKtpRGkcy5fKPpCflQd1kIuhzdWJxHb3jKA/aO+rMiCszsfwR0PFUYTN7Tx6KtTDAEd/c
32rHTL1iuwjcRkL7wpO107RY/UGNivknwD7chjHVUwDUrtW+w3ApGjodp6SnS9oeffs4yhb5op15
2y93Rl+jAAbRRCWWhi+Y8Ftc5gNkT7IAFEIcJpVbwGtQ1xt32h9ekAgo+LuwJmqxfd/AP2mdtaeJ
OKTX7Me56/ek8Nqj4lF+qsivjafmMNX43t2B5/0kGzV7xq19r/w6acloBc4a+AkNXOv4CdlHAdHF
XJ8gqI6/Sd/NOCIqxraXJq0gncuiiz/tITGNYS2GdXKP9UHN9Zsp1x9uJYHLhIpfzeyQ+tjfsfMw
N5/lncDn/80MIdmlbt9HhgIpxVtenAF3Y9nf+Oybl2C7zrjkoRJ7UjA0Q7y25rCZYGosmBYKKBed
SYVzr1sj6CmzyL+NJUpbp6IOtpp13twvB243gAljqM2lAno2swvgwP96vI3nc/vgcVXmMEvXKpk5
yO+7pAx+Z9+y5YZIA5/2hlqHI3wFfkZJTj8GfSKneP3ybZ7B8e1fpsFqH6HCKEeoPJ7YgrTJBiSS
zjKJ+3XqZijEYFXGB0sb4zer6cCq+vjjb7kzreuIIW1uWngUdT8Wgdn8qz1uZB7Vd+JCkeRQzkhQ
BHFXg21OgxXuASdnhTuJYhtJz4UJy5c3gTn7kz6JXqP8DLhk4b4HR9rZed6vk6qG9dR/tAn+xyg5
xF8SheWj/4cT86Ymwh3sUjfzukHOvRvaAQqclxHA/xuJxBtzvw4dd34ZdgLqL83iW0CqogFiNXiz
tQlehEeRP8cFx2w6Hw5T3a6RaYmhHC0XsGIUCl1d1r5ZVC6YhoQf90Dw/dUHibBJFuEffslXOMSL
MSC3o0V2vmW7QUv44NjYSoOyZZw5dPV6R1Hu7HxqA9mU/JMy7l4QA7OcWe011X3DkmMYXVwJC1pv
xFHflopYbf0VDqTQ4epJOk4prJR2H9JyTftyVwaKQ1pj4sejaYvSaM2GLP038OEVpZsNkirvx2Vk
V3qZ5y97YomoztNHpo1gW12BZIF4+BfCYy7Tdpr896Jht4lpwmrIUKi1NG12ZxEJuOSOaTzqgCnQ
ocILwTNNaNEi5vtLAazGNXTM9o8ZOZ7Ip+rSyqAwIqubvNBWIe7KIuVtOtjGBytwaUiKtTyrvZ3E
0W9DgPgKUMhxAiDyEKfuvKNIK3wVk+22iEkLIfZcjkVClzJDeG30IHRfj9oUmB9r7BTHUsJJeYXS
e/9x6k2vb8Mvllurl8XFL/DjTQuOsFDjMvniurQ62lsnFm4aXICJyCyLOGjblNZ6DPL6efDcNyAv
cR6bvaRNzfhGHcpIvwLOErXgoRSRIh18zj1zq2pfy3SV68frZQU64OCVkfetXblfVwigGJp2mLYg
h8ma7Ox2U4bFUc65PJws3qaZtpCci2Oib86K4vmz893balisTUAkHpTXJFXqzFmOparR8fQhyUZ1
YQXHU4EW42RyTaBSmoD2aXAzWKIsY6TXoJv81HqqCU6OitoBzthKWPLuCKkoTaKGeH04P5OQwhLI
HmEv36FrF4b7auXLZ0lUUirsQccYNuXOKC/+T9gNktRTj+rmatn4ymWRpBZUxmnr8wKYHDmKrckT
yf0v96a3wb9IxhRXp1sltafCQOIKSwnWyebk+9C5yoYWIbKwHoxGPxPZlWHRzpsGYP7KS5eubdmg
5OEC57nxW0A/Q5xecyAPIF3uThJ6C5okNJPvDlp9W1euLQN9tlBsp1CfQIHDVs+KFXJVzMYYDkGx
vKa62EnpTo9pjShCBRopMzW0mwKpihz3ZJXQGi8ytGV3rbS4uCXZ8L1vHMq+36nNHbfYJaNsCS/t
w5uTrOINg+Atz8Yy7s854FKsx7LTl43BlAFXWF6uInKE4GJIiZPu9FhoNjzMMB12caBYYB/CjpCc
eISGeedfmTpwbaW0jeqctN4drAVFJshY/wG7YzbHwdnUTvozmE4S4Mqq3YTBoQvG6BRTzpo1D3Ke
9ohP/F0GDz8JNbpgB+B5fRQcLrwk8mw1JQTfGRJL1P7VpErFLwnI7U8KJPeJBV3v2rx1ivcZLD6Z
+UD0eQX1kCIxlnUFvgei4GDteQUtI4YW0biZnQ+zYAftRL66413NEuY/rEEMC80fsWhDE2ehCke+
r5fINZbl6xLEEuAMcRdSizLhuiK+imp2V4xrmQIdSyab++AgR2CpjxDhBQ+9gmyvyasW8RGiy5zL
4lk9u2Lu0F0lPe8vMU70Q/aQUe0fR1e3Umzo0tip29lBEEYfhwJESYmg3ivvZ1BDcq+fTEFiJTip
rzZc/9YCpDICfdPej5QyY7rQmXnke/HJwtzpeF4GHJHhcN3eEB3r2WPtiHZAjDZU/cFAPr2WVGkt
94Pwu1854we6DkaK1gSc1GiU7hOw4WoI+H63wxBlIN9vqMjyLjqq/kffdA2wmTM9Iv92yiwBlo68
jnCzSEyZvEa9YaU38bYyqsfDwaqHy8LT6VTVkveA3CdtGmK1kMkWuzJj7RTtUZseGkj1XK8LSicB
gzTD3deSg1Le5Nw7I5Vjq3lxoAaRepFmQe3trNYZnkxpq1HpN25S80zm2vK59v4WMyvVpwfVjjYu
HyyEbBw94qGrj2/w1O6Sn3FKxcIi9HbYvu09HNPieIlKwpEPCTPsx8xGYwZbIDU/BJx0MNjQEaMe
aiPJgzBchnQptXtKDCET03BNOQHB3HDkLmCadIs2AQm/0XbqVFvzqtlMHx0BYVFQ7FNBTID4T71x
QnCRtOgZu/ATFaAzj4IYDDoH1Treq2RajLUpdMzsynF8FcXYGuDII3//3vCUEkw1gh/dYdm40wS1
55Rnd8AyDeTjVKoGSoM4khaYaWyn7k65HJ2Mo2n5n8uEJHoZPgjUHRpIaVA2/v/MzkppaorBIWhL
7fDnDOr39k22bpuqaZdsUju/+CGv7b7CJG5Q1kJxHLDxhrXonBEAjn4Hb09UzOTMbxTV0uMVWffd
eTiPVlMzPuUaYNjGc9X6i4Y7yXxbU5QmRhYwp5Id1EpCDM7XmHrZ+7SuxecK8ffZ9VFbrO9gvi1k
AHawF/++Q6Af05Kyp7ZLoxz6uaSiiVVfKN93IvcA5HtmfCglmWr929cBzPS58cdpuNq15vbcpxEW
zQsSPpt07RX5/D2bqzmjsYfUbJ8uaGbkXiK9ItzY2uQDbmGCD9Ah8C31bsRMtkaCKt9feCTH7Ihx
xMRaur6Rqcbf4O8VVLsee9zrarA+PjRBmJwzOaluHT4qAkvKoD3TuK888MRHmA+sUTQhiOKhVn56
ovM4yReykzyA6GOW+eZdXC53sGQGyQEHgh0S3MdlzAKl1yfhwiWC0A5547Lus1jPlKf/ICV0KJLX
Yp7YdKxRDZX9HY5JohRy3QRXAjscFyyM0U0T7xHMUskRZL43jkUeWMOJ/bI5uz2//EgTiNfMfAWT
yY2yITlC4y+c47dpTiVYZXrkrKIbkUYOiV3iEbF6s3Z0WYfBfOKJnIfjIc/41+pPbv5Lr6k0tsqM
1/0fbVKJ/strf0R1fnBvCPPy4c8PodAus3teKa7fZYJhdqTB7J2KaMUqrTFQp1BxTS7CQrIKsp8r
5waxHmbCYkdPEt7QPFaUKjDUHm2YmwlE1edB4vF1HCrf5j83vcHJIuHuzLS2j8X8u2EpO7MwA1xY
LjUNTZz9TrjKEk2LA97sXwqXUJN9Rnw7Yo1AP11uTS38kaBIZDwp92Z6qWbu+jrQTLImj8DAR8X6
lgVVu5gMTTecEmWT6Aaii2wB5+l+hXK5SsKVcrqVzkEJIv6zk5EcXcqWfDVl/fMsfeWxwACaCFoH
67FmMzGrCFdaO3eWO+jTu10W+ibW6jYuvQTnr2R7DDBuVColtCJf0IcGm1R4lT/POAVx11NkB302
LHyVuyrg8+iq94EcVFeUzII+3xvOlyssm6IDAxOe9O0CTBvuym6w6O5C3DY4n74wClF3WgU4w1R+
MaEr5Ih7jGbXXJdH7XG83hR9FdbL8AJPP9jYL6V0j5PjQkCn4az2QIUxanjQNMJxgDt9e921Tzfc
fTLlyalU+4MGXjPiJWqKYEc/XEC1RhzYPdgKUr/KuCMeaYfHNS32ieIqjnI7OZgPKiKhdP0cuemN
eR4BBdpEA7zommQ/ipsyTF7QT2ppG1yHvSwcNrkUaKprftuM0Ei9kfTu2yGEKcIw23HhvhTUfJ95
i7aOl4/07ka5ePyH//aANSdq870Yu3OLed7G0eQ7DX26Lv0YMylcM9y6WraU+eKalqcJ3q4c3cZ3
+1dOa6KMsFvJSkD0IeAOUHhgI27YaAOmlMpE3u5KCYKdwhsMsWXlVWRk0pxWl3aI1OHlFMTLRx2C
qkPiTvXx7mtIiGKd8vROtqPk4oXe7hekko9dL54TvpUaItI+ptMjlg7xIKOtw9Lq6ADvAdih+xVT
2yGn4lS40PLPkp5rcsVTW/NpJXHtTF++mmU9x3YQSI5AZ5IPQAR2SaIWKj715b3RVmd+0v7DVuYt
WyN4Ft5DtXnB8IMhRVzyhNmEKnit+4sceB0Y3QQ3nFo3aYYew7n3TQVNbFaAMdtC3BEiPHPKoS2g
lovdcxErq1ba+e6BfJuoJX61BvBnVjKn0mwR+2UC73hnO/eMVzEoJU0Unxp7bfewXqPAtleEa4ET
duF02VB4AgmyTcWptcvdci5iP23PGB5AANcbujGpjdTzuLcVJvbSwOTU78nOOWFMmZNVoouJP3nQ
Gi62JRXcpD7gm4/BAA2/BtL2FtktE1shq7LrPPW0guxxS/RfIo1vAMrwCx0NZpC2lEJDwRLvW30f
Dy5R70ON7XTmbrijeO2LgzH3SYqBDXZQYuA0ea0ed7Y/xmSpnTWpF2GpMDe8e9lQ/u99zPYZSldu
oEmD59VL88QvRH6W/NrbzYLRdL60rQkxq0obLk3RG3+lbetF57mpjv2q+J2pHiQLxFiAe+kxSrEu
Gke4w7G5UhhhJ0dRYQCt28kOFZZlYr6Fkxaw6OrqIjmQTb4uu+4sONM6qhvU2i7szWpAzYqpIWzH
utcP7apkOSp9pOpvWWjMaC/+UCo++M4PGtqUiER5fEBBCuhlG1ykSdUDz0qnZMQtGyFRDTCvLl4n
sj+m9f5JnNbkw394T9PMV0XDN+B9InXhJkJMgsgSLBIDkasPs3IJR10E2Bb2e0NlAr5kae6UO3yL
W/BClbjda5U2gxzbpq3glNg6Fjvjpbo/POtq+u6qDzS+jMzaDGhQ70WWov5mIJsyD4oah7u2kKXN
D3nEyMVcGRdlHdWeBy+w3lXUYnmPeQ2baFQi4uHPXgzl4ACQwCXOh/xl1XsXbUhitVhnrx+sP23i
Q1n6z1EOkHZICLDdXSNpOkipkkT7Yv8y194kH6RGxOYNzmpOdkgHHzi187m2olsuVmfozPz9gRZ+
hfQoEMtW3p4kb/z6EGE0BDDUlty/oOoWVvi6hq97qQH4Niul62ptnOvVj4fPEH/YpZR/d1iXvfCD
P6XhB6aFt1dS47j9BI5NTLsqkrKr+G59yQsF7nUE7ip/+WHP9eLwCIhY3697tQBoEmxuXTZwhEgG
4Pmam1zOlmAXnUACgIuXgwjLg/Kdfnf2o86lOdvIGNButTBTbkXa0PD68JuVxI2QKhFwUhzcGgnz
J/lwg9jxvUxMdoLvXvyWYbO+sGhC0xbdIPhVxHdhc/rbgCaN2R4zEx4BqbAjCUgVTdrEBQjjqjlq
/q09XdU2SxipHmkc3oBSwzuTNmhPMzLH2HHFxhaMubji82uD2OW0jLsBWKe27n/o09UMyquqolY+
jrF/tFP0vwiV+bYfrUjnPAr+TltAqKVrQ45owS+W3pQ44zEY9rPErR9wotn0kcqczdD5bM6XbM0B
miU0ZuQ0fi+66YkdV/4Ga490MeHZE+69R1eblHmfyre7bsL0U7zwY7T8fqCl/R13LM0eWgaAzjHq
g3+IjYeE6LKzMBv2Dru0NGTT7ioqziP5GnD3U3MG9jvXnf7nCv6KXqXu8T3DLmCKmHLMth2N2AjY
7Gzqeq/GcbTcJojT9fijh7c7z7V//9e7zuXMit8r+7cnArKVVu1PVjYRwQK8GdXatspaYqQuywuu
AAJB6LwUCRpPQZTWTsij2Jb/FAgKH4nOh6ryE7IewlMVRnxPpClbSQNwhNRNWMbE2hHQYGaCjhV2
x8ellecnYZU7r7ANaaJFpPGJEK6p/uKP1B0x+SaJKmCOQmeqYxkussrgzVppoTlN/AZ0KH03YKu4
rPH4TDrdWa/UegSJAGQZ5lwOzD92gtepz86KpN+N96QDi32jA5AZegmlYn+cZIYuEYvm9zp5ZNeZ
W/5hLszmxig/paR3IwDjLCz0Iiv4QtbtBpBfoATIs7Ll9gQJ6fihCkI0ZA/YqNCtoFnUDVKiaWJA
N+0EHrGqbv3X3M827aG3ikh7oV2YfHBpPJQ8qpVdYYnVJu6whuKgVu6mm0EKwn6WwNen4cnK0V1j
Ny8+BkToId5e7BWRUze79XzeoXdy6cEHSBTADsFwYny3kIMOPNKgymZos6K9Go4KomY3jGM4L5e5
UKR0SlAYaJ+VD7udZxXrZg2zUdaVTKdGGW26eROhfgbhrp88eoPW5gYHcMSqbEK1gJiXRHVepgD6
jqEq9h5lbLjVvWjBqvNSnprVOx17zL7LLe5Wu44rywa8RqTiSTBLJDfFPiODxjaWMCv079Bj726z
c+RR+2D7JS7y/WXiqmLAuj8WxWtOvMGFnjySHvzEAqs5AB/jsW+cTL8ualCmPzInPzp5S4dZS75L
EQB9nb9E70zBJepal2ibUszer3vfs4KPCrbBpNPyHaKKloi3K0rgrukyaVBX0lwXnPNDt4mf141+
YFzSY7kXdfELpNFS0WgizBJj6kgCznph0CIqftZkFxXtBMfqJl5r3ibx78y1GSfadGpIQVYwLCxk
8wJJnUvm2/5dpqHAh58Obniu2vG5UrekhtPdP3naTbBI4e3txRJuGOXscVHQEEBmOz3nNGUqToH9
U4fT9Z8fbWszXnxBl+grua7cZlsYDdpvKK/n8Zqcr5KKTtI7BmIuEPq/tYqg8eo2+DpHyfcg8Lu+
2vcqnM6+6YngsTp2LLF1q0YfI9dNMRdqKjta9/OfpWhs/H7b7Ip94KrqCdNQVT4esrerxjKY+w19
5GfcVl6gThks6qmPjrsC8P6rGgoA2SCLnqzE9ZcmVM4nV3ou4kPbrhS1l9mRfQlwmMsy+NDmrTji
Y/QPclDx6OeQuM6i96dSV/eEuWbzeiw9emhwX+Qo1lw2iwhzmfh3o9LNeKAsGe/TfhjQijstvI5R
TlR7TKTOIfr54u3JkoRRkkUm9AaMnW74748fWfGEELmMP2x0AX4IMS6BrKwAeNw/jPx4c1XdUkVl
Qfhfwilh7wmOGUdfkQI27HknoN2Eze0xAKAlxRbpPnmwLssSMjEd59a0q7OhNPX4UK6mWzWfgUly
3CTKYOGqrZBM2D3zHERc63SVKUvOyiGnntDQ2Xq6S4HBF+/Yt47RqX+FBMgZxxivvL2hQssEvzHk
Y59NKOB3/30t68LvbGSg4dLWEtPGNExPydtNBkcZ96zAKIta8GuQH6MDIdeQd7yPJvZyTmbwmyUq
jKI94N6E4LyJFXhW2gGYP5EzK37leGUyc6TnXpg1LErTq1RaeLy6Y8yYHRdJQgxiRZA8oxaQ0bHn
/6439FF6B2XkXRZUa0LLJx7gtqDRfY8EG9NbVPcgK4KnuQRFdITEUtf9n8xz5A6L+ncUEDrB2fjC
Uabc55bNINhQE9vuNJvgDTbtCVmdiFxyBqN8XyxH1/Tr6lQvcuM6gir7wrlijCjbk1QX34rjwCKJ
SU087BgnM5cQ9gawQsq27Uk3T0UbjKVy50WCErw/h4QMS/ij3VCESEqtjO1AeCBBrhIOrCxHHUrs
Uhm6Y8DABxKrX+W45DzPyxFvTpxNBJHHAU1/ruxWR9wgnAC+QBShnIM0aAolBOGjYftTdFXHYl7c
UnGQzcoSIaDFQxl7ChloWaMPM7i+K+qnzyFU7f53PJs9nd8N5RfL+UruLmK00GMO6Xe/+h2915wm
fA6dXu2LG5TqIEDlowqOMdlbHBOrZzA2HRvt8pODce/eGbbvs3xntsxVY1H9A7VuEYEW9esE5JTN
0870Ly292hJxgbA0B2sDgAXbofevD3E6mzuSmySKyosU78GRmymM0yQN1OEEWXw+e1sEgYHke3aA
mq5iMC+HV4+McqR6AT53HphNxrCwLJbpgkx2+vI20pBuKgT/irHrotrfgQsROge2322U2TG/RvNw
3pQPn140AdtYw2yG+Y55dS8/arqHjZXuRUQuNydDsaB4cFoqdnahJRvl6JWwCbUfi/CrKE+W+Q2z
qQs/lM+u5fGSWPfiRtaert7w0BzCfdAMeTlRhowdOeytHsiJvzLSx5SZB5Aou32gov01Hwkc0KL0
OATtMh+OFKrM7fKK8sR4r6eK/OEIao2/0jzjQ1+Off7N0FylMm7qYm+kHZmxEgMHCo/gkJno/L2o
1SajxE1g0kiD4g9QcVsS3bgW6XhjZBlOoGFJJ+2vP5iXg39XgO5XJjSp+UzuckY7g8GhsjPwXzmr
3A2TeFEL0nEvoI98ojaaHBxMjlAPg3eV8g7zzdCBRzUhoBUVT5sERD8HVZA40a9B6tFFGmB6qRXI
jlcZTNoodQTO06Ank6Z25uQCTICJXN1ZQNY6A7o0kbbZCCh/7yXboAicciWmwS1UqXsrmXhtmuL1
yPvd5NwMO6cNl+urOdMTX75gAkSttUVU8FX0oJ0SbCboKXoUlNy92WWyOcW7fK9dtwyt9OTUHp+P
DZ8YKXA2d99JvYO59iS60cENSrDSV/5Dbl04j9+zSHu9B2djNnXt+WQ78ELwnnGlcxtZtWziUe/N
Ae7lCJv/G8omoNYmp7kpX9kzfUxGHp0lheSjF6+SnnUOhY7c8fwLW0kNj3iKdyeTfN/+wFOBMQTF
DvfZ8GqOOdbJjCVpYZZFKKB6jfIholGLsdKXM02aNAFDj0JTmkls68g/j7Wqx7Sv3FCbojig5q7h
SO//zyTpUhphWqidCYgiAcOdj5U2cxQyqlnGxmKPNfIhVQdMWtAb2mgE0rDemQEBgjn3I3+eRB/7
Kfmgk3+QxnxUllPmHvXhVzTRhYM7lP45ttWvlaQ+Tv803qjY+YnLQXxjTfH5f6GHXeQeRACfgDtv
/CDnplH0rMcJXTOX1QINy2ZTTXeZlPtT7LLjo5EWlvcUl/LGskOsB8NtXCZbTTtjC+8MN62oxkag
tuVObII/ZP/ojOt+GTvaqU5h+REzvfu9ADrv6coCnHZARj/G69+STnGAwfrVsxdWnbV4knuVJVfC
ol1rnaHV2yhWmkWIh80dw7lox/9BRtz+fksO3a23pYgO97XYrsDb/X5G6rYkQ51IDgb35hF5DdOq
//NpPnMARWKqgmLvVqF//mF5llwNA1bEGnq93yQD6faFLcPXIBaKRxI6HP9boSWH7SefZ8ZAuEyI
ITFdBAZN8vBy6M0Z6YmdA6R1g8NXnbwiHmNHNP3pndJRx/5T9DmVCDYOYggbEEYQbHRIKOj9aBBF
C5YfoQVel1F6FN3XgOOVc2BgXHndBEuyrGhTK0pVQAGHN3XTLqCQR75pdVLHgVHWHjvZGYOq31sP
VWiqgrrnm6C0a05tr+XzBXTxzYJvEgmOG4ToVewEGvzpsCxos8bFhRSTAh6qQGt3yuYNFkhQczWt
C9vCHb/+EVx01daPNpHtRwb3wTqTlXy7r5Cg1VAOEcGRSJTfpSKFuqwKNovjmt72um0sEJF6J3ic
tsj+tSpV2b6yAeYJXImnmV08/r7yrW4HmIjRjvuwBoVUiUb0Z6F+WpVsgTi6WTC7YPfOuMjUfeyz
WoY4QYipvPDrkfApgCNeFoGdJPSfAHZVh1Y6xNHEAKyTPHZrIerrnpy5TpP5/JPwzn8NO3AWoH1+
T8hoFyt1LOev2eGnYQcYmYb/nUHR2bCYTSPp+ikJ9rlGJQ9EXIqquqoVOz+sWsF+oIMR9OCLrmx5
NmIu4OBA5xEariw72atGtHwwiNVu4B+tt2QO3YZKSk721qciCMydrMB5BpbRsDxNe5Bnrr6UHYoZ
fb9dz6Gh0qkC+/Jr6iPZcXZKCGr3hIabpl+YSbL4DF+388OKincJ9RqnMh2gg8xlaG4wzE8F75R2
n5wV/KEMtlNaGpglANSr3lRWRmL1yHhJFVadxU0OqA5JHQmoabswKGp7X0k0uHlo1EVtKB4YQ+R6
E4Uj9gWwMIZMTzPAM6p1mxoFrGXINDR8rBB2SUYKZQwyLXLrd2276UuPDdwP5oyTa0qO4TotUFC+
6sq77JKn4bjn5LPb0T+BRfLru1ZOHGTKHDAPZjSWyG6LKPUy1vmdpfKz4qoNVInxaGSAjrYkc4Cc
OFnwO8uyK8Gh1VmHf4Hg83oms+/QFERCig+vmrJnnHM9KhiR7eBR4kFa2ftigsoxul4wCNMIkvAI
DSRcf171Hx6U2QM4h6dh//DtnD20mbq3KKt3JNWGgpeu7ytuYCvfDrHtPhW+LRMsysrazYonZlKv
+4gn8zfg0l2KvbPRPIaCvmOKyv86AF8Bc/xSNzYdz2O7UeJLCnDbWKLrRs1vnOPHoqPIcZGsk/BI
7YdfGT/+4M209UIuowM887shGd4IhITFk7v8Vgj16Z61jA7VpW+XV+zoQUI+THjsjQeEL0J5Ir7U
wKej7QT4pK0Bl0XAd/mBxtfAE1EAC+7dkc2fMaXw5bwi9+POheBJs/UwebbJ8Cv84qk6Pf/YhbEv
QZ3Ym1We4wCxYj71RUHGKM26YiRlmC3JzN5qu5bmvIuVaNubFvurXAPDMbqoQlB6lPRFPsnOMQCS
dBmLlm53dPrsUq3NT1VulLfer7V5Lb4CnMyyms/7VJHTWKxyILOLrZ/B0gLSXCldyO6gzED++LO1
8S7VsOCLtPzKNHpApSlXA+YzFI6HNZRQVV7B1ohwREn5Fef+7BgB241m9LPirI2M9q/7urQW8BMC
gwAks7DPT+cVp9uAGM8zYXOpL6XE4BVq96ckljjFDzhZhXY13Y93x3lnMpSvW8yDkpU3ULV1YXT5
dQbDWYyun091v00ec60saUIvBXd/WfuNTYLoIzwtw2ovehgiM7HqqSv9PYb3hTwqRx1ubZSJ1ylX
Wel+lxW9QS6ZGfM/Nz5oq2oPBOweFWfV/8wqSCTpxKBQ0QNNQ8B5UY/+bxpApjF67sTOyCyTEaXw
52nN2pogBz4V8yn+hNgf+xg23Mn9iKWAq+Ht8U6PctXLxD9U6V7XWPT9TgTnfsNXutOQSyy6zm/c
T0TYsvCkN7jeYjTgFE4zzoh+jbCBaIsZ3y84DPwSx/RjhfRNF6XFA1/srLLl25jEtlrsqdHPtf2Y
DO1Xd6TkPLb+XTCG2Il0RB2asSGdKNvk0DBRI1giRqMtothe3iImTvJgkqKm0Kq7gfRw4JhqRh7i
jVeqUSns1m33P1QirBRsFEmzUpPJWlanEaziXBROxJoR1pKnfYgzrAeYX/8ICwliocQ7b1TIWRFU
QkurdgD89Ou4PKOv+DIPeXzwTqSWo9R3hYdiDLTnVd+f81VYokUrglCDivWyaE3XSIMmzKWgLgsc
LCps2DEMVdh8qTz1FgtCHFYPspv8+9NziFEjhKkQfA6zkjKTC6rHtBJq2vz3DT11TyV/nTr1Yemo
FqNidr02hhEcYje3LZa7yj/LgQVKcvhJPZPQ+vRwmP0VBPJV3DbsUwotDSZOJM/sJpjV/x2HqXMq
S6kype657Wu3TiG8s6nJ+um70MLFXhyxbWzM6/AJ8fASuKEDouc74rw8URyYVVLFMi+9gWUagork
QOiOM61So+Ko1KJ3hQIqBmE8ye4dp2BsyQwOLA7rGtmUxJzJuyffT35xSadeuSf8GW3cEf950sQm
mrr9357WeE8tpygAYEXgNkxmSbIVEwflJp4UHWy+bCIj+2QnZUlLSsI3CsjCfJj1ic+KpQaiYFyI
fACi2FMFEQ4H1hiIUckDO+AxpNZIjahY9rVNc0aT3Sl2g2F64WJjqjCxH4vnvQ5CQQ1iXOIvWZLI
rOR9tibn3gIpaAmAIFHEupObRobioP7eK/ksAUrqRpEwtR/rGhZlAP8+VtAdSulsJW0dqAvYvkdg
0dpCnN2eVZlVa099TGrGDa03Dreetl1By1ITM3gsJXKZViO1Q7m8nhHfpBMKTjx/KvWKz90MO8Oz
YXecNzC8AKmsyWavwQy5YHO7Yinj+uGeZAm4G7Ky1JpdLfa5YRSv1z3GTjSBPDwUMacPuqzSm1m7
SzY0Y3jMMosAEA9tqyNI9De5yQyhicf8hMzxGsRDGClbcv/8vn0bghc7hMvfr2UGfiDO/Oc+ly8q
SrsuZju/ZTtQcZBIuyTz8Q99vg9mmU+w+0oF7VeIM16QeFt9k1M1COGk+fW0CyZrzAw5T/hBd/+4
6rcLbxDhNT+3lML+1fcPeY39PqH3SrM4Fvmz9UYn/fmeOIUmK90T88eP37KV3XnEa5WEvq2Uzxwe
B5Hhoe2g/aq73op6xNci/Ywfh9g52g/l3iOq6+TieeidXb3xSqihyEmS0w7T8Zm7HToI675oxbPp
pzxr4Zy/ZebC5vTLLL5nu4Stnj75Go1a31s2iM1DZSyLvPZbtZ3Lfl6HLibb7k7dGklo2OCZ/y2z
q0Ibec2E3kcZRaZvOfuVey8upEqLCIp/kpb5s/STCAETyBaFUfePeyL33a4W+rQHYVGhFT8XjWa0
QsM3IOtTvhAfJQAxe4iWor+4A/zGFE7eTktO8wYUz2CmXxbG6cS6nhIG3GOuqkqtJ8I5RNy/rtnH
aFRb3xy3t/huR5hlQzGc77YhcGUsSEX7BhFkNMc6mVgdDW4NjeLJSferzXoz8mwdx+3c2mryBPdF
PjtgtCQM3MPPvyFFb8MIA/5ARCGvxwMX5GAbHAKKEegPRiakaPkL1Cc2i/OZaVyGod0y3YAi+S/q
ZZTV964kR2akyWO9/qaZMWt8M8kDPV2qHTFaprO/aClxypzOX28Tc/0+KpGGn7ucI6CriSxInEOc
S1JYl5YDdmu7FTFIE85MclMzyy6oynB/vmlxdYnxv+QhKD2jNJQN0Sq40aDWNJkl5USHrKQCPsBb
gX/FLVxza9evh+eZ1jCwzCNIusPoIBSabmKj0mrHQiqIIoxOZVyYOwccSTv5EWBQ/05q4sxBa9cP
Kr+/YQnmIhWXaILQb+zRbXTHiSLaZ0oW0MAkS/+l3jglr2SdwYXomqMxnh5GnqhVV01QsACpoiIs
lXtOcyu8osXDnbWmR7UmXrbIf8Bhbg15mMrHxLDGM61MNM6U570jGsee/hYBNURZIqHTt3nnFTZF
8n3O+jPK0/4CHqZus7PartMHpnIWqxHcOf/ZS3bIzM9RaYK8wLVF88CgDFoIsd0oT7zBSibb41hS
yNkooSRnc/rObxv6PxkJqlrWJUUlfkCX5BGlvpOlRdV0MFMsqoVF3zOQ2vGuv9iKY93iqGsyfoZl
HqX8u/AKxqi11kIGAcjC8L3izLoqIiGMe51TC3UPR629eQU1FnSn8zeEUkO/n6GVL/Aw1v7c4yP0
xGSEgbb6z35cUaVsVzmcbJDRLd3L0Cf41CLL/oZHybni33q2z+cooD74qxKnfNnbptztM30aISGZ
SaPFSQ9QfvrG/sdqMLQuK7qfklVRolpFaFv/rKKXYgOUIvB2aaeJv6BeiDlkjJys/cb6AHJD4Rzp
mpyA2iH/CVK/orLqu4KxNzkMm9yZoTpBE5kFV98JmokJYQa3lZU5znKzZSV6l90qKzxgUmI4W0HZ
aDJpqHQJDQfT9rzjXU+4jG4roVfluXehQcSSEjgY5LZF36NZmSRUjhZrNqZkvWLs+7I/5iFGP5Mz
EeoaMZpnNhj+xCfPnu+o+XC90KU3auvOq36QXvqm/3N5hJeOOhH8iAFYbghs6nhm3UDA38ZspYX8
LwLKoflJYSVXuojmNUVIQsdrJxqxKBDcGliLMyh+INxvIv8lQWBBYKtqlxemTzo8lBAb2lRfu5bZ
oKtZlos/+BQ/WdXsUwf8vGwQos82l8I1E4YMtlQm9wqGRWuxTTnaA51/mgiyYBc4RcdMMqpkHgB3
JcND4+m2Pm4HQiGJ80a90h1laMv8mgiNZfaOQCv5wg8zWJT8Ey3pt4KEnSOEZnrafZ/c+4eHhRv7
ESIZC+0lJaAGE1zAR8Lx65XDvAPuES0oN12quCmmZEnJdlai5UV+Fbl+MchlCdF+X47AVdymhFWW
r9TPD/CraTQKJgBH+9DSu9QJiiTEac8qWnJQA3ff2YWSeDBP1Kt0SlXgTIdcyTjuR+RHyLQfyC35
aXz6ArJ2V7by0WonaJKoPPiEQUIU7873bMK4MU+X2MAjAGVf6ZDuFZv4gfZPubD6baTbjoGtE/pb
mV/3Cm35WVeuVEMx5maaqxNZrVEcKS99XlSWTpyNcqQozImLn7M7wwjxjpDAyi0TTpMrABSWuxIJ
4IW1w5V1m4GdthdlGSBaJ/ovckNvnJnNMBj2SzqHkgZO/gwXOLqDpMMGZ1E1v05aqdojOGI2I/mB
mdKVuWFk7JeC876lyBDPQAzv79SKu0NdIecYKvEMaXPcx6YwIR6kQc/jQlhv067K68mp6B2KZsut
35QoZeZcakyAlJnHYWKAhoi1mcQ9PmpgoUn4WhlIAkYJWKPx0ckqsRai2QvHM99PPkO0VhyQ/p1U
fcHRGiS1u9VbB45HKqnCjzsROMc1jTW6QOe/Y2GCKZjOOSMP6pZZkd+3/7XaGmDQTlpX778blsoM
TSyEQVDYgjY9T33Umbu5zp8/qBuhV+OSX/ByCkejut+gQmnmyQ7prFPjQOjPB9Ntz0bKDw3dT7wC
LeEIDal2LqXODtLhB5tvjKZaKQ6kknPdRpXjqe7YlUsgcUZGz56bgdzNq76oGOakwmV/lOBr5F4c
jia4WbgmJaqqn4S6/byMDBmHsnWQRYPEbgcZZR+etq6zNQ/lY7bwIOSUtZ9oYbSCbUPBV6tdTY1s
40FBOw6whK25nvm0KIvKdklFXvFWPj3us94nDTn3RtMXqYHabrUhY0l1r923orKGL0GLmQmU85pP
JY1L881KSuMHKCwqCk4AFw5xC4UH2T6+PCFRGrz1o4ZU4ZvbwnUMxDg0P/PIPZcteB1PATXAS3Jt
5ByIQgEWGlMiPBr6KodDsK3JKDcwscYobCeWNjCu7ussbdNvga/M+Beu4yV/qG8IEWMX3uLnTpp1
8vJrgFMia8+MKCZOqGD+bZ/aAFXnskaBAvmGkyPb3DbEtYVMqKPrYyF9Ms3tYXu/u2vJKvj60epq
GbNoOhHW1YW9xDh+80rYzinEMvIGj2COEnDTx+Pun9LRKPtVD1C8rY84LdxzIE512cN/OsvHFETI
NFc1pBG854La/m4Bb5CQ0rIMoh2eDzXLVj3DgX7z3y/cFBKcWTDHywGjRZDVnMDSKgmKRETnX+6i
aZZKo42ZyM60nzTp2WWlZk0L7ayKgUMeEbTU2rzDQV8B8KTFI6Qfe+tIqIKtq1vEh1iZU8Wsvrlp
/J+kNAo6zlVDFBjuSGDX8A3/Dtmo1cfuA85rqTY+skfJ7tOvqaUmcS+gQEBvx6sQyPjbByBGMTaB
r2YaMEWnKwQml/NCmITq+GM3iQnyNKjcknG3kJl/I+/ouA7sTdi4wLBmvm7x1YBMB4Yo7Ds+OgGh
TrctUxa3p0KKDoLUmpbj0ef/1vB6Cs8Xx9azZqL4KQsBoxvChULj46odCOKLosuuk1R09Ew3vuW0
k+7EbJn/fGGFC4+yFxTQqUWqjOkExo5h7eXnEPaHRhmlpPzmJT3/lzpOMtFB3Yy1eNrKuq6xP/4L
YLRVTJhOik34dMh3692L+sXd+ArV7ZnkKQGFs4X3xtj5ieNxK4HybLgutHFQfXcQycm1d1XMMSt6
2OH/S85VpRx9qzqS8sNilQ2N4AsLD8ZUw2kf1Mx1PsF2mr5QzHTUp9DL3X15opplu/pkhoJifGn3
QxdenqDU9Fcq/8KUx9OD1aCbf8dTO0gAOmc6LZ3U8cmLQ5KHEC4N7DNJePVvcFtqzUomQMMO0COq
P6yhKROrFQNcwxN/gDB/pyWrZz4EMywFZ4/FxW9W9VRuhTKKbq3CBCMUcIyASheFucv/EcrEFpW8
nGrS9UVLpcpQMb3HzECo4iqNnnP9yemBfT6zVEW9jentclTxcqpCS08404QZm/+Jtw5vplF6j+Pq
TGntQCdyn7hwbeY4CKVXqbp4b0qNbegWVixMkcMvSZgL11i4fLIZj5LnpJrjkx8PHEa3jNY8g7t7
Ohea05Wxr1y0UclMPuJouQ0+P/5h5f5Lxp0Gl4LvvVpU38wVPSFZnGIZfEd9GOkHDI2vsCUN89DA
6fVfkTGn0o140+nqBOdwS92qB9fpVl2LfA7s2HJgjBhFFHb9fW9mtieM9j4skWomGzpuXOkRau0V
MPmVGE1PkraxcfxI54x22cq2mJPrx8SzY2K+BzyquFgoW1PxQRCQ3em1lvK6VaC5+wbHyzKRu3pQ
wqNvPgQiLY0omTREEN36urjBx5iLUC4LgwXc3nYIhzdTW8GT3Z/pstmz/skFSgXM48Ll45fE7aln
SD5wYT5kptcZ06qmTKpJ0BLPMGoN7kFw2YkOFdsxe6IE5vUHY5pQMe68UvJf6l79QUdhyGndP9Lv
7CoX7CgyerxUbJUgBY4kg/z4hwIrcJjqv/9oxLKVH2pbORNIICTSF4mblyz/zMfDmdCyAAnrj7ih
YPIwhGJfODxZ4xaex3Nf2x6fQV1BbxBMl5h+lauoF4u6tLUpuBJpjfEMX+RpEUx9+76dOaHH8I1i
JtVYcQB1zjv3/95h2OQrmEEg1e/tTX3SFgMESBu4Av0vXCPt2W+lWEZlH7SQ1Mctd/LjQ6a+K4h3
EyGr96MLOdj9bV73z7giYDsLKihIBtPsUOC7wq7iMqU0qf/S6FUK7aompI9FuuyZ/XPFmPYP5T5c
oOjAPHRp9XHqNxAKiuFscBnk4Jm4eqjjsPpZYz7L1ArShZ3Ts7hJb7usrIeShHcZcDFc9APAB9Ct
6SprZ30DyFs0tKufabL3Z25o+3BfeXHCXNwb9KkApOh3mMVOul1b1S7vnJMLpdbZPZ5IqTVASUFw
YnAudBOG90OEP7xi5qznV9cSN3Sb6tXZAB5HnprXeRqrkwS363ol71dc3ofskOkUTOigwTNuZOU1
TqY5VyrAVPrPNUlql+rVULCUpPP1YCtOb8iJzCFBu8fCgUyKsIVzrT2W+RVZAG1zf0OTUeUwvt1y
ZosEqmSgfN6A/4TWNCHclj3Kve39CHfJBOEPs4mu9NCWPtTE4HcklJn1jnV8srf0RX8iDtMk58R8
gs48q5kwPj7y+4wkV77P++G1rE0xsIwIKWHoZolGqTm9ZUaVzJc8xMTnNuk1Q0IS4BNRBiQjkfPA
Hp5/G4TXdx1JRAEjFAuHpExepr93DSD9XGQRdeuX26gYua1qid8DDXG8k6znj9fM2H9Vx9e91BsX
n8s3zz8XFEC3jxK6slyb3SLPmryEggdDeX8NXMxzn/XeVt/2ZDUsKW3te59snjtMdleX0HRezBvB
B4MFjimEt1JEbzLea9s0ij6LjP/wbqILD5YvgxUlvICB3ZZZZc4Wo0cyXuiKgHhwJK36uPfZKNoi
R+w78l0cF2qGmTSCSgs8MvjZSZ3LxOEWxxEu8doLrdpFV/RPcK6PxME2Bdmi/S88I0DRTx5gvEen
3/lZVVBw+MYFOHUf7Q4BE086jFl4LbkEFlQVi5MpKavHPG1qy/x8QZR1W7Uk9ud+WpYZ1v54T0Gc
+szKIJoBeBWSVve19NKKj0ebP5EUmGtwzfWoIB4VDmORsyI+TQRYYkFVHrMjN466lSORDvzA1bUV
lftkVvY1YGlSqapzwvEyXTBeToUrM+I+CDZq/QXFDd4jfZpw9UAhmIg+ZlyoQCVSANWrWrpL2vsX
APA7xEzCtu2LM1jEOmHWJpYgPh7dD8cI61VMb1nC/5tjS6qUlfZTzaG8yN97/JRHtI1lt+uaaGFd
TgFYXpbCMq+9LRKHCgqRUa3guZ1OMB3SM0EKvWmRh8X/zy6yWRfQVb6jREduW26ugZZEJXKge8RU
ebVkgMkBLOCH9T7pOzFafiYFHy28dZ12y/fyMPCRV+YHFTE+C7jXxZ53VBlyXp5+EUPtye+EJjcd
Bf6/Zpc8R04QAGaFAQ53omxiUhdLFuSnX6qdFJRDDC2A/bZc0R8D6PNtirNfmG+MX2p7F/X0ZhXv
INqZY8lb5360ObQ94BHtgwEM773U6VyLbnJS3zo2VIcGxWQgRR8Rb1S9qdMQgl6LL+mgc6BLiPV4
d5h4+rnXQ2JKkbvvWNjxGOYBXHhhpju8/s5HbVbUl6qz+Nb8w601vAmXBLD1vvuPErZEeidN5Mp1
Td1GhPsutGifekncuCCiWzOkhk5r4KpuyaKDo7X+vcYq5B1Z/jLqiQzPpbocbF7dN9w2DVqbUJ6L
NDWeOZb5ApxDSeUYIdRA/9I6DWMVWb6+BuaQZkwJH5gNoGXxUKzrlvJ3ZRk9x9zGfi0UHRZ6Z0Zr
MLNLmxTCqyp1Uookd+Y1v3JqH4bIymLMgYdETr1a+d9aYGC88i4MT//pBT3QvGAB/z8Zc9IkA2Nn
y0G00OtCSeDd3S7I1/vT5sk2sEShWf+ceM3ofBpJU5MpLsTjf7UXtNoWvdnGn2QkW5dxZUb0e+AN
z/nhtYZqNJN5Q8xIkQy1W0XLDSCJQSA+uWr5DG6RFQoTtiyPeKPgTirs2pFuwZ4IGW8LTYi1cV5n
sBK+oyazEiPRG4c0iBGJ5twp594HEcRDaA5AsKUUvOkvty+fyJpimPrLq0qYxff30ugRYmNUocSv
z7yVVJJax30t0MGHIm+4EX7Ho6Mfpw5uXlnkFo7NsdSdVDM5yw2daSDZ1nZuxM40iLbAofV4eMib
ib5ypvlo6Z0MrSS7lNICwQS/I8PpP9UU/FLE1PkrzWaZCR4I4/T6AfKN6xj0C7gMaYniLL0VjD5E
r8lHWKGAaWOA5W16IZH8F7jgDMQw0FeSWAx6S0hbAy694EYHpn4/y/GKElkWn2hvrvRhDzMqCAQM
xlL+laVKB90MHj5G/gMrVzgtpBVIMtPQWGQQRWuEXyyorgBHWPiqW6G4t2u3jnws4M5sbfD1tCdX
qs7iUs2ymlosvqrqAnqhJgYTTN15iBC6kdMIfT6nz2+Oqae8zzqLpCEF99839AI0Z27SRCmaLzgM
AiQBvGJ545rcKbc67N4r7cIRTxHXKD5D5/MRA6bPyYzP8ZPR+D2tt3AgS//TZoaonM3nZATuE79m
FOVchXc9+8S3bPbJQQqdoBIc1dsmfVEV/lPqOgYKU6T8ZwALi+hrgry/9uMf7G0xtB/TjPXKIdrm
TLT9fgB4XO8Q0a5kPKOVQ9n6VoTL5OsxUJmcASLsOFdgMD59ri218XMTKq0xgUidr/G+fWFpMOyi
1vF8fSDkWvjC1YKCqeGE7eceO4di78T0EhJ3qkKFziX+u+1XeJ2Dd+M29+yzGtv7/cap8xK4Dy0O
f2qQm/DDNLlAaNK/tLb0GBbnSJ2iivEdwMJ/A3KK2z6GLX/cUrYuopF44lpUqD+l0KxkbWqbxcOx
QxAwucYOy93woD+knq7HsyWMuC/D1H0HgSf105alJQed6ikD0UO+upb3g59rXZJTSKGTXIwK5zdu
QLmbuS/+e9WOwiubQYmHZ9HCJTEGF/oz5sbJnBBcjvo5OIka0PjzPvEYt9kFKvfK1uARdK9kJu9q
m334uHbgrXP3kOzBIBg+v/8HnxpogTh1EHeh5jpjG7LsSnEQDrJrcXXre9PSqhu/U0gMa8Xo9psz
xO8T9UzrXIJpVXxDWxStR7OINhQ9f6Ip86yxC26MeNaT14hPYDkX9e5SUO4kSNUF5eFaX+Slx2/0
ehOmtXOCy/7xjoO1W/rDEwIonwGt9w1TiPekJIyFgb0uNw2nvMRsr/5FDAeCmg8sIr/CDpv34dGE
dVtVRVB/lf4ulCD+3D7s8+h4bjNiDQH9R3QIdYoamnjDCfnJNj+VNF4/NqDDaYQISQ3WJh/in4B/
p4lWTvTIGMCGFQkHABhrFJrDsQ/72KQ99B2DEWcju8VumNq6RhphnZoYcBOg3DCgvgLZBiIQU5Hp
X3GHxfWaBrOm9xRTGhC7qLkoLkfGpa/8qZ4wBZkVEyX92O3mHRvDbm9J12jYoCWyHO73Y8mGSgYI
aUmllO/T3d3UffDi1AXP2PMyVEpyZhskffw5Z7WSOf5Vr3UJ1SXunv9c+RymMNFa/YtprpDRjKt4
fZtqTpEuMbbEHff/ccaVsynwpTFwwchxWPXH0u4xKyTnWOMR0s0wxjS7ZPpA5BOhvpfy3s7uKcV8
Rmol20aeCjOQFOUUyaoGjneZBFAE9S3ZlqjR2sU4/5QrjGPOyzqlD6Bs0C0pmDP31AEvaU8d0dSe
G3VcL0qtEmALmwPCCvkza9oMhsX/Qp0OZWxhrD/W9V5QVjiGG6RgT4k/HcbFs35SCY3VgNR/j7ZN
xE/19kR8irlrrVA2YpxN5uBncWcJLAevSOjGeTPElkasBEkoXIn3NA4y3y6TUY5Jrw8LZk98zXMj
ucTAG/C5PFc1NCWzg51rx9TEai8TNOqjeKB6dFBd6aZ1BpyS/vRFGGDkV9GmabWIPMxc7lUJDUWp
Pfrx1e445U/GfqIC7dSR8hNr8T/X2VqdMKpFAoz1aRydn9YySklEoT4Nit7rlkulvUkUNqSpCEyH
d71jfRmOVniP92B9KwXrP4tF5nqOxp6Baxx51sg/NIGV8XaB0EQULF1E5EF2Lmin/Je496mYD3xf
ZkjoPMfp/vRWFAlnO+9jqALPcHdBFmjSR9/kRw+3MZ3u7C43R9zVuOoTFC+hfGd1ZR23ytahf7PH
b8DDko0rlMB02hEXvHucFzcVCnA+huIuTJ4+JwuoZLe5io2aeDMT+zBfJnnWZwCXo5c9b/w0Q3in
xdN9CwipienOPV3+SSbnPQB52oKg2zlBB1K7MvrreLFWqBX+W+OiFt0Hq7CebUfK7B6QMc4RA4ug
cQapAJJ6wH3NBHsBSREeSBnUVQvfpTPzZcxidz0MYVJ6F7tZzSIvBZCbxMo04QsMq9hl49NiS85H
VH5rilKkHJXdu+KAB1jCv/rVfPaMTYK+pBNvq9flK0WZL+pLbAssDmsGoPuhmgkPBJ/a/VG3xLpQ
mA+5RltgnepgqPyYdEqyD3sPClhALm6URyZHtHmO2TY4dlIFjvLAuCfGABl9SDDOj+hebZTFIo7H
7bhSQrxY6H2Cm/hEsxZ+ttaJfmfXoZ9C4g60Fmm9Wb0pIDQbpTf56xfwhZGoVhDrJ+Akygw/tVLp
OzaOkG053bTZWYnFI6odYEAyhnHQvGtQtYtMbSdXL3dQy2SF1F/a+tOLBnCBzF21qjs3uV0SOIqB
DNrFDzlhuHNu2A6krdDbYPCr/TpQCG4Jbk6nwJbb8N+PYB3xlZC5sIID8J0UrF130ghMSfT1pmGU
dhGE0UA5GkfTuTp0lxqvb7YrbgCQCozXnYHVhzx338xS38IaNgKiQ8aGemC2fDxB2MinYsH8awFN
Yty1Al2PaI90otuuMq8f2/gIF2Cz/CDXhdNJuXtMm10/A2ZH6lcMW032tIPkG18ef11fdKglS7Np
xgiiK5rtuLgnMqMzLh/xSJn85pBXOk1traKXue1l9ovkGtpllYsazsfrqPd9oxrtPSYUdyRiV27s
gbTDoWnLxofsQUPvmEUKAm7PgWQhQRGzkkjNXuMiFfjZYkOKQSV6n1Yp1tZBjsnFMuzFSC7ol4GP
Vc4Iq5t/BXg/LyGfYhUrCxcFga1R1DoHgi1vVPaURaCeRcbhZK4OtULaHYdduu9wqX/xh5zbl+Bk
VboJbj9Y3xcDf7RjKfVtNp+ipaE0sQyXjAzg9P69ezuuQoqn8e1Dih3u8qgakgxjRGqLM4f5AoOb
hi55fxbIEC7twuFB0UGV4pTfPw7ZXfbrbaew0mVp6Nj9sGKwlCbO5VYw2TCXyZWngEJSDXTMB+yV
u10w3O3rrYHFFCEesCb4MaDgwiVzuLVocbVyWBXHTePb618czexevFZMat3/UfMv6LUcBWvj1SGz
B8pk3nmI41omrBnwGxIOIY4spFmJ3jgE7Rt/zR/bQ3oW0HmNkJl+f2KmpC37InfL8qXNPeUnE5xq
8iMTwKja8zcIrjk8zT+i8Rq3O04UYDvCoEKmG1ibnsEzHItD3gErJ460yTna++JB2AxbnRTnyqR4
jqPDIp4GPXlgTfpz4eiQHrLYlCkXYv4SuCQli5s4FIGg/LSTZdtXOeKP+3aB3yokJX8FkS86l47M
1ggHl2VppQmlusGtEbPrjnTft5imKuvrq9fcEUn3X+js2tUL15D67zmtxde8h5AGL8h8i2XGhpus
UAqysK65P+c4mOqnmL5TelYrwZdWTp3mHGxS2ZiUsQd9ADvAq+q6gB7nzSEDjqhC5ROaOQIMEbHK
ftYPF2glbOKZ690onST++Daw+wOhv7wDJyXePQheozHfYXtCYNYAb9f0gupDogXyA3+y5EeBZqNU
GEP91EA4AvdqdIRiBwOZYiGA47+8lpxFMrbw8S3U0TtSvB3ovD0HXQEAdgL7Dwt2s5xjUfXRM2hM
74FVx0rzDyrNWg9j7khRGSfycCcCKeLDKSBQT/oiLspSiQfnGQN0QuOKEOVWaTgF3oAmR/TFC6P5
Fg7zXEVDWpkczHIE0ae3M2KL2qeoSHl1myIEewW8IclLqm+rUs8pvJlk10ufXZCHdWNZluJdgYP6
TaS+cZC+fi9ES2UvnkbHLHjoU8Kahc+9PBUgiYr8EqmuYtL/4rJgICdn28nlqBLEYq916vlSsOL5
TE0kE3FoBX+ZAPYdFe8X0tPpjphYEYXFMxd/sXfYoAuQ44pXN0GAAYtLXhLPvYTpU3Je0eYBaD3C
hpHbkcfT2sKTk7ZSu69F1+ZxpN2/3999xwG8ykSFi54MUs425MkihGBeIRkV+R1TrZ8WFSgZKOGO
vBiRqMmtB4RFSP4CI2AlOMalX3+T7ReeRYZrPteUz1nazHqon9CS+hBYYOrqyjyPfFcS1zByYOBM
a3tOA4SsbAEv3HTKLNc5gpBUO4xmCFWBUvE7DMgLQVhs6vKs2y6tlujAPjlK2vW0BRFxOvGJoVny
HHM/Wv+xvPqy3lDgtt3rkbMu5uZaz4CHJLQ4jRkca2ckU4+SZx2gR+I5Ztt8TlDZt3vCf/0EvBUV
SCq3HZlVGPXDUd3TJ7S7gQpMsI2qb+zjXZoWS4zWDxz2B1Pz4owimdoJmcaVeRgB11r8y/taNVBj
keswQE3rCgADECDmq2UEJwrujMLXTyg9xoPBKq/kOpXmfRcaVma3bYc5cqPiGyDmroPxjHqU19/d
YnTDSm2sHpy+t+4OzD9gor6d1Nhp9bLlRbacRHCL5yfwfyP4teHcpCx//7zBmSFkbMp2OZliNIOM
YJwC2PVjCgc+5K24fteW7NfBZoLZY8Z9wA8jSNepMUy0fYqg5mAE5L0kn9WZpBAEtzurgDsxSUJI
FhU7oCs1OAgxm5Jxdau4e9nwKazZGOACVoBwF7ARA5krw/13seHgTRulbRC6LAhirknw9mtmJQ+7
mhKqXK46ANUfbN0nLghj5O2wKKTzULTxhzaKv3Dvni0oj9axYBF7/3t+KgsiYB8HrF40WrrpOOMr
j63U/rBRckqrcSpjHlUCiX0SVa3cUMrxXpaDS0oNO2jAEfdnlQf/WVe87dPQn/md5T6rW055MbjW
zJBYsOEesUPBGVqAwbrBQRD/XmlK4Xow7YvWVbO0MkfkC/JD2kWu7bi0f2q3WvNYRhiENFrzJwUw
bDhsKO1X/Db58DjxC1UeiFTEkYDNAGaAfyfPNqr8g/VQtcJLdcnUyzwuVUS5Oq/oA7ujV5OFl6lj
zrx/Hbe2mc4T0kwRd9sgbeZZKlXzW1kKDfJQvvnq7w+iXHl9YPE/Txug6l6Nv29qSTb4THlWfP40
kcfdSeRCLa8ZoH5OHbtYmQBDn0CVYEReCgem7Jm3P6CbDZgmEiE/acihOjU4CtUzIV/R7nPqV7xw
t2/5ygPaG4Ka4rbJseZ0iJbucpcSa1PFQ0CnFqzkEd7cc6R2Wcqr4+dHkuGh9TaIVCSyVymZVaTc
jBwpOCfJ2FnrHQv4NPXZeoOkUTvl7XghrR2TkDb41TqsFA2fgOuFaZhic3K26RCi+lO6yNhSkjv5
Lo5gq0voABW1tVcXquPOA5hCd6lQRmiW687cez1YCBw/rpKtoxcVxDON20Xh6pSiWtt8lTlxuItK
WB3oxRIznjt71tfq/2+vQFFgtzaqKXbpjdYso5s6go4Xu8wU16OmGbz5W3kLxEIVFQUnLb0LVWY4
Po+X/7hz+vQbwpBLVa5ILZHOLlcTlfb7N70P1GF8I//3UINOtIdHUmBmpkHYxljSROWa8NQqzW6K
3riIOXIcO/3p7qzG6devjFvT2ylKd5IJV4DOrPrxenkO0uBqidVBcLVApAeRaKLUqpcatLnN6kKm
uuoE3eApDPUlncZjQveeALjL5tsQFNTOWCj/3utVpueDMyMLcRAcqjHCUqwHf4H1/PNnN3FLwmrw
y8SXMHWLHnJoh7oVgq5nE5WtqywBQCivh6ImO4lsD49miVcQ1zXdQ8zCZSZ4MTZDMSngfL/I1Yym
V/4s9OhNjG5KnUcJ8ioIeNfwzznpNhF6CZMRcPXZdGpQ6TYmEHZ+CSnOtKJsO6ltGtv/ypbtWdcJ
e3zHxztaIl8DjdKezBfMbvUlTkFMzrbOsfLodLc/a/lBTMwzUWdbLrlA5G60TrnKnRUjDdtSpcZQ
9oVTrfScWWpYly6aqCzaTHemDzNwz2XAEZ2fL3cExJRCTsTnqz9GDN6H+8z+HaxNAJ2rCCMstTP3
znyhagGvPcTForcDXrFgGFMafEQaMYHm8YIby+cpQGSOJLh1emnFHFtfKXonQukjVGSUbsB31c/S
qaqxTMu66ZyNmh1rEyheJ1PUCI/fnkwJP0AHNRnE7GeVG08fSsRxgUo0E8SE5c9cGsqlSDWtmOx/
GzhPUjCwn77vhESM4cXtK8LYy5yNA369S8UoqSDUkS6cLtYeOBwF49cRNxzUzi3JlSAtPIxbEw2X
Jt0Ud4TYPgR1fsZQNEnVtUHfb0798YbnTZbEJQ39224bjaXB4njx6ukaJV54v2XEk3DsbrXMWGnc
+rxgLdSsPrAhp/7CVsG+XM2IOLCfid8nO59OZy1a1MeiD7cJkHGB7QUyQj6K+DpCFQa1dvPbDLhZ
03rKGD4GY6u26Jcjo5SR+FZfge9p74WPOk5q5NUIsMLcFv+pwl01Bf/fiDMu2ZjqWNUunDeU7phU
0sKc/Z0zxc6e/P5cxudXlSSun6mQqyn3WW5C3lLrj5o4h7mnnysEsHIlEWMomqcqdOU4LxCvYz7M
/J53GDAORERG8Cy2vbMdIYEwLFe9WoJMLLJZN5IlIX2B1mwyWBwSJEU6AhEStrxr1hU9+2Kp1xk2
ER1wA9bs2+Xd/y+zEpF+S1zMPz6obItwfS78/EpGVWxjXx6kAxyyA+aKwd+LDWSKWvYmDv/5wcwE
0bxx/kZkHym5E01CyLlIqgy/dQU1AmQUXfeqNFh3+zXdPVTpnRVTJ4rogPVRq337U1aD0PWvPeF9
qnHEsdkrN4Cm6C6uoBtP6pnRXxIxN7yDVWD1Y3Ql3gM+G+7NH0BkR9I3XJC5hjfnNRl2/zhAgkpf
AnXDwUvaZ47SknnNnQ7wIVFY1o7tAEWsH9Plj0on8+vOJn0lqqXhF3yCmW7n2eT1trC63e2foxpr
2aGraa7Q44Q/QbU8/z87p9tJa+qHbLzRRGx8lmWqh3+OXwIiiHl/qQCyxX9R0Zj6WY7xlDdJMLdO
BOwf4YNu+2r8xJJWPD6aoIMQlebOyXLwGMXKvaRsqUrrajGXi94t3LXu47RI6TjZQ/CK8YUpvAqm
nMHu6Z/Npc4OgCBqNgiiMmJK0Drlkvc/AQP47MLg+rX2x5/OTP3pA38HmKRaLNytD0h7WY4ttTT5
+E59nRV+bePqSX/aFL34zK7OIBWR0+Hg/vDDIWJOSyBSJRo62XvVhBc30VQ81zXX5Z/rZ8OfIzl5
tpmHO/Q5Qzzv+P9ckB2vImaR/XJ0P+qocfLY4jkCQQaONIpVgRWlignQvG28KIYklN62HkCaQhqY
eXilqkmNwoXyityI8NLVRbQRStF13JMv7A7EHELA5sJ5TyuwHsAUdk09vHd/czKHG+A/QWgioa9T
+1vaV0qqFKcteGA5N1k8oH3m9F1ONjBIFcuC9aJm4A0SMVSa0q8EnQ7IGuhV+ZNk3LQYYwxAd9Ow
vT5Xhg78BKiFPF+QKTJeF1WqgqiMYk25tzVz6kzzsf6F2rm8+aD/09OV63kC0MVG5PR7hRAZE7Gi
HTf8GGWk4tmPWW9ogAM8GCoaHJYKhrvQVNovf+s4cAFw9BixSSGd8AghhrOZPeA0JM8Ljrfh1+Ee
XLkm6zLYa1DlLE1JBnvnQyYuTN4oglY2OaQTTIYatWZ20NDqlzRU1yHi+dWqT/gqn82NtWfDdvPp
ejvrTsQ4303XGHrPwDyix9rIP0gzpXJfSsCMj+Qi/Ym4sfX69sfOfcvt9vC0Rv4TrLwNqGrN/kYb
aL7Wfl+gMgjSCrQReoGMpgIAJGt1fsnqSAQvmtzIWb6Niny4om3XvM72+4TYSuwPH+f0GHGNcGVB
ncEmrYU5HnJbeWnZG43dWzsNjKlx8y0h4sQWlyd5z2X2qK5eQvvztSyBTuD10bQCumaTBTkAM/ii
pins7j4SCgczSUXH5Qcob2CNrGsNCl1fcJ5KwskEnR+O2t0QrpSYM8JBECLKJ3GenE+8FCW9eG9e
5WqzE9sqsIMhOA7/bJrvIO0Gc0syyDOFDXMOqNveGYL1sDxeVTTc/iax9YkBegXOJp0tC9wX0b9e
V3C63xxMS1YBUOZMb+gLnZQ9qfe8aywx8eV15mmehMjiEJZ5biurSv92GIMR/nNmxGbR9u+ZxyXG
W+Mi0NIgrUZYLPxS6si1gn2sivPVYWvO5eVNj8S93kmHhh+xSdGYGU8dXkiQJfSwSv+uHGbkZflc
aV+Qg+P56OXfgPvWmGw3gu8m9rcXsUs+DFRYK9Fms6qGTORI2lfJDftlqFGBVOlyoLg57/3kFe1u
aq6a7RwAkyWJvq5K6XuTGo7Aa11KgpcMiGlLiVmUa4VH/XGgVk8tQvdgfGsien5532LbQh6ZuN1a
dbAXZqrBj0xZWCzmMfWexGMaBA80VKbLhKccCDCD7qUtpb3rfoNg11o/9B+qJ2Rq48b1Ujr3XGSv
iqbL9A/7GIVcQ0kwaFOI+wxkUNxXx/ldkdLqqYxuUdVN43seG3+phOo/ElCh/8O23atey1PrMnza
NJYVu8bXPKYgVNxrrAntOFWH7uIo1o/vDxPHL3a4Ukqd3iiC0C0CIJN4RnGqOW892ITiG28fr5t8
uFP8Wv/huDMB4UfsyWLM9CTZUVgz9NpKkCsRfSsvGTN9U6wB1hxfwCgonpzy/zNq98dq94Un+NPL
F4D7sGSeW8RgbtqNgQ+uO5OaNSg7qK6eTOkXIunZ1jX7ozaekJyqMgw8nZhpwpV8/0Q53JB3H1EF
dXb0ExPxRBkb9KxwiSLIlEWuUgQbAdfmZXh5xDd+cTucdB/x0WiIttNARhCcKfahPaDDcJOw4Wfa
ewR2qpwxEnOJnn0SyS0C9XHI6FYSEVdtE0WEBBUu2coHXIX/sRp+uEYuQsEDzPPubjmrn4vppmsb
Q2Quage0gKhxeQycVpcZt27IOe0u6xIqD+nrxffIVfFeYilYaP2Hy/m9gMR2g0W1jPFJDZQDiwdo
BT5KUYZ/Xst6IglwUP04pbAYToPrP1EvCj/Wln8T4L3GoHc8x/gH/mNGGD1tOBrLHCmVyiIHuDVS
4tYp7hnowWxikw1du5pn/gAOcstscLLAvQZ/pLjXnyFiTOC1KE4ewVUAC85h2gsqlr+jaBb8f7tQ
vEAPnq2RAEzaUiB3g2pz/tdtwVfWIhki7Ub69dIUdfMBRZKMsEcC5U+WnARHL39OL8hQvAt0nRup
St3awMutdcEnC7M5C50DjWeV2DXXmJn5OQHSNKOFSc0WnaJZsbG9H30Uo+FvsaRUJsCaTfHWJov9
cwSRPr00TtmzKugYdfLnBWb0a6OR0fQdrBNtnrr9dMhlJGCzBlpfqV1R0AkATOBKDdoQAntPA/WY
jSxfVC3Z2itbggSp/ekI01XCB1iO3qKGzsgrPCufzB/3mGzGCiC4Oeni31805tMrC/cQac0t9Dro
GZw/mJcI0PD5jlQeoj3qovhhbEQXjF4wuJcZ1SLPSv6h5y5awCP5JWuTwWHzkHu8KGOkv1KZTEBr
M6fTkx0DWNcwCU4xiS2kZt4BksNeiIcZJrXHKpD1Rd6d0SceIhQ60NKoa8qbZjdDr5Uy9ytLAEJZ
tI5aUlpPTHsxZqyPUj85fXQBfDr0AntsXBkjzUMuoDxFYtbIqRtQ3NJ5JJUyjP5gHQQ+IW7Br9AV
EGGZkzSfQPisGjUBy4mVU4jPkIKgvGp5bbqjQLlrIcic1tsNEhN3h7MlxtvtcIyGQ+LFtaKWxgkp
iByY6lHH5mQmkaUAEP0uZURC6ZJfjlXAxGyI8jbaFnl4kbZO0vRFbrTRUies5/Ncxnxe1OWOn19n
it7J8C2hERPV7N2Xv126eZRNs87XEWFCtK/JzGQYSyC9SykhyXNNmEUDtZlm2H0du63lH3ZQooW/
seC5wZZtsGz5u4VS6VdNhyAoaWYj153P9VSyEmGmlN2hzY6lS+teCvArOhNus4GFyjAtJC6pKC+9
OtyTgauFYCMU3Rbo8TJ+PxfYySpnutLVg1iNpaMXIqFXuP8xEa44IV2Zaghaj13THKUfsdYhK0IW
Ao1HMotxxTrRqWElFwIcXIkrKq4yXhcggGuNiG+33eodSrE9RUk3h2qP+gtkOPkrzeS8pKpOggHo
ncaiuY30KL6HFWZllVNcDwXy3L3LgAaLGj6dOjOhc/7Yoy93aEjb4/F33pdSOgSZEf+/tsUYbAhz
fLHHjbGvEFcyceK+wFqPWgC2u+2Oo9qShQi1laRFQwS0GdP+Wk+UYj61heCut47M3EQbystBAFex
J/sLpD7rtwYyJTlqBU0OWJVxY6lU9h+XSXCoQyr+mrlTSSCoCLVTMEoGQHqbbBiviOFcWAcVucB7
u//4HPXKNYSiVck7huLLJ6guDaUtO06GfKa62N3H/hO0eS/x0tcg891p4sy2M6Dptb14INV9LtlW
BoRM7zKf8nAcm5KQH6xvEBOA0bjHGGInXBZ/+4s9pvvTAC+nJ2TTW1dxfC7FiiHQWoCPO7w0EsQd
dShl2UrVsy90j+G4n5UEU1s60x92YFxUtVX6i9aWv08NdXWReuw3Hp6eWsZvh2aX82eqPRnYLMf7
890+2huWkiNan8dE1yqdvyVXfrxojXQlKL6sns8ClFDJyU9CLdoFkpERrS201ZWgJiVBsQ88Irya
FGnByrTuPitmmhVOJj/o31L0as90lIRyulK9gVuuf9+znRAccwXtzIyhnrFPIaGOwuwQAgGnSwvS
JYXSJ9hHn4af5T18cNo0IGum8faeD0aOwoHyfhreJ5iAft2mCHkNDayVDjhH5ssVJ3g3SC4AZroK
+6xqp7gRZr/Y3tJ84I0D7PRfGSN8NT2Gi7RxUIZN6K/qRbJBCOD4CKx4Rsr/Aspn2x1dXeMSqNaQ
8sfSbDmbTtEWB9WGTAyw8ZZamoIG5kA3yjISVXnfwdrEKjYCqFyb8eYlBZxSj747FEjfQeNamV/y
XP6j8awJ9gEAy8Vz34gJ2zo0BzRjozSw+mGeCXnigx6avK4zQfU0xEdB18tr0s3Z6p+oA/Vxr9is
OkD6fdI3PyV+d7EYpBiU8DcWsS9FRvpH7KPEc7tkqeXwbzoQ13kJd+UujR968O7C+1f3Z1oho0XC
7JzrK/eXQN6c/cs/FPQfSbOsL4q8X+4E/Z3e/+LxZhbNVb3j7ATF2hZfSNyD2Iw8t93/q3Cgf25s
BSTNcX0psLWggO1jPW6pYORwLkUGTP4Z6xGMNZUuByzk2G8D13evd23twI84oD8u3wz45uoeOV9Q
byvi0qZ8IwzxHohhRePEo3pjUBG5KIfXrhwOkri5sAWRqbD4Mg16vfYf+qQQgexNNwmgVrYawc1w
8FrmrI2Bfc1vui07QBXlZ4b561Uc/TSuiVxIIjJ+U0CRo0B12sWgSIOaWGZMpjRThCF97PzyIDAS
uYryBELWmF8YBAl/8D9wFxK24Hc8lzK1w1BMbt8IiFFt8jVXK5+sX39l7Qdfv7PpUcoYrpASUZIE
EUnhQ+H8JiWzxUpfn36LHS2tQxz4/4/zFJZ+uHdxTvGAKqV+iw+i3hQV8Q7oa4c6wicjW0ZRaDOT
DLsY2w0pg4xDm9KnF1+jlnSfaHjrEf897VdG+3M21GqsamJWQWLTc83FemruGYarWY3xZeCCHPtv
tDHS7nwzesrJyFNLLUfK69WJES5ECRL12kCwQxWtSQxvG2GJFV01N880J8y8xgkeyaw35kbaFuR5
3Y7A1OYZicC5YwjHAvejLfBqyjlWEDkqORNjI2am0aWfmKQGZS8pUYiVpFA2hG/439B7dI82lHoc
ziQb25jP6MQeVW5IwW62GIMYErCVX4DV+jY5rjvSFwMdj8HTTfX5MHMmWcx/sHhRIu6DX7gVQYRQ
qTqJjr1aZYgZyHJnFLF8XpxKE5fXcsjXJMFLF0ESwiTBZshZS318xaGxsVgD19/m6AF7irb98kk6
kg4g1yUApN8Uog5nrmMstnNiWYvqpoSTEM5+83BnX09YsXel08hLvoB9u82sl1ZXcsxOAeUGJXmX
4zb3KJ+x7w5NJ/+ZwjWyAd0kJ6ULgt2yGEjBrmqCZx8h6i5LUqt3BlBBpjH72/m7J2UYkUIi4ls4
HltFAfNtskm4duG4HxKRimJ1f9gOPV3rDh3/Zd2sdDP/+i3zZr6+tHAZcaJJN6swQov4rlFnQMZL
K+1tIv63Y1Biun7/iJzIgt/2vQlHeA5teVA0GnBbYt5SS6u1TXnBtuEacen97Fkdx0V67cPVQvXc
RrG4BLsT0mdf268poyuFEFmC4NhWQ9I5pipoDYZxOFlnOPMZLg4XgfPWXwKtlKXC0nHbYhzTrVYb
B9YBivx0xgkLFPQdtq4vfma8yD4iC0qq8W7fJNOBQpZfTyyjajPKagFhuaPoBlH3CQNBwrRmRWcg
SHLyePmcg4GUC/7P4uzrPsRz9906ErkmH52s4UDMFjbiD5YA9s3ZzrmEdydddeKRfNcqdapfmiRR
NFtbBV1gfop5Fpe/tTZ83FoF4XUeX37pfmS7EMk9AsmrJ7z17enQgTXWkTo5c5QRMYGsDWpGUESU
veTkT4giSjljE8zxN1ULQnqit3/ZrWBQnaNsIbQzSgkOAlC3zQjM0aL731lBkw9vCXNJibWp0XKr
HZPVSR/T1/pbj11sU1UD5AAaEF3BYh4NqgZwbDriMcdaNKX+vZwhaJWabkZr1eKpvhRDXJe9XkjE
pQK97wyUGFvSB6ApcetGEEd+WhUxxwE8ybrmJ8X72Ux73QjkKHCsnhpCpETY2IJ84ncKw37PuMLt
yE+ckPUj6czGSJz5KVrL0eu0MO0nJ8ULw/pnnPQPk1i5x2EVquKMk8XWgbg+UpEtTUX3UAMn7M/Z
wdfkJXmH30XLfCzz4Ps6djtoCNeRp0yfN0rgmjFDb4YTqd3AchlVkRAldyL+st2eleD9D0hZ8Tpn
rnt5YluJzvNxBdXQF4P+uEHYdOIKXGJS2XljCf9sx+INXj2Oq6QAbwhBiXMeFAipIdO/jeZA2PF3
Iu6dUqH3nZIW74Qe+Xjdba7nhmxqTMfGFcwxeUHPFoUC5qAQzHODniu976vhzS58ZapsgOP4RGsj
X3dwnYqSst5CZ4vQm8RSDJSMBxgdHYBwaDvM5fa+ahsPB0mhXxH46kVwCD5hFPLPibribLhkeu2R
1pKajY5GHfsu4olLbfNbu4joIXGDFOnd+zk+cgP63tdRzY5HXACCLSZJFKXgHpCPwpUJIrRe3j81
2MGgyVVqth3sMvEpI0Sz+VUedB8kuWSlbtZy54YAuZHtDLJxxoBO38Q9rmDiybAPTpOySRg1Gbsp
KGxFQZniex2pAWC5seaWlcWvblu6pcU8TyehQN9F7NgkSOxROhSp2yUOd/UkwBnWfckSOrsysXSo
ilUTOxP0NvTcPZbKUqC31KMs2/6GdgfP8nPVJD93wM9ftSmL49gfy5ltwGab6VUSNor/6Ikawf/X
GocLg08Umm7Y614R2WfZ7L3hOrGYl5F6TTyM/UwVJrvnCCzev/sTwsMinpdIP/7FMiqbCG/hRJrv
aNZ7/br0yWQW6pW3FAEjMkMl3kjbB7q44i91Yg/5eAhGjTJ4W08oVIT6r7y+ZtlsjdKJh8PENbuE
s9VfV8ilLBY49zHnAMt4XHLlOgtLki6VfnHZdYmGohqBik8SshM4Obd7s1QeqedE2PhLUmDWlJfU
5yDExCZdqPGFVc9EUIionvnI2u39qyAy3wEd+8yK8F6X+vvYr5C8LrxNlr4y2xs1fziwT69vpUhy
nZz7s9yB2x1AmrGhJQlWT4se6xDQwVTlADDbutU41X1A/7lijy8HSFZ//mw8FLTk4xfOe/z5IBZ4
pEQNfSfywK20UK6fFrvtCf+x7z6uTuweBgwewaKxLv13DmoQO9zLfXRRWb36eRO9jzQ1bVzqiC9d
ijguQfg0gmjay8TvujKyt+m2inbp+meucJiZq0NtmNlYN/uF45iQivdK7ovQotq8cMR4CprIRNob
Ucp438FyfS9dRqcv6rbGiUfCKyKnQN9kg4jk7SCmq+Hjj852ABaKs07OJxVaESX9x2KARjjtteGR
u3Y5kMYaQAQ232f2aS8iieT3u61beESe8MPLQC/wJXJa4gbh89DmZfMvwPtMzY5XYKsqf0XEYUHv
RHpGrmrtcXGBvz12rvndnWhL/AFvc6G0zYFpuuyYGbQSISAOFL2S46cqBUfwJh67kW5vn7Uej4/X
THPuifbraBT+znKaSZxxxmoHUEK3Ha0f2S3DTiPV0b2RzXDQoaSbbH1xvg4fL3k6oK44gbM3JzGX
VST9T98+i3MnA2spgQSRQ+rzOk6UTakuWSDnhD6HcZbUCtbjvsrrXGzKi89TpCVNPAH4E9xg8e4t
mmGrSYdqYBh1PhqfBAWquypKWQe15l4H2ocs2ZWAXzk6kx1ueetMjS4SuXDQCr+pB0xLf9RYfZ6G
IzJ+ajtkroVDk4AnaR2B58QwXt3JeqGbIsCf+cAW8vU4uUEvrv+3ZU/y+AdHo5LPYVO/Z8nhtmm/
swSf2xGCieqAFHQm57vrAET76mhFPZz2rcyANFBP/9W6cv5n0THod/S+jbWocnPIBnWuYsGveJsz
v5AgOK2y54MSBtr2pEuHu6C1uikdzBpNL9jb6gV6VLZeMwR2z4oi9NzGl4fw45tEXHZjoSppx/hv
vKctWYcqE3Fx/WeHJEteEAhjnaQRB7LY61QnpwAHtNr66I9JYhJNR/zWyyTAUPxjCVbcanJDd+S0
CPa+c+jmK5EYPJaK+aV2TB8km13eOvZdYkwwxCXWhyQit4XtYuaf4CL+jYLNlKLSNR5pz6VyLj8h
pSXY1oft5opQfMZFv8nMRbbUYIhrFnhXzbLChAfLJHClIRjXDhY/ZAGwLpu28gkzFDfYz5BfpA9m
S3wnfhzetHl+t5nThPp+qOv4eXW0bpiIe7Sy+kChw+mK8JD926iPuNHME4CTZiLcasw95GRDspdD
Iw2wmKhFcG1J7uTzPTU3w86aKilQIxzqtCFaArBvH+JturhiwNjJczRBIkRlnDcgqmfYDtdeTLiw
AnmIFRliwKPoTiTc0gXIT7rFpH2W5dT9OVr73MJYW8r2xKwC4Yt9IUk7Le3qDN591dzlG/xySNOA
OJcVNt4zsiNqDir0qoOXU/k6cYSYx8O1nOMbrSy35ehIgs26sHW8f+seEMF84dzveF5ysNM12/BM
0BKP+FQgHo0BkOZjDbi0T9o4pXG/hiStUwRsktf+a7nIs8bFpl9HqVVTCk1qIlrOytsrBrnC7AZP
BE3reh9Qyn5BxMOJhz+e2wqJ1qTn4UHhiH9/tPdy1hxfhjYeLRwIq7cB95A4jAw0K8F/J1uG4b1T
S0/IsGl6vi4uO+F4s6SIO2+oTskLUAYozNS+qr9WfLgqq4kj+8W5/YUCeFUOvI2gRCD0SKvUKPHw
j7N84jz8VsLo6cBdRjnofvYnv7aNL1oLdp3ux7QVbgqXpZyDRKH6QHoW3anaPbcPNKag7C1pkBmR
wiHYtBa2g5igCxFyeAELv9YUXwbFv9ZrndX2KrJNaRzpEVruzLVAbP5HKMkYaSD7OqTmjlBqspc8
aTbj8A1tdSC8toFlij83oNKzcYvJmsEXSlDt+nr2S4cak9FWA1JlA9gVDm0CHQ1KvWznxljT2mN0
x2LeqmxYq/w6xUpeq/o+MrL53AM3Tp3kK87L1INN9x1/WLKgKZjStdp2pehEStuWhZ++oPOsuATn
Z5Z1LmE0NrjdrRqAvub4n5o45sjC23h4ckuAYypNhYk1ohfSomfvLJDnbZcnM8NLzG+jUF0uqpOt
mE9wW5pnzC8DeNXnWTGPAUrHsO+fx1Ib8lwANIBHQH8nwYYRRzxNDzRS0wETcmCEdA7J0WdJ0R6s
Ds362V8ywFsxDgySgWkmMai5dmrHeg65LdnOEfYwd1Xzc5Dxe4dT3+fPhvg66ny3V5UykoL9qZpS
OabQ2LfIpqUYJIzVMXQ0SaM1HHUTF/VqbsQzX+y9hmQWsCPYI5Qkn8IL0QiGthWiMwEKT/aP8oev
iHx6jHQtz02XeYL2I9XlIS9v9MFCxsA5cCAzfo5a4JqPMYXQ/rBv15jS4S3G0f1fBPjCSqGcNZZi
dC6jN6lQFroTikod3clll4XkMiDwD+SjYGTAtE0nFMClHcR1WSz6TCCeeEq/7W0KdquVfVEa6twy
Z4rBW7mtg1rEpzEW3kGCFLWOKtwjaLUC310VvE19IaaTFWAoKXQjZO02vY/k3pFv/bSTiQat2ozP
FXvnMMu42wKYyveBYMGDezC0aICMhvUFIVFBbVjXl5hnIyNQeh3UQKTGp9ywKnA1FxyRf6y+u250
d4gQnx6Ue9iXSfNmd1A+lNSLPN58O6A/3zK3Y1J7dpHXrUW2G+JC6GZw5mxp0RHOwfjweDrBZ+fy
BH4SFI5QTw00b0+mQav5zQ4c1ADv3pSRdyLcoIbfuta40y0bVe7OXaxjCpxg98IfUSqUekadLZVk
Y2MzXtW2wvdtq5brerUnmMGcqGVKf9hfGPKGqBWxYTKFwfftNCZrQh2HDgFHvE6oo/eL+rQ+tnb0
DyPWosCgRHN+JWVjzwXxeAiNSywoykLmS06Vk1QOj7My0zk+3LbKM3QQh8Wg2P7kJ85vQ0O2gBUk
9u4ldw78vVmwH3yXcxC05Sn3cGTbLvYjqFc/C7JTxiIjqParVCbtVBecQnKYX82c0nZYkyZTXdtC
0JrRzfuOhX3SHH67IQFQpkzqug8iO39KgZmSADUK2tzR9m3f9+ag0jY7IVjnDXFG6Lj6BO6MKPZW
FzDmoQvh1V9Jw9+YICZ4he8oFYj2JyMIHCa2bkI99ALbyi+mJPn7m3JfPzGMGgLbDeN8UZaZYbPt
xxYlCCUt+DuTzj+QjDYKfNXiHk+3+JO4kLrbeDuswCLSQMwUa3omwFLStTEyFB3BKuUXoYK8el3K
dIwF/Gpe1QlN/6KvAnGNIzSEaBlDlZnnDy1BmsW4cVCSjej3Ncv421E29B8HsNXuTfgPoaNHBpgR
8ZOErC+HjrwHekmYDCyvTM7zCDKd5GkGlsblqECmDKUx3Y4xrzEc6erYgKaYWoignsSocro/zRkq
utGMpViHr03wV/I26pkv85gW7HLixWtWpw92ipwgBxC8AGJtnAHvirl1Gz8MOjqDN5cMDnkdVGq0
VaR5d9bEQoGLXLZYVPfogLsmHZpTJLXp5yXg9/H63ZERaG5mMndWXNhsUd+nzOy624SBE+j+sOOU
nBBT9jM35Ae4E2SklKd70+CVKhMoO+0VncO8K1Qf1fER5NyCg8gxIyQ9ZMGWt1cXOeKAeaYkI8KR
5FJD2mbVRZzzqNKdAX+FSCrEtYhaAWP4PsdwwZlsJZ1XXg/Vk6nDt/rVfpmoR6I6OD/mz1NWMUD2
M7bQKMbgByz+LADapQlGfFYQ+kdLet/EYIlDltHIzur2u7OLcGv324DbbcbmtmqlS7w4vL9OZqVc
c/CTvhspStaMk3gKPnIibUUtiWy4UeNNQLp6X7q5973uvywKD2tHdZmMcevfLqlW1uR9Qls8YxEf
o5ymifL8J9p6DvT2fx/AHpLHc5/fdjna0Qr+W9POKOkSWuPFzkPZapPIjS2rsozejpvXyAd3OdFy
H3s2hpGSDQ8E8vQ8w0SToTT3v1Dq2DMEupiXtXILj/tFpF/LZ2zNON+XxfsNUl27NmUodhsRr4rN
vaxvfTCRPxxHomzgMkueqRRh8a36exL4HLhlhma4/6umPOpDXJ98T/Z5fvc/SIJ0A8BqGbQQurPG
0Q7Sgt1wUlwSwaZr7AH7dNhCso7ZaCyZpKmdaEHjItlUT+EHXoerffbKt71ebQu3r0D66Ke+Jbou
sqMWXXPMnkloGBLGx3DwM1DKCoI0173TFvGa9RgDyuPozFkNv5L+YFHtpBq24H4zQZoI3d4PHzUo
WCnGyGqaVAoyc6uvDoKg5dsNFc99zZ1uKN8MMKtxkVgA4NYhLBi/L7afJx3uUcsR1O1Ikw0Icumc
atShyMzoNt63t/9UdBcpq65tLFdww4qSN3dGoFE99Q1NrNi/yuQPhSm27XYwwR/H+ZQkx6sEpfGp
jbRbKhbl2/qEOhSqUF/Eadkgy3nhsaL/kU1z54pYmB3J/Po1fMjNSlSv7yebe6cVBiGRWJHqmZkR
tksIzW3P7auulR3oRDhLNpTwVXA3VPUeFzw2qdtppzJ++C5AK0MW8+Ede3ELmn1/dS6TvxMtFY2K
Sz/wHFOtT1qpg5er8mxp/nFJdAb0fgFN7ttUq2bGVKAzcOa84dmP3KQTuWwPnHOhMLx3LiXLuo6s
MWyYrwoKAc1hbJDKmFcDWkhHjNeIe6rWuhKs49kJBcYKy9TMsXRfT60GZhUR+tdD42MiCTgICN3f
BhCvpCc7XwfY7W4nUb/CXeyaPod/j4Nz3an96qP2YNCZHXSCCnLjL2put6n17jLVDdVYeS4nMT6n
gaE+i8BX9zxI1KVepsBidUcyrqgXS+xrEfYWYuJl5GxttaBy011kXvWHrDO2c5+MrAGZaV/7U9LS
g55BNOnl1cSHOk89K8M0Qwm/eoUjFcz8+DKZQvRkbT4iFpb4bZiyceFWKRfu/2rLKjulOsZfzORI
8ex5+l5iNaNKEr+8eFFhfLF6hDOpZFQO3Qg2+LbkbDjM4jkke1nQqvI3y2IAtUhjAwIzm2+ZUPHF
9t9CUkvnfQrvjYMPFQptMn1uo2E3sdFW5r0aTat+HyA2ieIfhq9Qbx/wlBjvlWQqbcVTxKLx9Ci9
4BbWcDYWealMJ3z4Bt74TCvMgre7ORdGlX4G3Yb85pO6agiqfAnK+K7kQ7j9D2FvSW1+Im63JMrf
WcjCcK//1Enncp1/udIC7BQs/NV0G+rjGEDhim3RrqQa4/cakdsD9rLqKX+Mu/fY4/FlJjmMuhnr
1zSgTg6ybuC+nBb1WODLrQITPTgjUcEZDaz6Lm2NUNR2dn5sLm0fDClDAozsVbrVYFvQLF5UFDjU
Ji4J88/SqaFQZeC+DhrCo+bbIGGaPOi3E2wXD+Iltt1btjNA89ZL5wvuPEOr6UWs8pjdD839lNOO
x4xkJ0ZhbWMDVwS2nWgGmEuCTUMMd9VUlHnBE/ioElbFdzWZ4zHiFUhGHoVw3L5TQJEA8tdhj4iw
6+AByoe0MznyVUgEWtiAPcbO8wPIPNaOi3jR9TUn8DXQowh2eEpVv7YkmwyFrkee/FkIFs6+I/4T
k58FDCj7Gb6yKNdhuG4OE5Hloxub1tt1QGmXGGSBO4eBaKacSjrLI+qLScUoXOxqBpzFvVZ0r50o
LdFgjETyf8bj+mkFYfnysawBelOsDiX92wx5Cd2mvf1HyycD9PfyBizqMzlqI4hbTGO4LeJoimXC
T5ZPFVLTEDLhwnowQ76WI677XPqWVR4SYgZ8r2FscFBfkK7u67bXgf/M1lFvEpeLpAw2AGMHWPR3
44HLRzQNAhY49/hxpZQtRAuiulrcaGc1hT+W5H+U/yzYS/tUI+M7DEtMCNnZLza+HItl42u5eUpS
/Jio4sD5wN6B0qzKcxa1nZwEoqMU4Q8W8i3mm7HkjVpQxyQmLuz99HTB/jYo2i7yoc1P7t7kCNvF
Yo5EFVQ53O8+1TqoTgfZl5O5fnxeiFri3D5VPcFKGDF0Hkr6Dp400A+nxjftsIkp8nCRSSvORZ9+
UK2ply97emK7c9MXIqtjrmCzvtyxk71tVWSgSdbmCZ0lJnGT9H6nrus6zJucPws+oClbIw9VaLsQ
ATqN7JXIbYk4S+CVS/jM5sWu5k7Tr5XPPUe2zx5XsJMNjhgcrWhtzkOOe+XYFRZ+kHQrmruLdTJZ
fMPv0KF5CD1QUvJGCZZhPxsPIN3do+f9mAc9+Ad7rzTNVv1eXMJ+pN7CPrN7ZYuU6fb509kNsUS0
sEvmFe4IBUzUxE/E+qawpekXmV5vEVal/MVEqLAGzl0i0kRP2hT3K9nP/lTKwInm7hi/H4VOKRLb
e1lVpNWEdYYCZDI+HmVMzSFs3ImtFd6IB17bBkB/jNIrNY/d/uNPVAv5JTWJCMwE5M8q6v0C80Nn
QnegvennSK0nC/uqz6uJfbAXCqS0Tp+nncjvir8v354sGyi7jZvVyyy/iIVN8loH9GFEXwYuHram
A0ONgdKEk0rl1JJDT4yYwhOsP+nIkyZU9IuLKwJqFwUK5qkAej755FKvvcNoefx58kxMFLvNPiq1
EqlYSZLiJl1DKpXTEbheRvaPM/d+iZOwNUEzGOeYeZXakh/Ar4oMngmW7RbfJAc1PWo08n6dX4qJ
y6h+cszv33aRnkJ7ZNRL7fQmRey7X1TQoX6tKBD5eoM1/7wRQrEnrQVl2pnxO5aiUCIgPMvttcim
b1tVKwWj6N2gXgRFE+sdEUc4ZwPgVqB7oYBAq1YalODD1itj+o7tIpCbyee60LAKOOF+JodaAzrK
SGNwLT6tW6FdokuuqYw1UBEJakAc/fDbs3o5kX42mZsvvxDlMlIO7mRFsFSF83gM9enYw5my04xf
G2RzhnVnAbbPRdzbJEKTPtg3o/n1sSxlIneT9k6v9XwBwda+m/BF4jLvJ+HUfaWCHgTbBUkzheja
lGKC7r9syi4oYYtTqdSSdJOU0frfwRN4fgcDFtHeVntCiBHPhUruqcOSO9EYcsFBFJ+yXd+n3a5l
hC1iHPLOH9B3421dfBd1Vy+R9a4y6QWk5Q2ic8BzE+1q0V207J5H3bjVNGqqbq8obS9pkyNpqCWh
3wBdNhc2Cu9t1YNArOJG1rwqa+h9rkAsHeTHjbH3zcfZUJkgc9Ax/85Xy1OLB1jhz1vwp+Tx592Q
V4RvDNtvyiRN1rMDRtTzbzl4OsFSTKP9VmbzA489CsD3JwkS36bb/XmB3GVkIduLJPOukddc5Xa5
oITnzyXSYiV9HV5GLEn2yj78UOtZSsjVOip9hNjSJqYB47P6jkr6w9IPnO1mkaYdB1ToiZvo8ISw
kLH7KLORXvhqq+ok5R8Amxw/qzHocE5hwWP+xPQgGBLBjVCgLTUzTYMFSQc1rDpe3u+Sm+jlqOBK
VzvT1jSUQjw24O2a/WBKNmp43gF0CGozjqMCal8gJy2QwXG4KQOGMbi5ZfPXeRmTvzO2Ahy1iepc
qaITiuFhGmLqzAhxMY9B+AJGxYtRtcO8hOnG5ugQoPIH43GjZ4QdOCqpBCmeWCUThjVR0lSbHwM0
5loY6WXAqts0ewe1+2fvN4z8SumWOVLANCut4AMfc3e7hNvr6Yt66X0ia3+vThWzs3XFf7FGcIsm
JgiHNnR2vNXX+D9p7zSNmu49jmtq33J/jtFJ3SHnBaIibemuMN1AMDirXg4Vo5xUPQzedDg4pojs
9UDtsOP44FlP/aC9o8VRHhXHRe6yuxKy3qOo+Wj6MWDMDXleAv9zi4H8utj7asZWsSVJrICwZoDc
poPxzkJj6Q+L3j1Xcyz0hgF14TecTX6IUCPaqYsfZ2EbsrzYdnkoP2sERmsfVfEQX0HP48FwW831
d2Jh/UkcrWazXLwT256X06+k8GqW2ItzcifnWsOYOcytU0z0mEyw0Ig4xKgTI/5LCVrYT6YLYEp2
/2cNJrJnu9id9tZZcG4KIcn0UPn+tNBIsrVTLB2JUWKs8MAF+R1qFuIIKho00UtDQ4VBWJOzrOUv
NvzTbahm5ieN6aDsoIVn39glpVdVYBDVATjyKsdljOdPMpvicQ35wKyX7vmsHIu9TPEmd1Ym2fmL
b6BcLOVX1KnyBk9jH+LklWLzq5YvmBPKvRXgYRKHpFNcDD2a1ARQlpzZYdhF4tPEEJQGxKFQoc32
FpnF1g1KLrWU+1FlMyAE9QFB3tt6mE2UGoe3L2HxMj1/wJ4EzaKQ5OU1I5kr56Z03kG8p4UqyMe3
Kcz4EVnjsWcuDb3Ab0az3CWPatvJ846NPnDnY2FcdIzju7khjTkly5r5SHftpH0elc97LQ45s8sj
mtSL5w9b6/+GKBa0IftInu4zRCTKuX7ZiFodCdPj8/oSflFX5zfUQcOkcj1KwXqwpNcLtG/LMBo/
r3fBTPEJWE1b5vXGiSHpuuaA3PfBBWg0xjQPYyMLNIMmJIeWj4xxoExZETFSpQ9RzY/pSuzc5gnI
nBnDwuoYUZ3udsShRVgwnBT4a3eVzgy0erPCHrIHJRxtdmw277xyb7fuuInTr0OmCajraywqgwqn
DSNaKyMVkLWhvMGbK1O433UWZCmvUMViKe09WaJOT2q3OEkJnS/PMNzreCzUyQm1PLuvah0vs8QN
chPKNlz57GoYQw0O7KyyoWywavh9f56MXX7UHYvD6A9Hx11iGJWHEmS5KtqK6n+pT6w7MhfYmTA1
MHE6u4ByW/Z3K83XTh1XBDaIvSJ8U2fpZnfOZwL9XqSAHDO/01oF2bW+YvumLgudN57I4dSh/kqt
qFOU+K7DBqpd1vJS+ZnjzC7J4gGoHZcfLXkxNI18zviiyBAevwGx5IKF9kdT8EcHDMcHDiOSXtle
D3Kg467Mh2iKJf4nS6RkhdnYcHGB96/n0aSsexFTDUsmje/lh8qp13zEDWYlKOr1pqecriGACmaU
W5nPUmh2EcSKoyfeyOyTZCbn8MtW/UQ/WsEOCSQdoEKfXzYNCmzDhfFo+po7W8kvPS8u85tLCC1o
myKKDSXjegBZhawn46TUwOQocl+lBNbujSyXhZZuUtoyOzA9uitdHPCr5CnBNK75OhwVkRQDzm2L
PwGKioBVy2s/xrCzpFd5mxkeoLy29eW1GQ2YLzdlC6ucUoo+k1cxYLBtJXMIl0+TEXKstl9k4yd6
m4XHThHaY8xjLDPmsVIfbedWKKawiEucvKZZm9MM/k9EjWqLovuI3+Q3Q4xi8Ep8IqnEoy52rfN8
eiBkT2+30V14tHYZUrAhpZn+nDegkiPd/UQn/DdXZSY8+tUv7+s7Pf3dm4dFhKv7GaLnvYy7sJOX
oILoptj9H1R1RZ35o1TCnheudAULk1U1PkL6n8oFPIlQBmwY5+B1pHEbPVXlSczXgX3J8tOUb2H2
peBpkRTzMmIlC3gVFS80i6euHR+cfeaCkgCf3D7UoJ+F1Z1Cukewkkwp03zhV602/i+ZwtSHGOOM
MZLIOjJj96Gy+sUj0uFhiU4X12yyb8ZBiyMc7TfdG+AepzxHnQJD5qcY/JyuVskbzY6hutIcKSpF
N87UFr3UmcIuu4LAQvhOEd741I3eUoP4A9KlWBRLAhQ1tmnFGoQyptjZeQNrOnHC45l20+xo8Bvp
dPm25YUVsbSF9IBgbUwG9qKCTAGvoIChxcMucgUY64c9dxAWET3S5QUUsy5N2HwzKp4ZKEfHQ4Ji
sJs+9Fx9D/Npw2ckeAHLmUI5m66K7YaH4o+lCMGSeSfaBIC9/IzQgIaNA+qcmnT0eGCWol6jbLOm
yX32ahUDGDmtak3yyZJOANGzV41+DGSwWlOF1o6ZRNbn2QT5ls7OotCHhXfJVySIHVrOiG/Ziwbv
v7tlm9QCrgDYYViSj+Tk+673KRZGE2RmWPrsLPlf2sWDfrftc5QdjjbWcFejVg5vqeX/b+8hvHxd
0bAsCBjFnIF97nYYcQeby4tBRlf5CEcQbXfC5Jp16MJm/AkFAoDsm39UiECs1eprIuvwJRL/y/nf
LtCFczWSQ0BRADyWYoshyZXqLDCF7BwNKRJ7vrweQF9MzA6H9svM9Kb0TEfysseqmEVbb8PO6J14
vlFAtEFLPz5daERX0rOqQ+1d6O+xsCkolyz+Gyn88MQR96z1Li9sE7PxluKWbrV9BXUFZhbapAk/
b4cWuL9cNaEYa28mrC+WacMjNkMGkz8Am/K+sgb1fnTRpqQIoniJbsl3o/Jdofe3EDGchDbcSdPQ
rY4ewBecf1TtiCQopTn5EOCo6yuBqfY+Z/zHv4ZJjj6rruFYlHciupgFfwe8rDMfR1SSuT/zkif8
uFpB3Lp6xbmbtajDfsSENh9enYWVkwiz9JF2GulUlGBV7gGPpMicpP73ThIyN3gMzAZ7YXt7R03h
L/e5/+LC2+vsGVjzySlIVSIqBke4Lgn3meu+gxDIprIK/c97i6/jKz1An+NcwpVcyJZQhhmhF12v
Kbkyb3uhaPaIn4lR5m/1dEpWt1204WOx5ZZTMyWXdgWDuQ4d5aCq3RqJe4KM4orimTO9rQQM4Oxv
aW5a0YWF3G6xM6zQFanORDHg6ARL8B6u24M6mA34ONFpv1/cGbKhM1icyNh4+9GseeU3LLfYxKZx
a6WFqINefGl0vVwFybgPLAYbt5iwvVZK3d81VtXBexJM27aaOOhUkH/QrVVpsZrpmYVxyYmIz2ih
z1Xuk5wZPQJHtpQW/10KHQ5cF/wskzQWmbjO1lJMaS6bQH+ljPSo4oMOvSvzbsYF0Umz9PSSalOP
pA3BVzj2W7UGoA90s15ixYj9/j71fgXLhthqbiZQ0isoaAuYs5nHBY0GoqNDWM/8hEQKhvvUfQiG
Jr4OPlVK/fc0+Jcg2CCyL3cTeVKSEK44D7UrnkWwvRqhQVCbqdIl2XnyS2TAg3CYiYPGPQ8uVQzo
mMMUcadkVL6clJ3HLMTRMXFgm3SRYHhALdgu8mLNIq2/G2kwKSmeRG+1QZX8irV4YNS7mByOBkxk
CUMnDvXmvNmPuGqwlYcbrsYUU8Q4vTc+qjRb/dgF7O9U4AOSG2R1Sp0FDpehSPwJTKJ0mrvTTjGW
GpoAWwjvv+9riwK1z6OuYBHZVQ0UaMaeZZ+iWexK+vphpqdWf0ooCp7TFNe/dPta8N5eU6esmVNo
T7mO37B4S/6wPv+gMoD2G7tnqX8GXitF6YjtB9IIF8ycmnwfRGZYXkzinMmjGcR0vaOHJvFG0VFk
VeFNw+34DZCrfFcnBMWEVzWqeTmi3bZ4Au/XzOtzgGVWIn5vR+SwuDI2q2+RHYvGT/FLz9xd/Xy3
l1svT1SYZ5p55HntwGG5F8g5XZ58JdyNUrb9OXDbS1zBYfnjd2o9uInWaZT9vovz4BIZjIdW7WuH
3m+7h6OG6JcvhaGxQA4PYhM5IFkJZ2H8U3bCFrlsyRqJZl4qcXjCRlUcxs6GMe0kCknJXhkda/00
c2g2o4R9dQ7DMccV0gDGu+T52BUa4OSkbri0XJ2B1UdegkpMpUrWao48ZFIMWSdI1xF1NxvBno9r
CICg6oQ36TGaqB4MCo4oBLrAf1h4iNzlhvyjE8/Swziv658TiO/uALezY+wsOOa8yigOtOGUqvw3
Nw+Jch8o3rhHIoS6nA4Jwk1VfGFiL9yhNULsvEH9oMH9zzU67e10VT1ZtN5QpA6WKkQ3WxAgW6DK
/mR92+9N1Wgjik/3EP72E+nGUgisPZU12UKe+UuOsKCp1E1nFAEwe4UbM9y++WyfJeHdJj7h+30f
mjWNjbXCdpaRl+xpnqWdjMw0a2UfYOuRltw5S1X7b9GapTVT0M238wU0WYkxGBW43IEfVmlZAicZ
AcIkVtdPNIJ3WiImxa7YwG0UVmHtasYQ3/QNOLcooCdUMlBpJdniPHD/naIcCZMJerJB19weLvxE
rQ9kye+Thw7cC8eGjpxfixsMHluG7PfzvFJKE2E4e/5bbDoeJqzJT/D5HfOIo/w3p9f7/ijb7qqZ
bQ13Zt8LlcXuxihv8rlkW4ixctxtVvm34BLT4JCA6WN4VDztPUxIJ66+jUaUkFOnUjw1J/T7iL0Y
wLTucbN8vTQF4jL+jgBgUYEbY+RjHQK8Nydrl7BxSE0oGLyz2+l7cUOFyYp21qgpb8DWt8VwCC1p
RSoCA351GmOKeoU7Rd0YTeVDPbCICpocHJGQMBx35PhkhUB83erJgKIpWAKAUaOQRAe+Dll5PxED
ugQNaIUvYAdYgcuFANtbSNpHK2PJVeab1ndc0opq6G+hD03O49pa9cY8zNUE9sGUGGEXKvZbrKi4
WmVzGfSmldhQRHPpvzHjILd7521z3L2scvvQCu/13SuQl5a/zXJUpCyqKbGy+X0jcKvkRdmmHYM0
9C37io1f2k8eFjUzJjN+krjFdCpgjr164a+fhZsU2e3yVVbs8Csmm2In/SuU3vJvpMgHfg1adoR4
jVyRndRVXHuI2/AGtCnQgu9ZcI91Ih8fW8ZU3Ut7MPjTDIwGtpByEXMOBY/S6H41ri0bRhA3dSYz
wUOvevnmCHXNyh+11e2TlBIGCpx65ROKwvI17qp5jLjY1atE6Kkfo9wErAv3tvnAXRXaOnt3n6ZA
cVx8dkNkmdCbBQd08cbo4f8TSPN6C8fXIEPblCZdQFftSQ5qO98J/9/tRr+sThoNaWoM5mMyLzLK
y4opaH8NoQkzYVpf8kYB/My+HdmKQvZcuoIM/hSsBJfFPGbOt+No8Jj3OA6Id5lTVNaIHZnsn6X5
JAtR922Coi4Gk252jL8lK2Bg4AFmFJTPF7oAERhtf7A0wYiVResH7BewT7haDDqXh3XiRnwGjUHt
BMX6976vS8I/Q+ezgaN+dLYBvb22rSiwx2vRF1y/+AXAUoddnLL5TrMuljv6eTn6ADcBerukdUNN
RUp8k1k73ZTAS7q+hh4iJT7OdRCEC4z0vRDeU4zGmNI3QvvsZ++KlYPoMtiDeGvAvlHhZQkDDi2K
VpdWYCiJ6Sz1rYdNfGAwjIsbpcf5Xf6oaQa1DAep/C8trsTTIU3dTi9OFYErq+8YNiMpjckYenL1
0Jx4SdEG2iGQqYD3ffM3YX5v3+PN/NL8HwAhASifdDhj6hw6EZKPKGRISMGF3jzjKYoBQw2CPVp9
JyXhiuIT5kkYiHhSqniwvlSi/i9OxTbm1P8ILAa/CL58CJ/ci826mIwGrIHUJxev8CMAW+GUVFwX
qYGeIt2PAVKBsKFGlvT1n9ifoUmAMM4FaM918KEMmXKf/4gqNfPZowKDgGDOIh6eM/uizbgEkX4v
71F6JBqxidfjxCfCZ946wf5c9BjeaT9yfBr4wxY6a/K6/b7xHi5hPpk5MBYHyiWbqjGnvpuPapqk
/D+aZ4oRM7/rdGuIV6H0+Qn4OBg8uY2mO9K+hl9ktna0dWtzCpg4HdJ4+zv4nRCxsidiDMzERQMl
Sbv518EP1Z8Y5KyGePZPTdB09R2bDMuaZEeCWjZb5oI+FeT+9j+2O8Rwvx5vhaNY2/Q872HDn16z
9Qwqr312PlZ65siSch3Kz2PXmV6IjfQxBfJDjKb/Pfbdcl7agfzUT3B/BgURGGmRnMywxQlUd60p
dGPFOSg5TwzUI3J0st8OkFBPZg9vumsas524sW3Nukk/noL39RhgFP2agGjOPP22pq4UXp5BOnWi
Gznb90zAb5SDJIItpPZiKCcd+h4G5jWcsAJWvuAMA2yfj/rXvhM4bP7j03kdtFwiw2fn6orIRjlD
Jjl+RmorKu48ZRYl4bCCV+3n6S1QqkbUiAtJnWT1Tg+R17GV7UH9OzzCRYp3k6jzRpOPtEA8bKp7
xpxQ272mZ1gDEb3NBwvj73WCzoKv3Bjt/mh2rzQfQcY+K4eFNOekGZR5nLU7Jjzg2jE3WyQh9ghY
KbdEtPtiz9hI2v3F0dy18epQx5p7RhufyYVzZ2ipqu/WkL1CT129dY1AuAUi02ReU91usy2jq/lA
dCZIJkr/YyFMEy/m1chag4xc7guXg7/L6eZQ8TH9TPVXcaiJxFtj9Ey9qey7aBZ6DWxWJRAlq1XM
yMVlhijuESEIdGmkKTuodn4RUpOlZwr/1+3eVuW6fM8SHK2mPHTFFzDYYIr/oAZKKTwhgDr942G0
pX3bqbmqFxdSuCIh/dEBX85DwcvtPMg93NjPr32wQF389CjfB9KqLbCXTO7p7++CTJnsxyrWLVhQ
N50jTQXqeODIjglpYRQQbCb+d/Un/O6iFrmT3VBSGGT6+F+iy5WO/H8Ytqwu5iZst2VH/xoR6URu
+wCjVm2cGZK0Fr/iQGqgfJYTKtoFY7PkPFqhnW+b+s1XPJ7EwXI9+1fQEtIe3FuN6h69s36r+ZOU
hV+ufG7jmrTferDETf3TZ26/41FLnEG8IWUKZSq8bdoux5DCwCgz5fZwJPx4NioSu712tqIc5tfA
+SEJMde0Ggk4Zh0UJgniXP9lfunfefSuqttVwHoAej435D9k4cIW9i9GAozzrqjXdWNVYx8u6kgx
7kiOJ1NK9DTAlssXAgj78y2NjdUvQa90mmjMYCpfgyRK3L3f8NVpWRCsh06P/LvJeyGr/iEa6bcd
HJQgDQqkdH6KzpFxpT5/20t7QfTUa3SSiWW+mS3AzQbp5XOLfZUwDcZ9m0PFQV0Tn3waaQmRQAqS
71pm9+1VoSjAdaw70ao+OKIqzx0pcJ27+pfLNbuq16E2aZffas9AcHkj3dAQXFzetdXAoMMdL4kq
igBf/vr3btX3SlTZkvbPNOU8+sCNSvPE4qZlmMPh3VP1JdfsyTMIfXztSG0FpOLCgqoCupCjXdZD
8tM4uwRqRbNNjj59WDBBntv1gOW6fZmy4sfqCQsffbdGqa0YTdvzE7VvNtk9v4HYCr7/BMtCunsu
zdUSxayOOY09ujcpxw23yVhDRyjq3Q9e5ueZrge2EJFOvttTaXrOQxJOaRjKF2ne5yY+/NPVhdhG
w1sDd9ZXgcnub2CXMT9Vp/OG3uZx4Ao+rKh92CR7MJqnCxv43O2u2GWQtWxoGKN4ZIPweuVYTRPR
+6S6sj9uhf2U7umfT7CqI5xI5WaeUdVUSBnI7Vxlftv/I7va7QLsTnZAf6A7nlxFTMqws6mKBocA
/7GI1yJGanqtXhwGe/jOoIt9UDnkYNq35OVTBnIWxZFElEAQw8AK796s7LG4y0g3yc1Dfni81NUP
6gdjZxxcEYM9SpcpwGcJ9yNGw6Jre28pmaHPTgSmUaWAUWjYgjQZ/X5brs13yINkldzxafU6w4ve
2dqKCATzhER3IsFpSzCeXG0p0Y3y5T8gCz3x5Gzw7a2pbh2270mTe15yxd5kFHGoetcRscQ/wzdV
APLUGtOF3lq8n9UKE2rzaTs/OwzSha7apCF3JlhF9g88RyBTh89zvA0ci5FtiNoBoZyX7eklH536
a54wFtgJCZzEewZxuZwiYozbG7+1nUjxYV7dAktlBRxHtXSrLBy9qZkTc6xKYjkbrIGVEB8HDCnD
qyuGeqVAopO0gevvkcTrK6fwJR6CFfl61rvy4vstDdL85zuAPTXyy+8uvUtwt4QK4c3EraOnBV2o
HOdL1j0k0ZIQ8SfwI6f7IncxlTJ2ZvAIGSWgw/NN7nwzyMtCgmNPJoCU/fwHjpq4MB4hYqIfxJJd
5llQwOz/5mrlzAbHw198EAqUMzSzNwVCKkOuz8Hl89gdlVPNpX9HZvpIt37rxGOU2Lvb3QJkQyc4
yilb7hsevCAGMVAy5yVodKmUg1GA9QeNrz54wmMkVjzSt5LdXhezgDpo/WQ0KJabExQvs6vh4Lla
wTe6pKaI0NhfYfEpUQC1Uq2FcMeuIrBHb6MlJX68VMKC/pkSaFN8i2WeUAdlmuJgX/kynaZ6oXxc
suaLhRvvmB4Fd/kgeAC0mg+aW0Rc9K+6O0lM2/YN1pdhxLU3a8hrhBZtIo0H10sN4A4W6mZIMX79
RY6WaCGj4jwCdPB3SdGLIrRBQ8/CWolU7q0JhrUWqgRK3gegk6RaVWkgb3DCyCmNiS1vdMkRI39u
i6hZYXGPhK1AmZnQNpjHS7hgI3JoxBRx0zAOTp5oupZE+jgF/O7fACuW1L3JVkxu4cYQ1Vntyb5E
MKdfPbtOCa54iIMUibtd/q+AXPjDxCwN3IihfbwHKYIj2b/3hsv2CfAq7jYK/rRexpVfMl04gcsW
Jkez6XJ+JIfSfGyOE1n9cID6/QlH1O223SZxnSkSKACREKVuZM8Scb6oJTGempCU+viggpH8G+J9
VoKOJIs1rQ1YKbCIP4/5s0K9zepi9CjW6YiTCsCrcL5GJCPGzQd4hGrz6bD8AXzgfUglzsks3l/x
kHOFER3R/HqiyfdtkJ0DE7aj16eGBOCLK4NdDpuF25K8fX5TeoVfglD35S6tYjVMS72p2KznkMHU
4Dj6kxKh2ZryJHi+H8wRvZ0t72Oc48KPUOXH+LDDJajSk8zP/SBJHaxf1Rm+OaDVlScB/izzwVF6
6UCM2iKJGae351Ntwh8apONCT8ZzOyvm3y3OJj7MEPGqfvYhTEFfKxxTtk5wb5TEJpKYCZNwhmOK
qyfLZO116h6nLsrM4UuapJxaemUWsmsuK3z3XTWpoHjYUuM/s3gJTsv/qWsTk4ZOdHNBEiBPefSO
aSGiG+DwB6Pu713XnnpVCukIh784BMLW5UdagMbltPHsDq8LVqKOhG3f0IPbd5qFN4ZZsijJ4tLL
+MJftiqNYSc9DWl8XfBgkLLD3U2ZtQUkhhHfK54k6RfOxlfhBYSHtQb0B8EeZGADXP/TJQYo2M1+
/JrCCGLF+qfyrAFxMWOqAuq0YNJ5cF1f1sBnOsGfb0hzkRNL0nIlRqqUDKV1+0JbIYTpFnB3kx2v
M4A9QXdMNeTd1vmAJHz2rYWv4L5ZmVLFFRhyhdHnUWjoyswKvV5SPxx2XoRhvRGnc/1D0ZfPrdAc
PfmBo0HPweLDXS01NDAC/eK0S1Rmed4wdNpAJlzmEklT07BmIbZE8w3K4gfY2yYt9kUscO1lQFeB
KZ2PXUalY2k66kTfBoV+FpiftfqNX6L3ID3Gvazcik4BedMkUgnQKxsJAwnYqTueYyZYGBaUfCOC
wUMookIHJ6q/D/0ab8xwVUPYfu02Mq9Aa1eBFjdJFsOejDhNsu+CyaxeFXVd6em8Bl2fYjCtCwqg
IhzsnmURSWfSjUJIbzvvVJMy9gYGf65pNmH6dAjfNl+72U36K6C90jKzeUu2ol/feyN/xYJaOBXh
sdwj8Vfn2UKJr9Ldl9ZSUKMYgokaMrGqi/41G9Q4uRfjwxoCQEynipCtrXnDdujDruoG1UP2xixg
13Dp1ANfJujOLfHAQHruAgAikLU3PKDXnu+tw9BBqbdxYlnLXLmUUYFUpnzezNL5kIm5WkYAHb07
ZfK5zsLtSoDiK1+WsVbj2KKF7c1MD5hSiJbDXTpnjMbFp/mgmAGAFmA8wTjpyM//lUfSDSmoA+2Z
m/wq4F6hfj5pH+0OajfCTPaRXLuY/MEzCktTAbW08RWV/HD2lywjpliUu3cDIAwn7EfegrU/xRJf
t7YPdL2NHKkisipxoMnYfAKeY3xSMkyoXw/iHuMLm/xfqTMCnyayJxlweSERMMr1+rRVh3VvG6Ra
g9KE11jZbI4UK2tdpXAfmJM1pK9sWDCzO6zGz35OmCU2lnxF7TSdJ2nfRv8EELiArlUQs5+rCSy0
hkixp93xa/yyoTIPpGcSI/eEV7YdpzYZIySpGr3F4VDpoFyGPGM3Ow615+2P3aJ8S/jIgCMiK4c7
6wjB58jXmR7xnDR45ZF73WtpWBGyZlwWJvWHfN97b9c0xiLAobFGtGL6Hp2+lfkg2ofavl9o5hrg
n6ALQY3i1jfjtptk2cuS59LtPkzovNi6kc0lEZqvulNwtdT9gJDUbu5rZOZ+aA3QeBrJvn75yULX
gWEhSACowbLzolR5ZT5EQQ5cS0TF7yoldTXCCwvZImM2oTeYtV/JMrV2APUYJwIGneYWFMF/7Emf
YqMQo/e0woMuS6Rb4qiM7OF+5gwfNVgWKc4SXlNacsYi6JzvQ4eUmgVq44n3v1nuuHCM2ZK9ExcH
JAN6QrNAD/6jNZWiSvkZI9bBc+52htm2VE5niIWCsrdRsQrDvMs6o9T2qXdY0QcgolCXvMhqUbso
D6OGvCzxGiQZYeiEDFBHXxF93PJJlS/N+YjG9AX6fdbaoVkAa5Jk510TD6AMGKb6tZ7AR5Q6zTpG
PulWk3Smmp8YlqkhV1KpWgqMC6Y1/P2qP9IYxKEt9SWfw/ZvS5qvkAni3P9vXearf9nTim+gIyqX
I5q38gPTR50nWaaE0QFZ4nhWtLJwaYEimNLXyPzQ3ogvFvY4ikU/dqvLc2grLebTKHeagGDwl+RI
l4e0ZYUB1cWp6cemikd7oCKsoO12JA4ndYY4qlvPyNhOcwUtw9hHlKekrvMa6Udm644omxY+2AvF
A9M56vozoaNUQzvBpbz7PvlrdvDpb63HIBKO89T1fqQV5mjaWbE2jg7L//6c+OjUIqSu114z0e0M
VxCX1IBl6FqV5Eh5B+J+fZLAVQoCyz+dI4PI40OCb3SY8GNv+cic9kfnk5XWhGloifNQsCTZGBWP
oSCrv756cHpgIwR5dkBRwFsZ+RLcKm5m6InnCCvj2k9xTK0P4E5jUsdXtZ+txIVng0aFdfJ9zeP3
+k2LhA7A8dPx9D8GVPMhC6wYMmAUNfM6EXOA1V9GnNObWJMmzTG8388P45Rp2j2y8fUJyObfMZrW
2TFrijVPDLwoSafTb/uoiLr9BGVuLe3KYm8aUal9A1G/jAZcoUIEbUuOrp8IfWUoWWbaBvReulyx
Q55ww3Ql94H0Yq/dwjp2MKBptwQbeqzKczr4AnRtcCm6tLz1PASC5kDwilhcbjfV0LbmH1A2+5Qh
uF8HcnWCdy9TVhtpd8z+ryWgkK4/KvG+wOGphdG7jzxtMNcr01QxObC/LzmnldQHc0+Xmkgg0wJt
5sw/Zl7jKMnBTvqIXmUgaEAl/XOg1g+NNiLMmcIWDsf0NobsoZJpW5MyTQnzhTpZyX2hYvOqAoe7
IrZTfeWE0BsQ1j4xUWGr7lUHMITDSZLGCzsR32hwBPONxMVQEZ20gbCsbMTo0K5TnCYfoY3YAQd5
1RrkwPrnfOSiY+5QgtgEkT6//U5F09hnVMjdU4F8j1q/RZ+H2cghFkXLti0l12aPTGIVfZoTMPSO
MjJ2FLTXJEWB9dKjTuQB9YhIG+hGQCtWkmWy+qvP6DmURXrtsdtanjRm4bnY2R2TfmznGZqY28eu
pomTiDbtkU0skyt2xGFQY6WwO4M0AhoqwZPxwKGXT0KqhxPGBsj+WMly8MzXhPsN7ootJg1+MHca
X7Mjf85eOjT3tapOu0OJkyU1BHDqeBg53ffUlnGBL69RbEYZYyIJJtNai+HR0JsoFSXc3DYJir9A
aAPwJxTJyj/OAHDV4c4KJU9JRODiWr5BCReDeuAwXPPMDO4g047j8tQmTHynRrzbypgWib7nf2N1
uf/CoKi+r0GmEP99mhq+hNK4cVyQmHi7F+ToxxpcGwBg68/8gjQgxafzdnTpe3mcp7ipce2k/8v8
3WY3kOskvTW4AoObygoYUBmKGa4RtVvugZZ2JnRqqFUBZgKNnH7rkIdxuhJjE+aw/SOzcJlJgRNc
ak0T6Xdpm2yz69Dm0IQd6KWroFBNFH0y6hUmDcWoWI3ecOpOg1v+TJbmcytHrUlpHbCe95o/UYRU
K5wvfUo4OKtaNon3AFF04e+sS3FJYdq92+sqvw/FI9DoXsnUoFgu/7G2r4APnBq+yEleKFJRQ1JI
V74w9sO/WooAH/TvezKasgoJS0RIM4ElCNVC0Hx8lYyAQWzaBccWjsSYuUSYeyNyv9K5u/SqnjA6
RuIQ2bNjz6hoZiphxrLNHTWSZXQmBuoiZ2wtOtE/QRz2THJZgZ9XzPwf2sUtNFNXEa8dAJUhPNBR
efAHy40heUEn4Ku8ZSyIDHe1Y499Bgv2l7ri876DL8j41fKN6J/8r3/O/gFrNl6Whj+dIVSZ70yY
05rHVF7JnYUnpgTH1U67c5N2d54uX3AKKTkYsJj+AOgZLxV7ixA0DcqL8mEmJ/m5ujg1eTahjGhA
7ZeVhSmDzoqA3+0You4FA7tNDH6XKHJOvLTOQBVUls2ywQ7FiThG2iIAUx3C/16zV+MvWd//W0cn
yM8dsU/bkORzXFZHhyXES1U9egmQzO/zLUcKvVkyLE0SjOSSfuOfyuwLpOCix8287bKLUr1uZ9Vt
MV5nP4ARdCxqk8uvSYgvIdOxS78L8HodClk4YV31jiumbRhsbdCEsHC21PHreaIfsMIsu2F/384M
nNwEVo7DvOzA1hbTNVadD0RcKbY5wajO1d8pi2EAtlPUrapHXoyICJicZw1sIF7y2GL1sA9VbavS
5JVnG+M/71CPrBJtmt7Ew7E1qvKQM0pnNGGmmes0T79fHnxWJGOS36gn1WLeSHZyP3aeEZ0+Vxsp
SCSk68T8ii7IdUqUvOMkyom7Hmu7A3JruYKElaiOTAUXFLDXtRe4HP4UN/64hkY8nPvzKHH/KS6u
IOmb+MjO4N0iEO1ZuD1In+FUmcoljt6i12omzakq3OA174+CszRRVimi9KrawBUstRXACZJSi9p9
pPEz+klE+DWCxRE0+jQiv5IkcGnjnTmYy9NUcwkhgELW16ctt+IIKEG//UmU5oPm4v4ih78zta1j
rMKBWkWOY9+LetbhVFSaQ9vTgHesWjfN/+OTE7j12Q0p9VH9951+4tQfA5GV+5kLAFxqPRt/9Ku9
+gjNMTlffyhBanuI/ZWVsStDiePp4TkvrX/FYT7yODrLCmSpCNCInkmzgx8c+lJzNVB/JyyjsrKW
ZpNhZNgHQ5j2n8qbPZTzC4ZfUmH8Jt0HTWhLcoYtjNdTpKABoQBnRSMR89TZxWHS4BvRt6cpbmaF
os5gzxlhmS9az6Z5wdoHTsOeqvOFFt6N9rwj67fSf05QgpgW24dGafsQ7ULhaHl5CjDQTw0Fzx0G
u4gCPqbVHFO0cLnRu+03Chq7+nojS4WeweFqtniIsTBfe5f+CLFH1faM+TwjlqW73llv63cUk5GK
cX6u5GjTNCYcVcctzSGfM6ePh9+D0+l726A8/74J4/VCKrFwaiQkloVMx/s+h/lx347yzNaxPx8h
5Q7xAjMXKrCr0a8vHIMuX00A9NSJcUTSRF04niAxV9WVXddZLUAzvT29GUMWjVJhyLpQcfJb/UuS
vkyt9MZgCSm/6yt5pe2KhWw16VbKo6oo3GATHkJ81LqLHJKT5Z8T+jyy/siBxpCIwep8jN5hTvnI
Cfhe/8oC3ZX/YkioedX1JJB/DObbkPyMgEXE4vgLIHZf6uqxTcwmMmvExyCu7ajKMx51EntD3KbS
aIrOnAgbgbyg9vdVice2nAIdBQPM/z1Q/ckG976Ic7zRS9nICg1nk3Z8DNbB82vNjYm29WXcgXa0
MHX5QaQOvJ5USg6Glw88Kq8KRNEYbiJeAWorNr61Rg38vW3vqWZ7mN4YYDtNnKdNrtU++4h0Rqch
XHlNWOSreFmHeTmKgRLo4+Qa7LxaUK8MfGdZcDiuA3ixN6dMtE5HBYCkCVrIP/C63sg6zxwLAmA+
DE9PICBGw9WEjqFODBuA8zZGzXZ1IDWH43ItuT4iniFm2c79zkimRaJ47MHsrvWznR4RFJauX8oq
HjGpONAyKO7zEUzWkW4EG7UrgFExjyGtqo1ooYAzPRO9vAMvUAGoboGEGUy0FBp+kVvQUDrX9UXM
b78hZnl/z6FjEir+uwMCO7kRkrdCXqSFS9YyKkKJvIKL3TLRIGj0kHKAnqrb7GvekQYVtP/6FkYT
HAImECVeEt48PDz0GzhSq+DiL0/6hl+fHwA6OG9OEcXbjNKA33JXKiz3VSAbEuf7i1rAxNL5uoWP
rPjjN8rrOVz5edUEvFwsyHtKe/xuI9hsa/g30EoVIdYBAp6mFNu1ppNd7AuvShWE9kR0qAkaiDDv
e5mDnlPecDxMCSKCOxnzVowQ8bIhRk0ZKsud7C2FP04hD3QBsxAuIFpnuiAa0AIefeglc3MeLDNB
EqPJPkXhlrysWPXN9vJEVNYRAixpLVacJCHc2uimNT7EJQg2S/4rJivbV75ZoJKXisztQXn8i6zn
a5tU4gZdYMVwivyO2gqodKBL/UoShYxdqeahvd9C6LLm5E0SH2Yrdwu43d023GiU5WlfPs3ZtxJC
uxIRAz9zZZ+G/fQkmRE1OQov0L9RB1+eStCXhs73Vglu4lz3df+xRXrBkmcG+KIAQudaOKLr1Eam
WwiuRfpyJ03AalL9rF3qPjfyOWXzIfABVKtlbd2YUfGKvmmbY5p4i6RmoGW32EmxLDeESxGZia2H
3Z1wMaaG2yN1loVQ9faDxM44fYQtY6v7hMTJauGVrKjQzjmK1xJ1KwDFBEL8oklEX8Igb3iqiE6/
YdxUiwAM0Xa6P3e+fgq5wNxEr6PtcOHtRQ6iZiZ0NtstsK21fcUnk04Zn3b9cuzlttBX4hVt2FQ4
JBpyFmBI05gNpArg3h0fZHViou36JuhSa0uvgKFVf6/ys2pOJgb5jDbFxFi3ywX1F/ZuqouO2dCj
uX03pPvZDX5CcYC01LeSWfDE34PJU+cIodLg6Oz2VdwQft3OJZp575li/0DgMcdvMOJzPM5L0+Tq
arxTaogX80IMWo9N0pecWLCcD7m2LjoS35Ycx4n9e9nCw/cW473LIA/g+E6azcKMdUCwJ/NGFYkN
GbKYtUi+zGgwNyONdOvAvnNroE/VcGKDMxVhNRGhuuggc7P1h5zWpPCor/1HErCJ825da+AesJ4i
V+5c2hjp0QNRs7hmp1c81lnVvqiSxLBUKbRqfR3nr913/59ekMowZWrVh7nnOFauAqbcheVzNOIM
MjA9jzfUDMtOsgVijC5TOYY9s1CKRZql9rcAgCC4c4DAGMZpadDp/0vbZzCsNLW4HM6RSnL6R7YA
WP/kfo5zhqUvGRyAT8zn2+Qjzo3JmuijBzCl2fsf4qyTqVmbjBisotKszGCA1vRismo3n+78cUbl
AM6apqaadnvTcEKmVQki/dw67+Z6tOpUcZSx6X+nT1IPPrJ7mkA/Wio8hIB+nKk8hzXILu4Mj40C
UfQDN62e9nFgYb4ixiiIdyxCoPl66UNSvW3kMzwkEsAk4cw420DqL5HABPrG1Z6wugpj2RzM839l
/7aKJ6haPcy837DfzR7QVfp5sjd6CWgB6kjdrfpb2hduQQKtiLr3Gf84c6T7UxIlABeYLMJAdYgp
fh/iKSPG4oiCrOGGiZUWb9pE5+CmZLPnVlqL+U8SBWDUach3iWCgGcz8CGvATr1RT5SPoOStMFcK
rSDGbU5oG53wQUFgXIlZoVUzS9ySXh0yG+xmJpcpc495JDxtxAkBZkoXGbCYO3m0WshMNlqCBAKy
DIDJVzbSjqABjTF3sw82EaD39kqxx+0NR5s4C1QXRNasg3FlhnjMhYO5cvVq57+dPLejZKAbj9DX
iPlui5sqNSIACmCrXRk/5+aWAo0Cstx+zMWMxNPQFb/NMDTngDP6Q8ZWQvTDgevGG5+1ga1pDnMs
4yTx9zeS+JT93X+Nchrqp5/9dVok8rNwpSPh0JQRGMm/LPwJ6IqCIgqXN9C8iFWZkuMy0ZyznYgw
za7BotnJ5N1dREqnUHAkqBLssNgHLGfWxGT1NIUyLmM+sM249elu+R7aVYhmSU6qKn8yW5c5kK7J
hGJI3vuqXopJmAhBv7tLOYBHP302rLOsJWHYiCnH7+mlr+Y7NtBC9aEDbofyYCf7PAlWS4qXJYSA
dEX0Pk/bfCd9RW68HeTecb0kab6rbWtUmVR8JB6K76wFgTdmfad52jnhv1Y2XCWPsKQXW9VwNgH/
IIph/izPbYCTqIu87vr+Ml1Oth3ZXqIN3VQn81YNaWhhuOW7sAapJKrPtyIpzLFRPj43y72EmozB
jrzwyMc3G/BCdKjiZ2LNYOofRluTKIwpXbnmwX4ZrsJofVFP2xbHUy9SL5waVBvo3irL/dQ2qg9L
vf71UUihbPvIYjNy1BZcH5FERgeSSJ9Hb24LMZKFOsIGRPT0KkE822Q61t2pJ2g88oQMfzdrEqne
FPBpTLbv88yidEhjyQaSreBejRkmlnKjTgUtisn3OlnZjrW7hgqABu3J6hW45+dSVu/CpjDooVfU
fQURydmX+aSPfkJmx3hlla4Coezn/4AzQdoOPj6n6s+tpZ70jYilxd6Znt/S/jrROxY3lUVbXQMm
zvOrJfEFSryHYNztsZzx9lU6rGwJL6IWkzAFwzhrQh9xMxcfR8Yg8wpZN2jMU0aElc3nxFhVe6oK
2eNfbWIHpel0o1ONuHprvUCZB+aPDk5ercGHq4z/EoYfKWpO2Ax4QQCeLnEpJCadAXlS4GkJrdX3
+sfqgyWS7bMio7ZekSAxXLVjM3m3Ib6NfRResjde7DUOSo+tuo29erqpqI46FNKLHmZgveQCuxi8
IW5eUUZHElCGu2uoTdPGtAjfBHrT3UNQzSeoI0c0jWf7f7J91yJp9ndbUbNm65S9aVxUwpWksSU+
lBP1nIZ43rc5/Y4lYhr2xmVhMrZf2nZuoyAjsaF798+pc5fKmqqD/q5+S4udwn8jaYKUyTNR6JsT
ThWkhuwZL7whNE7QnmJSmQfFz+CFt4yOnkPvRlU7iw9hy6D4K6ZiPgeS4Fif9WzLutWW+QKrslLQ
whfH+TIwqns9XsQL9mxUa3LmbWdycvtJxlFm7dRWSJqvaf3ciDdZd48UEc5iPDkwlUv4E/vjsUFX
eV3iVLY1TNE89BlaUq0ZKGAb8Z+69anIBl/DwzhNZ7s17Akeos93ValNcpQEhJDfjJ6MaH5S0hYI
yVUDIrDcP+B3LYmJzvGT8jWdx94V8Jhn1BBUNQLMoRKz1UkhqF3WBhEB1fNtnMohf9zCIOPf9C6D
V/s5EG3NP8OLKRnTVt7zmLDyVWlGzvQAzbKyll4i/Cc6T+nJPfFo53jhrywrnwiXSVJpVIOS+uAM
wkRlpUi6HZ7ynqLeoo1YiW1gm2ItYrl9Z7pNCx4S3wvKlVYQ8jcnMmjLiONnZ235rK6JZWjYnCMG
3EKNUPro06qY9mgrEXe8UcdD91PnVai3uxdnWSnVi8qOclDwNNwR7zbGotQ4vTMfYcb0em2xVADB
1MdevJU4DiOUf3t1HrJgEAEtL74qe/fVC+uqEpLAHGFeFbJDmfDWv9LRizmyxy/BsfSekKC+9QFW
LyrO+EXBtAz3cG71cbULlnps8JFrj8GdQWBhwfzQdIpr2A377gLTEh83Gd9OPx7V2ApoFfY2GQ7i
ySCTQPstaNd8qZcAuhFd37+OiOtzR1k3XCNy3eN1YfWqyH3QuLspK7xDV6+v1LzkzSq6xcR6YfR6
l7+GG4bb1ELdcskY+S79oDgyF8GGHJWZTJEOpjMByAIgT+8N3/MjmAr4xFeVfKb3TdWXO6M38PB6
25HnaOpcPwLzvw8zy7VxDxDAttF0hOdcQSpZCy2JSIZ3Q+aJwaIBtM4CsFL9uab8x7eV9Ph/cDyn
tolbSCNPbzwskJGRCYVoOZlvvLLvwvpXlaPpfcFt8xgSQAW3MqgipHF22mCMppZn3WD2IoQDwG3W
pbnUErZOglQcd75P0wvgTUUsTBSirayoi4dRX6yvoY8F2Luao4dM5hBjv7E196xioYsM7eEOr2U8
4/rXzOO307G0SzPEIe1JD+0CzMKYKxo8KCElQZdrD1i94g2KGjNiam4lNqlKYebBKiOjZ8jsH/Dm
Lk3M0XU9lDOG9fI8QGVL4NpbnKiBBg1JR5zjzI92CnWXpG4cRxxNWA2yt937lP3amm4Pq4JWPub8
6i2NodAiQFZgz22ouC61L0kis3qmXr1EdFV2MyXvJ/mpgFepZNMDymh7mGhmiDcrkjLFnmdrrkbm
yThKaiv6nH4bABlNC4H6zrfGZyZCwTXx9P/yiopZBjkDYUr4bb9HRqDCgv3lkepF47uMCsbZQCGD
ZF05DWWyQk9iJ8cCY1R8FbSo3tyFhmd0aF15stl5pW0HwfNlj/E4jj9zDB29M11cx0XaTMjdU0i8
7G1kJokMnjEqq78yH4GLGI4ddAebefw1jCTCJVLFpBt4GXHY8YYsthHpUbsMLqJE3lwwLgLgF7JC
TlKozBC5CIR5mSbmqLvYDwA+P/gDIKFoJn7aCxqh6E3yLkViqoSN3fRIMkv9g+R1tpMzMRrmwJbe
/mx61v265iQXFejYxpbDsd5RYQG6WTATVugGXEwWxMfYCHZrb+6c5gc6Gk0xcwCjbhwUBr239II1
Wo3cb9UknIhWXsVcqzjJxiCqyAksuypSa0ILy2uHUUL6UL5yfbk3/h4Pi58nFnYsGeCAyKcMFytB
QWpE2SoVej57NqaVFRk4KU1XL/WU1MhDnIAB09n6/DhOvckPSKzmlZTyKyVLbzSabpzrjqUh6NOB
L246z/xrFMj7ai2HYepUYVHgKCcNLcH2N9mGvZwXOUk30gxDSumxLUQY+e8K3AIiuvrV9I5NckNH
Mx3Zn2uDYwVbpzprPS2+AH+xku4w54CtWFEg9GjpQIBDc5facoeT+JR8I2rOR3DCGr/wSGfVrLm8
XpcF5CiTBbdl9lnZ4AMfZjzOHTUGUVia/PcFpJH6AtlCvAWXYaG1pkDHFuwV5Q4iP5eCtc2ZGQo2
Qa6e6svnGLMWpOakccIb7LK9anuukDQVp6yGAkUVfCWLOUmfDZspltGiqMk766+X1rR8VC2I0x3n
Zu70uxFprx+3OtmuxHnfkgZOmctgk8FToxg20R3rsRSnN0S8dbRUXSKGm/g5PCOsVDatW0SAUriv
4wzIK++KIEA5QZLHcMHRQmUsE6wwYj2COB0dh5cVx3JGfj4fPPrqYlJ9xGXFjLk0sHQt8FyUFRHN
YTM8jarSeSyVSXJLNtTaQ15csBHoYUkIWzprUVFIS+9wL0EAONSgq4fgmjxm5Gf6PAiNcxlNx5qX
wt8AS0/RBiFu2CUf4C4bF3OJpH/qt9L4W9lMh/bBzMssIv+Lftsz4F7SUA8VyU8ECzbHwis8CO9B
XdJlwC1AQ35qi1irGHbR5opM6Zz1yturJXpb+pV8dePE+fSorsdmu1d/HSib/0sxUQ+m78Yi/1MY
7wEC+/h6/MQHkyWqag5mfXgMEwkqYsGfeBC8IhnEIKCq8vJ1h0Yy1ITHnNOr3lXI0wSZgYQhA1/9
/sCkSVPFgb/NBmFAmJOziEX8eZQOzcm6T7Lw0WyJZ2PoLB0kHvH859zqr1sQZ+5QSyKmL3cnNJuf
CrXKtsBj0+KUf8KgRqjU3rIywzuA5c9LlpE3LFEg/5jcXlKEw/3gKXaXnosDMfi9Z/pkV8E3AyVC
wfegylgibF85L5LiIODJI0xAbUrfq3fYSZVj82VH2dqlzO2uCZPHamO1ow9GSX33WfUCihFI/FEl
RqWDwqLXaeBOyh3cyDsDZ1as6D6nZ4+k+OxP/eKVxzDHJ+ecCHtfhSgLOCVX+//gJze5EPcbqQAh
T15ln2v+7U09Jy6jPYnLvpSLb0QrPRh8Ro3S+zkfEHozKO8M1ooFhgUaM1VaNWTdhx0du7xIcL/4
TrqHytu23kATMCQoAWViahRAE5TnGtpXu7VhQ7rwtB75DneiDLl3bKszOVh/2HZFFxp/tYVu4VER
Pu26/e7juZK1t2vX+3ZXjK8f1x8sdk0RJ+vuGJChAc8WpFmkN1jBHTr8tdsaWJHBV/LNwZQoX2UT
rkGlCkh0HpIukRMXV3pT3294enY/4i79v5P6wWl+prQuQ8mV5UzqfUpjBXm34p5J2fPolK+0rN1I
xCpVFgvkVNmYrfxJ/GmZVlQulOfZxIsBn/RAcJyh89TKK93HfTUUWp2QoR58p7znOMpw9ipZx0jJ
esXJZnoJB1cMTzVArTYwUiLxSwD8vM8A9WvmyNf804VLZNi8ifgoXXiDs3vP6RK6P0J+1UPHVi+c
myR/9HZXeEOB1SE1vPR6pbsetNQh5tl1bZlBypGVLJFcNDPKFVYF6DTe5ZxjJbIviA/fcL92USrH
7oXemX4IqWmeyAv/t6Zq7Ht1wKB5wY1Bt4FCMSosZcuN7XEeocksVzDPkXiq3b7hsguZ1Npo7Bsv
1gr0cNvkPNtKSeIoOOArpmyjh+yRJWJEl0Ozd/OPFPC/9Hyef3Jt44MjAZaCraoEzgoLsXwhXm2g
7WFfvVj3Nin9o8uPY8fbVWW0CuIiW8IjUNPJ/Mww56EeF0lU2Po1EJnOyqqWUX5iSrDJ3DnZQxoM
G0cCUNQ7KmPyhV68j+mgg/YaNUGeoScEdMhUInNTKCFoCW0mUTvgLbqvaBeg3JoMX/eYi4kunZ52
7zf424lx2NpqisitQ83gIQPiwfMZ+4uxuSP8OOg1GJac5YWspS/GcgKvFHV4JfVVgGZXapxR39ES
N0Jb5bxaKkDpz6P+dffyrqbX410Dpny5+lPreEw0jcIT8FZ8YhnoGTvVD7Kq2ZUM5lQIBkyljzTG
K0z88PImsDrbJi1GIeyX/0bYJVPXTaspshNNEwbg9YNmRhdpKN1En0PDjQoPnD8TOKihqiN1O3dL
oqw2Qrej6a0f6qbPfLTUKvTDL9dcnGtje8SnvdA74Nf9JEQa+Jd/mAGCZPkHf4Ag+L2RLWEuKTwM
C7ZRQ4xRIkbxZI3MgTZYhXAVK1KqPsuZ6e1A7oPO4B2Q+E39xPs5U4ZcvhYIA7gHRjkZP3WA/HQ1
DNo0fQ8AiHG2X+11pj3LMxFs4ucKB477qI2LaOr581bJuDDwq3ZqrCln6J6RtF4J5thR6fT2NZL/
J9moYWI1vwcrKH1b5b5qNRME1HhDEdsPfYtkZhbIcDnTE89spFbgThzQwN/LoS0g415iaI1x2xmR
wpga1dKA7tHA6AEQcjw/KtiamFOZp8Hd8hPIWkLIX0TC6+lLeK4JfO/WfE71PSse7rA8G3tZ56Jf
01qCOcSO1CjBtZWB4yVO15LuwO9vZzTRSfZZW2CCQH/THoXkBdbj0+UBU0y9jrm4A6KXKmfwnj4i
ML6yzm4uWU7H1FeUWencPBHdmhr7ztbIBmlbagmMe+I7kigud29+6wmRUUEjYRGn8/7ODrjXmP3S
91ktskaKwXVQGkKuOXJ1R7kI+brL/GqTfVIrorW9NWc8ZI3VRpUTSvwArpKkXzwi4OkD0QDyLzBX
GBAM1DFnbJ5Lhok3y3T9XTkcifaJusn++Cwcsx+h+aVmcOvn5YqRTKnicUmZvCNBY9VMik4OVq58
pb3Vuc9fG+7a4hK06ES4L53Dg06lvdAOamMQIkV3DD4WBb5NjkrZsbLb18MPHJP5+jTFdiiOPxYw
a4+WPp3N4oRjUIGjRKhdufYy5J9iow0v0BTmYE7vFNFJAgP//BnVkXaZzeh1U2tt38jQ41PQiTH/
uS/2IXzHATtUGKeQ7GGjWI5r2+o+6hXSngRvm/JCNdMHyrEDJSgjo0NA1oaGV9uSEvN/Q3+mkIT9
9LlMPOIZsO6IA6emfzp8Uoxp4ulI52zjTMR5c89Knz8+WSHhnedyX3n3skR7rdKmqfuiJUedrzVO
yfFUJCN/jnAskMjt3xCVvw8xq6iqtCFmPl3gRbGT3qXlNXRGXt8NrDlBeBTs1JCUzqDjgrJUOc69
Pehg7cLmJpyyXhi0NFeZG+QZj/BKeiU6M8YgbZAVWgAGmRxkLayFweyt7wjoGEINQBek2JH8HIyE
cS1jY9htSbZtRRhrZo11C9kd8HFPFtmsdOlruF4QQPtWFRkgpqCT/0jh8z3aKt33RFfNq+2VUb4a
UfwhbpsEtxuHqdiyor4m9r/QyzuffWPfxptwLtK9yXOD/PA8NYMpN034N9k20JqxNm/q2J2WEYXL
FS60HUfUQW3h97gIos2BVNJdYZc5Ckcnt3K2uta4ADK6QeOzyYW3Rskc57bl3mZCXjGaWZTlRMuF
6ZJROnBLReQuqxQGIw6+GuRHogd+T8MemBEdcl/JOnH2JiOxVCdkOa6Kf7o8kfk2hFB3k3SAIRSr
nJ+3OTAI88VTa6O65wQP7qMLocXwTjsyqYNVIXoKt02xWLOVxyT2X7O1JNW3LbSawohW8UrI4pE+
dOaYjjZLXDqBze2QcN8reJczxjFuqEmkz7mNBXjpUhDlPN1a2v7/Hp3J5q/ngzh9HZo64l8+U2Yg
ql98O9gRq4NAI40poS9nBWiIA+1dqRe4q8Tw8AoePwodEJuUlk/cliZ+Kt1P1gXHmNr3KnIW7AMX
p1cFy/yd2jQCervmJ4twp4WBqlLKWni/rgkKxKnkNNDNrks5j+fcJWYoItLIabXQxTz4kxy/1KNu
fql2oeRn2xEE3iZBX8QBSkyDQbnyI4vZu6W5p+p6XOZgnOY+Wii3AA1zE3Bg+53zQe51c8aG7Lu6
A2aiV/yIPj0cEFyH+LP6zMHbjp2JgG+JkNMEeIui51J1ICFH8GAJgvIECxEVRWHDFt+i+C/WXkZU
C2Ohrcl++MyEzMLBkN9QLP/FAzSelZbs4mGaPKTDfqxNuO7jqZwWd382dNglTY9cG20vjwE7sKNv
k6pTuscwe23TJdAC/FLNC4uHkl+j7qWVNBrvegOh75/+uIYNW5HFmtJHe5/phLi/kapOlqySig7K
gz5TJ9Oj368MA5Tgi9ntaq0drdX64ckX9LCr1cOgMbVX13VqTWetUgdGJq+75RnOTuRu+a1OPUF9
H8y5wryu0frIFrWt7udeMa1dQE4G1664Nkqi8BiKgBxwgV/SS8RDifVr/E2y3CUWOuZXoHbgnVED
8TWM91/KTF227RerTSnjhwxwr4+Y8opWeh/NUCMubyal4XcSh8xglvyk70tPRXcQgRsuyhSfvEyi
QpSr5w35ZtvmSF6XTg6hjQRkhy8vWQmurGtB85Hqpw0jhPQLhAXbaWL8bCoXPiaSYjSgAF/MtP5h
9fcbTE7iziHU8jA4dRkFAQb1Tt/3CmYVWXuT6rgCfVEFIkTiC0gveRedAwHL4Z8liRo7N8vh0EUB
YytImVobIAqxsnfkJassUAXInqmRtOGxZbO2WBSUcHp7TDuSX7OxfAAltQ1hZziTVeTj3vMaK2eN
WK9OXze0gyjouyMCYnFH9i8PrQ01Pft49f8kUHx6SpNoqoddDkNVqHxsYdZ/r8gYA0xcsIxKSARc
JbHlBEKd/zG/8Fsp8OhTocm41I7Wr2eBpH23ct86SlLNxP1SACRLrj5R3F1NBH6ccc9hGAkfAyAm
r3Eal+/dKxbkVfgVKrnXOBdjEbKtsiktat8tNh89YAAUpySX9ytGxVeSL7toAC8NwFkUTaUfTa+4
yqJVEOfXrU0kE0MbQTQDInr9dUZ5S1hSh54SVHuz7lsmvscIZKh8bxESnvopX+biNB6C5m8LuFqn
TR0f/viAYTdEYfUsEuuDakMQWm03qHzDZ9CPEQNx43Y4qUNN8nuW+0fzdKxv4MgMSrZL9sWNKaS5
6THiFYgBZvaoYCBLiy15K8v74SPONrromX+jNNF22yF6MGj6oLQJftOMOOb7od7AqTVEXSH2C8f0
lM33YECRYjzT+jyQIES2F1+KmYSCsPUAYYEASBCIaLvM2CGe6rTYaivkRG+VGg5PUEC52G+4E8Vt
DoXp65d2N4+EhryZc82+cgE539A0vy/Ru5zynbeDGs/d0zgDEwAthffPr7smdx/To3wpUw/J6Vhd
SwcJhG0+N+6YwJEMBsc0/irWQqsNhHmqQJzLGoXtgH0iavcN+aywc0wNCs59GCNEv/aDycOCL45B
TqMrVMsMveonXDbbOshZwVLfnVz/vuzbRlozijph7z2KuaRw/t+gZiMrX+A5Y3horNUwoexV/BQ5
j6ZaRBpB8CGjw2esiAWRZc1hcVO47Jl9QP1MfHozAA7r2FhRFTV4nFR4EjCTqf7L84QjSW5+/8kE
7DmZkA8RCDVp+isFRMvev4PWjT6gfcy50i1uAnm7ErpqMpsdnaS83depqQ+ywJFAHYVwiFhmnhLh
oK3nZRUT5l2gYg0rVHlCnbyNejK+KpNubJBkd96ljZA3PvjU1II3Picdtg6KHN61i7mxO7yIZIQe
U6v8X+QeopVAXjyrn0g7iBrTgKS43ooqFknf3KmM66hbCD+2vi/1JZh6mcPaPrXiTcAgqF50U108
qQW+FJTFI3EVOH8p1eI/XaWXhKwaPBfDdWCzBvbtunVm1n8RPULuUUuYA35AsO7tlrgEu25Pgc6f
6VVvMKu3V3APRK1lMJybCZBD0EznxQ4Cxf147PHGIOvNFLWM3bxebRQMfOETI5+FNl/mYNonXeCU
overECqXLKhXbzWYHeonXczigLIkyVIzrtEf6pWPSx6FH9QNKnU0gSDYBTkYJ0hIHQ3dan00nsxo
pj4WFESYAUtJ2J1w5k3RqO804vCT9+vYfuwZlujYu5kiAr10iZsO3yKDSGzgK2cghZ3sf6SZZl0f
zuf4UxBCKv8MkwAYHjKNnlCB169hzvjgJqgqCEs6g6bviFJ5w+N/d6mYGA6FxQHb5wLbHVtY1ZJT
eX7jRmpcauQs9ej2ZmBM8c8JHCO2gvEXjJ6+5pKQQFBa2oUSkK/vrlc0LrpsoP02Lt1XHsfNN+/K
r0tP2mIs18PV9LbjxypNiVvpbE+xWK6wig4HsHo9dJRDDVmn8pXx+Y8luHzIKKVzG34/UPISwXKb
txwHhv0IaAhEy01UcfzT8hPrwdCVjtZoLnPm5Fb0sjVZcEU7/rxtESnApiqNUZI4WnlNefubvnxY
KwYJT4Js1tsETYRqAQDGvUeFMwoONy5jTsncbL6QjVf1I/x4vfF04QBZMHTeyoTITFAAGi7mauxe
0X17KWpIwhyLK70jAjrO6TR/VVhDjTOYJYJ72hWEdTNGAS42/rEvRqjU4+1QaoDt7blf5yvqNpZd
AWBJbDdbHZfZMd6Ue8NLNvRjZ0SgfZtl0mXbOXpHe9hwctszsT8fqFNGVNGvDxm2rjGb8HPjE6Me
kAw1DRFFWa2U3IiGWV5TD5eQS3iBBrBZTlla2qtoNsFwffHo+U5u6zlZsodM2XvgugYAV9FdmOan
B9ukFvxPO9mNeMWCiAv+kEwuYVpUSScKUv9zo0RV2VLOsSu/N0E/GkD1JV0atVpVgfXkMDWa3C1u
WVGtuTQxCYqGuOJOx0Bg9CcUgWJ/sFGJhjjHfS3t+MSy2Gb5mrnu6mGtv+zyNTCUYAKJVTFe+l2i
7osxNxO7QZA+ILaFJmO6gKAb7BSqgutPb8S2mPkFwhj2otZmoBLm0HEmvmzGlNt0Oow4ES7O7JTK
C4ZFEtJD5dLkxyoxOuTF2GaVYAt0mK5kjDlCs1fzf5Y0AW9QAnXE/c93MDMCS7ypR9njqIVT/dAt
GqFvUrxQHJQBkliFaMDpfhQPPwiMNBFH3SZafgpiCotcLEM+kwBssRX2KFKTLVW+qlpLMN3ZzRdS
07txMK7Lt7JgaItr5dniL2zzo0z1RQT2yYwYAeeL634RY6gQ4Tyxqe42PVpLJtndZxE0YvxU4IS3
fWtgIfejKRotN7OEez7YWzOuibqaMLGdyVNyEnwz0GktKWyXgUKN+g/3DelvlZl7zjEq9W+P5TjJ
JHRmByEwTxmQ8l147vZLNEncSrWjoJrcCqIFgdn33ZjYm6+ZHhvOAZl4l+Qc417i40CjfT3lurgR
l42UW/mn0i3MDOqLx8D5LdDmWIO/pSzve9m8Pi7z7TtqEEnFWsFxWtbsEXqxJ1SapnmBpeA6qZyF
8ivjAB03s4VSimpjlVI/ifx4ZQqOZbqjXYkviIiSNGbkUhtIc2DJ/Yt77yQQSI7stQESIRIodNws
JlRYGuwOKxsCoCL2OUdtdqalEzuVV7QiSf5GfCbVXEghOTkvf78+yNzhcUHnq4DAnmTBs3kBDkop
2X8vKtaIyDyISYEwgIaV24YclWgP6/8JJFnNpRsw0RgSEIOkDu1I9eA/YctgeNyGyGcjmU/4grZj
qrCM6YAlx2zjEuGTqVyMhitQWJoEx28D6Q6YoAw/JNAHUd+4/3WX3obF6e4sm4ivv0EOf0NDBu3D
xWWpTUYVYRVfdZz/17crlWhvC1iS+xKWhH3lR+ty4W4y9QVeoCF34Wg8Sl27tKNgxOHlHan6KwDl
yCETkQPG7fkAXBlNXRM4LG6u+zXUKTuiqWlCvuNlTJFqEHRbdRKiLyAVuDIjJe8oRfkmExyzXO98
D2Z1MuZsEvyAN5hacDfl+m72key0SFUIajAwcwRVEVZDiQuJxCmGlD0Pk8JLgEuhu93IDVPjYO/B
jc2furMDTm3RU4CVkppQlnsJEWWpOvykjyANnWA/FfmQxPhJf2nKl+0chxVo5/VJWHBBgMzl3sCE
YYVzLjPRWZNZLdBjfuB9Jn9S7ogEdmwyOuHY4Jsz18zE1iaIIdtn3c5ST8ba2f9pdKWw6CYgI0z5
8fYBUnHQvEmB/DA1QjQyfXva/JMuSMucm4UqNheyR8AjcUNGfe8/2LkQk7UFXSJ2BD6q3PReBcQr
Qfa9v2oREjAyGCgO16VUka38HU0ApEBye1wmUXcHORliIrwrCSI9EIbha9d1FA5m9n7sTS4Xy6r7
GYknJljJgybqYitFaFNOZTfoOoSCzYo6U72fqYKAUwo8z5XOOoz2MgIVjI6SFbHryhGpPIQl/6I+
zm26Uj3bbjjCz0kEh+dX9pNMzsOAa5K+yHGUXeXNDXX00XNR1sKiJabyjuevrpBPn2s6VOTFhBhn
LQzwNHsVI4J766mMqxqGAzr9x3GnGmD4nsPPaxrchwj5V0jxK/XpTIOlt4ZqH8YTX2bedA2TFZkZ
8VnGizOKF9KFe4aVecTlVxvtQ1ZrcVwfvbAAxbYC9Idp90hGRNIdgNz5BKwsdB00d08SjdzTbG6i
mlPNVEyqtsgeBbGTAe6EUP7paIlPoicPeD7cM/WzRUe6TP2obXtw+GrqOFij6oenz6H/lbsmDeB+
Lj3FBmhJaAqIEORkH2oNw9QeXMpdS2NZ/IO+/ByxuhmT089QfhclZBnDG0XkPUAo3IVxndPiZSUc
oRFpf+00W1sqLndsI74fMVTdp7yjKzdWyCzJIkJTeqAgJP2Xy/ahO4D7T9uy56Q7BWU2NG9rGZaN
xZ1g4niyxbCdaHcG07AvyB/Z5tAo98rUi+7Peaoi5qpwHmlUUsBK2BAcm/JfbUP6WajwjN68Y2Dy
BaBcNh63LHhAgEa4oaJfoDDJUfJ9PJiXuRrid7tdpiOThdVG40UyS3yDw/8wRCS7Jh99QtI36NBN
4uOWHIa52dflBJqtPK1Rs5e+9L8avvKtbclFQm/lLzwOABagQZ0FlxYBj/mfulYLRUb5FGwXTe3M
vgm+mRiQSmUa6qq8Joz/E7Zt9rnRwgqbXvbq2hqWajDpiWY/MvwFdV9dPv5BtncvoLm/DnbKADk3
Y+S3tBJMdtrq9orcImyb1ToyVzAY7modqwq7AM+n46jWinYZdLM7AMNEeAm2C9ml0UlCsPNXShgH
7tDImCE00lUkBTCtsNaCs8o7TvKGMTFGDw9SSFcaNxCFWuTj9rksgJGiyMv71aiy4tUd4BihGb4Z
/vpRdRlbvzI6C+45zTP1ZjlBn137Rzx20wYmJaxaAHA09JdN3ypEvISIEJc1rPJDc7cVZvCfRTzZ
190bbaq2BKCbcf31qrR8PCVdiqv0N0qHsa7D7LWfgUtg4WRwhQWOtljdfcXlforKkq7G/SjL1+s3
+A1m+lqvN7Xw33CMbHVCyn503Tr8fMS+Nz+bAjT7l43uzASZaI0lSgPqe6j4dTmMh2SqI5LqLZHh
hz7rUWugiZZFqHBM062PKdVVsu8nKKhbw60BX3k+wxqICnqSGkMBlZCGmNyH6oScx9HjDR+JFQRA
nt5T1Evfgvo8/7t+WD3XuvCrhjgMLS5RYRFdtz2FvHolY/xtVmDz5s3xStOyBrYn/sYTv1sKnuRm
hLw2FdHLLtAamFwpHoA6eSM4xi8CGfnqBHuj3ntiw8mYDevyV0Hefhlqw2k5Y2tDr9DEV2rrYvfU
u78l+oTsliICqgXeUBi9FgVE4hoLkQGVuyIxl34T1hhzyf3gAs0pDcxUN1zVeizIGDiDCtWBjNg1
ZBd5v1JjI2b9BkaQ0UoIwTaI51QPT7xJSr9j35Un+f3oHvDERJ2oo/BbFlwX8SQhOnYS8l2i8zp+
ma3vDWDkP9aTdQ8qzQvc6cZuTGeJT3TjckeOqD8gZxKyIfD4YCdpmZS+fFjIUkJdFKGE5x1h1H1y
Sc3aLNqCPQrFfI7aqMqmmjKpRQ+ON8xYvI6Sv3Wkc7SrzLhKkBUEKojM7TSQXgQLq6VVoPZAN8i0
EYneTPYcg2KqWLKVpAxD5iNg8CYB+KaeJJ40Ljos7v4n8kVRPVrUEz5H8ZI/w6TjnonM8YePXS4Y
7CL3jK5TV5nHqZoEt4hQUtmBu41AKGcJFEWJ1La/mLd4bR3FaRlaRzrkQn3ozEWFrIQjAC32YPbY
qoNCeLQyeXGyRehFY2U31wweu84NbB6eJZELxqt884Il/F7GPdnZNWcRk3UH/mwRuK4ouV/zTXVd
psKbgMRU8yCJYqG0j2OjluQrgFzlKDvZInn11xxEzEUAS0PdGUg2grTtFeiAUbqyt6GpSfjAfim/
72fa/JM7Y6g/P6SeGP+wJr/mHwa/yeTy9/ssJw9ezCT77PJCpE7dLvCuYIw0DZ+AuQf2BrHg13+8
aAwUd4sSPgAXUlPvDbylyX4kfPW3FlPKpJ5e8UkKGQxbGA4MwlnuLVnMDhpO8rCryUZ5Wp8J1DiI
cIKSOcD/lnKTYHzpiDoSoFdB5RxsTIto4jLBjMRN7+KvaaVDZmUBfZoTnJ22i0rXrQgEDLCRSgWx
kBCKpO6pnvTTMFzszyZN9y0/7QehDv8yfS93+3/KLJMzlgph24tZWIeQ9BCzVhTUUsnguQh1ZKPV
MFr0kUF2yx7xkZV1by6R00bf1PsNRN7Yn7fCzBPStR9s3TsuvT2GKpD8Xjlv2tNARZkh0dFrMSzB
z7OT0bHIqsQ1sviEm8NGHaFByogMJk46knzmMTIAmZc+Z086XktXx4eLM28bN1J1ybUyiviIlslF
Y6IVp6Yu22DoxugQzU4zx6zWaew/Ykb2tEkJ/ZZYtu6OgEEtuLP4/BFm22bXQQ0fHcKcWdrUGOsM
mCoDf311EHBQIxQ/Uw2+Twg11FkIcQaZNvuOziE3dpdqZVZKFDnuz+9OMgIomZgUGfmNHy0wOT4A
FFqMYN2TIV+SAzjuGamzNCOwXqNkWsK5+nS96OP0QWRs2QMHhJipB8zCdACJNLlQRfERygkyiKyX
RY5dfkpM6K08m3tlxEbnj3MvTrqX9OOCbuyHnJWpY536qiHOYl3Urw9sQGWPOPVoHztZT/w8D7C2
2/f84PiicP8kIeq7rOWex+8Ei5PxOgsOoMcejqWpR8suSWqwupOO04Kq9xTsooBKdhBkUaocYZzM
JUjl9jauf/aiyk6GqPBbJwYVQh0kP9mVR9le93N3EYEDccOT2UCUeDRAf4tQJQ4XpRVh74ThFEQa
lmXyg+kSxtsfWLufg9cjv8I7Nm1YYVP0C2wFPQBm3srns6zrzpP4nj7DvjYhYHDHAnbHtwXx8KyG
TcoNmoFORYEPOB7taE9Hffymx1zVtmdH45iTDsqdZIsK63McEMaGN4M+B3YnrggsOBY61x1q4I2g
tGB76aCdoqXyhq9lSfrFqCPlDmfHgg8vp70S0avnJFgZ5JIj6zgO51pARSM0TiXUWiR3bPDTJEPt
XpkPaOw5n+NBEydHu80rKZu3+uoK8Q/puFRZTsozr6i1gt1Xp92rbGOsEnFsnpK6XEQRB+A6Tcv3
3VLrWdThSlkZvo7L8bJ3qlrGP5o3ulVk61iUrCAkJYT2dBt0ZXzsfRKOkNM+PWPhMIW/pe1H1p3E
10OoHUGtzC0ptTyu9rXP4yBGYPtHWcgb7SmqxF9oax8ftY/55Gyuh4Wn+82DBbLxeHGyuGYYUR0U
LA0kFDGF5ULD1xNjuul4vVYF9XRTPoirq4c0NHz7BKnZZkkjulPzMAMMG1Klbg+NhZ1jPJPu2ib6
sociR2Swal2l1U0ZIR3rmfcqlCS4EMi5dLAFS9uc3UzYXZZv+a44gTuUZEK6goVzwH7vbtMg3nx6
Tn3p4u5FCNLTuVLWGbfpRI0uE2D9EYPwxzC8nUEZSWf+tBtEokZ8DRMJnu4/ggy8f+VJ6y0Jxi6j
H7to05ENvZtmsb5yoWynNR1CIXy/bKHdFTT97Tk66mpzf5sOIiRiac7ND4rxVTQ6kl6LxQ1+qpLw
nZDNyogT7qvmBhnlS4d8c+B9zEIvHe1KjtUhAAShybhK/zSxV+HMlL5OGwjKI1m2rNZUqT9yYFPX
4bZux3Ss+HgqSssWeXxme7cZmi7osW2eh015Wr9cyzz4kdUOkBhZu6olpTYEZQXVLra3RUJTOJkQ
P/uzCQ+J+0jcpJi3H0K7kldfjSqe9jmw1SlAo84nBo0azrZucsr9crfjrliCbvfnVnLNhYH/9S+a
BkKnrk1uDaAOJS3w2ggDaOpmB5YAnm29co0z2e60KpnfvTI9VFsczH6O2sLkS/QrVm2Vu2pCRt5R
EyMIqac9YV+NaH5lJivUeOITWQO8ZEWuwnF8gKR5vlE7IJ/y59AAAdkkQKVzUBWDE5GERAvhSmtD
zk+KDLY7a0Xv1BwJVkpqwb0hEVgr26qFfM1Wtpv0/DqH3HtpPwGo1NUVQXii1j9QlXYfrT2fl6mH
DLuDnazj3ob6FkDMFUuvLkH6MFp752aLrekw8niYl0Nm41CLBvrseVmnr6k9C43FPHr/He9P5ooy
0qrE0R+53MwflegTEpHsmwd6RhneoEMGC0A5l3LUpVgQuMzQdzO28BrEtyv9KgZD4YuB1HZaQybC
UFM+2RvY2Kpo3KH0UOLsEAMMsdsicZ8Rf50oYIhF4run08pHdARp0zF46N0nLqIK+MPY3EUu8n1H
0FZNPSN9J7CbW4/9SnsTWRFUQN92ismQT67wA9Tco40AdFkEo0GRcSoItwJp3dohebMA6jyl1yFG
7vjqsUokTfjMYTkYJOvlEPhg3fK5TyjCJH4vXEYHeTrEh0KBDacl6EAP86Xz4k4kAJpV90ThczjG
ukHT6tzU5MvzG6CKnsJmsAk5fhEIy0s+77U/wsa521k3gfDnnA43REi6+84KT4XZaK0qUgjiJp1L
dGJRVlgh6NR/S2adakOyCwkEVe2Sb3nL+Jz2VwSZFQ1Vo6d5WbGkNfcBCYAwKJCmM/hJgUgobEN1
/2oG6xGawND19IakdyKz1pcz7pwuSIeXGYgHr0BbPO2mi35mEqTETTPXfPpYifEEfBBJIXc1ZcfO
xqFjKSYZWAa2QHPRRgWAOCtNW0s1fRCHHfNS3UhGQAL2NbnkmCqLdbaUAAMAj2JPiUI7efaUXm3U
SI/wyHR5QGJ4Z1vTWieDS4nI6szfb1hricEm24/CzS0N3SpMlrGb0l2JX/qEHFcLS/1gkQID1fgw
LcLz17srf0XImclbDfSJyMNc1PArakkdvmwvYchHyCvPc/QeG6c9FGSB3e9iTwad9C807sHwuvXT
LcT6NjDwvxoG5F6NuYSQNXbSBWF4Ni8hCiXFmdpDcQ2Sq9jYK/aTEksTxOlRx4IhDPNhUZb7Ouqg
n8evs14HsJ8kLQ4B032lQnc0f7vWwXj+Ofyq437p+7GS4tQzMkf9zDSU7HnNccyQX3WTdFc18U0M
Tj7h8IrDWVBC5M7woHOg5QYVhyeCYQNwdzj5ApB1zmmxl52kzM1EZmp9MuUlRojP4uxk0WcSqQzL
es7mQo2gTEJAEg4vc1UaODvaRWfhuKomXqkLI+7tLQLEvrv+/4G8pP4jBNv5Fb9nwnqOFC9pb1e3
TpipzfSVWs6+sL5j7hhhQuwVoZycJYgdzzqW0uiaF72kVIDm2GFOnuNEw/yOOkILBM65wlBBSS+f
Kq0eLSm7mHj5LptWZdi9cXuBbkgGK7rMj40V7OHRqpgcOwV07RE1Dg9ccM7pEXkmEvq/ovvRdmNh
s9eCfQgRX21IiTR6M9cVMarZ7NkN0RxGsKwmQMX1qscP9GV/K7WL14xVT5BW2JTdA2KY/32VhMQe
QBCFs/skjpNzp4o19wUN2QOUwr+rVFCPsFS2FVEb8YXZotipt4yvP3Mnc9jmfJ+yKgmRZv6PHzAB
vBlF6GWt4Hm+wubFYTwthM7GiLMjuSLVt4i83XektrY4FoB8Xxb4xm4YMk0mXO7oowqVkdaW5W9s
JZ20PLVz8sC3fgscao8VhHSosq4xP0A3P9ZvJvtT/JT/BQc9ujjRe7vym03hsJvUH2hU7qQrQYlC
JfBqcWTFXsNR0ntXP7ldWNV4N/FxU9E2hgPL28GBvgzClXYPgAdk7+dVRvsl60JQAilZR55f0ggH
rXCmKBv/Ze6CNEgz15y/OuAwBn5RcYLQt/Z/6VOO40Vn+RwsQImcXqMO/6GKH3NzIQTEx1IKz+p5
NWh4QqWy7yD/gnWDJ4jvCY+kvxqWn+UWozoBbYtgBd1UFoPBRFcdZHtU2PzEn8rymaxReXR3g5V0
ji4qrYbX/z7QdzjOs32+0EWBCKSqc0+H+wUQ4Q1s4uZeg2/SRINVL8QoGIp6cU8v7/XBdZUaqqF+
mRRbtj4XUCfg9QYqgj12s0LILh35tuj6ZG914/DWS2XveOHwB9sUL7W1V13b6e4ccr5Cp3ucjVGd
XFFF21TtZKl1c7LzxBZ9IyyLQKHoLqNy77aUIUZlU2rkTrXlMLzlSK8jRp2lPhtKjVlIJRYMHvux
S+SaTjsdKpfSZH19ajWmX8S1nyCqsbx2fiPmWPXzIAszf4tCv3cxTQwdWVQpm+tdUAijHJc6aINl
p2VLIaXjoCk9s3UtavMtzNQjHrhqapci7CN+cKyOCongtqO5msWVgJlTJT78CDkgpsCpG33cQqag
VxtTC8hVf+EOAuDiDf9sSi1bDDtJwfPuAS6N7CsfCvnYdnaj8L4jEUqrJRFV56p5e8L1K4seXMMV
SG3kOxcYDzhLirHvgzYDy1X0sdTYCkyKxcpT5a9SWxH1OD5om++8xZaJv/X2kP4i0A9aK7iu8lzA
JD/2Mwuhyh7m/5BRvjm3RJzWEimVoTJ1RJtVOd/obNCdenezmBgWXIcfeXsYhgHMXFqmsiQZWqbe
6+dcrqrVn9sDZssE1fegRdIimbAtc5cd93D0lowaQJ8Edxq05BUBNzc17caRDIZgA18iIvUoO0xP
qptPJrnnE6FqT9HUEUQmoq2/xG+tXWNw1T1eVaaGLnZ99IzB3CJw84QtYp4Kho3X9lQxFwwWiA8H
9rHmQRB+McCcC58HVoZl6oxVhtjzWYiw+BlRC+/xzW73q1bMNyrAuutQ64SnHNTFMsrpFWRI6Cd4
AHyCm75vPedGHtZoaJcucULqZiMwAJmYBoKyxL2dNCjfdIFQf5xshhzOiMyWhOZFPeAH7WGZGnyS
uF6VWDijRGmdSt6oCF0uMPWbIKcjp+5jVgV387cpmotZ8RE5i4thqlty2ULx3utyWFYRpGZmwMgl
h4oY08LINCCE4grI/I+s7Pn3KVBwASMsJfyo3FvfJUg+r33Z1MPWiQ5JXSw/NJBTijxMT6ouuqLl
7V9fi5hcwa96FahqZqbRUeRCUd4SiKhtOm3FdGdHmQcbtKjJTNvp507C1D7QYQekBsM+hNIgSa9n
VYbJR5sh5PrFLx8reD3QnebUr/+psBDumqW4eC8qI58lmL9+S53Oub6+Fh0+wB0/TTAwsZ82YObE
Jb9Rfnr02aZD1Y9MAoWDeSB1RWmBN1aFbravHdiZD0sGUzngKGljYQfOwuklTvhxQ4VEndZNDgOz
2BaNbj6UFnciQW45iFUTJg8VgmfyLqAYkdasikYimrMxsH3zys41CSg8UADLDfCgVytpxwOh4rpZ
77/PL2ptXGVvYCI+1WhTgo1ijWkXx/CtScf8D6wKr27KbkQA8unW53LVxoFy9YezK8yQs/9McLv8
uMPqoWldFUhURZJ/nxGoPcYDyPji0oe1Ae42MyyqTCj6P2C/nOBad9+1AyO8KkZDjlfC90FBhygC
Oja3VOZSR9fjig60kDEc2PDXLSLjSOsrmELYBHEkKgAixsqZAR8w9ENB2bIpM3tFLs6CHOIY0QDQ
znRZuUNyUuBRq88A67pldtJN5yMGUhiAg92GUs90ti0K6ru4O0c766xU11/kglNqBn+LPXsk6gpJ
J6G+R60NaG2EQMpHQXpc/NgcInsrLX0GaZWvNUV0wlti/5n+P8v746OXPo6k5JIedC3+avmHkr6x
ekLlV6E6SziDSfiMRh0c4Jc/+tmYgHnHVMAyHWgsmJBAuyxDrEaxvuZ9B6FtoTkN4UnPFye9xTlr
6UtmBWfYjWr5PjGVjgEocx2HaOzB91i+PPiGEYxl6PVqFastwou3ygg4d062xRNWZGlVdOu/M8sa
+hKFNKoZZ5DS8Pd/Ims7SxNrzvZHRmGbdzrgbeODaGhPKMmXq4iIWlMEa1L6XQlMioFZ9JeHkfva
76EQflbEXkeMaWtc9/8jTifPJgh9Ao377b5VARxn5fw6uG6c1OYqQUsKDT6/vyKEZ7aVfOURi1Ra
wQUqL5lFD7RsY+r37OuPlfNg/bd+hsumW045U0d/PDxyIug4fcWpr/jd6w4et0XMEXnN3Ty0XC7D
G3QQU6PZkmduJeubgP8yoqToqlLwZXWy08WbDwFkIwNwl16qyz0Bsq2gpXhWLrjTRRZbmVFVaAxH
btjhwaE2ZlgJRRhHp1F2SmA/jKcE2sxWrMZTkQ29hT3M+bvs7i0Gt1Dm1UkrRGNLhLR7M8/KMl45
e0t98RvYbnCq3/kh/ZFFEp7CLl7yS/iU401mT7VLK+m20t6u9URbaGzq+t6k9Zlkb6aw1ZUTAsi5
mgwU5J7gmFmO4vlat+WRBduP4xZFcWycdXRvDLDGlNWZ6KAoKNt/K9QB1/tTOlG0yPzqJq0vjYSc
Du/k/bSi5smYbOq1hRt36KxpaRKFv6sdvcciV4K+qj+d9DOtAG+IgoVKvgRSlssKuuCSQvaFcbyC
Ork/zAzDFxSv6A3RvjIUZOxwniF1QmAu5Dy5jjhKKYugM2rIQ+RJQGIqRc8XpiqTrRqKmvborrl1
iRE990VBwhWCFBhqzf5MwNCpHcQ/I0TuxBepos8+ARVKfR33lXBW8QABRbnz2kWeDU/L9yZnzVAR
fTqEFp3PJlkLjX7pIr3JrhM5+RZpfVUcXSDA1DsRtJ4Bb62F+Crr9pml0Zw3U3j6xT5QOIW7sPYi
z0hSm9QjeTv570s6gRSjKevQov9L1NFRzhPoyNNDygKLhwGRtDTmK6kRYNT668AR4BxYNIc2dr0W
tHKeTraXSgNI0hLQyTwrEwGk8JPtYfBl2xdZIT+1mjNLagA+n13s5x7dun+Rl+1LOmdR12aE5D3e
T/g2Bum0QFEVbcfJVcwjaBD1LGsfXy1ukzuxzbGuq2bQN9jy3LVo//VK3lDYpZjHYdTy53Jbv5xM
KbgeBBFxH+sLvv+qczoLDwdR9LAu7mt20now1z0TSIYPO63xRFmnQ1oLxp3+b7kzxTm+DCJJ2L/c
BAqFh+5uQCWfBD5E4hs0VrHDF4ylpRqnDZrXoTzsnIiRp8wEM5X7y7yY3AGTvo1dK6j1D97R9s0A
tcIeFYJQot12Bom4tC2iR1R2T2s/ZM2OZhB0vvzjljfv9Y3nUYK1NSrQGxrtriID4ExhXGaxSYBK
8p2UP8uZ+R4QPDtoUuavu+xqmb+RyWqq5TRfku2WuUPHlQAZEXKhkOjualCUKUb+0zhbRIEL28bI
hsQu0EQ+yE2UcmLjIKihrczoigkVKZq3i16fs78ZZ1q+QCvZLX31arnAdq1R3MsuKXs7monfZwaG
528Kb4Z4Vld8VgxIn758Dw7zO9k305YmStX0jNe3yYyBmiTZvZfvv0vS3jx2jiZx7DvSJhD/FTJk
x4121sn59gCWkjjxF0Nm8Gw/K4yWIO3j0GzQIunTQS4nHmcTpl5gpJ31cEqA1qwMPOJwnQV8RZ5P
r5OHOHCUrQb2sClcrt/0FckWPq0xUoSsDsd+ByEN0oZg/XJtLH7xDs8DtYJLMsrPpUDSdTIkLZOL
cUzl6rwIMI8dXguPqTWI8I7g1AwMQ4NYcCqSf4NjS8WLH0b9LXaQmTH/20GtccuQhBRBiSNyP/MR
vWOLQ6MT6ySFAnQuU9HvdCpq9ENP5QZ7GLUwsOfWGtxdA2nmlbLE4Vj7A82Lg8i2vi7E2DhW9HV7
L16Q9TZBd5jasDuAlni8nCvlAoXAoAtdZbQsb4tTgcQ+sgEhGvpKqAny3pUGOvvCRJMqHZiWI5K6
nGos2xR8Kuym0XylyJdDrsDHinVuhpJnQ63RAYXfatg6OdUPwSMgurE4iIZXyAQ5Ye0kaXOlvB15
8j69aUJbXuSindCGIfq7SPX6fky8QOe34IiTsMg8eo+MWMkIWZKPxMebTdwO3DVqTxEotBxn7PMK
9F43bA7Flgho4wOgocT7/iO6/cgOHXhzKVCkIRhg7c1TQCqKoVwOQdMx/eBPvZkkKB/MI1eC1FNC
0Cn7Tppvas+vaHW92sywlA2RtRppjPjnb/K92f43DvujeDLSVP+Hx2RqKdEm+/teCFFyUpwa2FAW
n5wVFacLoJXyiabT1BCl6n/sUaKVxM4oZb//o58ymxkJpHAJb6ld6LCBWb8gbCYp82WoSt8bmC1d
Rhd/PyStJFR1Ctt4F3+UtVOXDnYkBxGko/73xT0E5abACYtSuBkU4sBx08zjWW/SX6uwLlhBiu6a
1qVXpuao5fGdD2pg7OBhgLOeu6eR4BGjVlxt/MRGtXuy6UN30wezNfh1tyMEjrH7ED/sSNuNPz7t
nHOxLfimPhTKjSqIVV7sj9uHjpzjRjs2RU34J3uxIJJ8aafNRKI2TyTZRU3McfVu+p0vrqTkrqMd
VdAtvq0DiKBMTTkAcqDXuS4z8NdtfaXPhJjZz25YAmrjXh4U8gh9PG94YjiRXfZW04YioYyaFRUV
bGuJhbU6+Blnh+0I4RpfJZuXMC3XkefidAVeC/K3sGOkJyPnJi3qh4FG4vdxtqFhvm6MXNDuCY3b
1S5DAPloXJnTB0HPOy4fkDOOS30sGnpQwc0Fd88UlajiwncZ/Dv4F7s62BvqXziXE0s89b/pHmg1
XDQcEqIU0Y6NFaTlAD+ZNVGARiCVidMMbV4MPatTf+5WvlZ6Jcz12Xk1J6qr1lQ4q+StTjZxSr/V
EWgx67/dPVt12s1F1cIa6wjZgnf24pzK47XPcDoOEGlAMvHkCS0JfEjtF5BwqQP29nRYqjCMombe
CjubyuNJOT6NkYA636wyOwubLMAXlS5wbkeM+q558EISLk8ttNQ/N7U+617QGnLHJLsCnEcsr8Cv
k6zgfze7h2OeyR7uA866Ko5De2lq5PQmnoNAnvR7B6XgztP65W2cSJm3BBEXpi36wGejeFTO0qa8
rE9RIHFvLEKQiQy9uRds/xOKvle32eDm+2MuNhKNLoXHahUV+XXBzcEfvssC+YEmHRgFCCYAXXtu
CPI6WtOzRl5nbXSvdfjKPVCJStXs59OwMZbSYeW+V3rvCxiZRNfTogl0EXjq8ezHNpySOKRXUnwD
Ki7i9r98WiEBsJf+Iu9K1I/Vgb9MiLRMmaWAf+lYn6/m55TvkJW9ft+NgJO4fTQogeH3EwY+P+hu
0JvbR2fQKw0Q4QmngtHZkxwFTYQtDo6Zie4Jta7PP8NggY8lrdBBmrfgb308KHBHVTAp0i+IB+Fp
sA9mKuON29Ns14BSHQXpjCWCsEnl0KKaq6sQQ0jpLI9VC/vyNK5Cj7dwPnBBsv54DlIY8pcDCLvF
SQ/C5OMwxlwgcYYGLvAnLPIpeVuU6krw5KU81Fs5E862ay0dBvSd7PinwqniXiZV/A31hlAFikBU
EzxSUq4Uj5sbtdyzE/3qCWhgV5NXNdevbch/8SbHRjDw4MUWUmqLsxPZs48NrdqluuS9ziRZ4BCh
tdGuSaPvFOSiE6eFtAOwd5RYOG1n3GDgWnqf91wMCCEV0Htq6lnhaKkTt/yndkFuT7u9AqHdpN0i
YgbYvafawN38DDIl54WRd1V2mnLdnSTf2CvWUzzPGtuNeR428GP4DRHa3KqBBJ2pWwpXAu/6emsV
P+sA6cT3O1qPQAPeH+LhbN54K6Tgf/IJBGOHeJclZkG1MPfXQyVi2LfWOTQqx1pqWiev+4vvFIBg
JUSHf0QW35T0PT/XasgKLX8x17PptGADcfDZMpBo0X+1iZlRCrIMJZ6xkPyGqirnIrZKIwp8sH8t
Dg41Zht+V8zBNvCqvLD4W/k033xxGAwn2lHMCb4oyZbYhwkMVbrIS9m1pOKhCLEOKTGDbESX/4Ic
SdpRiCuXEIlgxoXRdJ2DsTjztEPh9LtOdykzMe7bQzQe+zYO71g+xx4GXsMEQB5pp69Xu2YVHgLP
7w0GKnojzTm8aVLkRfaVyDBtQef5teikT2luSWolrMnAziGqOufDDLh6co0e2FaxK9on1wEODxUa
+/c0CDJrtE5Em31C+TcsjYKPoaKNQp2D1BgnVzUm+/SeLXQi4bQeX+pPbOEPU/MErotwEhU87YT2
48dvXgrHT4hbNWst9Bc6Q/lb2zPtvI1iBPRWTwOutiLqzNS0rsZwk98wGb6FctoW5SFdgrhwygvk
RHt2L5wVIL0H9/7wqSs8s0AW026lLhqdZAC/m2cri+2BcsG/xY66RJ+RLKXMjf3nsQnLefVGXqV4
7M9WMuLOGA66m3xC8Qispmeb9HcOvetXHagYoh39AF+lQ0aaW/zf8dpdFH9tpgiKwGN3Xj7oVw+W
krgbpUFeJgAtgmrd35OSWwAgCkCm8oddpyy3svqm0vfPZPiC/mb+ESQ+JMCjnnZ94nEXXvuR3Dl/
8PnuvL07H40EDwLB7ly+ZsV1gJcK3Nyhtxy5l+/jq6W7eq3WWijxE3mbZIPjvZVRjcT8PECDV6wN
M38pDBZeDHOiFszlO1hvy/h/5uZrUKCLcINSEE30KmkMMBu+r9BzEwy9Qz/MkZW/aak733IIVhej
iVydJTfFGk/R6HBk26erBkfZLhQfaPQtDZtgEqrM1F7FQ9HBaJAoc7WP5ozUkGjZmr8hGC49tbwu
URRvJr2s1p1RnFn7D9w9cWVhIVrg92NDODHV1Pkmi1OgR03jPHWaQxUPEgKr0NPJfgzhcm0N3e+2
7LHd71GFw2uqcW16TLSZF3mOw6qx0H1mCYN3YnreCIDcE7ZnByLBDD/bWiUDYwcfylccc/z1YzFs
A08EsbzWxLnFQC/LpbK8eCnzi9oy8ns2wsfcfI2ekkIs7+44ZlAC/pV3CvqKkua+lsDPkQ4WSz9f
wOKQZyMamP6kVG12Tg+LSpg4ZT1n9ivkhsT81F3CevjMmAhD2dnE5YuyMCvu69Se8hWOt0f5ZpVf
BtD/+ity7uUh3FhaVM2ngqZpvGSqr6BZ/PHGpQ65tVZZ9RtKrCdY6fsqx5hP0Q66EgfIWCNi7Mor
FgVeBj5M6ayAcBdlYde1Ukvdm0vC6RvITuDOTVI7H/2Ng38REojHjcrp6lR9QfhF1/hYvpF7z68D
73u0j5dwhbs6ISMgOjBA1FTRVUJNJAHryGU9x6zJbs3683IYgklEQtpAScyXUor7LTpbtgTdS2zA
ZQVINu0/SvylFiUZK/TrS68DvSnOjYgpiSTl9Ck+IMXYiHiyuxdQfEN9gYBasalWPKhnH0Cxs6zr
2dmPejKNkwJZy6V80bq35nftaz4lbjgQsfNHdCJOeIyskq4oVvs5aoewAnb2gCVsgu+EDDUaT+Ok
479Rfk0q67DSrnv5xKeiOJfqxkla9BM+lScAHc8aUX4s26Q+XETZtu2IRSVcehhqz9H9PUvaCltm
7YqQHyDINyT0fakaaWLmEufR2jN8pPB4SFqAPzXwXMAvzrAkdpv+M5CrYic61wYWtyZrYUAxKVxz
fCzRrl7rGUuUKs9kwAL/PZvZBwgP6km3Um5NGtxRGE9XlQRbKAu4d/6cTD/GZQ4UhgR7KG28I7/u
e37maRRBWXbEhNSrcwJTHDCbh9XORU3+PzMEmLyWzOECmrgJxml94w4N27OO6dcOrph3uEIftqjZ
8FI9c1Wv7hpRgvdI2X4X3MbYGU3Z2QhW0cBIk8kVCZb+e45mhPWvryJ378zk4o+iYOtAkXPijzs1
oKvhWFN4TA2Pf2w6UMhE192ja2nYDhT48u4p8XdZ1rY9G4N7bVl7Hk9hYXPmiWqL1U3Kp+AKFlu/
upOe5jVgXk74K3WTP9SnYul0pDVF/NYpPMOfHkF8/hd2xhgRiXmSnuZo+7T147laX8Y7beUCCVIm
WNAqQS+R1V/R/AEBRfJ3y0lBYiaE/7md4WATR9iAq9X1UOZorS7ZL6DVLFAGkP7KXJ4Q21BlFqN/
2fGIL0Vt3EFQFrVLhN6McevsO+xnirIe8OoLzK8TSRbuFES4qRvlLGOVGXEbSZSobshJvbcBX6FE
KBcYjvUuXSFPldSyrso+yiGkb6h4nKHorRHPQvFODymC1n9BfnWya8LwXqxdOY8sGrBJZKJb/Oum
Gnrf6T8St3FqAYINNvTAxJEaj0Qw6KU3zWGFR3M1Biu3+1nbWzWtcJ8JJKKogePvd0aYTnGHQes4
wVd6aAgNDffFmtmlmLOEDUZGNGvRHC139Wvn3usIMVLSjZYFz2vh6zdGgF/RHz/TQjeR4YutxmIV
syUdoC2MXpkhiRW9QEe6pej1HVJISS37lbbbfY49zJBLnf0eo4blyXY5u6vqPkmzbPkJ6EVs6l/f
MXUJfVy8oqYTOywYItn3DM0xA3umnEm1zz0bFiCBDHbV2p89PuZEzqqFuWJtgdAMr9z/MS2wAeI4
iqjQnLm50JRrEazOCTT4wMrqyUldAyGmFdUiiAt1LZWABghqH7iGC6cdmzclDA7a1/LS5XeAvyFd
tLFAFKrJ9Ixw8RMtl6opd+/krdrYDGJlaeuebBa11iox9PFrncal6jqA6FMkXiHoznyhb5CcnqMW
Mn22bVKKPO8d6NyoOlGV93Rcw8z46pSdJk6Jgb/pmhlSekIV3bSOeZg5ysp4EEqMTjZNOo4q8VQV
bo4cTto1EKWv4u5fdr3cEy+LS1775RetMX1QeAw2BdFptpBhJk74YPmPxshX/IMTuBXdSXdH2dsz
57j1lkCtlbUSJKhxZhMGNkawKKuCFGRYgzD71V69upJivwEMq3MHCZk9X3Al+meLRlTPzODGOhp/
6Ol6m/3eVPq9o7dDUI9K3dKAN0Y58LrtMQG+8tzQfMDmDARyJKzhkSA2TjBq/4nY77Uv0Tggc8zl
I33IR2Ao4+dJrCe7DHwX+QoFcLAmYDnZwc+p/Bh0M4MBOjA4NtLmIroYH8ZNCwy5lf/7zdG4LyAG
AL+3u7N93S0PbnCD5U3Tcv0ZeOcy9cYxkyHhH2HHWXhsBUFpucJXLIfbq8AaeRcIvSHaxm7m0YpR
AQ5qNEmKRbIweaJ7mLYe7NKy6ClogDslKDoBVUMbwlg07iV3YaywUZfyj6oxoefFWI12TqkIGZMq
lKWX073kUfW8Qonsuw3oEOcOkts/Dpb8JMRnsm1ROMTI2JXw3TX0kWVjAjh3DYTMSWNEPim5SR+H
Icyw+gvaFPyw9ubaDOz+4pw8MWVTQuV1rEOrrdKZGkMptgVfOhNHBzEuY34Vqa1W1MYzsI4aIUWo
zf8CKB5O8VwC5khaS6Bk4e07suJZ3qcPOrGw7jMrEa1wI7psaagv41GPfYnLoW2fCmRzm67oQFb0
TrqujB46M6OsMiHpfpMUuafbcUdV0XPcwbmpgJL6KDVulqllRoxk3/ZfGpzWWn424nF3VVEaEKK9
C620WMX4JElm2rBQOTOAmT33X5gqk6vpysv1krHcCdkb4zONOtcTTKqprMNrKBl4gB07wocKzJAD
1cHWKCP++iC+vMA1DeveYpqrFmL56urzlQsNrXyjcpA0ShhpXXIpCFtSoi1YnYKWVdYQ9Oscj7aB
TgPyJWNCtOu5XLMkGY8c9jwTiNGjbPgFpqnPKAGRSlU5yUmj03IX3Mo87Yw2lSAeFYaCbs22g2ku
T9jJAY1WdZKx1FCD3mNOqnNm7YZG1APZ8rJaUsLUBw0LGxUQRZAxBinWShsb6qVMoLZyd6D8boSc
ReSzlG0PqeBonxD4XpBuPGIq64GfGP9lZ3RI+fzIYJLgpY25QrixFf+RD8rD3h93ocoEIiO0UqvE
pfU7LckhOv9sO/sVUL8Pql9DTaD9DF1aONitMQ5+j5Nih86FbK5V1JaRuHfaxvWiJLSyg6SXkSCR
9RM1qX3StHUE5C3jP+TQsNs0iY7rIJW9Tp2roJEM1CLDkBX+GhFnI0hTMtpyBsbfWP++h5kFKbcs
qSjLJBND5O2IUOBz3oOGt2s+4HrotljywaYiGT7RECxYR5LbdLS7ig42MnJYGN3xwCH+FQfNXF9O
5uYxwvhm7Vd8k9uTsqDcwCYMuty3wzw/senE5PWvNXjtd6lXusirCg8WiS/IMoLf3bFeKfYBm0eZ
UCuBCPZRsQrJhjx6QTFDNI0AhjNAon0ZIvG9LpLMom+YkeQwvtB1XY17JVI4IFW11HZtVwsNbnUF
EXK7jGHlq9LT641F8ktIjjR0iK33Dta1thcChbohLuU+FVoLdsvcXDJMPnEqRomMnpVUHDhmpV+Z
U+1fnfI0vvtOdWi2kXbmTWAVMJ+uidrEfdRdbQnW+/VRNZmR+uxPfiNjoyED241k+YhDp7unOypp
IW6SJ1YANX8ueTvIYwXingUEQQid+bwunJUFW92GN+HMfilsDCGkv8r03CHFt2fr17327YBbJaFP
P8njyboZI7lhZL2rrYDOgmmy1xOyOBNswXk5g4YPQmboJZMTkfOLZmeFOjoorRg9YTkdRHQ/J2f5
1B6PCrUaHXLKPsHu4v5qv8cvRaustA5Bi7hX70GyOdWbFs+a7fe6kIb1wvD6mVtkS6t+D0UA1/b3
FpMZDGARhjs9XTxk+lbBoPaonPxgblgihs8NDEYWT8bNlFNZYnU4UmWwdkILnSALVEuIG5L4BdDn
rvxob8yXawwRBuVZd59NkbsMNrIMtXgVwmi3yBUPl6hSevhb45KeZd0UrrZX6l87b9gmrscommsZ
3jlnMYZvM7SiBtJkLry6ELLUuOMNb2awQK1IHcLrmz6rnILqUeEsu7+FISChPZxMVr96OwE7dF0w
8BrCh7eOm+/kedyZlIxT/4ODe4PRcE4rhhG3HLyRipVD5s4PDRaodRwh1cMT7Ww/KDIZuGjBDe2P
lMueWnlh6tydvcunsdw6KEpXFR3YfaB+85e9v+k9HVI4Cw83pRwHtnGieia0uJ0d0zc4Sd3Hu8jl
Z1eRONIeeOFVsVPaUdv1JbvJCNkN59h9CR2pK/cIJJ3bmVutiZmQTrAqGmQFZeKjiubszPe7wwGA
H+y9bIHkwWGEKDquxRdpEWBvaPW7dDWGKjUgjjusHzi7yslOjxz18mgsEAl0/7GE/+7KICxNy7I/
WB1dLx9NV3PAFuusJc/fWxdtXcubgUrtgLu+lHifpEXq0rAHyFw1rAU8wbBxhMVhb8ypHa2WGVrQ
SBJQxEHSPZhANwL46JNlF+0PalytPEIiQqD9CJt24cf9jcGyFkQzyj/5iYE/mBkgJWb7uVPJBAOJ
LGRddY7P2DRe3Frx4xXwumGRXsRTHHlwpWlo+7ilt5ycWakOKOPzkLtK6EHOpzcCG1hpPoz/NrqQ
tuvXPlabqkftnVnjObXvn8o+r/nfOyQKwjhBl1bWzxXnwGRclp3U/mmBEEQUlF5TT5yMlWOkpOAi
iCzadGGRbx/dPAA+OgOmiwWHD8kHLKKSokuI105e3LJ22v1Kep7Jj40VIOGlSbfdm+Hel/0cA+99
ERxyiXfU9a7a8+fbzoJUQYBDsbml+SpwA4HY3gcmp7b/+b8p1T/A7N9Duuiz2JB4h5RoYRpJph4I
4g+4BlajcdQbAIVngqqBhxWr8mKve/ti7zBCoM5hSzhijKZ+uCqZeRM0YNhoY3unT7GXCK75W7xB
ruoNp6PtEQ7b3e7ILKnK1/PM3FWyGecbYVUpWOe+t5kD8X3oxvY0HIRz1gQabopJZuOQ3whgIjYE
HhUqLkAT30bkZHZAn68bRdR91ubZWtx86WDgNMysK44Sn3OiEr76JZiLzCpMODu3WwkFjwKil1mf
H1NoCEwD9alN6AKRUBu/V1rIT5/d2MvF724Q86PXUxXZmk6LniW+H21/Tz0lweoy0Z/3jJF0+/he
iiK80XlivbIsn496SlS1MtxULSbVhoYpV1LxZ5g6nrRnw0/eQ78gIVY8nWNKS0fuQtjOej+GPeQ/
VTLYHApoDRH7AncxekUad/HS0oOuIV0oqrO4hyhftJmOuXLgx4Oor4Oxcx6m58IDueNTRrvIvgBa
cDoxKGHPcO11njsfunMFttZEWILiJUdx9D/0rcGXqvcC7jcb4cLcQU+5jMy6HogApewsKkU79h4Z
2Er387qq/XpcsdYUNTPourlzVHY/w0NOhrFej0CdUdd6n8xSMrqK9rWKPGpVKNcd9CsxDNl50Ifi
0ZaBI3psSGhpkD/OwQphmRit+RFhlJgmktDVCLffVV0hQoWNwTv4XVlTwbyuHNl6xfTSbd1uUkwG
r+8iI91Js0AfzRC136VFuJIFdVgz+CE8dcMN0o1G7qnqBuBIDtzjx90HirsVNNpyz7tMl17+Fp3M
DODAd6hsIJfe8GWv7ivcBm6FJNZfyzTHEtsePrhtjW6bOeRp3pNr+eeaZ6NL35HyZNT++kSPpG4b
DB/mmzHSz2p1dRS357A1ttVO8WF3awXI34UBTDkMPekpmN4IWQYGGUvlzPabAdd7v3NAydp2qsQ8
te3tegwaanoWp9AveHcoNuBf+9bcOvpBAT0iwDJoh7OI46Qb1mJlnQ7IRVaFOdxnly5e4LMorS0i
kp91CUlorMKJdBifmwbJtetGj2+0fIcz20oJbsFTIOpsDmBtFpqdfGNJ3NbNrsCKh4dZifoB5wfE
ImZyLuvs6qqXQMZZWBnsB/kVBhaRthNkNK84SSGMOjx6mANsQ95lPO3n2X1aCP2doocyKKF7cbZW
QSgemiG3ZwZLnqyNFZR54TwScH/ymTJebQrBdkLJtxB3i+Dx52fxZ/eOYqPIZCwXzwj6so018jIO
ek3sBH/uDNXM4lgnz62hQgUcf29scZsmV27rn3addyXNz5E8ZULjqrVhbFka+r06YhZ4TtReJWhm
wzbhJ1Ys6GBL4X/YaFaG3QMqqOBV4qiurtGKZAVwyoDnuYkSXLrEEZCO8RmSuGEKkgX8JAuCVewf
KEwYJHE88iurdXAPrCpRUmx4lMBNIEkOosr+dm+as8ZkAR5mE7zqpf0fCY6QlNkCK39N6dMdNKvn
iblYvqdt1sAbJxdSBf8Djt/3nVpdv8IiX2y++Rt0xxNpRMrNo+HKyhBA+jcvc417q/PYU/HNKvrM
D0JiuURgHC3jqasN/Upo+UCetJH1O+4uptHzt2Mr/C/+PiREcQj8Fvck+dN9DpKeWcMtNqoGaaOQ
xO55GyYAtFTfN9FdeEsP31nXjgSnsoFc2jW/rxPp+7Q11JG4f1u7Otxb5Thmg4aBoFfV0+FiihWK
aWLLyOx09ko2MRTjNWjG2RoH8SbUM7K09qo/oLv8LEV8hp2GQY8QnNkURyUKhIqxudzd49V4mh98
2/8qwy3DX84JdlEDacXFFFa2txHy/KrKDwhX1QjRlPMKTF6nOi+V/fKT0wcoFhT8jEh+WSskhhsI
8dcDjtGhDeB4mQ5cgUCivLH5oAlIlmnwUigSo/m3e9YJft9TaX2/efoIznYTYbWHSimubNWS+DoK
TCXCSJB6mJ8MdUV+dw3et7Q9STHH4NyqKNog1HvzDwxxeHZMcX1pn4ye0MFSHTN+4YwrhvcaCmhZ
xOpjiv18NbKTptjkS4K9fI7vrhzDx4zcVGyXK4g/gTBqOhjPHQ7Ys9GP0jv+19Z4Y3r0jyvO4U7G
8B3Mznq8GlS99fSdZbhuv1TKBwypRMxNMQsndhDbr/RbQLVN7vS/yfgWyD7YE28oIp84Yo5l/mXM
xG8kW9QiCfD4nqe6hdDWkchMce4wxbEZg0xPN1f1sStiGNyRsqGkKGZSeatd445GZPxwfqwepxjG
/HIA8rH5izHe0DEfSoWiyazmA4Is0iU6REPGvt0dH4jNS+ILeJvnqUE1G8TjoIbB1/h7RhyeowS3
2sV0/BHfL/30asaUeYombLwHgAhJqB2bMzkO2zGC6iHkeaB3qgBRMTbAW8zlWybZ8YBZa1lbxtVI
P40XQ2Yh0duGY3qP9lEFBaS3jEZYPlC8GDgpT6XGGOB/J96tyL/sascAuo/p2K0hO3b3xYPzLG/F
Faw/9ktRqbNcs4R800CjMAtIO0EvDAioJ+pgIpprfeQKn7uy+Uaql/genHgvexRBi6QHba0BObcj
JUWALb03odnNMvLb4LZHN19lewfUXddYrEleXSVpuMmT8v38b3JebvhmQJMlkQmmZAoNRixugWar
k7cQA+UQbKnbmoaOttfq2RWFz7jNMjnxhgYLSKKgzf+cjwGsXuNJ/LaX81smUxfkhMnivbOhOyMn
diK2RROoT722o+dCEOoTnNxsIoFWt58DKsQblCmLIbdL+Qrpylf/2lvSqb77u5lIKN4zoy6zp2rz
505nNn23XqyQq7+Qu0urF41GR1ISClKGvUUNZ8T/PsjBscAVO6moxtBAVcjZ8nCfbQ2lg0v0h7x2
S2r92alVsER1A1KyG8gDp30QCFmUxvriAHqxO8bO3a69vxFjJ7cTnkFzXe+xUlMM3iyRNCFc/gWO
ZRto8WpX350j+cluVDnGV1wdcm20KsRA4hjMHOxlzJG6bXmqxsoy61o1JQTCQagppLaUxowHaNxp
lgKkqIqf2YRqpb0MalSdtUhd/YcvvL86SZYtF2lbKJp7yiGYLRDOa9YeRxKo5yf1xeR2AeZn24tD
dT9m0baWjJvW7+8SkVex6EPiiyA9iFu/VCJ5+0ghdFEs8koK061F51cMyG9sCbbTz/pmu6bbqyZE
XAD/IU3gIMd1pfoaHbuQvwCXQhJ7oTbYPv7JZ1tphQduGlltb19FTBJrD9WdAo9FDIjqvszqRQ9H
sgffoCgR6aFfKo0M2MMuo1fTHYi9M0XtHyRg6k8CK9aWS79yLmY/hkoZIgVOrs0i3510HNhbBBMm
BDf6cp/afnYP1Cex26IaFTs6MuchhvHA9uCFz2IBMvPV6GVuwzraf8FHlBfpX45ZotmLpyb/D2VV
D39QKrhn+zv/7ovFMI/UGBslDHiIwekoqceiOR0BkiFb7ZW4b93NCFwZoTOUKooZSmRdjUjhwig+
fq8qC1xCdxln1aH2IRsw7F4yGZFGzmj/wtYItuZUMFKtUS84nbenZIARdeGiXmzleOyv6BWjb1n/
55otKLq7BF5si3mIaynXIvrPGs7AogtxRVgCwIqc4ltvojy5S1jOexLDWT2XacW/7lckm3WiRmYI
dX/PHNAGWDHBbjhiASui4eZAizfswftPH/VQ1u1jADV9nQn0RGqDYTTYlbLP9F//VaZPhEwBiy2D
EORsP6xvCWwFBCl/+/U9sWLapehy17lOfhVTiGRJoB9VS5/N9MxzvwDCSeLhCpPjhXTtSK4exNe7
XhZXllPc86Xn0oZqe5w6+IkPEwKJb0NhnoubHJdp9bQ7cmTTOL8bMLA4CbpXMCVQckOd4IxTSjAH
SnLwjIGZg7Tq8F5u/Z6F5Yam6bn/bFiDSy6iGKZRL/BAX2wynpt068ZDXAZDBpBKz8Qm5zR3kxH1
eSQhTtSDihho9LG2HKwYAsTTO2nP938ucqXYyULYPZ40OuiMuJtkJTHa1snigRMHu2R1IPNXfjSP
mAX0/bss91Ah8Umu0C1Mf+HldYdgqsJK/X7otVAf1Q5hwsYscw1+jTbXrCcUxyVL3r0GmxxBHGcc
KNu/fhubYwsGoxRo4jPgRE/eaMgrPLddsO4HhSgn+1ju8UmxWSeCwFW4rrLBFjii66Z9cibhBMCe
MDzXbvQLNta5LyjY+avkzYWElPjuTo1U9jXHhd1GhBBaKoXduIaJfAqB5YDxJG5ccEOwdtT6Ghts
4Ta5OMwEQoYvg7bxqTARr7gIBh+uVW2qBg0yqLce3UoGWcrZ1V4RENP6rFct5WDzgYFPsKvAPR9o
6RDdoSShMEQtD+Aa3qcnL4Zpt39J1/aDLO+qrb942/yqOSohdFjkrUCZn9EVGwknJBo4SwnxHs8/
XPiEV8fwtG7Ep2L588LKXKfni/GDYXE18DiQ8CyZG+at7GjAqdok/WV2xUY4/2HAWy+sOTR7PBVj
tbBYJzA/91MyhZqxAJF26J89F+YrgOoyGpgFSDm45aKZpLdO9M6DS7BgSXsN37u4PYldq79xZwjB
c+bsDJxJ3k5AxQhoCUYSQU4N2LGx1aVxARMsjQzZLxYJIo5A8i2UHXRd/iXtL8vHRowkTSWBiqV2
GFtUcuq9ZW+2sWsruNczDOHWGw1ebganPgmP4xwxPaaytZ/haDAwUwvoJ1BKYEzBOR/5c3dmEWOa
h9rp/gGqQbbxbO330TUCwXxdr10MeVyqqTMcfTG5/30MqDe3rl68wPQPT54ID9XG+HvWMHEws/rI
ifth999IzzM8zLGYLM1bVYFHpRmAUi8Hplzz/zgaKWjAsn03/xHTM0P7ZhoDu75Wi/yvFiX03vbD
Yb91cog9qSYhdYERgrbcr8dO7MsQ9Y3nAYolSkxn4HmqJ3gaP5/6d2twi8NwvKywFonCEZ2IUQFN
0Lvy38mwaiEQTTOKofdrZ88XqKlsKo27kODNd+jQnTHqsYkX8oj1frX7Lz00uqJ4LZyWapyaqRoF
aLYI0n8Fe/EPAWqZ/lHvzAfBOa3/P73KGAEDN6t+N1rIO0Tbe7Te7DTuiEIYsJUaWhDAsTOnFAt5
n6Jv+EEHw7uSp9umQq4Lgk8o0yrfzLyqoKvCHprqLQJ+dpJyIX53M45tUA78TwYMqSdI0YPEHXyQ
z90UCNBMJRR0FjtA3XN2lz3eUzA4UPtGfHT7Svvo6L4FeI72ZAd2RvhwqEmf+hV0xQN/7Ryq5NJK
ZSAmp9MtFazLYjCOsppA33HOXiumqGx/z8ZwfjtaaXVKdLyoWwtvudaKVTclH/mt6iY90qWhIkeR
AuBjlnajrdJYEhzT0/50oM4kHHDgI7xQk7s50/6aU8r3xYwFBMv4tPkTDufAqFQMHyHqj/jRhgWD
il68gv9c4D0mizLK/zb6ImGqjtXmSbhHlD0cCBReJRtDXIdMLgclmJeyIRK63COSIFU0BU91FuDj
bd/OcksfXvG35YE9CLQJyTVTILXl5ag4lIK1iYNdutnTtFA9MPJ02MZYXoPNyczs25nX0v8nNHik
0XOAlFNZ/x9hej5ClyIWowedqLaOhPNuOsYv35PDa6+Lz8dvclyt15FXFq0gXBuOaAVGmx1dqkBk
HOr+qWSVL7OlC6OIieEHe0T+qbMY96D3GMsX4ycTJvjiTcTcWwpqEC4bjLmQWh7OoWIsAXS1bJqd
mu0XqcMey0Rdp923GhMb+MfaBVw+MPZErBhRMXOtZ0ggUc9fxcEs1Nr4zRnn8bL6tC2gzVH0Wd33
DpAc1r1VlPOjtdJDDoFwwxfFb+JfLiVJ5hUQGnfL3g2RgV74dUZ5RRB43Nsxx8gO8UIYUCX413MX
hVpE0hbcU25/1y9JxnkAy06xo+4g0UOta5R5IHPh0O7z4baslB2Eoj4RKx7jl/knFJncFQ0Qfjb6
kz5NhIF0FYVsuExKoX/nKaScZh89rMDHnubNx2RqI05TuD7MGAcwGLTIScbQjZ5iU1KOOTdvxs4D
LU64+AhlPH8DGV7B9uEobKTmgh+sUwjxj0bwek4mxQHe+Gj8hhaaFmAGFUCTQfVs8objjBY0kTi9
duPC+bw7EYN7w5XGrlAyQkPrkhGiigH/Q9+j/SJPo5+rHHWGWZfF8sA15Gx/aWa0+sxYSsb7joCk
9O3ZikynBezDzwzQjEm3SwmXuTe4PM9FZlh9R0RjRoAVrHLgZl/33luhE8yQA3nDRxbHTcqLVppC
8ImdQfYhdieuRcBeV7M/yNB3d5GGiX3EsFtlT9kfV4mpGbJuJQOeSeajsexIegZCKB+jA2SQuDDn
/FMVXspcS38mzncoO5APPGt0RGbiC+vyUzneGk0EQbiZG/KZydGChGEH7YXf8kpBTy0Je4gN5kb9
OYavub6FlLZf4Bmzo0ZinrsiU7MHd+I1kF8KbUabIqk6+uoLkbSFW6Hn9Z8BFdM2+eNgG/7ker0T
ZrJOHO3zyfA+JZhtCND+ilfyxbuo5BwedkbiERGndEGo0HsB4f50srwX5N5y6TwioHxpPzAGa/ea
5DfqxTUS2nz6F8QRYEc4pWaNdF40B3ZtfCQockA7mGWisqUgKWjTZQZdLRz+8bP18IUoX1GUvRzM
sSCEj+rPRSNTYa5kW2GFD4lR1Juux+Ka1oesyo6TjlxoOSk6wQWAVgOjBbFq/hvx8xCO1iibGAXJ
TR9fBf/9Vc1N5FIcINXxj5p9ZiFHGOPhjho6efO4bel4GWNbL+ZM8+klOyjcZ8MO7U8yAfaRpKA2
d/i8ehrnbnffT5luK/Zmt+lx20NSOOJhvki8C6j3x7cS2fK4z7lR5F74k6+0coo93SuXaTwbuX3O
MUtuC1Yzg9e25MS/DH2de9CAKuv9XeghmPTkXiJILn4vn6U2NkvqLM/vYFxkCRApTokLhOFjsIs3
/T/8hxM6KyQbLRLl6N5FSHSWri8tIibJ0sf2oCWQzzdwx5iGNaS9cbkNJN+I1X58ODrifUHSsrEq
emdWW5YHMLOTg/KfMetg6M7n4fJIxjdQQr56BI47qSKstE173ZnBUjyW874layLcH8dAE5a4g3aG
E+eRKGKc24prQ6BRlROHO0opl7A5vmcPsCVeP+UeCToKQBx0+t78pYF9x0YhvblZd7DDAEStwELL
reQ2vc2mLX4VGxv4gdTEGOkGZxMjBj1AZQBBn5h1LhW4mCvkBTZIgBQgcr85J1o2Yv19s5QW4oG9
OL8XSRRLh/FlGIXkdt1AndloJA2AhBpUh2m6IN3uaQwMLGexCQZfAaWACWk5PEKydkKuXD8LvsUk
/39ZXDM6d2jjGNiVfsDMHcGjlIqESf1k7X425YnyBbWu28ipPBptqPyaaqpsnaCSX8b3NOgXYQOR
SPj8zij5ZeASrcYDtXliMLcQKq/gUCNlrtgCWTLikx9axRd+muSV8VpuozAxLOzSXa7VXldu+Q7P
3KNsl/aNthXptbU9nF/TePIQguko4bBCFnlVQreNqr01h8p4ag0tL8R0wlCfUrr+HGiP9iUGEJ99
XEPczKpUi9oLRsL39JACuAGzzVWwZ2ZhseolaQyhej30rGV39qtxeckk3b9ZsanDzaLzNCYgheFu
i9rJcuAmU/cfeQSRK5R34Pn+Wnv17HcpilpkoyWgl7Cz2Y7ZQKKKVAcuNwuPdA7LRhMDDaFMsNSe
hlQEHHZUePo56KCjL/DMdlTNVSBQyRSUY6FrBa0mFlcpgLbD4ji3KVg1jeuftLuyhTSNDlrOJiiV
GFWIa8tSaAX3j/BKRXGT9wxDGb5q63gbcJ/ryWizGh7f9SSHabZFGI3oZ9AZA6bV94/BVhaJUvbq
YBQjVNudjEkqZPP8bw5vtOnloC1NzvlVtlk8CV/Qtuz2TQpZT4rY+Ei6MqB4SGWalRBym7wEBoVW
KnKh7urufmZ2NR7GF1JenzyqUm8tF+25MID2pgqsvleQeaJvmovYag+q74kLDy1a7yGLSg2NxySq
5E1L49X137Wd2c2YvMoj0qbGrya/6t6Q/CCv/ITemw6gLhJU6QWytaUa3mRuREph89AJCAN4jTBe
Eqe00MRLAoK/UwMxE6MMCTEX97nfkvNlkNeMh4rgAgJXNPdHdbIV+dWyPQ5XigQJkeDEWB9FWHsQ
8ji/8IHya3f22JNy/iD+m0AsMMBatVqPo4Us6wXt0WxPdPoBVbi0B/INOJcGIL6i9OlCrKF/zcLz
ppwmZphAkxJNB5RvS+MfJ2/oo4SNPtUyyeQKTGuaTFh/NPjtC9ostCj0PNycbqWORQVYnj7XRLIF
9LwRmrf0jplypmkF3oHcNdi12ORsXDSKVoJYSSE7KotsCHKR2C80rHZx3a/8obiClugxdDt9TTAx
GFWvUj2hK2QIyPGSDF3g0JfZF35ULeTDVWBwmLSrR7c+h6THEN2xTB+zHuoyoXyF0uwWUhkXb4NQ
wjNruiMHUYd34xx8qXqP4LPXS1Mt61dpags5T/QFQINjUG9QSdiFjdMoZkMo5V9GO0tm16elM2gS
bTTYzQswamd6ug1cxuhWtm5ducD3qZQRT5p9dCPM83ot7euCS/+ZJ/LYcbKnZHJr1yocbXi80kVl
7S1+liLUo35IPhWxpgyXgsu/MctS31NuV7NH83ImUHXWL//V9kgyVzA0N/k72+xJQn/kyZqLY1to
RFOJknm2MPRiPq49pAVVOXJ4KqHFGLRd0rIXr+1f/meujOmxBa2Oa4f3g4tyO2eSNKxO7gEkV/rl
uKGkBzJLZDbs95kj47nwXP833C2A+reaDehAIrWjYdBoVbltX3kOxZzp2ZQUkFYlVxz4fPldLw5i
Iu4p+/4JhYXoaLJulNkarZBbwpNWs6ok/7V2LxrhviysOhrg/I2c2YTzFGj9vwruIjqnz4nLNC4r
R+00lSzjzw4p7SX8015+B/o/Yt7z5W3i8MI+yQ0IO9kvXmEK4DDCrtuPWSE/35UrYagfoMd7HjBw
t5vyF80DbqSXnoDRJoPNlg1m2HLM5O24pv72r9hEbXU89pZjNxbhi1Z0RB01w9znzDKDBU4IpO3F
WFcQ9EijzhJHywoDyUZH+q3vh0XSiAwtsp9V33gaMhe7Rr3b+QabmOKMeIDFbuGd4Xl9/SzNEMfK
z82n38WM3gYWfYQWuW2EJ8dFbCsXegV0ne+/jIWBf+sYA5OAQQBjCAh22muSL0p4rhoXMGNYaH7l
O0dF7N/7U4yT4uZeryGQtAHKM4BILar+K99yncCs6XcCzhE52+t4QWLlNy9ogZyvV7oHYovaRrDE
o+s+As74fFRsVh8MLTa9XKG0pWNb0h7ODcxheSwReqsKoFdveK8kWrbL1B3KpdU3dC8u7tTnvrJL
WYQTLc4KmK6uATbR9b4SPrYV+33LjL/+c/XH9LC7N9ketDT+6qI4r6oJfFnnrN9b8wKUQ7K6VSZv
n43bOZPxy+TJtP0fk3at7CQSWTndKTwG/ez1OuprEagqjIpuirzB8nt1csSWwMQ0tplWPPbyzznk
c2Y+FMFpmh4BPDoO/L+jUh1k1g6ak9cchZeFgu2TEw9WA74JLHWQWTnRaDagOuGYDrJ6dbe24Ldj
EUCbiC2H1D6bEt9CreUhS4JDZ4DcPYkapod/TRUtQEf/VopP0KgyFFiFeZf9QNuJlE4vgdExjHtF
vsXnMiE6EFFq8WraJBVhv+PQdpRQ5wC9UtdKb5g74HmMNKoFyUN0WRLLn1kpRHi6hUOFYRBIH9q0
IPxUnQja73MP57r2CSJLs6ItPCOD9BAzWfVsDEn7hKtPXEFXYSS1zikkYVkDXcmnZ4U+bJ5EUCOt
V66VT167nr+inLdjUM3XnqiOhVVwnUZ2CuV8tSTmD/ES0IiAwyffhY9a+Z2GLjq0KJIdq9hcfll9
uNL9ElCPHK6YlaHX5vZw1nLmXak2CWGn7rTH/guuNW7teCFTOBeXgKK5Ti/P2Yg7axQuUm2pfwwD
7KHpfHViaA1n+TXBJmXXJDvTbqhyMCFTljKUufT8cR1E7rfF91ERUZxP9aMErpDyxgXuq7KtDb6k
jGQ972NYq9dvl5vyhLBoB9MjzLPjt4u9IIsglm9mD+YfIsrRy/CjG9UUTMVqpw54rVttOLTSpEeP
w6TwFJYIcxYwC3CBJBooyEvdU8I94R7GNIQ6oBBIVExepG4HGWew1iyX2Cjv5fVcYE+8s5deNr7X
TjOya0VpKgKN7YqkAosN53ICQoC7qGYBA0u+4K0gRrTtet+oYpEvEQeERcu3Z79eG8VeLBwQ67k2
GNSI2XAK+byGJPa7QfuX/1vFD7DkS0C859H0QAjo8+hgPYngBvW6SblczlXFJHc82Xnm6Or9uyfb
5hez295x+jpOi4NKZt1fvly7YE5U3DIjhuAKs/haq/kgMFvKZwEsnZyPVlLEChbaFvwkJgmZLZ2C
2wFtSDWVCUWeVEJPjoKIiZFtF1O/fVqmoTFnOCH6qiJPaveMoeQQCG+S259dCq0PAc2YpyGGZw8O
Z9E1TQComdc8kRvsCwK7JM9GLJmsK4XmjwLiw9rtDjmUC2a5ngkyloS6l+EpjXvaR+dmu290pehX
NtaJMywW/nMEL9S08psYUG5dmQasks3D+H1Kq36VoPNRziypmHggqfpykITJqxLW8WPHoIglQ2uc
2w0fZcHPVgiRE6SNTnmo8RSbTuTUdDqvGyqUzmHDqHKLWh5Yxy1YMZPR/Gpbtb1hTfYNTJ9RqF8D
DuNGtpMcxSPK/onWOnHoEgi5+5eTlItQkZgg+1GoA4HSO9HA7U2cHoONSbhxXn8brjl7oTu5qcJd
wSn2EWfT3tMGyJUBAL7sDUh1eupnQ8te1oZgPoVZ1nHYtU/v0xEr47fEVyoMMqIQUHSJ66mhJVex
ReoSgwCMWShfAWpTlan0jgs3Lv/f2LQ3lhGQXc2qWo6yqc1ZMxG/GRa/GiWq49WPvTBceYuI1niV
tnkggUSTfsz+IyDpmcG8uWYyjD+MmM79eEnrrjwDgrrpOjP/saTK6dnG80Jz2mDUJZYyUPmU4JEW
KZbL2Ol6u0JmPOugN54d6Pt9JpVQNoNNatAZyFqgiVu8dsRP8U/b68sQO2GlciH+zc4VqpLHD5HL
Cp/5iLOCqvXRxjnQ0AtxWOe063Jj2lpuVNMzn/3F4fJVHAuTqSJ4cnXVFBvrznuuVTHhQQdAX66K
D9jjqw29DQ2cfr7a41FbkelQIsMzLj9RODUag++efMY2fVy0Bh7DiRhe2hsGarl1/48tD4GnodPc
cidqizAsUT5l0sn/0szprDrXTO5zPbYmXQeUiCGOHz+4+n3Vz1EzRjnK8ootY2TWa3bXlriA4mzU
3p0Mwo8k7ECH2LTkUoOZoOTZII4iqHO5dtAoEdQBj4U5IDVR9rWSgQL9DmxbIe9k5COWWSfkS4Wy
wSrV5zd5Ixpy66bN395KvCE1NyGCXct3bn5gTcAkrAU5HqMy67QB3LaPXrz4E1DBy1XnE2RkHjx6
acz+1Vpu3gdZvVNvPlrBQsP+5Lc93rFiUCOaHex1wqpbd7EAVz52ryBV+QsYvNeNdhM5/lDQxoii
xDUU9u8JaIvzUl0r7C8CyIkS2Llc3ltpqyFdQ9KMBqUsEV2XNUyfmWSM65DUjMWX+chfplKRckFW
7hNiiJFNFElJJ/ELdCPOoXwC6eKEmiSjgg+kvApgvmOyBdvd9A/RDSDqATM3EtNs/RvXI9lbk/wf
KJD+bmC/D/b5btGHaEJnXMyVvNcH7moORDVVQ6gV+j7qhmoe/E2NfhbytWaXYQFygWQ5rNW8yor0
C2nrjlt+Mgegary1/7uz+CUD9moNBDVttimykO87nkJw5Yku3UraTI2++QOPKd+tMM9zWH7sdF1d
7n5cjzHv+a1zShFWDTOt8PejQVDJpenDe450SgqHQUWyjKJ1lZxLuBOdck/P22P2NHjw4ezDBp8H
gRrbHup5LUwsMyrGq/LaQoG3u/n19QqGRP+mYo9m4ChO3srdR9KgEAAQ8G7d3A8opKIBv5jEdMhl
uUS3XMImXyJVGchB9tD7k2hg4L4Y4yDBWZ39YApEbHKmTu6NJQwo2Sk/MyHnvTXVoB0d0DNqY4Pd
it3iB38ho330g2LjzlWjHzkLK+m+DisY0yTYxV9SsbI3Ut0vNZo2pN94huMSuv2j+hunVzsJiZvL
bEkTxGwBg8uFbU4DrhDtszD3KB7AHwY1VTjEkoYZxL5m/JzGLkz5PJ3Ce4tOpnVvuVXkdIXEga/R
vY5KgqJloW5jNmwPJh+kDGhCVW8s2LQjCz/Ms9YNvDUTDagJmKRZNCwXVdfR9UuRdtxPlVMNomyA
4jYMnqCXj4+LTmRXOo2uDOr+TY5UwvOUPT78yShUfZhS85KJUM85GXrXgUIIEG7eT8/Nu+WnPIoj
bkfy2i7NJSfZDKJxb51Hqdin0ye5RMU6h9NbHtXvj1i1PwiBMTfUkjPDxLMPI4t3h4X1ObU9wV0G
0iqxFVb90uPvCT0NQ1aMJdHFSZcIxSYHVQ7DnF8XQKkd8YHyoAf/OH2noSexvvZBT/6Vtv/9+Fc9
jWKhre9QVQuNfTx4x81SVLDdApT3bGIUW8i8GmEx7Cb63Dhc4Dy2Ud33tdIsOkY0SSkXpbkaorTO
qLLjjwxWkghT+B94EXKbjwqMg9U4ZUf1Tvj029PqgXK1FGonukfvC+h2VxMWxhzW4uOpyORK2wMv
2gkllb3gSRN+LzENfjBK6hlepQXuRTErFSOm4OP7Y5WTjgz3AzP4JJRM/USihPmQ9VeJLermOlM9
e+hiG4s+s/Z2SQk7dMH007EsF247OyD1ICqhn2FOwSLx1+W/7dPZefDKuyzHdKS6CjX/IKEGh9eI
R9N4rEjncz+kixHhZQtXHsjnMCneu21oOFBBjr1E9KsW3USqgiHeUWBJkU10ZWbDm3m5YBo765Hn
9GGdt8SrvTgcpKORecz9560Em3g8+9D4zh2baqTkuUQzM0clVQ8E6wauu3e4j36j3Rz9lVNR8U4a
UIqwbNVFPFrDQ5joVf/1RwJsZ0mfj8gk9nG3C+GneDPQ2pgtZtuq3CpYQdUSMV3xnVOHwup1PCg0
UY5rZSdu3/P9UGyMPHuyNQIk0jsCq9Iq6MvvYprSKM9DsNwMNBXzvKaHguB59Oq13KtdtTrvOgnj
G1CE5kbCvwzPYhhpkWShM2GTm2pqKR9f4yyZseEvWTTqqslsupmvkyRl5uUg6zGHYeFyvCksBmNX
S4X6R3evXelYahoeapWtv7TQ+gVELLYs47+DVnZ1+NDnCrheJELuyT8FU72b8IoiR+X9JnB/7Sjw
Pgt2D4164GBExQNFSoqmQI5sBSoBEVa//9/5Ul3Zxxi4Fw0N7FThVfmDjAOyPDYaMc3R970ZPGBa
js7Yr5CQ9psPGhsMIJXEf1jPscFS1pWd3t2loSzt4XUE+d1zsdS66bYCg6gIyylFnfhYW19SQiuc
b4Fz5gXtmZj1andddLziyjIGlbF1qwD/uX+gOc/nK/iI/TbaCIkPStn3T/bTCPhrNDASw3st5+nB
qYfhhttnOV2onUr7kv9JU6hCpMzabU7brCxJC18G6Y0NvfN8lxg170x4AX4jW7rtD6j2QRuhfIZS
GGit18mlKYR+bP6O50kfnsMDMCGEtVP5j4xfFOXnkrL6lsDsevZKstnsPquo6l1RgwStMTXHS/99
Nwsur/EMS1zrdSTXsbxX9XcyBTxXbEViv+vh4MirH1Pl8dM4k8PpXJfCbzx3QkVDXO31CuN3uW/O
pQ7MDdSC9kV6Gb5kuo4ZvU36sy9AIuACa+YaccoPj+cgLUymrUq9DctCd/i/7CCQvNwAxjmYC0BT
juK5ufCmA4colqFstM8sDW5EnEB2uWJ12uQErAc/ZOry7f0XQ24GEIYu9bLCSZExK1Xy0oMlHQLb
0oA52Qer3buhp3nmZ7q/G3Xok8phzQEO9Vw3IwONn0CkNwFU5iRvcZm7k4sza5jFIbb3Jsl2XMEz
b38ab+4ktvfc2Z9pvW80ZFs1uSLvp//p2tRp1d4wwgarzcu+33zxA2BH7ju/xaULj5A0M5Ly13e+
J+N9KVH0W2QVPAAA2vL4MHlyisPYlaEn4PytjUtLeOvgSuOmQfgNcVThvRt0BVRH81MrFNMNBMpE
pYTqZ1ClLkpMlTEw/87Wzsp8cNoq5LrN+JbWylvrKeW8bC1a/2c0roMvyy9Wt1yVrthMbRD9klhU
N46PqS/YZP2CPUbAxhDDxWdPdAYuFl1V24jgUu76ecwxrhW5s5JViRRy5bfvDw+Zx8dKvlGfbbj1
dW20Jsm3EI3s6uoPXcGVlwqvBOebA1a5w4wgd7uhBbS8sCGH0U7M8FflGlRnOLQ/9YjGsn0qY12k
Wk9rLBNQdyytYhvLHstTCAy8W5EGs94XC4bS8qmMrOKfNW9NCVKGCGkK31+kJbAS0KfsQjBNC8g6
xjvjtQL29waAkN+oxRTwt90T+2MxKZdctKBcv3wROq1Zt6veL2a5wYssvc6eXH+GdDxy9LCq1ys1
f9GOMD7nZG+AQgqdEgpfukKmZDbTqKiTokX997txIL6ZI1xDlDceXWWzGb+ctmZVgVCUmAbRfSNH
Fz0rjdc6veOCAXe8XpW2IDS6i+EmUrQlEfkHyUVthXp92TWQp+B+rrtTw+os+xgJjviJhS+4Zyl7
Jt493ulviShiXxy9h0voo+LuMbkOKT27+8OL2arcShedl+ZQho5v4d4Nx2KAFt5aizVmVGMlAjhZ
d+wxxnSDqO4HPE0xEt0HyA3XM8UPrNbXUu9SO3yllhpfjuizWErUJV0LsNR8Wu36fYW76s54qTkw
WM2ke1rq3i74Ug72QVHxvhytCvD8Mw9W0TYa+UJohAwHOvNoBDYFOpn3Le3c9jqwGOFZOvB0Vvtr
6nbgC3ctDd+qdI9XeHwQCTvSzKJDBx9eXWJoGE80aBrJSeertAfCP6oLb7oMRqKIsMZapmUS+GV6
Th3QZ/Mirc/tWP8G+TJFXCR1tLphrVvLp2Kl2HshPdS8h4CRbAMpwrVDAb+vSO/Ae4qVHFVOeaZD
BXM4RTo5JgmXTGCuXnmp87OGrsfN5hc0+nbCD/ILCGhciMaOFvgnYwb7qzU418ugI4sOUbiFUMo0
qZrYbjRYLv+nOp1FIUMxO7PqkPra47LUDFWnkyAE5PkIFFkccNxWIpoYPZHMP6gwfZ8SKey/E3Ca
UBuKpwsz/r7INsJIATF0FBhCHCv+R7d3ICn1KTjLNPwXwssiwki+zz76MWK/rl0O81rGi0WoM2wr
y43SsAwXRPXVrRaLKfWFaj2hMlio+tcs/NYVqwkrVuVQpZF4jRNJJJsHPlFJZIArVA0Q5u83DgQt
PjcmjBuo5ImZthmj1kx3P/LTKvCfXTfxsOcwRg8lJQl4bDi32gA29+2jEXEsNITzebKUSWcNdlSS
LpzmndaKS8EEQ2bBZm4WZvq1zAsGtCS9TvfhW51JwwhobhwDFwoKq6qZUNgPYYstPJMY25/KDHri
G71zKKiF2I/cvlCWV0TBerDeaLwX9ysfeWlw2Jhq8P4htK5lFsHDPk6T0+VrugiFBbFJHfKd6ZBH
gqNDPApENH8sa/8HGr/iI0oGNprL+0ySNKjTNOSJYEGwASOlCliOXNiBfVIQUzAYEZC/+ebasNmJ
hIEQD76cV5lFsjCdYee2A57K+Xda2piXrSzSMUu1ihrs4hrW8bTyPcxmJnTg+k6+jRNM5QlC1+3M
b/9Qem/q34f2dQR2WxlCLyqZH6ZdqiV4qS6pdXT2qk9WDUhucM/0a8OR0mrayaBG7lLRZs1itQB0
ufjpBkT5zV3nQCVSCAlxtEfm+g38/GrhJRgR6xcBKDBlcJy8j+PGMLZoW9PxNn8hKa1mNOMa9P6L
FLfbbk+vUTK4E8I6tSutNvAcx+3PncUk82IvKRgAQTF+YrieO3lVW8d8qSUobSbHH8JDmw678dId
QYWP/99JF99NbgIKwD6ezZcbIrxKDx3ijL1dR6h6Gh2NbYPw+3Y0AuQnOnJkf2m/qv8BEGY7Lton
46mjqezlvnSkhL1/PWKF3Gazrmxngc5uWg9xb5JH2BO8cOy7uf+ZDVshUd0Ct+tlK4TA6LEH6VHJ
sDXGD8E8GTHEq7v4tI5cSvd76o5dnhMMyCn1ZAO5vhI3VLmvjIW+VLNZR33ZGBS0pX7laos/6eYs
sQkxKPU2CiG1FzXdnzBZGZXF+eCFOsn11FkPk6ejKbqN90WBc8G4arZD3cqgVvhRUX22poWbmgwK
4YbxAAOTzvZSGWJESVOhpa3yKXgeljFFdsdMzuhzaobRJ9YYSJkvpPRrsT7is4l6K8JR6xqSH47w
fBwKhliopEHr/s/Is7+QUD0fDs8RKexjIcuQwUTAenjMhF6Qd/Qf/aErVv9zQC/Xckns2+TQV2gt
9NgaDqBDXqai/8iuL048sSxxS8ORbTpoQZN5Kjq5a8CbcPhxVDyTOjaBBxTlkEvbzJb6cvUNcO0k
ILDjWFBtyAIIe29Usa8Mja8Jhktqo+MfzRxnJbIeAMhFFyX8THwcpjnH0rpGvoQlUoFRuutkeXk2
G0eallWhr+ca1cy73E725t2wD1/tmWxDE5IKlvn6SLFiWL93+RTLsbvJqNkHBvSmR8YIcUNlIRub
lHFW5dXqPHYIUWa7gYb2a8RXouYrAK6IBrL3jqe5B+mV/hLBAMMfl5SEaOUioFhT3AcngEbEpcs0
ZE2IYuxQT+zBWyMEKF9nw/5YKlcafZLewhUWMjSewFbMJWlTDpmaDpOQQf4uva0Hmghiv5VrTx1C
1rLXfbdMCI/xLXRANxIv+KuPKwzd6iEV6af+dAaDW1R8Hf6LM4dORMZzVX6F6Yen8hrtq/oNDLu8
P9p5tDYH4usUqv0XI7irhNfQRgn/Ghy4CBqU13lzHE29u7JjlfDuA5v7TGye77dGSqQkiNecYxkY
V15ln4BTVpXHvu5MWqXwaPneBXlO91Am4grX5Dk2iEKOD4XgqB+UjsaMQlu0GBAT1pLX/ErlcVAp
AP2Ugw2X0uPClu1n11NcvFtKawhyvtQFXFGaudCIf9hPMnOKOwvtiddSRyV6OkjZtIScPlSTI1Xz
4AjSRV5iDDqPHATNa2l+cDsLCAV5Nfk7lknhuYOuKfasmWnkNbCIRm+C9n4FXa0X9OvbL/9OH3Xb
aNKIJ74KFyeFaTEZrfpocwmhCXofYOxAijWoC3qsyueb1YslCrQLZokjYUo+mFig2knxeO964ivQ
buyQVIWcbGqNpj19JYgHSOAg6NgPZYCEwoX27qaJ1FxEABHfKf4f5e0+OyMX/GgxV4C5p34Qhmxn
tYhcbxzt9uRmjrO6LXckjqsg4/g6YQevMijknBCYEJeJqoxTeaMBBKT2JkpdH/cn8p6EXnqICDrQ
S3IV4JFi29L25F4dhbmx7YxdS88I9yUiYfpHb2F0EIp6MOHYvOi1zOf9wfxIkZOGCFXGFTqoaLFa
lTFa3L0MJBjE96iiWDX3TDCvqFXOKXAfz8Vj4QYO3DvM8qDDseyqjzA4pRN/jE3dGPclsJVPTgoy
i9aLOwCQ57GMcAUmfJhIUEmAkjCT1yNOC+3SV3leUz1TFOghY0CoISnNz6M62uUmO5BBeyxzd0iD
xrYhJwxrDjxTSvx546lf/vp4OAxzFULMsn6giy4g0+RjcfFT5ykdBHpO8STJHBt3uDuX/doL9e++
CRRxn2BKsmpabZKnklTAARbVfWc7rWgn0aT3bYjqpjuChh3HBzl2wick0WE5ZyCrVDKl7j0L+Yve
EYnspLUh0uvCDMgjrL3jS5rtSeZcA6SeZH7aKDFd+mZiIDLpJBmdhBGNGQ7StK/+pA0QFnthVz/F
Q1YvIB3PPO8sTOvl6pT1/wSHt779UgYXRyYIxsGSHvqYk6xB/JQdhUpfTGNtlCnVu8pvCOiU/uyE
hjxmoNT8RK0Wp6C93xdozBkzZwX2Zf/piOVSVuanx7LE9kJfDv4M02scfExjiMKr4qHQf/CtMUdi
Jt6K1GO2ENVSXsYf+KkYWmaLqzj3Lun+/HUlhm0G8YRKVPNBJ0Edat050VrHt24XPz5ttncC6fuW
Mt+x9lUUxXv3dmVPpJYFTm0a3uH3PkXrW7qbEpGI7ZGA9i4Q4Nti78QGsSehccG/kuvLuG2Q6Fnx
q1Vml4pisUdZk1loXqPzZtC12RiZijuy27gDiWv/1ODC7EHdyRxSvXdOpCyyjPrHs3mlp2ngJ5AF
AuQeg/Oa33FiMEwd3U3HdsT0i3+oaLLGpNXc6HV0gOU06NXHACJNsubd322+Fo8V9xP4OwMtvH6e
5GuTHoC/KIzhSqQYMVAuk/JU5s1uYBdb0PKwEM7crWbmV2VjvvTWSTEL8/G/GtD+skabapnGjbke
E+xXX+RLjqTbqzsFZC600AQrle2sO2KMfb9TPPV2zJydK+aTfobp1EkyTwjsUdbD2HEV5XpD+1qD
9guHZKgXVJ/cfQmob+ZlsgN2Z98p/DInzvXnLrMVrb5tmwNFnyBznoXHJrW6e6cQ0P0zeeu7smQc
7+QJEKoe5yZ28A3bMYzeat/k4aA19aAnwFSHRXx7+qUkzhP3OfmB8O0i8nOLaYPStD42IDHMZ0DP
dOPjDy16vQsuZCF6Z166J011dANBzB78cQhcx7r4IvNhm29GooZAKMtW/Lb81VrSivX26y9K68vt
AX5GgwUHyEm+L4tzDHX2C+omtqPXFXRH3PUhtHrnfrbJx/oPxDFu1kKa211z9jxDkPhobf6PQyvm
oFoFAOvcppY2YdAEZz1x50oUOoRQ+/wJKBZ19IBnvgVOSiZFFweVt68xMD/dLWH1xKKgUqrRKAeC
mydrXxe2Za3fzqfQPLXXSVb2MuSxT7UHfKJphzrVdmYb4li5R7sj3HGd/VvB65Brld2reIOruhwh
r42whsbXhR9o6/nyla41eMRlK0iAVfkQuaUDE6rg0CNMFo1P75GnAftAFNDMXvyZYvKLG35V0dXm
6hlLzcAYEIrC73xzLJrKRpCIHEiS3hjqxEYDkgIU/6EhnqMRRPpBMlOXLz7wJybF4z3KvbY9j/7G
21xm8cEuymnirT6ALv5LuSpRSr5Xbsup6LbzC+e0FGPgjO0lkneLtzX9x1e1/6JBbOGF+b9QOKQg
5PziIbs4nvAiXZO1A5sfSCUyQFCwv1KJLBQ97PIG7uNQQPWNN9NlUiE6qZT+m1z5UEOcaNPcaH+x
aXbi7m3L31vsDe5zidTpPZVDzKvqyWl/rWqk1RyXNXa3KsV3UC629WmlX6eKklhSNQGGzk4SNxlp
4K21C3Ww62ANfro/PlD147T4/tn4vIeHzXZeuBvdP+L97YD7P8g5aI+pbOMz32vLGU5H4uLq52Ac
116/bqQnxrJSYAxVkCVZtRykYBbW09Iy3BY8j8uLMxDptEqns5myh7FdjTZddoZIFyDBtXi3yuIx
QPQpkInRyDBlGspyj8gqpHKgf8cxSKgEhIQF60HGQOaArlrUaJ5QCpv5JU1hUAwGgC+u8zUt4fdo
6HBYHlzIQUc4+7ax0bAaJmhZywbDKn0RE5eTWDlyULhZklD7jVEN0Uct/NKLj2Yt0LfNrIj9sIzB
yLfIyN0AUmNFCfdvzYOuaHIoWMCgeELbpCU/OH4jwjcoeAzpBgnJlVWMzXRjMkjpuqEtJbRAEqGV
4ttxEVxTBjrPCLo1Ys+YNoQ8hQDY+VBs+YVtv2QYEZTXp2XjRj6umNvu+ZX73MTnewkwLLIZGUf4
UBcqxJ83ZozsppBc2ifqc+gkByajAH/Xrw+F27ZmZEpN+PdNpbGu/BPkypwaDwtsoJHaqXnQqIXH
GV6BYRDzQw17JAdF+q7k4UDR2VV1EMn3bS+/a+c1NNp6TOBJE5ObgCb03GPl8q5xFBoby4Y+OoLD
l0+k/yt6SjJiaafez3I307ip7Citt+/2a4B02gwhT1TGbvxwxulShphuUsO6LaXhLgLZ+Ps7TyWO
EwcwYOo/dJ7ACryQvC0ekMzt4T43VKcYkV4jPlCnycHeT+eKOFywBD0Wl6Wgp6VYLA4nm5tTtxG/
e8YdRPc/Xw02BMTT9F62lK20hVqgcV8nZBiJkQxkeSCz777dFbRqwVPEhQEWtK8elWTSHWIFHRms
BqVSEKGCyIfQhtzYah4RKTujKyEZMW9ZGufQHjzTC1pEJzD0AdNS6bxTGiev85HSslUXG6rmkBML
uRkYZru9wfjgX1I0DujU/QZkkOG3osjEXDv6Gbm7X2DOHZga/ZbmG3SUVKhSfYAvW7BJ/GYckuxq
nw6tb3z9XpSFexWuy7kmMo3uKKmS7aeFydp4VNWtfNnAE9CN/j4mU4DPItiHIMoKj7PyyWXiEDxi
22w1A4wwnMHLqSddRXA4+V/HA+oNxC4lgn3Z9ufIjbnx/2HdX9KfGCa95F3GSl1L64CCtwbh4u8h
XVe2quS2kGowh1GSMRjzQMuz7FyOQWnAEEL9d9W6Bq7sImVH5/m9cPBHKWw8bgg3nw7uqbn/u9dl
t/qMdx+4W6OAIwgwtueZixpLyLXnaN29Mf1//uFxteR7bFVYgl8JBsWl9tSF7qC1dpYUIF1GXPGF
LeAWScIJbhxosQ/TViF5VecN9Pxu52eki+4DBkduGbMErX1nQnNNldXsngfEF0AiEH7hEajE46P3
3/PVaCNO/+HV5ZGirv72iHgTz7J68eYGillQbIGdlUCuLlX7udSj+FAN1tVMW9UYWFVcRsRXvkWx
N1D76AvPxD4dXqPd4dd45ViVF2U/jCynROW/XRnofuzHgyEHrVyjYgfjE7P1FnCtKTDAHvUHfP2V
cdfKGsGvIn+OEt05STMb4NicJMFk0Qt6BpUXfAoQ2Xd1rPswBxFKgoJpe7lVqj19SERkfJmQNk4/
W0KEmp97VC7X4LCsjvOECL/Ubt/gc26L0HUajcrTNEo5cXRf6TdzUVPdci4A/rBmFssVAVbdhUrV
xFvTJJ2gNHC25w/VcNMH9hXEsHvC+t0BWyphuCKXwstojvOcGoSBv2sB8elqdxeT1fb9NH8a9wZM
ED1jJc7QzfaaiH4RkeCsShIAn+9FD3GuuGkAawPVVBbcUHc/G67N5Qoa2ZacUMVq0ben7zSFT3cm
2hMvxGzkwOuS6XMoVvnK8NOkHr7rE8x16YcNCRmWbf7Za27n/AHcQVP5VNYMnJAVt0d75O8XZjNi
6d9soUyV/zx2Oxgdab+9pau2J+N/UG3FS5bSofkQySHmr3BAh/alHuOUovSCfbXlzZ4sZB69ROK1
R05QHGBA80ZOdG4jHfwaPVjnKZQFXtQRG9UX9QHqto/AfCXomm01PU0UdvhAPX29xY9QaNiKh8Vx
nll9J/LT8Z84h2Viehr2atL6+wTf86j3M2+N69z3rSOFTbuB63rhniHfNgS2imMkLlSATed5zQ0z
hyyOhiDuOsjXqulUu466YMae5jvzSyE4C0/tZ/dw1VcMhwN3pnXUQlxjEn9Zd67IDQ1ZruHZ6cq1
Q3x7ZSU/AFvl60Pyl7eLmMtRZES8VWs05dHgtvLJIYdh+zmqi5cLe2+LdbEYTKU8Nr8kmFfeiQya
ceFaeQqv1gFYvuDylAKTvvh7Z/wOOvo2AMGm/PD7afzK2ekB1JN/mD9pYNbjdiAJ999VMH9FnSrb
ygyWzRLgdzgLVBEYUfu2jfYFujEumcSn3ebTx2Ei+8xSUevourB/FvGG2+ST5qNiIj3MfxUSPdqR
iFFTZWoE+m7+5dxpnixu1yNFwn0eUwrgpOr7uPu/aYfE/LdgtbpTy8ZjZnp9ZFoaUxV9mm53jMap
PKt+FZ9sAqRr9fufJr/lcit8Zs5yzlQk4/VgmSSgy+P8Z70qFO+R3eqI6epeh+rLQmrnU7FL+5PX
Pc4BeB4b8oHNYn2r7TJWYQnCQGatAujG60fWBi2y4mPBCzYbi6Yx+x9+EXErHBXvlUJsAAjx2ie1
Rh6t9llyP35B0xAhBVHI9txgYxiQBbx5Fcg+Xo4AlDPD8vp0e7i+fnezRsXhlGYM5xht0NC8M+p6
AdUt0brhicJbm2JyuPE5/LwnesfyX0Je1whBIPVGIzYCeB7sYgZLPFziJSxkLbDTuJV84hHb+EUg
tH49oa7cxmwEkWJNP38cyXB0Jqld+HEjIx0aLn1KZMISicgUnieVmRcgCp2tLCEnSsXYSqT/yzdp
/Aro1YqS7YF/YJAxb/X9pYfFCAgP2LKrZ2xbvPDpgedACsJ4Bc2gHc6hbWLiGfUy6CiBncgcIhPm
WXbOsUBf+NaLwhInBLmblOYzWan3xs+vO2/LnEdgMKeng2QHppomt0K5+parz/uJx/Vo8hbPFri/
vt2T150IMGsY8zvliADfG+UxEk/qNgqaG1xGIZnsRz8AjUBgKqY+Tqkt5D7L3O42EYSFTZ8hb5rm
PZ+VvHhKmSS9cAFJUGQptpEMgtrGIslNE50VjFwoK96dLLaLIOQfjIqiSTnCf2L7su0L0+8fNQ73
+En/DNnIDWE1fxBP+0+vzGMv0etK7ucqNj6Hfyz45P22U2yL+mbY3PO8dD8KBX8SsbV0gPF9+Rhc
8EFZmN8plz/ZK6hqzmZbq15hIiT50Yr7vqE6VXu3s+BtGaHpdaZGmBGXj5teTvkUasAUiIZwM/Zl
+1gx1qKhhviolENQafpRqhhmntAmQbuPVSBQD1UxM3sk1v9S73lVegZj7DSsY0PzuXSqfS4hedo7
wMY5eS/WvCtH1uMBTzyfPtrl7JleRUnBPJFZqewIxwCNlxwUOjhHah+kJYzBy+6lm2y4tenstG+v
k4OYzZvyWKYWalX77JRzZQqiElXaAohrDDfZ7GMv5ZI/paOpvIq11+WzPWrw65MoMiJ7NdCM6L4J
aA8q0ha+wNxvrM1YRSWV4jA6l8mScwqfIsN31B8403uyoyBr6PsZhV0VlgXq83euiokKfAD4fRkW
gVlbDYz/m8TPJSg0X+ZsZ4Mxrgml85v4UosxJXoQy/EFc5j0yKfGbeEJHUhon9meqfWTwE5qKA2H
mxYfnUgfig82GNsIhjjbe0Q6Vzw36D1PgKlpnX06wwLvsq2WsTReZPi38TpaRshlyYTX56EWDuNK
LHkXoKE8LVcaubRQJ4Ob0lcNCHmhiUlb0C20Erp6vltIQXj/3PYB8g3OG8CHKWdqhmamYLH38F2H
xiCOj4NkEPNvXaKcxgMvtt3QU2SAu073rbfkzAAJP9kx9EBPTo6wyBVlALG+AKr0X4i4SCbVZasO
Nwsv677YgmYMttozmE6xuEExn44eRbxa9x35f+yeMrqp2c4rmEFcCyl5TIq5MwqlV+Fo+DoKJ0KY
wA8JmRK/uAWYiAp4yTC9EYDMiGVRs7cYhMOuIMgR6BJr2vZJ/v2ZkXwOTksQzFDQn/S+8EOu0wRu
4TAJV0+TVEYmXtgqvgMhjECU/B6zgTbyoTiAiiIYiN/m7f/l9IsSn2vkupOTFJuZGVEPKyxnxhbx
9FB2o+gQ2xaohWk5QMbYaH5m7X02MwgAjRHNFA8yB8aJF+NLglzMyyCSNUYC4g36PRYY7IqZI/EW
NQJKqmwgGrtHwecx0or5DjjBF34tibTIGshjHqIuk4V75dfx2ItOltPecfpOqjvIkJhsdiuYKlvb
T7tbsRraED7pEKEYawnH2d2ivoeFAZi8gjXh4nxrenLjbhYRb+9KyywTKQZztp0GAOpUweRvbLaJ
Fj/WBMzV5HfvVjwleBELBF1Wd3RbYdLz4I1w9xkouIxotArhJeXhmgTpc78Ihukj2bUOZCvy0eRu
N2ROHKhbqTp4dOMiXOx0FDpsV+M1e8+5NtVibtmCrYhLFwwpwiVCUevmZFof93aB4g1gRSGOZr/Y
iiVJgqhNXcOXgm0NXnMDjRO+7w7vxHtK+8py8GCheA+Bbqx5jOw9yTb/WHm4uHsc26CYPLrc7JiA
yDluU26JR0WV+le9a8pysxqN9aHUHs4CA4tJUnsmmtqiMArinhZqu8vs7UVmejgWflY7JQNa2Pen
VulrZRYMYjtKReNJKKhTS2uz6291rsp1+V+zwXjTI9YcuNl5kbNlXa/A9OmQbw1j+74iISxD07E4
7kD/npkUOENiECiDwf+4hjm7XS5xW3bA36Npqj+7U6Ce5PXbsrzBp2d3wYIXoNU87c1rcf/ANSZ2
sg60qA2ZV0pEOy0LjS4hS4y/7di9XbxNhGATDZeBbiUM2MzF1rmog8omVKNPmssK6sOUKLkuohzH
Jt5B2cotwMT3gAE4f74MdAVbRTnQWAs1VjIsz+ofCAXFD9/ZRV9j2p+vpdQ8qK4UQIXxWOl1Ic/m
EnoFVYYIw8Y3ul/731QQ97NQOFgQczhexjrbuEOI+MCWpQWge5KUKDdnnW0HldyGzbtf52D0HbpX
cH38obRpjmeVcnEA909BEyGa8caxZbLVh0++k9ghT/N5RRAj538L9iBS0d5geCYwNoUjimxPs5Gf
CDE9AfPmPUaRFNZdCy+hGax8PAj8qcc69vw/Ov9KDLGnDPYxQtwoFQf8d4VbDwsxWjobtyGmCNga
NtIukEK/DwOktk34rZncS7AhEpPucF55ozrs36kKbKNa74qwzYRI6g+UBIjf7W+ppC1khTb9et/G
4OyAO2aSBgJO6B+4twPhmSnqNlaTA2Gl08biJdbXiQFmrQCz8aQLzXHLZl3dkKVTzlQ+5dlc1btO
bOnE1FEZ6GojNRR3qiVRS/mSq7bWe/Ld88YqWie1PSZ8HkeEwyunFbtB4Fza8/uB1VwmL5VWFBLs
CEhCALNDuSGmYctDB6f4Nv7dmxqGBdSwwvqVklVc+LpQBaQzhn+icfNGm+E0xY9uPSOchGqy/spm
QjyEpyguS3v852aAaLIei5T+4MO/t2fsQAUqHKV+zZipvB0R1ekL9fzoevwAOhL7l7T9bJUhZGgR
c1lJMWw37WYZWdze383/ubfv8iwmN4zTT30th04brMXooB5bP6o1Q1ykiVt5ffnO4iv7PXc7ujfJ
5FMXKmn2TN1SRwZcAKUkAjs4N9aokjZAxsVi9THJnPoReLdq/+GyTgYW9UgOpRQN4XEIjlFSTK4h
ZKFq7oRGMXLA3XOlAMLiuwMARx7eJQG3pqQII5FrQstBS6x9qvS77cEjSKoAXy7slL3/3Mw2BySA
EfopufTlN8adVXp8h3wAQw7zSmpLOb35VzU8yjPNUcll6gnOoR6wQYftN2iuYM0Y046GZzgO/Jbf
XMFdjzoV0dyxUd0EutHZpTdN5JjeZGvQKZYpqtjfb13D1StuKOb2y7kNrsoim6oexNvk2wrTSWqn
l41+af0PdPiz9g8TPHt+MoIpwDcupDXyXCQJw+cdLQ9A5A0FeALcm2z0VF9jJTdFhXOYVKebNqu3
0EtL3Bz9HvTTudU6GackPrA4wcNPk7+ekb0/95aSQw5v59MkbTM1FCvXPX+rFmb4vamYApd7X+VF
lE6bEiQh9YXRdQDUQmVnscrLN110u/UhBn7sdeI/ZhRSHu0tiLsaUkmFObGthMJLJ0oMwAweLmSU
m3I2ZziFwPABTiyf6QCgW4kbrQXtlUFy/fXHbS6is3BGvV+eSdgLvmpB8uib/Kz5RFdA7DGU44/U
LaztMw8xqBGfcqrrf7jQA+RGBhTi9QeuGWXuv4I8fTbH/JXrEBoZiNMk2DIWZqwlsG/RBkrcuWfT
7faaND2K74ruYjBGJDYv1fdHEt38XI/V5bZ9g3j05hfKV4bsKOSyjKIyEyq3cNEHpfjMq43n2Bi9
jy9pLOHE/fOv5nqgKH7uN8qXOMQDZ9ufG1Pw5wH9oXzmW15Dg+te5kLM19V06SD5zMDLP53j4wKF
dOH+9Glk+CCR7iVZ9MT1KFpoUJkPUKMrEAnflc1FK+vFnRxz4H9InMu0dLuaHyQgJTjhxpWPydzx
L2O0DNQckBpp85xhe7ghZscNd/Q5dc+OVpoTS3iL6kdTtxuflajfvLbgPBR0yoD5+jUt+R2zb92W
YMA4fJNfm8uSo/wB/fBUq7JdKi8DcjrvTM5/LCefFiXtoeKi3XHBv+sPbg0vwi5TZ94sgIBn1yfD
oGT8JFx81SHQbEc+AHU5FOOh72edDx2l8eENRMWghGwxccxUfzvUh7c7UjD5IJ5618kzuJwQbniD
hJW7aJMT1bVJYpVeK+n+suhTRnx/OXjwu30bXW26lfI5niHPgXCLVbDN2yoUgs7X90unA9ZkJp32
WMse+EO0+t3be1Rgs/X0mjN7g1a3NJVLQgVxRwespYBY3VyT5lr69l7H87/grQ8iBoeykTviuCgz
ZvdgvUmkddk2fAHlB0Y5vS2l32xO/MxQhEd9oDByHQlmOts3eEl3PuKPovEVq7sC0TqY7E2J2Kfy
aF3yKrYdClW9C7XtHBQtT5M6SHjxTA9hbykYCSaXeiH+jvpFY3DDRHvChCFJWEw2l4a/jsiNN5WY
WfbISwoskM8HVYcEYjPEy5jFIKxB7EpPGsBAxeKEU5+e2PBDlubiq0GTql67eUF86bc1L3/T4lLe
nZ1KeAiksfWEnkcCQCumKegnB1O5nRazCVwMO8iCpikFUU/s+ATwRRRRVdfu2xPqHu6W7IF9skNi
GZeW51YmDNa3NmEIKbr7WkS3UAd8MY4dBQ7Rgvx6hqeeOqAdHh3Y1sb2TpCztFJ0ETpiWQk1+N2G
872AWsptzOFfKtNZIcKHFZqdtTisG1zkkK//wleL6fqAZjVXqNErRPja1LmSRkAKCkG6Z1OSqpRC
glb+ALJEdLLgrkJwPAhjEL5MO4nhXczaRP02z30dgCy42axfRoG00EmLCQwXn4ipyP1Xk/OZr2YW
q9NykNdcYeiCrg5+rKUp2c7bjs4ySAJSUaL3edNNxM4Wym9pURanLj+V/TUz5DdDNWxiVPgq8Rj5
AreO6oJZ0jr9qEveOzPlPV6B/zF+T1XEDQSfMQMFKw27jv9tVa7VJLtl9ltfkbsRUhopNgksCDMF
R8+LWRwnFaDInZNx6Ea5072ixbRy5gwaH2MF6tCHHlIKvhS80op3RXyWbudvtHeamaCjosRpx3aG
MJu9t6aDK/QspQ+VsqvnLUwVnwWvsBOni1my+tykmV+0JcafQDfqWnrIdrPjAQZ1XaIgFnpaL0d5
NVD3th8ZFGhS7ahPrX9n5KwfvlAv9qodfLOd8zcd81ppZah/NnIZFHyAY6jdQE0Psvv0vBR/U/QV
Mmb+8Um9ubgDilBK4KivTCNJb/FTjCxIkeqVvKrwodbU8952PTSykQ6v/vynd8d61zsF1uPITPhn
HpDyg4GZQjTMKYSCIAs7szd/XXFAKeHkSXNUPs/i4e7hSfXGvsGz6NjgEozwQhLWt4FaYtLbHe7I
91MCBcgbIduqXlK3ZfMT9Up6oUdpwAhfLmqXYg+VEtnKqe1XpqdkBwKzibj7oASKN5jZKecSV3L2
lps8W3/6Crhmj7ZYR02OdKvAyf7PTQNok0gmMMxtR/4LPlfi2OyHM7Ne1TKJQqi/a2qsS+4shVUL
b25JQlFYT/chaYpVpetlxgfjntEgvr1xQwU19KnGJBawtqE0ViCkNIDthkqd8QOnMwvHt49Rt7uP
vD+/HmZvOxWzisDzod7SAfeHn203LzMBUZY03vv8n421kOagabtqoYYcIf63IDHyf8z7HO/lkEtM
lfnwzKOz5UKK79nWfcF3CzHYpO8jIFUddCa9m6zKMnHXSajaHc54TXqmL6vAkQjIHwghxhN/Z45q
B7E52nqja9VjDFexenaSH3HnEyphV1zw7js5k8sLpKYwke0Y/erKlI0SE7yPhcy3ZIHTY4l7ZEsQ
074dGS3r6a/evAWy1p5hXsfCHxzWsLbVlMO8YN7Lk/hgspX/nzO80HMgaENH7U5+sIRjJBDFxYkZ
FqCzDT341LcrGxK5RxJmZbwp4IK2QOGWQWpRQUwfmz9s6zC91hrtjaUAZhGX+vSJEowsC8fpwr3R
Otokux0onehcDMXHnfEq3zfIodX8BSVjkPSuLKXNEODlQaLU5BYBExaY+EnngjmZLTON1l6oScAi
r4oLC558dG3RpMTrIcHa1MM8PZtDlzNUJ4jjePuwaBTJdKxHJVo5G+4rKCA9rRhYgmzAoY5pXtUE
zyCxqR+XZUWFvY2X5MsGAn+gjh6orblZqKfI1TFl8/hq3wwFM4AtfsnjHnpw3832D8zz5BTqsTyj
lGDS7/+Nom+dbX/BPaMGun8krGIZ40Q7hTt5eBq6lj0MBUMuDH6pi+NRTq6e6dGDZba5s2JguaRo
0Q9E6vtDiwTuX2UQprkbyF4Sg2yb9Pjzp/4zuFqz2IWF1wPWWJp0qivmzRdPy1JGeVW7LOVVCq7L
V5vCH+S4nnvUEbfVTlyZR8ja7Y+8swkZLU7TqrEP5B8Am66qLdzHc9X4BuvH8Cjk2bunJAaSCGBG
XjXgu7pg/CUFbUzawLHP6IyrnbghoZWy7zHSLy+oi6Bo2XfKOQrdfw37ItbKJZ3uizkRx+sJs1Qy
Kub08Fl0TyE+avCs1/NNI0PU5jSEezza6P3Bv4mRmzSZ3HeBvD1KXb3WX0/XyZVYnQAx/6WEjpRg
Hrlenbt2cXvLB4Gz1jDsmTd7n6tvckpTPAvJ9skjTYkcKuAtFWBqZtdySP1gU9TNs+7PAr5N4Fcf
Thv9Flxsuiv94GETvbzDvaIxNTZJvqJX2iZQJRojUUNGXoARzIKz3Z0cNW0iA/pBXq5oXPszfWoq
BeNONMneNesTN0/2cNv6hLtA1Co+T7V59IladuFB6FgkyqIIHRbYbF1wnP73l01FDtdayjTim5av
pFhTG1+UVnIzRo8Hvi6060s38BAAGMrkdJ+5JrfsZJN1FDrX7ZZXvE/L2BxKEXgdE/qqFxYat1wQ
+5w2aAl+mhIHycGEkClEaHGyJEUcvNjkExw8FEKjiYZZHCB/qwoBmBw7ZLyxcWBj296ewHIUq2BD
3VhKlXNt8i/S8A2fbjAHLRJVbonBp+aAffZ4UfGJayu/w9vLlSe4QDsN1CF1f13kNnQLwCaZLqRS
o4RZp+B01SkU68JOVjTSiqb7iW3P+FoInyYtqoHOpfiPfWJB8IcPxwzxWdPuWrTvOhdR9Zm4wP3F
9j16DoS/rHrUwn+yGDYVo18N7AFHscsHWK9AA1HVrLJu4GNOUDIUtyK3mxizo3EUMMUQvKxjLlpU
u4X7qYrO2dk0L7O4tKHOpLaW4lvyLSYGtHJoGx7iyNzaX+KvFPlHxF9q9BuWJ+IqP5AuhMlniSmm
++/HeXdlJIbmW02+pQ8Ib1COJzuZasbEF7fgAWa1QYUEQvfm6TE6Sq0ICE0eX87fdr1C3o092iAb
kZHPDxcNKrKG/uZl5itH84rxXEy2TDXiwxgKGeyaxombg39Pj/sf/ZfpeXfdlv544LUOt8Q3dVsL
WV14U95Jh2rB/HowZO3AnkAYTbN3V1yH8CVpGQi/OZV7TS9ICMd80M1UuXtRP9M8ec/TkXeNmPgV
Km49qoYtXrhe2s4x4r4y5c9dxQucU4DcUC3yR5unyGzP1Pj87HOeR2dgUN0GFs5B/QgPQFxq+H83
0nMwOzrkPbKeSO+4YvYWFArXZ/zcVm6rqWlrVOaxLUqEvMMLpiz8P2ywJXDCPB3asqAYuw7+4rMl
0gMsB+53NO3upgpU4DTj/ATdBX0m2DFPRIo5rMHcRl1acxGtH/wWpt5O/N6I46o/jFy2PhGyiSIM
0zUJ3ESeHis7TczKAZFU59cadViVmCmUIyzAtr6q0L+bJHep09YonzFTVoOZ29Cg1L2I4YUVk+Zl
D1RukAiEm1p2qg12Ri1zDaYTR2qTBKfkEm2mXnr9lfiL+7aCajp4n4Hqpyeej8VnMIgNFxJ1Yd4K
2aHzvPhmDtxneqHYeACLZH6fw4CzwINA5gciyAZK5wmYrzUklRIrjcEsT8IGJ9NlZ1nN6rI1LL8u
vh/cf3mq3LCGTCpeElWO3DO2Yd4euWxQbaN87Fl7rB504UhAN1IBJ8KVtm1kB9h8Zqj3DZp5V1RS
rQQST2+Cn16jSvW8tDOR1w5jNKWtl2gUljbL2UaG7p3bUXbIN4OCLDDpygCP9oLI3k5dagKMhEnv
4vBF28ZsDj3O6wOxyd8wP8xSFyJTMLZNhDzDEjXVq1HnHuhyj9OFxRtlBnZRDJ4oi5OJolzgCTsB
+pkQt8wuD/qa3jyOhySqA3NkiO7r+vEuVg2fN4qApaQ/riGmOf7ALgZBdSXweS7UMrK9bReVhdTM
GdQyf1kwZHuzhIDcwuP+/RIDcsWq3FcD618KidOHf4ilzmbWliqJPyg+DLqbwuXNJRC/FvK4WfBx
2Tq1Wf9txtnwtKE/V31uTQQhgYVUHFXJnwBaxLKdO72tiaQ/pPM7q5V/rd0Mh8V790zn4YfdAmPs
uj7b8S+aTp+bai4DkBPJPB4i0skhZEZKumauaIcyq+9lZ5p7Ejbr4DSPbCPVzsWZNUcx2seYpMp7
D2ruOUsT6ou2DA4lKk/YZKGMlgxtdtRLQZvWN8jTD/Di76wXjmqmawUw7jrSBIDaw0vyivH4tubC
MrxarZ5xP6xjtaPtIZ0sdsUIvLqh+IuSgDOq0U50siO6MFMTXe9zGYpDfmbps9dI8P0mR+ppx7IX
cHSn8WGcv2L4rDWmCJAsXXUP9kOsj3m3rBiObEnmDUie7lp9hoCOpXc0Kql2riwq2JUi04lW1IU0
gc0kzmyrvtUQFMfNCZdV/JA7tLmHXRe5gJCA0p6z5kFE2ZbhHirSKbAbLevstoIYTPhWanUDXq4V
5L+w9nKiiwBHUZn7670TYN44VlOdcy9QnkfRBWngTxlPutlys5D4YOmb2wu5UlvYRMALNr7uOhSs
LDU4N3rCGwPXHjTSViAIUgJM9k2gYAQTD3aJ2Culup9jdK3jiuYsyPAtPrMuTBsdnefUVhtdalsu
C4S9MtVdLdPHQG92Q5lKtQlh17jQMf2mJqwVE/DlD4vkTwFT2bxOIlr9KNVcdlTr1Qcs3M95uBP6
TYjl3WTFY2tyInZpbHFa0bOIxhi8lFMHP40sWSThXX7KcdSvNduHgZEm2NISLn0Wen/MHBVAz+ye
bQesyRM3nljGdtoenwBtbPfTp4ZpszobwbuEGoMLtrxtxztOSIhamvR25n9jrhnowuVgKMLsdS3r
EQRCMSGxHf6LVFuAmVwFB0Kr6icDGLZIz/mOyOH497FWrcgkE0HHpfslqgZroLllklbrYuZmqttL
7WyA66BrOiW4FzY475xgmDrRodbNnW0xXF+m0cKp2ZazlJbPg7rNv6Cr45r0veJoNR5gppzydyfR
l7cztX1aqKUApj5tRN+vEXvnPKhHIQgC0Mc822Og7VGmkukuhbZni0tMxXnUdTws3JtrfHV+cOJO
zuKmLOIbmi0xMvUjLpY2RfV0CPFQUucsnNtv8qzbo5fB8/vJkMiznQLnMQXGALDXw8dtiqE81pzI
laVivVaAQzdNrTFGOyo0NDrHg1PUJjYQFidw+J89t1BRyIMskU3AEUMg/SHxrsbrVQlguFhS0i8D
LXwxJf0V7c0UBfupIKWOCmPfG+PSwMmunBtiaS6haowmwFGgv6CkScMYLFM36ZbFAtr5BKJAzlER
E/1X4OXTwVmahtlraDDXRlEls58qVfV0mUjjG1k1upVmsfJ7njyAPmOP3vIo6l+7pPGMNkBMxPOd
vl/kI03l183Ndu8n1Bz1uGhdbRu9p1NquYUbkGnOeTyLetzvj4Dv4wx44upR1zlEZbxpRQeRN/ZQ
BJd3u5dVDfv3SSz0QMKgiNdc7eMX7i6nfv5PncRHpfYVvyGSvspOeFAFr+ohD6RSj1fHBrPmSpbN
IK4L4o3Dfot0gcgunUJ4GqH1ah/t8UI0PWxLj1LTe9Z7Gz9wk4LGMXN7iLm5gYUIvn8s6OAHqgUh
sOZGmLFC4qzwjejVzWmLJLrRDmMYqAE3GOqFaY7LYQPeMXFJg3jeSIt+eekc25oNewhe+j4HhmTy
pLLsiM7bGR9w64clcT4udO5qd7JrA0Y5zhWEABQuO9JRDSMEe0sqgsp1cETk/bOd59B2MV36lOWS
f3kkvqtp8gud9uLna2VDmH8+szNSCTntKo8UyYYme3DDeNfonOzeDVgjf6CTgurLO9vJjsO+imlY
NRG5cRDimALlh4sxKHwPdiqhpaGnm1n8lLX4mVyEwfReco1BNXPcHUOYXAX8XAgeTOtZU8qb7JVp
kDgWkpF3UY/mRQJsy9+Y5lWqgb9EUPXMcKtSc4yD8odqpRCbDoQoUFflNGvGEhTo/bIa+thE+ib1
jYIYhWvLyuYGUsqJAJaGKeUpMgfXQl8S8DaXfMT2SsAVAOSrxqn1su2XAgeQIjczHztb4OltfOO8
yVwc3mEuSCViwT2kVhaMyJ0tG61Nm2zxHlgdCykDcwIHRT7xhcAtedrSOAAeA1S73ddNzJdRhegE
7UIri7HbKqZlUHHhifSFI2VQmXj6z3O9888kHyoxaBHtEz+pr1aV+FyVx3ehdJyFzJ3BNk70hbc8
pwBQrdSNAOMOOCDX7XQNzMVG50+KIppzgaq0UX2KPU3jAJ7v/ro4HSL4wRXy8kyJ1AY4t+UD/+QP
pBeAK1dQhRz8wVocdTVvkToCAv5LpUKwTLzKpXFWesNz3hcPn7rVgU7Kmn13uUEWeOg8WXUAoihe
cgyhx4oeA1qF1RTktqj4l2zY6qBJ1TCZ2pNcuPpaPd04VaLlFf59gSP6U6OXizYzIVGtJTd3AMI/
6ChE1c6+ehnZ1P7M2j7rjiTw82Vv3t9GF+pvuG+eixtKb56YVtTqV2zWu+gjL664xeKIpN8hey2c
xbbTvyT/deSYkQ7g0pAl423Uo3MOR7WW+4sZpFDJRiXTv7hj2J7ZSnkZxmkUVNYbO9pD94R4b2K4
n8zSGgZpwhVVnOss6+62FVwU0K7AZKupk6AhqJPvg0o61EbAFFy4fj3tBXXqmUP0LB6Q9CoIuc3n
mh0eLuNlyC8xj5YVMUXK7Ztv6zrM/aR0XsMWCRLEWntUiA7XNHvs0ZAxzAO+vC0oMGeR6s7o7C1D
MgZ6S0LwSL6nTk4LNUlkyJj8qBVUHcN17SHjlNRY89Bywtitk52ozBo4wgc6VNpMRB7eWRXB9IqO
jX5ZrJsvbTu0sYyPCbErQTdD2TkrT/mnNT+oQxwNl8FN4TvZlfjDpgUaaAWrr5uKqw6xp/gJgmCz
Ykk6Zr2X7fy3FDyAxW0tiYO9bBk+9hXFu7d0L1vjnBGfKY5o4U34JO3O3THh857qqwyWWxO0mhzZ
JbZ97yD0ZZZZsOMTA3eyK6j81otg97ZAGsrrQQnyBxIbeBfaBEIAkYyg501NX6+2Ic6jPbmUAhLn
UuzalU1zJarZ/Qq75Al90PT+cgND9veS7jJ+TnwPE7Zd5tS4+q4UH4dpfKB48nW6weNPZTTUiFUu
RhB7xPq2s8ak435j9Ozklp2N7SqjNnkV/gOCeX2DxUa+XcL7R+rPJbBgixrc/QMTLl8ixutL2ixZ
zGiXb+U8lS7o23mcJt7o+3SKh01TBkaVLNgTlPF9+LoYIzMiPecLkniOx6YrzO27JwGATi2ILwx+
uQZ80+sXb43Q6WC8AHpAS9hAMDlGIocMy14oVb0j0SyXh3o7cvBaeGn2P5Uj8f4Yk3g+MOG/UcaO
cHE0ZGweliZCwBhWHLMm7yxCN0ILZrT2BZRnVJbml/xHilWSXwRJVkkmhnbbLw+bOJPw7v3eCYQm
Jcw1FeeP6zHBF3xWiewbcVgqCQXCjOvPP9usIziB72+jN1wcDxSLEaYrsOvdi4z+J4Cd1z1L07An
2BV6PDCmo7TfZg8MQbRLipKePjda4NwaafnIrd0TmzY8nftw/MkKgZ/+r4Ow/hr1LP4kgc0tCAr9
g07bFVxoq/wZHe6wvTCe0s8kUUkoUn9q2Fhf2rFWQoR3zzfeqzZfxIW7xSDDeMpz4rmFosmE5uhe
DhNe5Au6R1GqfO0pL5U4rATVN4lNeiAHkzkX1l/UkwBuXkM6lswYIyUFinoQh7XAImt4GkJSkFI1
ErRQQiI8kP7mX03PFc1T1Skane55EAkI7JW8ScP7Z/LPC+UybO0TNtkzjwLjOalY7p5KDgTQP/di
Vp5p4IdMF1yObZZM4g/UW5VF+dlqKtxiolZftw7LR0Ixavjh70nQQDMyZX4buHgBrB15+QOuICGZ
Xc9b71B6Av2QBO6r4DB15INTwOVNcWjg8uyCIRuJCREVU3nleN8fUtk5T8JD61m2bOqyaRfmUAmQ
bLqx8fRf6f0ECehmwNZCjAKvXyY2kxVNbhdsYutVMp52N67FFJq8Cb2tHUaxKQr6Lm9ZrCQHYtbq
kyju9hsk4JDRR3nW+jBWPzHe8niHX5XXXtKajWl5sgAyQKl8XsQ/ODKUDkk1rLyyqscV9SVMYp70
7DHflCHla0uRhUK00GCTWik2Qu/Ub4L6mZBTjwhMHj9eY+cxBKVA+YqLOqhEM+jNun9xQHeJPDdS
PlMx5QyTwItEScFLn/Addlpv0G6l6tOVaffeeEGaBe1hyVXhcSMM1zU2b4re1euYNpHKbJuHK30Q
J4rmSCSuG2EEbxcSYCqCPO3t7X+wfUc2ScSKvMkNNJscLdmqEqJNJKvAO9ydEE+3unnO1FtnH689
8+Av+Dd9Tx3ZH9icHksv2VAV4k2Y7PRIoHIqVA16BFZ3eaayIVllTslE4KSpWvkNjFYBXKBAm+8Z
J3tYUvMmP4SjLQLuocT6bi6uEU5xIjDJKe3H+rUUDJ4sC7qsXubE89navu/4npKggyxlegbut88z
jBl2u/wDNtBz8T+SuxvO34Vv4QgMeWtbpzh/wOmZrFYubeyZH80BALb30aNCW7RyIk6/DZk0E1RV
bg+2ETMtCmdy/vNAAZ5v50OVlxAVcLKPuiCc3F8V5sw4w7h81U0qw7TCV5gn2uPuphKyMtcqCqHy
UB7at8Azh2aauq2nla/s1FUNNOhlqtiv7FFJl5I/bXVMhtTgO0HlmOlN8DZYl2eJTsSLP/NN99Q4
j9fA5lFJDz2gIi6pWpdMN8H6+tZ+0xM5K4O82Q36HRWp2+0XzubBWsD6Un0gGrrjEv7mIVXTYZMh
Ii745hu//bPq2W7gVwZSx7vOejuIaXmKnZyfXkPXfikghyG45PCAXDVK81/Qi4x/zGD861Q6cPws
syLmBr1kFXHts6xa1JRfFVN8O3v03YZJXWFlcPlPAohRxBiYCCS0bfaFewhtlMGzhO5AA8kaoSVc
DKlTjSAnBTcm8FOtcuC8c9Wv5bQq8LWLLuAS5+BWBO+qlSuh+J1MWhoGao8oJSaM0yg4IFhByYhM
qehFClw0z45TaqdIASr1qOnGu0Di5n2OrnJm3gqpUBwb6j6CfKEiHmhx3bJ6rCX3MTR3TLrAgu+p
3fUFhol2kSZ2GZ+NFYjcXHfCuN5Jr73y7Ox/L0Qz1eXuJUOGUCqw4qZdzaXgeHlW7GQ38N6stLmN
Qvyg1LRCjO33OXZF6vsbYLaXC4rKH8NL3F9NuR60duF0Uacc7Kbjf67KrCyb0m+xcdKOBk9u5EJL
GZJNMtXd3dW5AO8pjLx8HJHQ/QTAdb4/hKlQ/O9CuVXM8OhUaUT0CNRNY8F2uS+yz+0+fZM/hvOL
ACl3bMQy5Dc5P6MRl4gNNe8vV2SZznW1lny+gaBVAPooubvyBDLH/AwEd/SCF4SzUldS+2wyo5z0
9V4fWnQZHWzCfHe/jLDoNoqxh3pvCgJk9WlwjWBN7XOn48OQctMF+yVaxW5BL0hbFy17mPX3BTpA
EhFue28o4CpoxPTXB6RNUiF30vMUTZ8AaPFuvduYDgl8LPwnpy35BH/rhNtf77wFEc/32PLcxtJF
+FrPJpWeUDaDuPYT4D59NihChGCc8gO/M6Mj/buiPm/wRjzY6y2q+lEhUdfcclRI9anfBxOUEesF
Hqzjixhy/EY8zJB7JwBmomu99KDILNmgDemk4AlJv9gJIgHxs2b86SP0vCUuAhllUMDIhWjQtORM
dYbqCU+Jj9NfIASXC2iP7zbC+6qEuQz1z4C3GTnusnGlRb40nnmzLhI1BW9Db0Kv3RzKDGH4LLjh
boA8s9FDWlg7Hn6KAq/nBl/RuXlZ1aLytsLHuxsqVy7x1vYjFpGN784bjxOdHhPzsRvBsVjRcIPu
XkSBQ3iSue9XqUf3rpQ3lmDGZtu1ockWi5/iMw409XFj40D2ZqmV+zouWnbMo6qbWDnjgzyU8ald
kWAK8UjcJzFvOx397AAU82Ohl/arcO0Dxv0/t3PKsVeZew+HUQlwzKK08pQfpI4PTFIPGP0SajJH
KCRNCvL4No/6W8u8APBtH5WpBz1iBsev6sP/VWp6HD06B8ZsHNKfo/WqOcnmMby5ZIuNE5pRABXL
ZD2XJPdPwA4DM3yq69iq8BDJF/Byflx9z35d11KaY3j07VPQPUme4PnFGgitgi76wKODiZbU4Pke
w6RehHDeNbmzwrRRR5c9JwVF3ZJ+U/4hueQJZSPXI+qsHe7gpiKisKdxCcFbyWBW43y9GSAM1HjZ
V3aoWyGjIiznM9aoss6FnduwnhJF7lDn/RRzu32Uwb8ShVmu4saM6ml6DPpu+DSTMycZs5QyIjhO
FLU95YsONbFeG+Cv28THeYw4nsYYjiNWAVmXHRsmy1aoalnKuZLXuGCh4OW3S61LIo1v9lRKw24R
Lt8esv9J+ALwegyhki58o/HiqXymO6Lund8HfilutU51OS3zOrWgNehRoRFCpsqT2aT1kd3HnHZr
iyqpeqsrY3vcZwJ6LAl3ZrO1Vdd0W1V6xC7qEoOjadfRrI5XR8MPc/u++hdWQ4lHb3jvd3sg7AGI
18Yf5+70voOw3bls/Dx5G9kH3z+YrMUHO23B7TOxxsHE800v5MtRSwCiz5wG6yNYTPIHlDwtngCv
BBPhVARYCC/iOZ13Bry93NhG7WqujP193wT3z/dajfWvpTxWpVfLtL1QGQnRCy1Qb/EnErJ9rkCj
2DHibFO927/2qvyiVYmeulgW+rMAlf41FtrAxeJzyj7MZ/6bo7IlCpipgtwBuVxpWXTH+N4EhBOK
Fks6V83PlEN1ch8lpIIZF/BWlds335rFSHFSiAeAGkawFkcKon8+P0e64OJrpndCpBrxXxO/CZMp
5AGK9O7PketGxOWBfk6sBZmrhphe6j+/BFExR9/USMxTa5MSYDlPdY5qb20GHtGp22MFyERbLC3h
VbByDMKnFJ9+059oYMuKD9ormFXNQc8HXiOMBhndzIscxTwlPbRjY1XhkbaGE56ICd/jRpKpfDe9
NqNs9PhfmK1QM9CL10qVf6PMMHheAIBUKjg+fV6kAFPwlguL1+cmCH5zS9HKS6UtajaBizb6RiHM
TelkhLUbQrEiaE1KJ/ViN3NAItKowfiGPSlBrNNDvz+7b024TyOsbr+06YZpMy4zZ8yNdv2BiRrA
cZNEyBMKt3mhMcYcCERXeRfOpLYkKADXNtmd7564wGPEsVpbXvJBVuuZAf8lT34iBShPNAGjUq3o
8+gMlbVeBrlv/wRT/JDOJQMqmUZE51w3PtwPtwWUOhg5kWhe6dAU95fZssud+/HJdMvgiTIWwVLL
+kRqrL+26nUFKkHZTxodcGTcc1JArh2FRdu4I2dzdPBDUeNIBGa5NRypAt1GrTu3mFmq6W2vDIep
RZip6QLp9XjOlY66ff1+FrgdaID4QiSS+HHMU/ZirQZrWBTDD7QKhjdkOHalh36t5OrtDu0oUDUx
g3BDVAOM2g10LQAlUeYkz3iHPq9zcRA/Au5/GcaAzsjoXgMN8uO8UNDQ8kg9TE+ATveMRxqxnhOc
LrtR+DDeM9X5gUJ1FtZTF/v83sLeatRPrDucYlSzmMwm8PQTgKY4yETB7fccs+KcsROl8ToVKklr
7CgcjT3VGIc02hJsORvenczxPTtvsRzUBnwI7z0UgNqRQlNwunat6CUkX8TCY/xmGdPMedH6AVzr
mMTvIhWnfM1svoiDix9NzR34Luk1gDiRW4uOsVC77wzA4tF4O5Q/jS0IharPO8wwq+zoaSjJlgOo
YchorBDXZsvBy7xvpk4bk4aa9rYZ/duOgvIgvOZuFgKazU/5f8Xd87QaUMeviy9K+X98nMHVpsgG
Uje7LFnNONJ7SY818zabkZ+x6SeqDudLpv8u/sFQa6fQVH8BLGh9SnSOvSFR7IhVS++u6VSfarjK
O0xeq93WVeDtyrYYIxRatD6I8yMpBB6Qjj+OlTtZACJmPf0mjbaNp7/8L0y44HiK4ynMdA9s/F/1
snsZUL2T338LYHi42MzrjG1P5N6in7by7pEDvuxcVivvK8U7Kr4ei+VlPm+H59phmVJ3mzDerORw
530SWs0ZjHzAdoPZNuUX6bkrtPOxPJgiEXVO2UjBmvaR/oFeOimBWsLxaZx0YZTgQqi7doxRsrq1
yEn/3ch4u9yFfOn/P4ajHthC3xR13JMhFc4f+Ewi0zGUFwNrGNTZc8OSYbU4rZyD5z9n81/8Sl1c
9sLP43vkus+dTM5HCLRmqpdQUXKlluWCJE7jon+ERmqWBVtpHcOq366SFD/ScLYdruwVz+3NYG6/
wkMaEXxFTjOL3jzK8CtUZvvFs1DlV69b93T1m82LmLSoN9Ygnx9GNTIY6lksig1/HQHuNgmGVlI7
MjC4B5ltRY2csuO01yvtCvHnk1TBRfT2Jn8LcTXjty7tzw0SCxfS2AD3ogvQ/3Clz0X94rpYFyj0
3+V4Njg1XYmG9gEsgO84ikOxBPbix59LkzIV2dmmYVX/9UXAzGlAv3qN3qq6EVUXee1GSJ4bR3Xn
H2AT+7N11mOc5/1PrBTbM6stenPVYd7cCl8tPJ8w7lwkIXDNo9qt7/xd+vgvL1IDGhllk4IOu7Nh
MXz5BmG892ev8+YZo/JAt2n0Awzk82f2PO3Gk/ivE3Kf2IYY7rdA5rzhNXLz4DDxs1nsUkrdtEGC
ExVHNEXP83aDabl5DNNRpWhSkfM1wowyhH/fPbIJf4LW9NdPN9ht18ftX3M7cLL6KMSKmE1wi2BE
uN+n5M2WYd9N5ZnyZ5Jy9nluhOgKX+EKjDg/0pK1wda1WlClnBfye46PGomLnqJSUsnJa8jINZZ9
yn49deyPEHVg3QzVc7YDjUZqT0kFUU72V8rRdE4Gpi1kE0RXvuuCsFQsfdFcJTxkInaZUfF8dxRI
WMaKFfewAqZN7emVl/39ixmn/roxAGJovCOscemqUltO22qTDIiVPxfvXDBaE1hdS6mKGUlgzvey
kQcjKi+tjdVA5xJ6gffyRhc7rEjNOb/Tnwr5vqcFOwkjLSHS6/ZxMo8U+zqCKw+QxSrCgN7ziyw8
ItIXatgFdJXNDgVnHIkqOApoitfbaZAuNagvf/tRxS6h4i0Aji3rD7Y7FsdeExhyv8MCUrXAsmHc
lUUk36T4dZJaw4QhxOkCl6rdBi5Xc1hATm1TyjiRxdlrf5TTVbv1qKrVe+RIucbt6xeRsTWZrlKv
anN3CS4/RgNOQDG2rSOGZvN55Em3wvEzlRtk+UjMvljiG1jMEw2RekCf/numWX0Xx8oYGc/W8MHQ
8kC+TRgIzewpd7ga41W3Kz9K7kVK5+QArEREgY6GXCkY/ShE7pkjOvMgkvGs8Qk1UWpeJ1sMiZUW
8p1msWM34eZXC9sgrsorlUVeTVIqwfqbE/y+ufKLaKrUXd8W1pRH/T+VLpl9Syk4CqZIjkhT72c0
Ml74Mc+GOzQ960W4TwABLyvDCXh2pjOnT8Na8xfa/nD8VAF8QGTMBkXDMcw5UlOMNG2HEReyx1m8
6uZhOoJhXWTtgSduKcaHo5uGNtP5KRd+Bm/3Huaw/vGkG9whByCnrg7Htgrc77SZLjA5x8XMiatO
ASeG8Lv0m16Sz+NgqmP7blTBPyFyHcPhYA9b4mzDPZqvPKTXoaQymtDfmSW7cuXPgOFICJNEbAaf
0wplXy8aPJe0jFfF816TbTAps1NrdqjPO1A7gmJi0VOqksA6+uWAz0m0aUHC2akYcxPFuqnd9uug
oXswyzJb9t8K9yMpbZvJY/DsMT5FulFNRdSnJnMJ2zvVqfVUKcD4p8Ocu/1uA8kr5D7XNfImbvzM
ZL2QtJdGoh11G/HNTgAHehpinlZxotXOW3uAi50BEK//wXOePZPKlU+r0oWHebgmk3x2yFd3eioG
pxNJUNyLzM8rgMWMzzsON8wWI1xDpICZAEf9/Gdbe0V0q8W+++vKZobH28v/IubZ+PCXh5b6Q69a
xnQ8VDRj/Iz4Rj5fhqBCCIH9J8ckNNIjcWuoztfFgKTFbB4TKJhbnCmxv9whOSduwcnw1KxzHZtl
rQ8v0Me1yLnnluKb6Z+hYUd9Sk6GaEQxJkFCIfto+pNjtPHJkNsjPyNOlnyruW6osJ7T9tiWFkRo
kvnCp1TJSG/ZMrgDXmEcaEa48GX48y7YkoEoJ2h+EZUal2H6z4m6xV048YCVgTEqhG4skdKOf+mY
aYi40vgSlvS17C8Kl4A4T3agazJz0aaxjG057K/sYoeP2Z65jr2EaU0k5mmh1p6lixxmBWcKqGfF
LxY5l7PemuRVh/LMAdLGx0ca1yrjOOnXLpwIel6L32gxurMLIUmtfqVffb2MCCWmtjIiQas8DlO3
0DTi/XzMfg/DktIJ8AWbRJo/UHuNQWvMBUnWNj5RAMsrMoPTz2oS3KVbhNTQqR8X8FSHtGA1+/G8
tgianw2GVJ9WSUwVZyfnyOvBn0GwfhptHqi9yYgft27wgy25pisOe91ciPEGdJyr+L3QjoZmAkvJ
SlQ/HzNG6AyEnsDxlroqYQtEm5OXk4IeQZ84QBNyc80hbnyEMQW6hm6iHclGef07Hn4/hb16zPOk
HzvWa2HvOlIzk45eOO2zotM3D/S7RrKnV67bVgtJzIn2a4LPEO9HLjNLcdr2MpT/8oGFgClyt3lA
u76KpMwl3JcS3gob5M93Rd6roW6qiA3RbvWifnmqeZ0l6bE47+xvxRUQSSL/GPHdmJC1wELZ2xOz
j0oHh8zqvRGFyEsB84OsMJYrkvFJjQMe6XIUGGKwNVGS8Fhzmnegqw5X1mHz5RLSgY7wosr8/tsi
lqWhAUqR4nGOAv4jVla0ZRmq93lSD9PA7jnDHsLIuUbIoSlXyvF8PIGGRtdm/xfes0gvYrTQBdVU
viIUOs0jA2W9/oUVoGl1C+U3RgrDVchQ14rbud+yaGxbbIdzWHdGQHaG4ZJpJlQ0U5dvfq7qT0XU
PpXAwgGUNlMi1IdWTk+5HcvURCXDYppStvyom9nCnJ7+ZGqBOiIG3C90iQnM7ARr0NUvyvKdHIbC
6G1Q9qdDLZ+de0cnx3sbYvhzgdFq2BjALz7coSW4oQxUIC9KmTuPLazbzZbibR0Axc7IKoQqoFq/
o/ycOnhiOJtaa7lkyVfB3SSOcX77FpJ2pTAKKwaj1MTiV3sbHhatrSrZHH9JdN70R745VAblpsf3
7sK+47zCujQ3xlXGnLI3JoqlydO3fHsC/S0pDwiOG8ibMwNXR2DSScModp4S4bgbsP6pizoBSUvP
V2whD5uNjgKDUUT47i5TigmSrLLT+7Hykc/VaOXtNgNPoUe8XgPE0n2vrqk4lc7uB1y+2MUgZLVN
8BEIlz35ubxxj1vlU9HqZLyG312wlLlcdAEq96XhkpZWRJPdrGLQ/FTmZXuqazx8branIh2v8vHZ
nwSAvy1OhxZQ1+HoBDJnTZcXaRyn6rSfErd1m1VBVexSOmgQ4LnrT87ZRF8vuRZarIioV9wG9JEP
SCZCdL0FwELMpna1hzLcoB4WGufvJlRRRPjgQi/muwC9rTW1Ja3Z6PpVLHgctEY0pz1ptlAbzUuW
zeIaTbPk1glM/J0PtVs3ogQA4rvrPlky5kY+aZ8S37RjTqwcqpkLJyBZt0wysdpkJ7MtXWBLKfoA
fP5/mjX5isFBFXuafFyJDVS1N6mTAhUer+39XPCCjAWKNUIl346xbS2qLWJG9snYClo/rYkIn8aa
Q6rfil51L+Te63LoadZca54S6Nzz+wFZuHRL684d9cfFdZBtJLcrcsx/GvT2P1zlTOY6IFM3tG6w
Lk0O9BqI7eaTcyH5aX2EegGAOTXJQsXzdG1VipWBNq5egnEXwqjzfkz3zLC7nC+Q/0Fne5D1jrAU
XHUOxvkh1/+i0i7x6NAolTSpDsJ2QzLFBO2+usokcEu9QrFGANxa0mJLyNMZmTQRVIImGG7rvbh5
OH5nUbcCuY2tjBYbv/qX4po8Gvs88NHGSMvUYyzbzFxlVhKrIGQJt6O/g+/gfJcYMq23OEWmqQB+
gfHfFBPR0VmJXS+0OVhvBrhDguJblki2RP58Z/QI4AUS76fMa0BC7euTQhUusUqnC2IDrAnKU7dM
TpzjfJ49zyDzSrwt1q6V4tdY1e7at76Xwyad0UdpWehMl6MN4dk+5GXy5I9pUbqiI/i1y0kOyWot
YNUMqkAC65k0YK3exmdksLVIsLUstpgEa48joNB6neVIIIjtXTRR2M5+4Q4QF2nHgphHXqkyFeZP
1dE8glaPSzG7cHlC3mMv/4yrw+dQHcpNWg0tNH/pIf0HdV4HgWblB4oRqy13hS15rE/udg2fVbaw
L1hKaDmu3XDh37IzyUlXPBE1qIqPB+Oe9Bnrol8zwhQkG+hRdUI+JcKk8vYJqWCMvAMd/Z0wYvYf
QkiTw5x/UnyTOoSEIviS/s/vrRWS7v54tWDS0dmLQmqLKENoC4lahLDSsvrlYhbefMRp7tYOYEAK
HMVj+mQiBDEAfGuZXUODDyq+RO4gIEEYD9ZuF4iRlU6cYrnJX1g876MaIrYRMsltIkUBG8xOXwy7
tYzd4GQ1zJ4Ly62CN3AWZeSwB03YJI5P43aGtalATq/NevVPhbePV/za8Gg4yUKIfsosjkDmAyx1
nI+l8s9G84eCqhEBBtiPv0DTdJPbOXIkkWwnqR5Z7QAljvSV9m5KyJB0BfeZ71rZx7v/Al1eBFUA
O3oqtQX/yjQIDiQtYxsj/wie2eNFvtfV3gj7f5NZ3C1qAmLUnWLFEHCHgCYPahQ63p9vVl1T7bfm
D6L4p9ovvfl1Nse+3OkmAA+Ag0x0pvct6I+S1WTd4x6TT0cD6lt2rLiYt4fotQjTplrbVU8gPnZJ
LRH10jD+F3megRvkMQew+BATJ1N/QX6Zd+9PSVX/fPOPFMdzZH5ADsDQjYAtpxUyjznznAykAd9E
+URIaSglws0bSm1Ny/pmCKj8LHnDERHhT7nWA3vn8Ex9Ub3YasDnTiaU9MFmxzhqEM+6G0jIGRIy
HjF6QSyBY/1m/bH+z+hrqUqVIOBwRzugZ/lPShxBJg93lD262pSC3w5tuUnR9kFanuld1LSVX7m0
JgHhZKqqmL4HbbFg+2p+YCsiCesp8tIZijDQOclAIxO2sqxgY+FcrwQvX8oYH0tdCBHllkq0I9SO
aO3ol8Nj1RG9LBHKVfBwAV7Vemb5U1H8HtGcxeBA8D+YaSfZvrTZm/7Vg4/hbTR9jTV61b7Gsmne
ST8dBotP3FaFE9Lyn+Qc60hpP/OD4riAY8RDqIqXIzQU2/espGmPdGuWmumbBb7IYp2HANO/l67P
ppwg/ZsBcmi5CbZ3MLD9OhpknsyoZZTsty+eLuiRAVOh08D0OFG/5uB3/BOnN8DiratWx4Vdp/9Y
Q8Q4phWwLSmFrQ/l8WY14OPH8PwAYQ8nLCOrJj/kaL+bQlPDKN48ilKPoB7nGDW2UEeXaHPdTBn7
bGAFPBhMXV/9uorbogMZkwsMhLB1cCqW3gxx4bMkqn0uTAgK3JwIhuCSDSkryb3rzXClxPRhFhvV
ie/uAfserCDjHeadOB4Deg10P4VT3c8sIT3q2OsDtSYgNJoH3ljo8lBSYq0DBDk3Oi+ric9votFZ
T8aMTsPNMnsAfK+1Kft3qtFuhFGwmpEmnkYnf0EQ2Ib91hytYxy4ylNLQp5K4o9S75jN//zYuxwn
PWpaWnbk/PnmBV8iGoUPLhn63tEMDYybejER1QUGOHT/hb+dJuNj0EqDdoA7jaJjl5nOVGk51Adc
rYtBl5jWucTHhFLqIi90FjLgb2xPSNJ6lKbYVkBwdHe4gehHx/n4KBhH9AD2rLaZPHA31WQil2GX
oNkrynBYOU1JXDI+kanKq8Up2qHIIBlQesIoj+NFJR2KmCriz7ELdnR+8sEx1zamrIbBmjt+fRJE
RvbG0tEJwyONw9PXDTGbJzD+LFHwy+ui8J3WC+39JCRUIXkjPamgKvYCcr4n5HEaCMF4Ly23OjZB
oHPxlfktNvYxRC8mQYoUAn6u16/2Z3UnC++NBegMLGFbHq62qc/0aez8itTz/TOJ657l/iWm4sFP
yuZ5NVB+FnOs+pdSOJum81QEpPl+lnwcN6wk9VdOiZkbtWVmfRAR9eRnRF95E5dxKNy+Nv/Q/WNn
RvC+9CASO61s++fqBRCXPMWcNQvcfp3aZXkCSDIUbSEHLvpfN8ISnc+K4Y6bId9qS0wen5Pn8wsM
gnoSRzN409EUOCgb+a3lhtYbsykGja/lpzAnJjfqKM9P0rgy+Xctx1tFx7CEpIx8Lo3y77WthS14
gJZp5WgqfLJlltMZJWcGEl/YKVeKKZgT/RnPH7LACkQOZW7zMmdaTPXYIquWos2Mhaj+JRgFNrJw
rT8bSI7pOUmXYLrGW+byeb13Qqgj6+FWO9m+JIkmOJqYsE8j7vu5d/u1CEEGDYGFIaeq2llN7i6g
BPqYjhpjfZnokleFHqb1W603TnDHVi5qPCxo7tZowQw0zh9C/QhwDLxyyuv38HLnO+27hvk0Om9b
evhaMBCNMTf2icoPqrhjnzRelJGOleh9uQ/oj0fyGhj9YH798YMRPSo5ZkLJ6z+clA9ei8t8Z2dH
XXerlQfllP54WJ5YRhJLC4eep7T6g9EtH0mEsOwBn4Bdy6eTE5dRM8voblOKgs04wqW5DSJ7Cspn
AhA4xiop9R4mYJq73ub3vh7Goi0SnOcCfJFQUqGARkll4ReGxRFjrGy+oa1DelCJZjpgd4w8fYrt
rHVp9M6OaGBYrCO2qBU7O7JTHAR2Qynzuh651z1XgiePr1dcgx0F8ylrLeIygw24cc4I/Yl8BQ4b
xH0bMQmwVfpB3UCBDXBj6lo47vmk+Gg5/sSoIEtZafODkFKjNC2WcQHAWZqmfbLzm3dw3eaNufwO
RcG6H4qVGrrzsQf7xtz9z4jZhjnlBsTc4GY3vzK+6GlvzhWrRMSl5KBL/sjtzbnSCl75or/QyExw
qslTrJRMx7WaCnJAHkhAk9Zik136lp4vS+C2i5lOxHuTx15+zScIBY4L1N2fymgE7bboZZdzXdzY
P8JcDsJgEsFTAqIOcG5QvROF6NpYKioSVKqixm9g6rN+FfFSgfcvkNRAshUiVRVZF70fBPjitOfC
HfL9GudRbxm+J16pWFY+j1eINVWlL1KL+XNh+SNxoaoY2/S9sl2laNNtPXTO4RS1TA/4JzIii8P9
v0q+LAKY2GqVqYPCnduLTugI83uM5uU+0RVf8wXLATA+sxLgXlqiIKmr5KesXQ9/ciGJhDzWD2ql
QDWUyZKgYaK7ts8FSszjrSoVDnVGdmtMQFeDHK9wbajC5riU7dBMV9X+5N77yNbJW6E6MVlhXMVW
hCUVKhh5I7TdwQ/Z8hTx+oRV72sirDaksZd6UXrAdKP9+RluNfFsBLdGyPzJwRoGm82ccEwbwuX1
H3wKGar6czWdfwTWbpExWZCXWxozMtqAwmmEIMkwesrSsfoEZCfOKnFmFe7xOACiv5EJOwD8LiqD
DBOuuSllHN3/E0G058M1bxHTUhurtzmF/SySolhXrOWMsOS/6Q7TByq24q90C5eWwRf+aPjmj9WC
rAxUiiIhhm6lNYk6MkBGXnoGIydTXcQ2aVXbpWSpnfgOYiJyAa46To6b7s+DqFYXSbfnAg27NvyW
i/KuEEtiCW1TRAtQcVfODyYOmOiU70OW6S38kSz5hp4m5iMvb6KAKAzZ+9s33I/JR6HLqKC7uhbi
RcJ5NuuS3tIXeeuhbEtt4fgJ6qKxYwSOLw20PR95DTTt3E25EqpWwV0fgK19he5HVBR2qq9ES/dO
PEQbTm+fqrcAndsjEyKVT+/ZiBL8P8nsjYv/RD2zki/SN9u5C1m2cF1izPT3cXwt+eityMSUBnLp
tNpEbFxvllpwbKvZmm/QXLqH643j/F/HIspDaX3xTuUuaCvNSFBkmpF9I/enCITWvljWWNwAF2g2
pOTwMymtlXeKUZUXrC2EvUbBlEzysAf0f6QEYBru+K8MSuUXrvz76Og4U2SrXFx0O/xq37a3Su8u
gzNulEWEce3PS24F0O0pmr5zvxUL3iiqS86uXxpIMtW7C4aRBkEIN9EhmFIGPuke3jl/XoGkoMGw
vWkwhTE9inB1CBsB9JCYxuKEf2NTdxDX3ovdcd/8LDQnB+8VGEwMsqkAHg8SK8W8oIjy5bSN8FEY
LrY3y5wKqSeHxfjyuYOh6EOa74fbWY+7T7GbVAZaqvXT+KfuAwN2NVT52NEuOC035NcINBTGuII1
M+yXB+l9x5BLoielVZsFomT4+cFJboPhAxZbES4Ch1IUb3J8KOx4ZCw5IgPwPShHwkf2xsqP6u64
1xAodLSwGIXcxiCgGgQumNr9V62/jTganO1Mac3fpCXdOSoZaIy7PCwDK8+n7m708tp0whO5ZB6Q
sPKqeh59sm/4NFSFqEiUwzD6osNmsk9xwJpwxB6uKKxv+JXPbHD75/1qMLeE14oqrYh3QoWmzxej
8xZOOnWRfWBw/0VvgaRC3k7M3wx9eNCK09rnCoWZmg4QsOJsimENxIu+TGw1TB6J97MJWu+91iRf
QIkZaRC/dWzsUIP1zViRxheuBQnlOgWo+HZ7TpkggBK7Pf8B1IRPehutXHNwjJry5YxTNDbFwKmo
b0qPQY3iMy++INZbewCZ5pB8xi1HReOCgTrgtFSY1/mBT7xZdNTHqfyqb+GEMwp/WzT/XL4qwtiw
nueL1997xvc1gwfSTm9+z1pmWntnDprQC4ug5JBKe/plx1H8KdD7IbA9ZyXR6H6YsPH6/OW4X8cQ
Sw5XvxLoL6xyD9r4YQyaE20EmQZIqBwjNYB20nkyTGVcovpQISmuHOiSx1UFRHHhGsz547ZfQfRm
QQ7Yz/3Z1Nnn4xib/oJuA47CBozkhFZNe8PkbN9a3ilnVMMaWYJHlpe1fACZFpAuk/6S/tfE4Usy
HJZRfZTmrazaWBunsV45/LuSj+S6qIi8I2F4Sni6kQ4k6eo7pmcuFRQP65YHYS+xsMIjDF0yTX4V
IufGWJM3lMVQkd6AC3vbA/Rpbd9I5+LjjSaaovm+DTNWTskdrjOG/Wvg3ap9e4niCraQaIYhJNKg
FoYehXMij0M7j1j32TSPeqTgoQ1Dv7YE4b30ipm47KjhA/5BpWxXEvKifRuLel0zknLuzpVkLRGX
reh6HEAXDklp5mJAHKNKRxcBej+FR7d027nJORUiFRYlmIEEaI72zWSAW7QvMos0TaWIl3wpADHH
2nrY50kquYmgGf+aES7CJjhdCJNwkD2pYPfSPF6Yqvd6LZGpBvqcQ0/Xn6yU4qaSdTM1KWOIiAL0
YQwvtSBZmpRNr9A+Vh+IlO+MW+/MVYiOGczxHQ4YOmOe/jnTaU9yexUOboPP6GIfcD7gscygSL1W
5m76MrtEuhfS5ev4hcc8R+pwzyAHjTa29dKnTVkw8p7jDPUnz96+BuQNHIFhGbwkQtgDomHlO/Bl
kATlFvEUnZhs0RMV8N3Nm5yR+v9XV6n1UGPALqmRdjcMvbNk9m/d4MB7dTjvKR7y7KtCBF8eJ2H+
LbLsMYMbJ4wkO56SP8tbjf5MPVZMT6v6rP4ZvdREvAvijiyZVZsS3EM2UpNRO1vDOlCc1diLRf9B
p89MUn6x8JaptjEXXj9DzvChaI0NlDbdUpUOQGZg0p8V4KSRBa6V23ZB1Kmkq5gCbYlSk+C5VPjI
foZrOOy75DoZeYAmi44hSChNyOPU937QuaJQSh6Yf5njCSM3UBVRguCcm1/uttA60706dGPgzCQc
QTskOFMfil8/q/bOg0RpKX8nYTNT7HeMIf8/VpzYtbC1Q8roCC+BU+P16YJ+wnxfgrQMs0WjwT9N
A/8O1RUkyA/VyIvzcHG0RxN8os7lRKrn3lPd5Htpn0gVeRuV269tyqIdPK3ZiMfQexbogK9LnaO7
A3T/RWUKEo9Msc7d4jRenbPTpx4N0RTNJjvW48UgqYuxy8VGfT1kgJVta1Fb8gWixxd3yPJARgSY
caJn5SwSSrOtGo6OrqMRzm3qIyTC3f6A53FYR1cfSNAMt5FrPCEUwnSJULCI87YSgQnfWZ9/voDb
2saFvoz4wcFI0krSjgGZPZOl0YK0fRSeV6k8/0fVK8V5x+2iNP/5Dpocsi78Lt21n+yqKi6xDHyO
GIHE6K/TrEXxxiYCmrj+7dbcpk2/Zk9uyIQOSZqT7dUBBUYBA0jk1iV6sAs2OjC2h2XnWbi+LYkP
gMrzoW7GzlhUpVihm9MUg5cpWuqSgNnrVGwd9SkVIzHi1MNcqr9IJNcSvWudvHUIjw4BJP0p8diJ
EA3aYK4zgUY+LRPlFX/dAfl12EvDsdzPPTMBo50+28a3YEGu8sHwwZd9gk7zz33sY2zGdD0QeDVE
5mUdIZaDNNpDnyOPJnEwMDoKYIUE7Kubd0t4dOGxEpopS04M3rpFGjDBj6FSwsC717fwwTJpW9Gh
QuL88l1kJ2V+jxGHj1KGaf7uRDqMRFUjDnxLdBr+5YSL8fwhTpitg1G/0MiF0Ao9Z1CDSeFjEo1H
khzIFoNN9uFQJgV5uiTes39OYT9AK7IxZhS1aPxJuQEOpeNt5C5+A6aWyym+E/txsShToQqtipgQ
D0jqEHhNW/l9qaX4T2TYMGYm4S21/TSBBg1RVE2h0O9yGWO2FEVsrseesQtNcRGNm1ECzrXU3H5B
5t3uN7+1gLU2QjPcoETk/K9s8bRivim8VI8OxO6E+d2+fB7u2DJQVBy0f6Stdud27S63uMFy1+tL
4EmyxL4kU7ZfPHAeYUt9SO3eVOXr/HDPnPaL6f1feAyOYhcqI6coVo6Q47RnySyRBMfRFnvekkiC
2+IzctTEYleItWdVjziejFhRJqECjdnDAfepv0IQP4Iq27IkmyX1MzFNSl76v5//ohiJCaIy5ntR
n37bSXVD01+wRtnZlUSjNuyhK9I5nKP7aEiIR0877pd7FxE5aA1SIj4ctJNY0uS9c6HZDo3yldNX
mzEnxu9BNXJhk6Oksn4XukB7N1Dhdl4pS6bz8+zbfP7rcl0eJ1RCPCfzSNql5My4WGFX0b+XthL9
jOTfdpFiyx3oOL8z78EGwkgeqYIB+pkWpa/YMJm/QSp+pgKcdK3xioG4RVPPyHGGH3Jq9Us3g1gE
Dud1E2gkcrcUwbqmSFNImVaNB7YfKcj+rlSIZU42QtK7jTmjYes4xk0rWu22RE8VGgxYW85Wo8Nc
f9v1hUpJ0LaGDB/xgyvnWWaDyCp4OSBYrTBxRl0t75NaJgZLtBM+13SpQClLnjfOBUO6qdeF9Utg
vaTn0mblSavyRLoTVTtOBDgwyzk3uvBQjXAhzPN/wi2A+bK+usGyvLCs8V2++D0Y6hrl8Yw14fXY
pFO5Ww18Jlm5u2zPo+PEOis0vgqLPZEt218ZUSPFxEOGTm9ssY27A5IV+y6i5MSykJ7iL8mF8IE1
sSTM0yQVzKijEocj5Ko/CmIKJXYtu0fCBewbj9BBVq7QGoX5/E1NigXN8oJrUwOHc98JFvQMMAUr
pEi32KRohA9vfAth1guVvozpRf0099hJERR0omUTr1ivOWdmch9OKZj2Qy4eBmCzt4M+eOUwlwGF
lmKAgkDSVGPWt2PuHniz6xmU/jYs1FHsoip6m4su8A25CpkC5Sx1MxKVWJETFDcKyI5BHPT8UgG+
kVi9w9BOUspB8lBnn2XUn+6bhdUEJSlqOfhx/LQSGPFPe5DUbUsyHczlcbr4/1mfxScIuhuoNyw+
12QLsoUx68G9/imJiRbj3CznHxJVhTbSHjRAeGGbYpi2m3Nu8WEvJw7m3pbXmnasrfXPld4lHDtA
+p/C6GJO7/cw5anqrHaT6prmf6G5+yMBSZUWC6SOKAvojIB4iuB7kbHLzVhOYdZXcMECutO7PR95
714n7ZKryy8y6BU/cUIm9rlxlYLlgBsDpRugQgayRRlbcbZLSNfjSWbecZ+9hQEo0w5OnlqAZg2Y
QxUlzxqcFoLyDiKsnQTqJwAXEoZpd32pD9YBNZSAIydkKmUa8r+rluZwpBbR7fUA7piJSM0SulgH
zHmpwVzJuUKzVmZm84fC+ZnJjNoemrk6d1OPCWfc1nYH/cSj2nD2VFdMolETUbWDfh6x49jpLbCP
IfnYIdZMDqIfiE/VcYfi4e3YLE54qlHNcId0jGPKQVJ/kM1k1F6sUft/+kyUowqmQ9xgo0yuGsjp
8nLoO6jsPPdPlT2K8DN9P0P9GAYnRb1KmY6IjwhZf7MuYslXkq535HervxRsQJhc/xLg2q8JK90V
pZhkNsyNsGaw4GdGrUS+7R2YNSTmz4tsFBfo6czifOAMFHXmvDHGpoExHqDh8q7ZF/N867XjrNBI
hV1bHxlMHdNSYu5GFuZ5izM23Rb7wNogsM3q7ldWAHJTDwVhrmSyeEu/9NHnGwiav9mrll8/SKTu
zkECKXzgGWY8NNLybLNVsnra98v2p+9xK0v7AvsOjBTgD6MdcSnr07NiMRd8k6ZkdfyjkqJh983c
6+MpBvtKmpFMr4+Cp6XmvNpLbc1RatkGE5vVOtlNQrrxLoGWTezHFipwRl4uP5pSc1+jQELHpK4Q
f0i3EzCfkeOwZ1aXg7AlnTB+eMzzxIJN4XSZavWjhsuL8lKNcNUhOl6r4pHRL5LX9wjOZIYc7rR1
jjk8wicsJOdeSjbZUI3sZ0H6qpmjePsBuRNIWj19w8IFr3xzoIOwtIBvtehDJhZHfd2pc7UKnh0O
pczINMO8LoGAS8mAsgLAuvgdha2Ob/pYsxbwDWN8NbY/YmzRg+3RCcXlaUc2WAkv9vjPwQ3Ws5tc
1LvLlprt5IA24JGU2uI7gXBDzKojDs2LkIpoT3QFLW9hyz1fQ1YjigfGoQvH11x4cpZwDtnnfnxd
qm15bZi8BmNnzBZ+nbRDUovc6c4kw8WIMwmymS/hEIxAAHcWsEURQdisNvx2DZkSRlkdK9ZdfnzM
8Jg55rRCjRpM+KFFfZxNxrYJpZl5RU4gCyzuZqOzQ3B+SnnQxGN3HNM0gOwGPQISLkTDTpdnHBnt
2MXF/QPE5dWnVBaRRh0oqLbMr2SaPgWc7PYA/VC1UZa01tcy2Ed5kW/i8awBhE4T42LWBpWHdtyB
c+g/knTd6gHEh8og2VqPrvX2jvgpq2F4cPuUWdCtFy20FkLPb24OBpECkp3pjCtEzfJLw3jVsUpM
PtKjyXSvMla+q1uMAWJCUnRPKkV9VN6HMgLiLht84ajClPjws41N/6Kbw8deafX4gcld15vqEuTS
hxcVQyDwUQ/MZ7qkJmiZf258oye96ScvA2qLALy7cupV/uET2rt8oND1ry/HTi/5jncO8IDXxMwR
5DzAs0umqYPbiOpjOKT8ZwoqMqH6zQcK7I0VPjqq3dYVU6O6Js/tWCwmaaLOIcYnLouP53rcVfPz
0e/vHfHNo4nn3gr2xvPnCn5K3Pjx8mi747elBKpfJFPiNL/smHVo6e+5JhK30ZXrosYt8uP3Cf2B
EgvH0EYUpvzHgaIb1hH5CymJGy4XviGfsNrQuVuX48ivhdVv/iiQlqy1aC+H/Q4Ra/+h/7eCZgSj
6n6q/jjXUBMGHSApbObVbgxVp1DtRAtvn4LUd3f54ABp8l6HnEv6UMyshU7yeBCOZ84nt/XwzVdi
HiUqqAjx1Y4u56WQ2OL7MDdzQz+nnezHo5IIKqfrUF4jPB1v8Gb3aDUeNVjwFSIy0P2gkVqLmRBo
l4kikoL9JCK38AL7kETFcsQavpxJ6iRq09zL1GOX9k8Cmyz4jWbAGRk2KdEHv2nntRdsXuev00xl
SUP44sqzptJb6iQyzvDv7EwySM7nUIRzNfHeIuIEO1VtdDAuN/SL85WpsSJ3iFVtQ/HpTWqGkGz9
Ni8lzJBJQSTK5qP6NG3Rmo2ZiAMnfHbkfdYPZWik12eY/pftfsbvJjekYfj+R5WuRuneEOcBYeLb
B1QXm5SX6L56Lm2+eWRosA5DocaVO0AkqlqSNAFYXW+R3M0CJhAA9gjjb7JiZxXICXzPad3EMHvG
w4TQhimdkSRaKyGWxOvd2gKF8s+cKjHkO1lpMj5ZWpoltp+eWXoEx7TV7YJ/AqEXTzjdPV94OYAW
u93Wy9MJuFCcL2Kc3j12dFNLkJG9G/3SBbqp9wJ//NAUrGYESQzicuOxWVK88Kq2INbiC6Dl0c3L
4k/3H7xpVbSiuacKekX62L0qTQnjqaqtrGJYwQaiFUIMcN5ynsz7ndqVcxQyi6adJhM5vT/Zxnyz
NZs1yoyhSuOK6Ep8GCwC6BkqBKasHefwVKHzGIkDK13RewJLS/oqFDIHwQawTozUEJWwFVvX7Gs6
+Qmm2xBTRLwWBz9YBmRd3hBgzWu1HP/hqUxIyIU2QHoymj2P8PfpkspvfxlMWe63SCoGSDwtmqLx
lQcbygCaioBKwArRxofO+Ox49Y4Ece6EBhkeOlMUSZGGj4aUEF6z8oKExI+f9JBa1jSo9NazWp91
+P/CIxuYfCqcEAdD1DczzBGDicuBL26zeXo8HpnB+Z6b7nJpFNHy6m77f+yJOnIWLnXyOpubcuBl
qFxPPwiMqY7hb/GtncPaKTYAJwYanVQYe0NPG3JM+hyTOoUjuwjSTZI6e7hamDqXA0AVlKFwhwzJ
2x0A9IRnHE5tjGhf2REB921DMrcdDBoCfblRwPZo+o7LaDsy+YcVB3tZK5v0s7YStzR+1gtl8V31
PrehibInHdctDiHYuayzClS/nQkZTW4TjwOvbAkrpLYym3fylxPJkLBtA3gTzwp6fnxQ6mkD56sn
Doo2QmHWXByS6HpDarcp/Sr9eaDNGcvGmyZnnTPxaMT477SSSp8rAIdG3FugbJbJTV2u82lFMgge
DWUKJ7YWqVleHiSVnmcf8kbEHr9hK93b7GZvPhnsEmxhNgFDX4nPqLzy74wUpA2iemi+unU+zGyD
oWRi0tkvralQHAc5dxfOQFh4TmijhYPHsk0eFV3TslzcayLWoD5q1VCjzJFhHW5zsHUS52tE+ImF
ywhS+jXeuZXVIwjuYy+5MFSJ+g8ZPmvf1fiXoys+xu31HCPbNkTaRc5y1UuO7HtF2lauAKc3TLC0
8tDD9szrqmqj0zqHllbBd+pdIKPPYLLH/ZXWzCLx3MATZOjikqxPs0CSD+WgI5S+vmyDopmhJrzu
Hr2zdQO1nU8+Jz/2FmivlCpMfa6llm+ywH2To3tHbMOj3/unFrJW1IR4K1Afh5cXYEweikAyv7TV
b3RO0bMiJuxhe0l6HyZ/ph2tekWnMj4O0qfA/S0Q4ibOS9+9jzO2sB8Vw3E8i8DhsUquYzvCAkXd
oyN10lVZaSC8BsLtdS+fEbb9faMIeaPjPWAxygh32+elJc6ZEoS+Gwvfp1Mhim0Hl6rf6V4TWDBp
1xkSlw7fMIEIeRD+F+Kf6dF6r3lS+X9jJ65MVE5RsuALgKNeeI1KWJOwfjydL2BCKTf3aXnwenY/
M7yklqwTXy5+TZ4YzYsI3gmbK8aybkx+RYIsf8/evqAJH87qjGV3JALpq943UjrX3Tu6dF5+zP1J
5ktRibt7mN4EJKlOnePLOB812nRdi1/NBrtiFUCrW+peH1AHpOYmC/vNgEy9BHqyiqr9QWP3D/1L
Umt1kiIg7Wig+KpfTdJW2JdZEpIt/RlBWtCzAuIk6FpHX4EB5YUfuXvjb+bb+bJrcf2cxuq1z9sX
J0cA2RxtyQndwS8pZ5j3KR9LhJbOOkOATwsLp/xFUrP/Bh8p+SRcLRmmsmT7KHisOR754xH0axPT
oP1QuVsDqfxg1xeLwzqtv/lymhnExOiC5qGU5NfssMYrMygAsMSJnonMS5lSs1SnkTUoz+2WJUy0
y2Pq/BLwZy55Om++JZ+d7Ym8TP2iQJ/7Ea5G6C+buw7SU4xas6g31x8iogPMV7zZ09Psijoh2Rco
30qB95frof4syE8ZWPmp/x7DRLnUiiLUOcZY47puuNtTOJ1chPEPFj7xNIlkNhtk3y3yfgQ0OGPq
cmv34eONZP9Lm4Keibnj+eUu03YLf/rcbnkCoRIokShifWj87/NvxJDksEessTW8LN7eFKOnH5Nl
Nxdt0JtVQA6CkVbF89ap9cqpw3nNKC942JeK6rSktHT/749YyQZkPo+8ZhnTGZJOQBvD+8ojctB5
TNa60Cy7CpX4eMwBjROMWhWU+sL4uZaZBdorUq3g5WDzB7kmEOR+Dy5mXMx+xDJYbgCNY+wJ0DRI
InWhbNuUWQCzHEODabo7emlPyigJ0Ce3fh8FTTDOWzB1YlQLw0ose5aj8xXrsVKhhYIDQGFLtqb/
MNDPNKJ3VM6a9Cz7WgCbsC5LG+krux0NQ2HE40ktl4XVfwohVhtyEvpUomOF0WPHuGupNUvBoEag
VdwLo2Tl1yKnGRsACzX+VRQa/rODCdfnDrzJPUI5QWiryrr4QmOvHzovfVJkbOqO3wHKx/Lx6o0T
TqOUGi78jCcUulVXyQLXkosJdjtoygeJJYA81Hi8QHtJ3Jn50IMiHA5FUbgO+S1ibB8ebh/1GjkO
lvKaz6C8ELo6eriXQWUrdbFWvqysxIACsbzJPKXxaf3kq4u+gWkJRfIsyb9XPTGFemp2ZbpSEq6r
WtMvPMIkIkXTOxOrahDezPRJgWtdgHVXOZlPryNk4eoZ7KPsaKX7/e0le27NtdQ3Sxsip2O+lHTC
DUmbE+cNbZYzNsIN01UwphMkTcrFFToLolGGAcxPTqVoTVdc292aCyguY4swuazPZDmcOvrAKaax
QkL16OZC+i86mYSJAaTGBPy3YUFgLg6KAGqApowB1usFCStOmtTkmsyOnKuYG2z5jma9k8wAxYnm
+fRfaMEtRWXXYSRHh1j8i/s+FzSxfqhAkcfoJlnFO975XHe3m4PJhQGUgGHd30A4ChyzX4P8HeIr
hemPFDEnZ8GQBDUyFR8lrcFLbsPNVNdRhO32dXUypIbBr02GyRjwlD6sOyWFVvfrdqaSCrmNSt8m
gxLxmA93CuLu+0cutdfBHOgJlZl1DL3JH1z1h5DjG8a0MFpg3AU0YYhl+lVyli145z5X3zF75OjU
g7224RfA49GI1GjEQ/t6ywB4Ya6iE7xnkG8DY+VOeiTyLsuP6Rmf9WMS40ixmTMqTFDwy8CjvBpJ
qAa541B+v9GEzpV19MDDPDDXwintYs8lLKvTBoEPfzfmlB0UPB3SiQDAOWGjOguQgh18d2aXl/ST
ByxWP+GzQG6E8QTfxu/uwHyXULAgrV2sllUq5MCghgQasuia+IumWBNpnwcUXtvA29yI5JHXg4OO
lyeDMpYugaYfCoPD/TcflsQeYARSnDwChDXOwfDgbhglsx7Wcix+T2oUZwufbsaqFZmDxkNfZlwM
5P5p+5/AWyaUAnyQ2A7p4/nZAUNers+DUbwJjfomUk0MvcL6iebAo3go9BjScfSS/G85HoqLxbxY
4SoCKPoSV7j1decVNP9Lv0IIAhEHejkzq2c4Mn79fmMmyVlLo2IUP7hhXSOmonX0tWkbWsgr0VpX
OZTjcKC0fsqfKd9zeZusjJMqltzKRLAZFDU3oG5PnWRqKGpI8yvF0SW4P89dy53/JBZsy5ddRkY0
5GvUfmoAIwzFVgQ6vZk89heoCXlBKYeVkzw6HeaGy+0CxURInC1x+ppNDVgmYTm5pDQ/oC7GKCCf
22Thi+SqFui7TCEj4EuuFtfOIE7DgLZePwtPrZ4ix31ZwO6a7zVrCijgsX8S+j0zQwj3B7NR5XUD
9kM1wDeoTilRtDLfFZ1gUfpWwWmIveYCIEQwZJ2NkfDTbfiajbM9hDcHG9a1qSGSt4dV8c7GiHaL
bmnPU5H1VNch8AmIY+HmPn5uE3nXMsPG0fvNws8UN9OsdyYWhCGjwRBkk8AR7UFu93XV1RqbZqaF
cJ69Eb8b9RRl5OK04Ka3RGwFfAPJkCJj0zEY0cAp5yCZG1hk9hQvsUZ62lKlBoHMEfd2P6qP7Ae2
PH4jDw7mWN9qJ0v9H7WvD4g4DV+ovPZOp593NRphi0hv8Wdg+1BCcVuRoJgSW3nzk4ETvWIig2KQ
YWaEtNwokThzcPfOIptZ1ELSDE7T2iiRRY6ggVRyWqITWcOpiUB7uIP3UoRhpxB7CoxeWDL73YzN
8A73ZguKEnBKH4xGM8Q/gcKkUnoFZhthvnN2Xr+ukMeAImlAOT5/W7uIQWG7XvS5xM9vubcU64mQ
biqP6gJcmpcZhV+iX9Pl1Go4ENr9Bp0FF9z4DEfs5OspH1JY123c5E19gNQyEhwpahpmP88LklxR
+5tkJjgYkg1pI/a3BxRmYve2FDnV4sr4/ajqMgpk5m6N3aEPAc4d9ZgvogKwBOt+PL8CyFQpCuYA
JokLy9YC7NEpbcqsfSzCdE5452RtdG4EGYDxn5ZVZ5FmgcG4X/Fwxc7ZYv/kH3UoEJgAklZQ64Te
f8WCAH9/q53cuopUwtWsO4RbD1cAPwoGzP1OqFIYDFd+EmNm6dCWLFMjpPhszRvFu5cP/5OzHjIt
IAlohph8YyxxtmCcdzJQqBV2UkcIKU1tj7T9YGiQda1pNwsIyr8xIem32cRUIW23ZZlURW7Uoqpn
0oGO07GSwd6rVTMbf9lQQW+7qX8bi6hgWQLHIlgvwZ2TLSGNm2xA3ocKqm9OZFNRGE+XA5UIeuT4
I/+DfTfIBjTzIhHAV0mSU5bhFokBzgHEKooVrkc269wKpY5WYR/rkiYTwfi5gn/jjPXNcgX4uxFK
wtyn6t0QYrZ9qHe4ldB45jOwsyV/FJDu+/Jk8pz8EscN4YgDYmsOPZsCsrxeRi/ffnOzdnjYQVOp
tCNVuBJZWi/htZq7EbiEW9YhZKHnXt372mCXCys7535Gj8tKZ+6FumFfUyppELvtjdCuzKkzHXfg
d7m3yvEgRjsmKE45mVhBz1DmmG/Tc1WanFwo8x4ZtF+Exe2aUsS6WzsShD0CIuoikcaRkts6WWp3
qhvQYA4xuciIdk2GV6QzuV1Lsz8Fe+uJDDCsfrzPmCStM5S06kuQhlXr0Hy4+L8Q/DljnDEe7Hld
TCK+ws9MkS2Re0zQn+5SU7lW+Q29WDg0GrOowPWw2Kz0ZxQnMgE21oaR6/c0ncvug9PgyItEcARM
fFhkFD2Sxa/59Mo6jdVSB4BETuimG4tgcfSYe7OqJXmC9xekH16gGkYPov6ZYMICgLnH6SuimiP5
mifbcqf5SopYq4nuIstUBO/4b+lIQ4Sm7nG7d3LOINCqgrKJ4kSppCHbLl2jhrBnDhWTP0dXj70J
XYv7TOjtjjp3QddrJ1wXZ/Z2VmJrp9rv3RIgrqQLvC/WYfx2s0i/CdnMYfSV2K39IDioxrZqE/i4
veZ0ADQVU6xBrxXiJdzWw5za+Xl/xuXzesMNScxRvLNmL7PjhVFR2liGq+NQezNjyIrPZpJBVr+9
gjgorDjp5nwGAT7vBpY+XWLxJl/lsAS+mjT3ji8Zpi/fPRyv/4of8OUo8OZUddFqjdz5xP5gugBt
3OHZ9wTIfnnvUUxs7Wuo/xL05WRr0AXe3Awj3v0YjBBPwnxbEs0vAboIoBTtj7jvsN6nHme9JCST
xCU7jm7VvZBGlBCOa2xPA9cf7W9xfH5ptm0ZQZyr4FjjlYOS3IY8qEoQJoq8g1qEtc36I0EARkLk
mg0vSfYhZblaJ9qhuxsrEYrDbft0Q2SGjdo1Y5M1FtMMVaGdrnPtXWk/Vqj7FYAUbdSpbjkAfvLi
gf0o018diFf7vpoOp9sJDsSWZP9caXr5JliJJfSXu1vpCWUiprTIjqPL5pqkui8i0bI8oMCg/UMO
G55/udb4qGZoJg7PNkjTsYqeubp2vx+y1g90MYUM075FOcmgKgTiZhnRhNNcEc4DNtFnCq1ViqIm
lBqS5enNRKi/8TLAs5ltuEM5zuddNRm7hHq7fyg2S+phERFw3PyIVG2A0TwciQ5W3c2mSwBQ/JiU
uF1rUruXOtk90DAQNtt8iWkYEv+JlB6BrOGes6fV772vJO7q52OEs+Z2o24mS3IBIu7BAi16+UR2
5sbLPxRxbIH09KMDDVSUCiAKDof3q7JHsqH4n+7ccXqd3mEG7z4VdVpQF1gBnKHJlxkzDjazkhsm
Gygh2KiuweQTiL+xvJcohH1u6zXrI96u/3UJzWi79D45TDhmq/CTmz5DvXQ89yv3GvGbk7eYz3zj
edx8KVuEHbudSeRCBJFR9dG9cdUhasZb8833FWctga6YfUonFK95DinHFFfVYSknXXoxIYrXkoHH
UTuVZ9EIFZAxKtunPPAdIt1MxnKyRD6IjwULI9FZCnrFZU/no5uPel4izpEiCS8TcqMmAcidYSEK
y0YiSSdNriwWcrGkpn23I325ganVaYkcGn4fJzhqf+t2myrf9tlxlqJu1fRH2twsgeM9MRE6qiCy
cgBPoyAfZ1x2Bs1TKBuw6T+EJFeivwPBa7rK2rjVS4OnxTort0FZ31RdeUEOKbXt1vkEEAu2hqz0
VnXnBF+CumZRZTTy7Deu47LuqUlB7qkd66CeBzTanDQdrqbiLqmZgDkLnplc3iTaVKHmN+uymXrF
d0TKIWId3QD5U9h8+3eJecooI57KNlDTB8eAab81X5q5QKEnDevJYC7PI2/AKeqBqOlWJWHCCLsX
+ECiZdAU/OhpzH2PfPImUu9HJlawNwaexbadJmJdJ1THqrIG/v2178lAS4sQ1G3Py9XKlXaMtFSu
NsTvpmNuck+4qpj11mRKIV7UFW1Fm0UI57UJtGZXbC1ifJQ/CWZDGZ+pDihKE1ps0kzN4w54+rIi
ZCY4VQzdCdMX9kJNz85USq/DgAhMuJE7+kuD6orbUzmNKIbqydStYkO8D3xfP7kIMLE/XlCWK4r0
SM2T/XbPOIkC5XyJ+yeN/aa5669Rd2aBb+B83hzrfm+FVisupwPATB3zYL5lRi2sexAucfvGMhjE
4JHaB9RB8GLu4qNq5K17fPWGVUY2n3aAArA9x/2ccxWfaFD59UDVnfS/85R2z5nHeM4UxD/nZ4o3
9vYEdDfx4E+v3pUVYvX5j5eI0M4ICRgePuzCXyqKR2RrIQikISN7t+gEewlRhpMH9caxU/2yDlHs
2n5BihJbhfKpUhPKT6INTYS9yqy1EK/RT3/VvC19862suB0JCZyb52Wd6QLudstzw9rpEBB4LNGx
CvA/rWB94C8pLkM01iogwMlNHQt9IGpoSkarTgDzfsLsKn695DaTF53EfUnpbCCIBk4WAF73wuy5
6MA7l6x7eqQxHhL1C/a6FqrYdDk9HewtCNtZYwoMgU364mLlA81HK1nV5DelredSLO6J96gfhmVG
4PXYZUHCNTtcPFHPPuurpnvGRI7NevtoPUYg/QaXryNWzEhc96MYf8QpES9GubGuWyF21ZcEVCQ9
zdo93C1v9QIuMsLWUKp/Bg7Ycnk6biK2PZHIDUFSHinQYkzYHi7psGOlmuZEnNbRX+vSGQd0feFL
VsFnNEJtoFB4clApg6tNN67EF2u/KsWWcnPqPlPNQ/qiEMOVVT/cMwC0wDrJUhSq005oj8YlFfER
Wjf4Qdy9YDNOTsqKHyLJiXFxB4feUCUDGNUOjaOzjiR3kjjSwIDrSN+wlawMC0BKkWHi120Jo+zA
/CRlZ8bo6koAN83Bs8ZurH7ab4ieCPBtv6Kyyg2b6LERn1m+Z4eqEA/0io/SW1yC51qMRmxK4Dft
PxlDtbae0Vf0owkw3bakIOy6ifwfP94h4QRnPEiAExwyDWti8CGLBkIrlVOspki4+h7bQ5O+X+/z
J4nmFmpHe8Tf/EDpDQQwREppPz5ujlOIDbGurbjQu7Zg1j0aumR29vpHMdNR5+XArdkH3jFphM3X
Pa+UbJhIqF5kunaaqtum1iC7LE8o6LoA1YK2POR+PBT2NCJAqxU6zlRM4pUH8IyhLA6q14xEc3ho
IEbgHa+sWAWfOGFqHwRuxXqK6RTmLZHN1azGZ2PCDAwNoQ8BPTrTUJdT5Bwp4jHJqP68dE+Cz1bJ
cW71iiO861+weLas3L1vYuKcr4e1LXMxAD/Qt7WgcK7Cn4niqrgfPWQ9krDuzY2cnks5aur1Qv1c
LIHQzppZeUTDabDVN2qnmhPzoMZ9V55ExyJ4JElNPhKHy69yvTKwJZZkWpwtRdgmBeheiHUX/qLp
ColLCsN0qsPyPQldeZlYoN+0VZI9aIzOwJLTGdQlDAnA+lydu2X+yujWM2vGQ7OHBHNgDz4IuYr0
XR9f2HJ3KGUQmJDQxbXXav4EphJ4MBIwuFOyGDD/5FcH56rTuRuxdiEznWXmu6RmCHqDw64gZQr/
DC31zUNxD/uH8TB8ymXCzpPap+09uRhFbiueHSvUPV63TycSeTr4Dhn+UfZz0We47vHqc2+GnPAX
4dcRq7se0R7oOjSKXZw2ZUuwBiPhT9pMUD829j1+DfalT7l60x6pAVqYHd7Vl8YgiWOZ0DhpB9us
npTtHxEnirHzMNycvOBg+vRI7QZV2nktRX5tNEoqwJ5hBqJPStaIkWOVio3ap82m87N7oe2NiwSg
u2+QJQuWeI7kyeys0l41stmHOYiVTZ+MJW34iA0RV2K7mN02gVvqfJ/mwpAiBMjBjHZOiMOitZJr
HeRh6uYOPoGrIeqRcfKqs5C2EvmYVqQQ6bTtUgAkD4hYj4wOKQxQtqtCHAukQRcHsXRmllK1VMM0
by1xO6yHY1pJ/W2zOVYCT9WouWqkSvPqBADByzaWhwWjpG3+60kSFRk8QmHoJ0qbI+it1L4iGl0z
e6q/rnAgpLTsEJLjEC3E57wzNzYme5QTLv9dEi2vy4MvZcJvNSGYz/kDE5mMYkHkC+4FPWPQPf8W
KCBFQJ/D6/uxiu0EhRLozibTUCg664J8AwnuX480IzS4zDVrzcBwH/DWdI+YfcoqVCPmIAz2Bf3u
yqxBKhe74Y3fvf/KSKt76tXDV0rGdZP7a8vtojlPI38JD2mOf3E0RguPTBtDlF8CnX+a936zH9A5
FWDb+jr99VsoKmbqMontSymBuDZcFzi9cRDxBhE9AfGXrT+kAf94bfQjRyK7mbOAoGI4wyfEoZBK
oVFLXb+C7DzZj5iGx5ssAaNFgZVY+xy0EQVNdPDe8paxzteNcQxzZF/NgtNyRxHZnQ/sknU5zjg1
pSbJ0yphIkG9zN3X9IUMSenWstBfUeF5BHkjAcNOmZeqKQ36AetxXmeIw8p2DSX+iFoKLO7z91eG
stdmnhnSUXld9TWdaH+QeQyOwmv5wgRSsKsnyKku/9meqG3GMUdWTzmwj5dD5jXE3qwGqEzZq70H
HNcKqIcgz6GyC+z/4c76w3q03NTxsYpxKN+qqHKLl8EAjQ2Pd8gnA1tEwrhPhLEuaJYL60TaYFcV
kcUO3RKqEqDYQSdWuT++NdVHxDgXcUPiIeEklmUsSBUIITsuw6F6GOQ6GqVbpjwwK5xvvsAvFLN0
QfRiloCc+dIDcGFnllBs3hbB/Mi8vJfYmbKJABHpe7MJe5Khv3cD07OV0bJ+av1N9mxA1/3BYLlT
gMggmdj0LVeEFuFve9hhujvxTROvt0f4mfHe1Op+KzGfBrf+U03LG9ahJDYinq9Bz7BXLsOWRRXL
fOe8sJJoNfTfp/67Ys5ubyhWY9DtIjsmKxMnt/5vkBQqBPa/na/Ilm+sl6YuDaks6BwoQKqWSuVM
yvJM7EQAuaygj6rFk9iVSENr9Syj195NaTxWCGVUqNoUab99KFk8yq0uLyX6UMHGlHnpN7Ampwlb
GJxXXQmgglHZKkl0aGJBVlUlecUFvnn5bd2Q8hwiQQ9cpmibZZJWiNp7bFhix6oXZh7xl1EqlVl2
bRFQlPpX/W2VEYqUFKXoDtMRnDHz7HHyY0jvD/GCXnqCh7SJmcQxMmSA7GelaNsafIkN2ivvJrCL
kOy7EdMJT/1gkhlMfbgR1VNkc2sTsZb2zAT1nFYNMtqrM+fHWy8mzvOQHb1289J1oDv2FDUbbaZ4
qlh+WugP7DrhS/qPNbHq4NclpldYojbb6lSm1Gctb2lbKpHAYs4TWScaiCa+8b9txDNhxbWfu739
SNSGN5Yo6Ac2ceu1Ks8QIeFFM4/AqJkNM9RyVChIg3uLFeRpoIcgX4s7nm0YkYA5zveL4OgFmkJv
2ByD4liTV5VLwl8LABJDdurms4J02jrqE79gsk03ywb1jpNNQGtvaxsYWa+1sJHrUaPxECo0enJL
2eHI8BRXko99Gp9Yd/LsaTvpibDzymeajrthTkxq3I4ElmBmXVscAGjdHOrDb3yCiTWozKCVILf1
HTakP7ydqC/oN1Ml1bM55eMEbJIPLOIFX/RhoQDg2muhJlFeVizy64KOqIZ6rBJeAsiC4vdAazkg
UO5iH2gQJ0z/eDwPPnEB71OoAYkrebT+rPaNH8+3z9nVpLTsSZs++dJSp+eQBO1EiNwici8tckH0
flvMpCRf/Rd2UCHrwmHgkXkjSrRY3wABxij9rE/Tqyfb3RSmeIwRPyFGGeZpOd87VMo0Y9hnQrFk
MweBmRsc00jro+WVym5UCJh9zb6qjLisAQa8pXY0jHazAsu20Crg80qB3Bxgv+G9bLNoZU1AQ74F
3Y9IXktX2DLeTsLrBt1MUHnin1yNrUtzqrr64PkSaxkCoNJD8TQdaAw+/o++GQIIVohlhpcDBAK4
hTlkwtZPRKY6KOvjdZTlziYM467oax43yfvBw2Jk3/XB9caZykw+a611zeMMkUsv0jgUtJH+Y6kk
6cKwOYIqQkM8b3/LKWlJ0DP4Ux2r38prqctfhCLT2Pw1e434aFhFG+Rla86/kl/XbIr45ufe4vS9
6O2vNn9B59pUgAVK9zm0YldKPX5VDfruGDQnWDWzvt8Ivdrj0pLRFemzdQc9cfs3j76CgjUCovIJ
9Po3IJLZUNH62e1yKHsIkIklTidTwrD0YPtwnad+N1qYlmKHqaupJPn8/UvzdyF0L1Rb8Uny8GLk
Ty13Yhl7TK8pdBXhBktLowdnPXqtakIwDoCyenpNXvhDO0jE145SPw+rpoviOraIeHhbs46BTSCN
hqnUjpipR4gQpw7hRGEq5hXtDK2z6zzGqJ7vcz1EwTP3bBKE+DUXmvW+oV5piToB8qq1d5Qi1uMT
Bl61ampB4VtvtXqo3QDHNLNXsKyx007mh3sbAMCSj7h6kCQWydAgrcwX5d3lezV7stECiLtGYnKC
AtTFgCYdVU+0zMPsWG1Q5e+/r+E0tzJ67gSPCQni359kBbxGIpVM7fajevVNiEH9gwzYitTMbdo+
5fnKEvlLRmFKCydwVmRe8zuW5VS94vrPgiYSBeer/KxxeoKwYe3WRk5v0BSeM5VLFgnKT0U8Aaro
28PcGIzAI82RWv9/76SRFKYM6Y9YJP0ae2imbCDw8ie+880D6q36p8jfcOBZiZFH+EfgDPf0LfYF
n5OtYjZc+5SUX96Gmd1XJqKUbCtrHV5kn1D6MuBP4AaRg7H2Bxghx6wyMVYpl+mTB5A6SIMG44t4
JqsOm8w7KqBjOfsaGwcgHFK+P/mYC0rXK4vmW+QgrozJOofq1YZkytXYT/WMWGcUi/LbD8voLQp6
+4p1/lhoR5Xw8WIUA+qiAAu5QYr+aiJQRhncIJDlSvB6LU92RiVWOSAYpVjKaFi8qXK+OTmKQy/b
Jxbi4x/JPYI3Elz7CTEocrovljk/rPcBIfpbWejT5Gigz/R4CADKMLSMYIF4QsET2/gpUDxGnW+p
XuGH8Ri0qSGuU6YKoNuxTZ4jIwSDA/jt/Ryt27KeLRTmuriVXwvuO6pUle5VFkqGDN19UcPC6b76
H/JxQo7xxqe4ziI8NgLkcv241Qitb2uVQv+vWmG3sK8HotdD849HnTAoE1yGf6GEx5rtQlibToqa
BckYu9EX36KO3o/LWo/ohfZb3btdJt/UOAdfIkkeivn2I5LGCVquR52LPJ7OAaEkYORQhpPgY9A8
Rs7L/y86UfzEQMpgLATJf1ePObdeap5gL9fgp8obnzOT5dLyG7nTgI9NDqgIuZHfwrutLrV8VjTu
C7ThmmWdhWC7wlG9eS1pvqE80oN10snVJ2tUfcqe4lIXaUQEjS1HDaO0WQQ/a66szhECd6Cqd3du
bb7sO4AlxNiICs1GWfEmPQKM42Bum+tTdI6ioncuurriVRhASjLYZ/4hITknUNlWanajZ3FiTdXM
qrHTWpgH/wtdbzLY236u/vbZAV4ir6lyhGYQPF8vJe+AA8NlLDGQUQaEtxFL9VCl3gNzU9XG4qnk
WcRuu2gAvXKmKilEnOvy+E1r0qEbZmB4SCUvwli3NK+HEqrcQRO2meXolxTFWQzoTjyfyMqAD/Q8
nJVjBTiT6Mmwu4PBi+VZDllHDUb2D9dXGUxGhqbdEo76BOjg0PnCDxna/rkiwxvDXiOotDGkm7GE
TofHmh4vIl7JyTaXu6kUvk/i5wgnLRGj0B162g1NZZ+PnJUDBrCWBAnBhZQbgFW9Joe7HapIkPmx
B1nLYGRnYEwUeQgEcbq9iSVBrAntrJ9rKuh4nokrswqUncGdL4mpSheBpzMfHm0dc40EVfKO9JY7
Vfnxg4pw8ev1yfAvXikCGZ2BgZZ00A6JfEOBYuhaF+metPiVjpTcw1BrBVPYSEXWbp6GnFZXgH2V
GpiBYd4/YUxNkGC+9EmbNHfmchvYVSOriY+cT/ED9QOGj6BE/eCER4lxqgUbNsptGm3FpbvkWODh
MoOnpzT4fFDXxKMMogD4NRrOLl3Ko6L3P6iQqGBXzl7RRVFh/zlW6f3y3WMbYrxoGzK6vFhGTcoY
RS/Vp79MxFh3w7RTi/mncYUFpK+4ED4oWqVp7woLZqoyfFBsVnwiAtn+t7Rbhnve2ABTMePyJMo+
B7Bhwlu/iXfGulNysBLGXxSHD6TuiM8ADr0TjfC5gPgXDDn/HYMfUs2cqPn9o7IWF3z4mTj8oasc
0YJlUvU6HOWe9fqVj/jp79fdgjFBbCG+s9hs3iqG8hkgyJnzMEvIcPXrG6DDGQ6xOA0vLsfuztPa
bw7TbD9548Sngz2muj5Yv8R6XZ1Pq29l7hs4Y8+4CtJRuS/teJTvYncMyO2oBIH4TZz6u9wAL+ky
qUU/DDS4if2u1Pp6sSYa0KQzErvCYkcx0pXUKSEUc3beh5902EjZpWJrvpupVKsskfKasRrZUswj
zTXKve2gwRIEtCArBrIwmfclQKVGmsf6FSyUetr19sDX0cSadDCZwJQtyLQ4xzWpTT3vIX5tPSlN
7hOwflHOzF9Z2j7p/Z4I+QsxTFhg5/aaTx9n3CBmvx2Rq0RjLSn2IplENWRP9UCT86dOZeO5f2iq
HXe86zDFv5n2tebTJcy0pfFI1gfOPb2olB5sUWX9SvWLoZgl913pxrYlUr0jXFvFdjEHpPvHFCWM
J8SGngHzyFyi/uzr6ZhFNQXeTombQ2zYWXIVtJuMQU+MRrL6p1rawD/U5m/FY99qpUF3NmqEjxGs
a/wR0yG09D6e6W/jgeiARu0rPGtvWqSDJnW2NC6cS/8YqPu2DeFkvS2RU3PywU5VtaCm5baoEXIG
lj0m2GKU/YrAENEEJpN1gj6nKtcGLz241wpYUBfstL5LkwJIKVJInoYU+dpU9Ve+lzuGyUuAUXTz
XH6Nus1/j/skv1Lzobr9absRWPkCRm/I5KYkavdc9j57ZnRplFmFmwrBTTmQ8y2ektAaf4fLM8ou
0rZMiQ16VZJe3cxfYNeP35olwkfHEUNqs4EfjjFDCVUuYSVxGnsubMUG0vCRRF9oBLczJ+jEGi1B
mXDfDUcIxTjzzrVURrk+C6JyBQyUYpgWYr5Vdfgk943OaQXlIQ4x0mRA0ruRKkFka7WAclg2Sdbf
MKztakY128aRA3koU6FHOkxMBlebyMhrqQvm62VuP1x9o6gpF5iAj5a4fkkPFTiZqo8v290gHTGG
i6TkHXh8LYUdbMUh6uWPXFJZmBXnzbQJXpknNnYaOzpst/hXcWvGn7VFa5OzXgYFXCuhX9qffmY8
T2nD/DlT8z+CiLUclEuEuBw4jiQpTsTtEWhv87EeL+8R4Q8xwWFgKpgViQKskI9xc8ET1olc1t5B
XE0Adsg8gSbSrIcBWQ3l4kp1BJKzvFMYGBXhKHHxoEuWFkE6ONu2I+e+c9ytPWUjQlhppGNlo6a9
PZhuNOfKPC3jPQjZWvou1nKxH4uX3vWhnlFPOpQzzKeYi2uzXE5zY6LQMvLPUa0iECWv1vYayia4
XgB2+hd9HTsdEgMGtPRu9Hdlq2oiaz/ack3mfPiwLxEeWMF7cO4qTYHCbvGgwUTbxTVmS61FEvT6
PSyENkEIrqAFS43c5U5zqvW6aEZtFG33tKxnaRcEJv6/TKX21dO3/c0LblKoIeth95Rpjfse+ihD
C0WwNuMZ5nixnm6rRFs3gz1Qfz42RlN0lEtQepoX0xLjESbfg5GnqkeMCVgkUwYbgif+aPkFmToK
ntfodHD2kan9ioI0cP9AYoVuv/2kCLTSwWdCy09L05ECHhPVFu+yZ2sJ8oXqiuKxW9Ho34ndFVV/
bTCHm61xQQuw3fquNBccQSJZKZN6arr/sOAqQTqDEBniNQTnrx3CBa0Wx7WhQIU/7FmY0bTg0YbN
GXEPSPTADCZwvUeqD13ckF43mINd1dJbl4V4/br9vys96DjmPOEI5dVZDsH0x2c3f1t5iNZ2Pc++
pYUm4n2n3Zvxge8/eGX2MUDJlKFpAKj9G4HzAo69++3PetRs1/NSn2jzKISGWZnIymXQi2YHHhjV
CzyYuqVKGFr+aEh9aiCdtKCgNnhp32dqy+pYTu1hainKTW5IGPGzB3xWiVXgqdlQpj0+28rabGE+
7DU1FsuR6wlWPuJg+pEJby82uv/gpGb53ukiMzfYW9vEQaTi44i1WSMMP+TaZKwqzRdd4goQaYL2
mBuU/YPCXPJqNmcJcovtgvYLbAkRJfLuI8YoHpc5gsQGX7d0tmL5pLXxQxASi3dr8ATeSh/nksx6
LrA0HoAYyAmBu9E8UbbcPnE9eN53jKn5ycUiWCbf1yqoxurWWxbjZVBV22lUUsrmmQZYPvKScURG
o9SHZIwRIU0DhWnf/e/oRKeGDLqjP0Pk5HR/jUvjuteFFRY0Kn7ue8ciNegi01nfx0Jml2dN178b
lWc1LBGO5/7Om5JNu0UcdIc1VypTO89DLd7F1MkD4BhPLAHKu4AskqvXMySawPA6sdHYN6pzM+IQ
7y4Jd/MWeFAe/WZM5ETZdl+8ZeQbXdKy7IjgkcmhFRxAw7Nyit3fCCVm4BrkhJM53ED08jU6AeoK
OzclN297yn/XIH9jmgDFI+VW0SGfEyBq2MaaaZ1XV0cBDUpT1fGfv2BEpdWkiQEuE4h5d7tmXHDQ
Bhv7PHPTnDDjc0FDzZseHFVcf4BmxG8R/ilvfR30UT49Y4N4zscUaSqbIGvhcaXFBAq4JdOp39ow
jlV+TGiq3IlwKgk9hvmUPVhGWYd5g/ZI9741zskhsvYEmnVJOlAbm3uof6ckJPfNj8cnhOL3L2E/
/ql/qs8SgnSmG2oiNG344+9BqR7wtqnDGb5Qt4+l2bKOXY/jwsqzyzesf1rq3B05bytpaLakfKX+
1NGegney1rA5i3PQ6hZdGOdUbs3yGuj0g9KWNsmvBzwsqn7yy43s4iQuhC8Lj8NDyfC1RWnZIIje
cc6AMuqhlhAbSGFvSUV9dnwW698X40/cr1EJZA8XxUOvFMPBBGUlPJs9xRNvBSa3lneRGD0Evl8V
efqrjUQCapFJu/zyseHIaGX/e5Ntufv1pInoJ2oOBR/Vv8oE3xRogjD1Odu5tK68fWD2bw7fHhc7
O3WKVqAP5v7PiFeHijvq7VtYLWgdohlFMmYun7PRtkSyNPpEg0wdHrzYchcagFMojr351eoVVmVo
fxlxUbMrp2bkQmP9dA2YZJT9WFNFvd6iXNN65M5/9PNWee+A9d4qjGuECRQ1ERg5Xs7jHnp5aThm
5GCPLeiv6U26Y8IqeiYsisneltewLJATp7XGTEsgXvbJ7b5bOe8d4r2e8OM1AN4OxcXJTQhTvDH0
HakG1Swr0KhBT7BlMy56WJFlfcVY/g0FMptu/qGqhiID/ecCkcr2oF0n0hwBNqRShHkWuJhHsb6c
mtoUZJoTdiOlLhiT41HamMIegvVKb4UUPLTh2w1oPHmngxbfOYuknMvJpEmA9zPgt+jQNTuUPkgg
l93sfBfREJtrzDLR0SspCijW0wsnTgi72PcGv7ZcVfZ8xZEoYGz0lAjgtRDsQjCA8qG/pQGajlv4
tHiLFaOdmKrqwzDt0xF3BOd1Tf2RedPDA+7J3K52P+NS8kTYDdF8/4M5pDBPrfJPBwHWLosX0Iql
A/WNtJsEsmEnTRrKIkS6t95zodLwz92iMV4fdkVqOFd///Z8bgHXojeoHalH1zBszh5p2ZmkEz7w
4ucgX59nYU8WSRlq6LbA6rDjxsE/4sikVFx1OgPAUTWD02/EcgAcYprPyFGj5qmsZ8XccYwhWSfF
Z/tTWEp6SsxpHz1vG4hHqHKoq68WBR1thk0IRDbK38/Ile6xRKhSJxWJA8hgoCYO9tLCcjk2GI+E
UMSp4ERMB76T41qChPxMdOmuMyy/AaCnoIquOgMn1ujXmlP3inJnx57l07NiGgN9u0ZFpFCIsbuR
mauCi2zrRwKcvHA07B035q3PHNQfTSebX03NTpv0EpV7zQ4yhoc6AoVsM/W+++JH13IjYhxmYzVe
DyNfY6uuxBp3Tkiiqsqlpdem3KcItF32qXs76A0vSJp0ZFpbX3JP7H3CKxDwQ50vxa/WEnlEBaWD
I5mUL+0560o2j0zXK+WcRJ9IKORfeKcMruCstKZXJtVAddrcLOj5R4LkaiBJg3W7PgBWn/++lXi2
YwK1Qw6qBmNoJ22mUP3Egf6guYZRGVLpntdxvQyPidAVtk0OkE0gM2U2xCDQHlYcT+I4HCw4wF2R
WstpSQzFIoFeE1PSXpCPoLtJk++tF48SNF5mZSDwCCUGmxCq/8/WUr6Ec4o1Oj3f0JJLAgZxDrCD
qjqNfzLSTvcb12w447BxNddXGe3jbecZZghYrs2XDiQmGKtTiJ9w0e3Xygv/GtkXGi/VJwgIRKc2
45Wcb4GX8l8w7Cw5tWITs1lNKDPe3Lv3LTe6qJk6DpUaqMpdBph8PZ7MfkUBS94Biscp2iTPqpKo
+DyclmIWErztLHc5o2j+60oXWsRYB6rqqRGYjm4PgDbRTP7F3co3TQ+93HNRNuVMN4bbgNmam8u2
BTC4S2ZcBiL3wdXfj06EfFPNgLs+nddoM3MCFEONyYU3Y7fDhw1q40V0A4MXgRIFPkN0C1uUz9gm
vFPFxVkvywf+m7ejMWvAukA5YNTVIffIFPbV2WWBW2mGoibEQV3VculbqL3iW5IHTC4IFne0m224
kvDX7n6NJLI0AFYNFLDZk95ZzUnqYDV6lCGI5IaG0QoDW2K9Bak35ys7L1eI7+ZrZJdehZ0bKJeb
KJWFBEJWopPgBEv8DjqfKuOx9amwqGJQline1LE/zaYSzMtKTj9JpfkwFB9cSMA31VdL0afwNCVA
LVsUXy3lvLcm8aQCpRtYcoP2zKk8oWe+zFImErVfljw2CUXzyqrzn9HDOpAfnC/u53vpU3oGSxOQ
/W0CuiWQ7rsYWu30I+psP+dLkdi8S2nwEZQGkNVZlBBrvR9UJCdEe3QxdbO2Uj/n5OmC33J9GPO5
KeSTMdUihOFXAdsj9VZywinri/09AyfAC4W5lUb22BUNODhZE004aec4v4xNYdqya3YHjynKoy+w
x9Bvg8HoMC92Gbh90QeH9QX/RssOj5gwIY2OtoJuaVewpmC/slh026+bGJUeCtUa2kq0lUEVacDa
CW1Q+Cy5elcor7SDlMQb5zqbNFfbZfUq3ZeTvixGVh4JsIfGFMzXoNRJt+rqidgMLD1s1qr20wMG
FIPJA/If+mIgbG1JzF3NWKlIwDC5B2acdz0ibf3tVTurpciZpHT7mkiYJIXolO0BwHl4Tw3B/Tjj
aHMwySrFIwS7B4k52uDx4cdtCCyWAsYxqoHht0vGxlbVxFdYrI0unhxW4otaNhzHZESMOXCSW8/o
erlZlpUe5Vj+yFc6daHDI500EmofmtfJ7JxZvkI/TSSQYt7i+abj13FH+mQJvAeDV7n4o0hrjP5a
m3wC5+0cW7bedg8tMWheecw9WyEqOzff9bWrOjHjfJM8tAd6AGL2dtiLGakmXx4F/Xl/+J/B9z/G
t2xjyN8VBkNSt5CPaBy1UTySzW6QV4j10LzpesNPCEml/Yk+OoBYsJryEReJQ/lLCeJ1zMGoNV4m
UmPPI3g+gz3/jsCbyXZmcmDsT71/aI2yd3bgAfd9M/qtJ8IwZrmgOC/eO/9+WEXyZ1cJi+LKB4+M
AMXosBtBo334aCFdum5Xty/fRYWl3hvDnp+6LjAkYKiLmcbThPPlBiARZsEzkEaj8KvDBUtZn3Qy
ZNqQ7Aymlk03l3E+FkEQ2T2QjgHEE7bJR4MdEStQIN6C+mEMuJMx+hf/jFrRbo84810nDoVUvT63
Ro3Gl8DFphaVoJWxq4Fe9sxnDrfZSRHBFyieRGaB1hiVugagAe18u1VYdzlbFj3rG0OqQDiMDvEC
hUIMlW1qBDq92//BkKzh/1dmDBPPLAq7z5qMX/AAaA81szoWDv3XRWB5nkMVYQWjQn7GCCcA2lsW
ZfdhM3BKYpsg8N079/lEtdrgIOG8B90cUX85RIhnLQsP6OphK+W38ap4WcLeKn89Y6gv17P931R9
hslcOs6CsOWsIchYwxVqkqPf/mzMU3+7OfVJIwY8ArA2isUQ1Mk/TlMMSLumK91Biln9RUqYsONx
Te/BF3JObjnq5SRNw+50YVON1Vz6y/HxTOT1owktf09RC4eKQaccbekQuxGZC4qBQLepJ+ZN40g6
Erjo4BSosYB36rXYA+MXOn4ioq2IclacR3fY5EwcfyJmJMnvehvMxrbT0f8ZXKSu/oxfUuEYTAOa
MiM21dWpio48MrOQfQv8lTFseetlXnjENMV8WsGcxKL99Ub/gpnMnNuS3eJq3909ePyyztZ2B+q2
0l6thifJ4WmivnS2QHQP+aYSaFYvF9xwrZQRDvh33P6MZh55UUA4THNmAEw21e6/L1EC2ZkwtUWF
/m+ff6ybgds9JmtMAMto49wOG1Oa/6jttdR1JiI5Igvess9JEXh591dBq6qEqR8zTHrktq/XrZ2W
ap4fNk6Pa/CPtlClNX2a1gfUOZqjpG3qRqH05r14rdetAy3H9ljXu49R+L9cCALq8nmkuWsr1yJ6
OOfLuB/LUGgHwgGCdf2dAh22+M2RiAS42+fgXP+4teHCvKMbVUb/15IRglN5wHN91u3r/pqPzO7T
/bVwFa+SUki1Rxi2nD77AJdZTyzLacawZvih6wuTzqpebIAWS6ugf+/Ul7cWPC1BNonlcXkTFBGr
1TLBebP1yl9rpETMqRbgPwcroGJGiCW4oNrDgLRYzXjGk7flgY040PKICDMor71aaX1vrVuEMrBQ
waNjEBaBUqkGEmtiMKYZvEpaGGgWPEoDzcX1vbnVmOvLEiGF7rqBKG6SVnXVbQkOL+GdVDqOlhex
Sg88G79kMkYKykAkj7ydMOXp0tOEYDxbIvI4l/pCdZEcFhwuMggBTN4cN0WQyRCVB0iwUlIdPVTt
QyfRfiaJzqGI6k7Y0moghS2/vxe5tfCdV1QObXaP1heGY576dAc8liFKqoTOjWxm+l2tbqecCzRv
3wcEX9owtylFrg7l8jy+U4BnPNQRSxdl3IWmTeczhunp0PwvziJECMXa7X6VLfQg4ilqEyQknJd3
/kt4N5qylTdQ5sDl/gKkvbVQ7bpHwxtj5Fetv1OAKJksENQvhQiteXthJrWGpgqXf6qPwQhuu79t
N+8+ZCAbMmiDfFTc7yK8pYYHLfRn/uHyqmfflSB8y9gcu8MxdhthqsVXPHEamXnYsOsor/ECHEO+
x/Tphr8eaG0sAK+dFs7pdj7teW21RysKm/jKiuate3ZA5A6R2NeXti6f3IaYGyLg6wpY4trtMj4p
iAHERuALw6yUbvLNV2mHW+HWuje4DiHtuAdBLxNYXFBIaxePPU/GJrYX9Ep5CUO4SYNjAPgdhSvS
+qLB4U75YHhoLp/T5+ZDEDQzQVbhWK6a9JaBoAIPRDrC7F/EcstukfxP6QYFt+LWAS9LSVbmQgN4
zTWlFYLynM2hFciy1DEnRMyGZTQkQGQ8chJg6O8w9IGt9+MhJD6xEWFYtsXLRQ/nztyzoptwchs4
PHuDWMYszsIK8UvPqPzYw+OyUfbnzptpvuafGaqqjpNGKrOmL7BK0ULtpXxLXnDhyuZbDQywnr99
OyyybtVzYWVZ7+5LO7sb8spgDOzZFlUe5O1hTxyVw3GCwYUS349OsUm5DiLZegTc1W5I1EFrj3pc
6XjIq12DQvGbVVkQgF+6Rafv4wDUKbe1AARUKlIRnq7P/wqZLMsJtmQzFpZvRGvSiCqzQ6x+KsWX
p7CWU6IIpYUEb1QrYSRu8lhelolkv/7GOkeTy4v8zqAeHaxnx9HdSvoYj3uAqJN/ku0C6rEXO0o/
1iPNfonTxin49RhxxkLDBqVRR84A7mMMWPtfcVYRdWYkBhJvqcLjO8Xm6Ul8M/THIaZ2UBg7scUB
GxZM8Db7xVQ9iFwIZdTE3phB6Ol+kSDj2mqCacfv/8DT9ls5lqAPIb1XZaYnjG7+zpueOlDBNGi0
YFUlBplWVJ92FOm7FiwuCN1aBDzjjQE4gsG6HdU1DHNOsg8nJdblKUS9osXpnprvFRTXqg7iYgtU
OAhlRvLVG5nzYHO9hB34vgcJTRRQESLhBvz2CdTSEThPM0QgwFmdt65uEAoKopqlndjpY8i4cMC7
HBHsJ4lu4Hzw59g/ksoLHVVp9RJJTX4STsIctGtWl8CVdCuw+wcHe64o7tTJuN1Fuyl8VV3+XHNJ
3f/aklA3PGBuE1redphj39Aont76Jz/U3I0BN2E03hduyJf/GlsGOdTnDpAx0bXhyE2lEmiikhIv
CQ+6kkdR1ln+fubqieHdbPXJDZ88zLACVtnnAW5ajQYWgBNQS1veFsLOraD5enUuyCfHgnCyRKKV
3H0tFpL1iMyBIXCl5R4yfntFpbm6Vw4gmWQHTdY84kqFUb0pr5Oo91DkTNva4qz3nvw6ayFj3t+m
30ipgpCEPDFvm2mlXt4F12CEdBL8yklfPbcB7Y4liu5HbaWZMgS5MWwAbYMM9kRWMr/lCZc/0N3t
LTBg/JKU5+jAwJl4wkGAzxhzw2USBtY+anXMNh8ROP9UqE5xc4ll8YFmuNnmTiTxCyov1RrzkQEp
YE1VfSXLSrvUc2BDH+yQE8Wzu9OF5Y4PhrOVWMpAPCGmScSZ+VoMLXiZSnctAUv9Uba8y96BV/kh
qVBp882XX1GebKcLPyUm3dGQZxJRpNLJUfrw8kaTcNEI+KlaevhmfnEY080IG2wWRvuLX6h00dLB
rgCZW8Q2IVUZ3c0E3mY/Z+cUoKFnJ3k/a7AyLxAHcmFEBDYfH3IUAeOXHwUhjknT4Wn6gtDETTpL
j96MBlqpNZPzSbTShUGhvNm8ZuJwlrBuA5iqklFJbVxkPI8V1TGGpk2LMjLg+BQFDrD831LqcOgq
jxtgkL9+zo/yVpSPO0APS5foqmH3a85BZRIUmtn8D3JRABdchmOz+uZt+hfio3/BVA+AY18or4w0
hNUph01bZBXKAsvsVNMZYKIAIC02pIhXeQpTicUlJJdH5yNnekaqG7ooZGg0TEY8rsqdm1TZxHWD
3jLjoLrY5Cv+GDtLSomDqUSdwR2CuA1Fw0YU2DhPxrcj/IBHYCCVCP2Parzvd1R1tCOUJJ87LILe
OXtdCgrYIw2PyXsnZXC/Uv2tWxervUSS3ZONRYjTF5PcF8MULWyTiNCBOQqYmnkkxW/ACGTdB7K9
07Y20qdXiSHcXwsFiAtd63CudlAAJ34nRKuw1EpOgHOc18jRmek+vQB9ZE080BJeHfFSBcbdDcZg
kE+65lVw3gaRun5/DnceKOxVBHLiU4J5Tr4Nmub0fyzSYoR/P9/nLjEZpNaRnom/wPs4SGRfawJf
7Zu23eHZO1za2fLSXbNlawh/VnceU6nn0zGNgYRsKEx/giZoPtLquOPYUhEdEvGiOJBvjuDZXoDL
Go1zeBAfKG24Z1IcxZKtQ+dQy7We8f1TG2JneSLJ7z5yRdgMWBn+nH+W6g3k0ohaOzDO43yIX4yj
kUmFtVULtpTzGdiPwTkU1j15XJbr4N/F/DLNHrLYoX35KYaZ6OEVnTDlNWa0M5z28bI25YeaUZ9Y
HeUNCsVYHpoLqAOw+Zweks8EhRrgdJKkpXFHb7DtAg+scTqs0ZoZf3wX4nw4OUBb96+cJ56sX7mK
KdLHoqbKRnCxyivfmPv4nMDgyDSWBlh7rIOSJiqxS7xoctIkHsIliYFXLi/DdVlT39UVUb8PREjM
xoIgsAdKB0refaIKwhb1mrJA+MLMgQMyyuQcvPI8nv+Rvqosnnr3I0AsSLj1a2hPFQy2wNLeHjLL
oMeuKUcOeK8kUpTlPuVK60zLPtjuzMU0ptAO+71VIRQnplDitCp0VsZpQEPnonT7mTWs/ZPwkW13
6ho4gad1d5qo4+zMr3DffZPSPIgvW+xaZOwmx4Q/cF6nad+6dZ0cMSZw/Dpple6SMHFiGEPoOwau
gHmVlMQAtBliqIqJIOdf4Z2BHlAZIzLF0Jw1+/sOgXGtF7R75JQ4CUb1ybDFh6GSD9PORnHeiMd6
4NCZkBI2dbTQtLunV6nmtgKCx+19xAGtIEcwnEmFVga1g+/ILovhX4A4zahaHirkgvAzW8t0bek/
oGysQ5Pl2FBWW7bTHy1FgW3L0etMAbEK6/WVrgzwzymJR1RVhaHl31DLgvpWBJaP8KMsojDq3e4Y
4qB308WJqfn8FaVudI6Sc5U7wKoSyejBIIpk0+3BHQzfPLlBdQ/gQOru7Jj93pwRHfVgaLUVGCtW
HlUXaJNPz9dj4Z8IsOWDX3yVUdMmrjcxiV82rouRDq4pf/qU1lzG3ajrWgvywybpE0LSjP0h8HBU
BQRVMpmllil79Mv3aU/TMVl03bCrtvhpXEWhrS0puveliskUjvXZwoFoV2hW0l7Ql/G1Dboxzi5K
YXFzr/20Zvim7X6EE8qNusneiIzfsuTdDaVUmKd691J3itaB3QZLKoDu4dbCXbDsHe9T/mKirboS
CHBQHA4Iwiqo6a3etNHkOrgi61T0/iihhMlrC7gMzxtvzDr56SdijmdI/sPOPjWorREFWcLgV7w/
d90EcTN6kFcwROwCmmFf3zQcfn8S2xfNd18vAYkSA0QTNe2x2dJv3F6Q1cZ1bB2AipcHKk2jsF2w
X2JtbbWK9RLWEj+4QKXKRyIyIZtg0o9vt6aEta/HkCo8Hm8F/Hnm3i/bzTLxwmu2YJ/pIksof5AD
3AiiD1qDjKLz5D+/fP8X8Dx4s4wLauEC+kuM6JqH0AEdWR1NfUU6bvKpHpLp7z5X2SmcxKoXVYCc
PV40K/1448BYqvRgdFCuF6MCk0iq/U/MCi3q6GqI018K/FTD/B0G7iUaCZ4hkbM7dHxk2DfP4/dV
l4CQpLFlNfdHMN1tUAjhGyj2c70lLiDCG2gbRY64bvEcgKQXNTRgT2TLiB4zM65nSP2a+ZO0+Ljt
5h17Ourcr30HWbkIwXtBRoAcA21SRPmli+1Zu44QK7xpmVNUOEZq53z2yEOJjsdhNiDqzgf7eU6c
gw5WuInd5DUsUSsVXdpe493JpLkzPDlKWjdseCg2I0X5/h8JXaaxAJutWPkejbX/boTgrbRePp+J
kMB/iDBedhzv7mqVOP7vi0k5RSIsK4RYGYgNMYffuf9+Psw9MtG/s1+DaHThxCCogdKCXB3wh8w3
AmTx3NC+h+FaPafJtvH93XihZmK57PFdi2yABEvj8wedxzFDgxCdtwatJhXcDW+7Mct9KF96hVk/
2I2o+zGXzy5iHGsN/Q5vpLPvU7MbaUWx/ch1TNXv+HjaVejjd/CkRxb1oyh0LXzArKDNv3AzSkE5
ObPoJxyWFc+2xde7XABhDvUjTgm8oOFi1PtXWp7XIKzMAKvKD+g9+RVmmeXt5X8wz27RG/fo5GtU
FQdOPnV1L7wVQjEaweeevsBxeZDg4MHPP3DY8b1pU0Oo2y3xMXtKCo6qcdBF0nV0HQjbbn/yaD84
0bPyKeLN2MRM/z2lYznOA+7w9U/mj5AuOfwtXGXP0o25FrHZHSfhnmHQqXKLA1ndrWPmmGpmeylP
077ByMUS/7wBD8fNdFKyTXGJLz5JVxBqd1GZIDbkSz8GdShXo+rbi5emoFBJru6aZhIugtqVQKGq
1TgK2T3sHHH/e0tMIXVH5szrp5pKxcg9K2bqsCtKNUtMlKMFsd+dEMmsbbnGRwA54RwvXG8oUOwv
ERtHaOq6Eo1jniPXela36cM9bniAbOiwgeS243CZxdyXUjtOZK5TugIlshnzgLH2eB9uKHw0M+Q4
lMjUnog6IAEawP8zYE5lKeLAfy9UOf6dJ8sv/4CWcfRIWvfrPdMpRAg/Gzr22qxqd7PpVwg6EGCx
qf56KgfUCLelP6Cm0cuEAMxbJYAuaVVD5tb7Iv1tciWcZpcDwpJHRW9K+uMGGyx5Hy3M98pHmQ4f
fReDz3b1ZGDV1KsQAVVM75iqKexTo589Dd40+r/VLDUFldUWRHW6O+j/s307ZePQ1BYtB7D6kfrY
rex3F6z6NX6SYqrW4o9AGtQvR0XnLyvxRrIkLXajWS+E4P+qjdILUeQMuGsPxpc/dEprhUr7KdLt
eFemzMIByf81vAgHZSU6xUtkxJRLM8df8zobjl60vPn+Lliziqa6Iks4PcjIZaGQW3R0TvXigJnP
qWzqmToehWJvmPeXQPyB6xox9Boqq/D2QnS1CkiaVKOcT8M7vr2ogdPlupmBIL05uiB24mWFJJbo
ELEcX98/M87zFGa57gHHiHce1mKJT5Ya3kBVeg29gTknZhbN0UMsVDagDhudQN8DJXrMvgM/hzI0
QfZie9Fu6b8kuptD2INQtaUR5A4Ww1Y1ajNfcCnhjDwmPaheF6+CoowZ1+3G2IrifaDJmPyOUhi+
J8gjc7BokIeeFfdopaSmTEyJKNVH3rFdY+fSqRrQ5gYKEpqXrk+AjmSM9+M5S2ijEP7odDyO/j4Z
Tpmosrf1B6CWB1J9RaTXiujblQ8dMTL30ooHg7GQEUsNkdj5kCO/ukdV57vmcMyERbnkH0cfw11p
lc7F62rRm35ugYhfUmlDRNZRnGADdKefhwjCAkOc4AcUZzc8U642eNH5wDTZrfZ/kYbcgzJ3YEUk
mCZvVWI6YPf4Bmhg7sTn1H916v1bWUndQkISzmeQaCUv6ec5l8FJnhu8gSP0CJMnHPdcuQTvHnoP
Bwzm1wTZr37LFhLZ2+OiQHy2oPWQC0vEBfBoS5ueQPutbKtm+OEQwy87D4MVQ69t5R6YSvum/n6J
8PL+r1H5So/CWEADuviVBgfRky3u16cJaGDzBiLB7KnARPfPC/bPvaH0AlIP9Y7JC8AydXzQa4p/
bZju87ZFZjrIdfD4CFpd9KSthL5TY0OPJmuDOHK0Jc05EBK5E8GyZ2qVkXn4y2HL8t5ymK9Hqlsj
Srg3RIxv2y3d3rV65fiTxQHIHvV57/rflRCP6IeF6MU4Ko76ATgBUWI3bIgzRWr8MbXPTQpnk84D
Qtv0K+YYVw4CANmWl1w/fkQGIecPWjY514he6GiG1Y4SkekKj7Rvsj/iLg0UCtA/T+LEzwj2/0r4
bSTHGfHXG655wzvSVidEUdoIgSAi3FLwDyuZmSGwTfGc6wjGR0Ut2oRPl9prAMGNWCEZyVDjsJDr
/0obAN3/thkYv3cnQ/f6cX5aYmyc1RViMSc/cJ+styLdrp1XNRr9AU4+usuZ/mOhCqkRleBfwqRS
MaVMAXXtNfA1Wac0cPgon2b9aFgjRrO/SFmdqC0Xji6ZiTBw6lBsqT8Ob1XFn3JvIbq2uPtLRCim
Ds5oFr9vgM4RipFGEJW43pJMs/Wjz2Wi48CQx9LdBM4JyIJLp8fP/FM2i/eEvQHhi+BlVqwvMH93
sGfPWC1OvxBH5gUNcHSM+RYUmg3gBAU0OAGkkY4tDLkDC3D63IWbbv7LtnwNQusu0ZAhjoNpLtop
rVvvm0Qc4ilwCHYEdArP+1tfM9FH+A8y3m3Up0moGzBIm2zaH9K3MpiqOIUp5n9bVm/elhi0+nSN
/KAmmA3nuw9JkKMvOlL9XCo/jGr5TzlBLoHs2U/EEkYuv8d7Eu1XEDCVOAv7M/OXTJK/7PkYE9wV
tXmvMETw7E1k1PvZrGO1XxlPsoOeHwrnn0uJQbJqxBtL1UDWH2HPYEixpcKtn2awzTdXrQuIqG1c
Yz+1Hlhof8d0Yf33XCOxPhHTWStCm4ig5+BQUQmXqfOY+7t2MbA0B049ahL/AfFyH07zpwJe4ity
l/vHnwrRmVpdAfIXkAahEs1AaPJfauqLBh1KMi31uYlJLvFxo1uDxqb3U1KtEIeIKc2fUfKEo9qC
sHHimG9Uf3F26bBcMs/QD+NfiROr6B2v9wjd4DIz55us1Cm9iM9zMvnJiYNBqqvIw2l1aPlNtb/C
DCqwbGfM6cwVymxaTnl1GD8JnQEEQtJrCMHD2+4NtpJEj71b4t85+CLxhVLZjzzP50IGLcKlZ6By
NUFaK2Ue0+rnbeyQt9X1DY/f8dih+D3rmz/uDFzaC4xkWyCeLfjXad0XlIikgQ8cbp5McVQLiVtu
Q5xL5g6rFVFqOZFlMdQh2UUEJavy1uMBurM/UnQJjaUsSQ3LMk/uOJPOj8Vejfl23mYFpQndzvkz
dljQUOGBGmIDYWqEXmOEJyaKcTvVugteyEyju9BjFlahjYMZAIRX3s9H+qymyvkKF4I0UMh6O4Xt
Dq7poFgmA4SNZg8pPsblltUAxbdOfDrvP4F+lofGw7bAWWMHJb/ZzBlSChpfWyvRy14xn8xVc8xB
ASDCseeXmCrs/FmHTa68jyK5DVSc0cbijqr2yQJlYrIxXYI5ZkwfoIGZKMoZofdwaqE7gO2SqaQO
4xelMhzY+RUbPlrg1Y5dQodh2vF3RLZLHaMEivQbyVKtMB4OYuSQncYIrAAyWx9xju5xiGyIFPp3
0/scP1eefG7ICgZgr9MgOtsA/ytXsXAhPMu4OAihke5v0tQcgJ9oY+4HUV61tP+PszAlnV+qWPDP
Wx3yEuGnfAfRqPuYoVVPesV59ILC6vuE8er+v6RhJc5AjwF5sc1EjfA6N+comqnM8qzvmvVdluJ4
Z70q6e6cJ9jXwl0lf3QgrDN1lwa+3unzI8+rW11XUh53aUDCcPveI2hR4TwgQ2TwAc50BObWZeI+
UuVjl86YbFI6E3Yeu/zdOt54lWXAQCGZ1cyltzDpgu5KSCbzLcUhcrm5HbhCNS4rV5Pi2JW/+k2L
6FpdJJX17Y+SzisEF8St2vSENfztyry9OO0Rgxacwn6JDGHA6goyWPAV+lGzUHF06Nc+nvNfuDaq
NEEkl3xxCNkpAAJMGVchJ0WAeEstOWZhB2th9XP5DZnsW6+ePXryL6Z3ur2+AbUfHDFBGT0DzZ9s
a0GCuLe2wUERYUVOTFilKE7MK0lffSVtT+ANcCPg/2WVyyEdkULYNenXvX38eWjmQ3aZ2sMXrRiW
OFQOnxxt5aE0E54RX3PeQ8ZAm+XyNenY4pqF5Xq2836A8n7c+q2/PKpTtTT5d6z3yAKduXsRiDZo
AeJb2AE5kLa/jEU+dvfIWffCxSIzxSraVBGj/W+Dg5bcuGotFoFdgYg1MJGS/tHQdiIKWVwEqsG0
ruZH0y0CI3eAToqxbftOhrQcaH8iUYGqawUZqj2hkkqLlnfRJN/tfSv2Uhswjjq95I2XGEGQA4op
UrqrT+JtIWYpPgZDcluGjG58ovZcum4QINlljfqWG3NcBtuJ5rNi2MKqX1IVrkTjvoHDdaEtfMoV
oup2WhwUKvodBNaqg3WovM3VdUPD1OWHKbkB1Vcb41Pz6+FqhGtiNU5U9e2vg4Kna68qWsuTpAI4
DohQRrCAknRHupJGbsvvvyh5jGk57LjfmoAqYXGqgLTIok36WtsnrqUiZA6SVlj8siTcdFWc0bA5
aYbPqsC+sRRZE3lbK6dFhm+pQuhPUmz4rjzob/CO3I1Niqjycdp/NRexFdQwva5MXoW96on/OFdp
67Ty26VC1LD7kq3UHScvOxW/mx+pisIA2p2OO04+v3zBAfjFc06kx3+fb3u+ZSh4je7+30BT6ywC
z6uI1r4Q6Med+QVjeG0qsJrc5vGtw+W0hd/ElmNfiI2Fq+s1uyM66yOl/qiBa6bPGOljPA0lupEE
hVK5STZiAxAS/bunhgou9q4spusKOnJds9RXBweLcP2/Ox4D5CHa2l270DnNwMXMP720WJgcPAEJ
ZtPqJM70OMhz583DZsOTWyr5KbY/fjINWY3ocX9BlendP9eX1e/IT93TRKbS5Ht3lZBynFix4Rhy
9t1q/q/vZdBm2cwSGavMWeYT5HpLCMJcgzDl3uKin2qnesL0/HMG4+r3RHL0zKT2nNAbXgR2F8e0
cWpj9ivyO/LszAFS9145dwnofy6Z4aFxdhwZY7DRTFxMBfs2JQU9viAar24i3lkmWlfDEBhmyvuy
NAxot47eh8fjhs+mcLwpmH3lNvcw//8XNstCIQGidmM85DUBC2c2t/4MFVfCNWqxh3iYMfngvpyM
WffqJb93OoT7G0HFlkND3QEv0Yhdlzros4L+792j3gIfu0+ndu/2PIpxCHjWDH24VL3KDbdm2yif
QS8rn48fSE+7dZSr7sIX/V1xWn/sJ0QVgMmJ8KlQJn22e2zrE21wbRyv46EN4JnL/xBcJWNQXaWP
yJPA9+dcOTpHT20XRmUHfkp27Hi1+DlrSJiQZ6EQBKWpzRaKGYGJval7i6SUQLITkl+rQqBPysVE
CkYueqvUJqyODwnyxsav2YClG4c2vwmkZd0CUlY4+qv8NF/WwLTX5Gps1h84+F4YqEFX7CX4/QJs
gWG8DpoUBxRJocYxkVb6EKd6YRibXNC7pX+oqDKP2RtddGPOTBp1Az1QVUS8XhnW+juyksLECdT7
8v8/hohYx47KrglYRySrK9uRZE8UtOG/uPYUhMIwIGU2RoKg1VaM95X/ol/gLyiVRdlwPLJPYHfz
WaBFH3BYvahkmtN9WFEODrw8OQ3F/Rx+k0j5gaQz516oS+2/71hofiWmvoi8wep0c/Wh7Z+HaDaV
M7Uy+hjhOZZzcXsbkg7OP1MMBZifFg9eMmT3vY3q7G0QQarJoHwdKHr4DJKg882jPaA5a6smIihG
BI8cdMecUCMPdG0ng1/lytmg00SicMB7/k9Njm5Dsly6R+3e1/EtewII/3yOBd5g31K2sfT7AMc9
5BPd4PQj8x6jLxyt+5neBn8ruLJLTkTUU6q3sZ+nwZINNvObtDKefbtcIQMKBkWDGve4U817Vop1
ErQ3eIm1P7e9FUPqyl4Fio5UhcFNCXfQtB1jrGsfSn6ccdgYhK4PwlfIUd7r99FxLFbtzpii6BXC
xHS7mufA4fUMYGHW0psEq+WiF5ByFgzz4BsD2UJIG32d3jUq11pw9rWAzg/TKLVQmRWT9Pp1WPIX
JmEDtEJm7lsKg+/ZGX4QaFqtAG4uOPq6hblY3CkrME2ioLUPslinMj5Ptc7ObfRPnE6HMiTf9p4E
d2iBznVAxDV4/v0d7jsfRVXNz8uv9mPTcQoKlFHKYR/fgqtAqxewqhKwd+ydKocKj1hLKnG1ROIn
pYFRiA8LDrBic27V4DfsxHNmo1RkuOyrjrOHPzNrv/owfiMkVM1vB5tIyteslvEn447nGHO07ak0
EbAOjOj0dxrtXUlt8tM6r8L8Y8r1Ia+HM3oSD1TLVclwBWUpgKUzlrq0suOnXJGFKRvQP+5T3j/J
YxGzLQ43o9p1nvCQtoqJJsywbJ/IlfqsBtTQB+emOfREai55pTfniYwrZVSV91qO2szUw/AXF6Xu
MDnAoALZiHG9zMcDw0R+aemchTaHlVcwo380BnlzxXroFuCsrd/RLte49IEH0utPOf663DhKrspL
onn8F9KQ2Lx97AIgkKIuPb32DlXbN2yaItKr9N6F9R3PrDdus+S7mN6JvPRh/tK044Amxm2lV6xD
knNTiru1aGK9t1o2Z3cAcqKITy0+TkvzFwiDCmwyRePPMCrFP1lT1W9Obg1gATtBXLEL55mauI5X
2VSbAnt8uDEYorJM9nE2eidhMX3ZOSgsL7MrmtygILyD1X2f6s+0S+jlALzSgMk227tcJdAHwpYO
i7rQPcjYAIEPbttpfWrby5jsjjsxkEbMieRoUzXN7yQAS6x+lxWCC9bGEhb7lFc8HcPCDFo61tDk
8FlDmeVFreOGfpP5jw6BoEXzbZGeUuU0Qu63m0AFwVYgsWLDcDvmUqp8ELF/PE8IHlUiyen7KQ3X
raR96Sp87qrnlWitLv4EVF12I0n33TOWLePMqy6lN/dVoxLULABU362YfAWkIRiIlO7F6Gpuhvv1
aaaxVPAJczKunb4E0p4ziHj8AlXJl430VO1kSDu9KrW+rNuOvIY9xC4WvKf+xgsby3c3uZY6o5+I
xcSOfS6Vo83OvDvA2xgHB3vWrw7c15WaNlez8itH4bpwGsryVgILi4v5/LPtymkeU6fGys6hta/D
OsDsaVfa/LqwrJwczVbjw4L9cvFacDGLOvUDFJ8IRlUFmi8VEJXhdjvwRYVii4qsmaUfgBf8QL/R
w+D1jfzS7w/uSSt0OFdcujdT9It3L4eiAqH+bpyBW8ExjYJIYFCuMONprgAhlHJDKCc1zHaWpO7r
gAoRhThV/pPyrEkFMvEN7eUFasf7AQ+ltbFtePfNl3Qz1JOitSQVGmF1SqIIBrKCAkXclOafiiVh
WkN9NC6JFnvKwmh7k0obvbVqGAXZ0N5ZQHLCHt3zZku0JQk1PLy0l6e7xnxKOGDaF9d28Ukg88e4
9WX6MnFlhFhSIDA13sOouXzhzq4M3bhtKSwD2JbH9QeElJtoECyAS5GW9ARYnGloQ7hi1Jtg4kFX
r0wRwQtDzvMWyFzm55jW5AP0PH+cVyfBDoU8ynaIgjG/JfEExaRd2Ti1Vw1WlLFhNAFoAYQcWh+B
KYAtVqx6BfBMdVc1Vxi1Sr9Yr95ErzhhMyIMIWTX7nyGqOAwJYi1sULI/uNCrSqaPsHClsas/3OQ
sBuLsXBUSDcjl1bTKgzK923sCxlMBhTfP62BH9Bza5l7rAP+lnGbRS27MzQomlr+DwyNYzHXQ2Nu
54BSR6pvjBkemmKkkZLtMLzi4eKcGmlSYCi9ExuB/MDHiRfXV4TueWK7iAH8LYj558O7RYiVZ/Y4
RXDene6RMDnL+2QTIa6Dag6bET7SSxvM0QXth5ztZRytTlkJCDH3WxCy7yhArU+jw4sPMPEj8n4j
HQWkXtn8OA4EAFBRW0RKZ1qvntGgxh3TNgQZiVhqolnGSUbmcxDqgLGZfJbUsdteT9H6wlXuzs7A
UP1lkP+NeKvW2ZNiW/ctrOHfi4Y+9sD6vY039tiowFjC15yHK/VshvP1vNtBQF3SQGMsYHZVdJgy
IYcY6HNvar9zmCfIPPlum4KXtWNv7b+wDBXJvj/jgQdyCTvOA3mmrEyNu+HZw80sfehP+Cajy7oJ
SyFE1I/7fFNyC2aPzWEONRfKz6f+Qm4gNbEFy6IOPZsO2mxi2JgcOP1RV/HGw4BJq+SWlOOmbvK1
Pf/PL+pvAhZnvbcbixPgM2w6W7nwxcaQaDYBYlkwl7p2tMANoIDXLNsaC4pvdaF/KoHkGjy8oCcW
AtETEenT73dlm0Ae3W/o7XvzNMJO9edNBxvtkUKBb2U4tpIIPe3QIk1r+Zq3uSxdxViawk8FARsk
Ewaxfp8/fgywrKCCqn9q8B4irxvnwur41YgvtMrP4buf/rpaQEkm3VJ1YleM7xtZ9oykj8EJaK5i
2LgVY3Itkp9z1otDqHQ/NaWmhVkDGfAqBzEHOd1TRZfhkpEQbJ3sEL0/J2lTMMpEEel2M7GIvZd6
hA96OTasjhKzgPCQYa+1ZLFf7gxmHTZNMO+4pFN6mdLwUs/7D1ZiDDGsQ+c632HbvIBUAAYlYzH/
3f/9p8WCcCxtTjrS+0CUAl44MfqJQkG72KA5+mdqRqPEvaTe5gvla0Z6Pn3iE7LLBMPGbS3jWkpG
+rfIL5vZGIqKIxJSrzof50Oki/lxdqUG6X1YzcrvStgmgpZo/FRdiCOsg2tz9b4U5LC9jcFUwqH3
laHZ3t5f6KmCFRBKahMu8yBeystn/1lJ0n96jJNGmQSangjD4LitCTztyRP2ALT19wQBjuT+n6lp
SCSOsveQ1s+1ox9Cery1V2u10uqFCLmvosa1n8i67+PuXUssA2Zk02qV1bj7HyOHdfHS+zz67DP0
fVj82IxkIYxAiKB+nMNl5jG5X93jpm0kM8JEAggBxAg75bPLt7cIQRjbGdKGfJOSQzV7SMRSwrf0
F9KRoHdMbGd1x/gW0D+Dhq0rDNUt7ckbyhvkMfjnGOsxXlBJHmddHe18qvmXUmRZLQ7E9X+Er4zc
/tCwkDGQyBgy5Wrwxm37PSnI6AhoUphSQYjZ44Lu8PM0gEpMImV3zQNsoeWcaEwQ51HuYliy4NPI
UxqxXE8Up9O1+v4A00iHv8s8nRTlySE2rESNFVikNApdn4iQEYhdVk0fGmBzV9gzgrv8/y7wMBYF
uamCy5Jn8POLRDsyUbmBTgLSuNeOri9yxFY86tbrfUwnJZ+gsiT5jA1j5qRaHlkXHaftQpJBpjGf
igjP8WSHESuxvQWkZsV/vBL79jKRtWyhsZjBUxiA/rLbUEWwx/T9+dBr1nqvt2SHuoa0vv8YtUhx
apbzvs13iFgRODjM6mNSKswvMyg4nY+TEGiOzjbrokLxC3IoKv9CE6S4dfwLT6VwFziWeEc0C+BB
NCDAPaXidGMqeWe2VOMq5fvEO2eR0hmjfdzBeZ1VgxUYlc0wCIDIimEu0DCFbej0hr6guDvOPebD
5Jx2HpgzZvwIh8hIvY2sgEPA2nCvKU3rr3+54vqmFepQTwZlauZvxUr/prs3BW0J3LrubM9u5h3x
+h0SMddggjbMtHD2ZWi7TaeflSN44ImMzHl2Fd4aHDp16VUgk373fJzwULU3+ZXwNIvSEZL9NDDG
Pgo0VHcFG0D3xpHqLRm/Ya76oK7R1w5GlrFP3EjvuZVZQchYTJLGk9sbd1tFfLROVc5q6J9OVXeH
vI6RyR9438Miaqf/pYye0Ypi7gtPlUIuJYsmQxBTADZqw4ejfZpDak/gDlTE27JMJ5/cxk2kYX5d
yd4ZDCQQ0+Kk/a6h3UNEnFT1DtwcMJHq3sLQpKJGHCCwt5UsdLIKqQueLERbozfZYiKgro7ut027
NMBDYrGkf6ScvCNEBFSSLapAYfz+Cd7j76DQkkChL3tTPzAcGRrkrqn0o547ySPqMwyO28Nx+Tyc
Wh8bWv3D5DGWD9AXiWg2e7I645/JG8lYGMM0gZsPpXwM3vfAmJl/4CceCyD1XgtMTRsX8mTRYJIi
aEWWVpa5u6rCqE917HKAu/3+7tCMZeiwnDgDrwmfu/aHvR/f26efbXNdpEHYBYwcyuZXr4hNkdZa
QXyfWOINxBZmI6BN8wKUaCxj2nRIVbIlR1hR9D17HZQzx2JvCwMXMloT5D7vHxRlF+XHEsQBXWU0
C7jP31dALrvuBS5VdFbIKfeiYVGOX7Fc+9Y8fdT+Znqsj8JAt81BW0CKACvMjBUb3Geqy8yuiRVR
uY8C0gIbUnSO47rNdG8HOLXiUvcXv151S7qZE5k2Isj09nrJSbkdaTiEmvS8XMQ/clSXkbphrGib
/IA6/JCAH3MrBFIOC0dvbFfst+S+zajKjQaQqm0iGfN80PcOI1W5uctSyFwjhVYxzfIJhXiYNdGp
sEyv40Ag/LJZx/rDLh5fVEvanTYmsnaHlvQLPg2DpLUvclO1PNPtE3rSxVdNcD89I0YwtUe3PCiF
J7RRmutObURjv3WrXfa7z/Z8aFZuC+330BxURAwip/+ME1xYz33hvsI4Aycfjl2WVF5gCTneNYbX
JUQBEcb6Q2OME/lfkAkkML1uFEP9hXLhmNmaspyvp9Zxdq8+q8dQg33ed9CWDSJfVKoBaycguFt+
7gQYoI6NOIQoomHXOpIYd5cs72Szh5uziqGEGViY2NgntAky4RdbP1CUaihmF6KBJ3q9HQu89946
MTIL1Zps6U3xqssS7yR/MKEpCDKwbj+93CA5gON8LqRwWDDktkUQl/+G7y1mKzqQU7AKopMP1Wfu
ro0Zx83IWkg02LyLz2y4tmb3RhwXh7kUNfGvzru3cMf81bU7uINm88uATZP2DQtl3xP8CLJRBezR
+jdN5yingyEGkpvUxEEbl70wtrHAXJojR6mRD+dno1SLHDFoow2YnP/pRiqymagDQ+U/XvXeVVyh
ENy9+I3DngT+hgV5GcNVyMPRXiAZjsZD4Jfq9tKt/NzFF53wgfKwhKCnuCUMfPcVwhqUMG7IJflQ
DlKZrSc/4X+x8Iqi0ayzVmEDNao9Im5NWUhr2UHPc4BGCXvuBUxF/JXoKBw20bQVFVXg7OcRhQlB
CYdGlp1HnrJWYKAJK5EItye4sFi9P2P514Dwp0Y74xzHETTL5OqN+nLHWeNzors7Kqqb5PM1lcdi
bwpWqoOB9aHUGv0MrwEObGmTrn3pXrCDWQhXfT27MBh5zc29vTpPnhqT2wOCcyPOHh/QFejccj8z
PTAknu7edusClBPzRXtXC8ZbBho64txV069g2tvZuoZr8FT4YhNci2C2FvNskhlq6lWb30MebPQc
0c7tLpjEt38RKU0yl+7l5psvS51ao6Bwr0DGbuzBciBzYHZXvwBrepDsKoB73NpMw1vPuFLJWDlM
DwJv2XKXR58R4rzjStbQKfKa4Tm1rUH7+99vmO8wWnW8UTt78z3y7QmlILw8+J8sHdrdK2sb26DZ
Cs+7KRQNjDwG9ONzCbZmcSLmP5yfFPjZVfCinbbEFSFLK47YiMF9YWlha/IjHL/fvmIGc7osKz/x
HRfTpnulcwaJMsgqc68qXlnR647GnMiGcsS61N0f4vgT5oPpsvxIA8bJCFlwB7PbVsz5E+rLfUCz
vgzkQ9o8psTgfCVaNnwE+NzT0bb8ZdNL//pcFfJ0/heYr8JrMMVUDFnzHb6zGLKAnTykKDdl/VYR
5HFVjAqN/VT9wIqsDvWJElcj7LtLEtnpljj+YT42Oq5kjt3PBzISq8UTimIq0oEBfQrpgvYOmvjs
snX+WhugeMDY32DJ7IddeVdxvzX5rdaCE1tObXtws7KUq3Tz459YtNaIKuBUM3laOCbS6k7EgRx3
s0FL8PuprMPAzfIQ0KpyV691up/ehzDRjSauF9dwmQDLz/Cr98rmCinG+lCMZSV9CpE1k5HtB5BL
c/yoCeo0zR1tcHGt5YHUQpg7Sp1MLuey6tnkOm5F7cND09gsdqZ4h8E3meEiokFUgfQivCcIf93o
sFdELTCTk06ZLTjB5ZjjAw0KgiONXwBB3XlTkndl7GlgLOTORgcSm74nI4M2S9A5GDhGddo//Clp
cJFis9bAHJu+bBmGnfvQaPdVqVSNzmHPBSlrkdRs8MlVWOtoJFqc0q+mT85zVv6V0O8T9kyxGj+J
yUpMNSfSA7Hec2kG/Ewe124MXEfUp3UcYR4ra5kzji+7RAGEJnw72p96aGkQsLZnHYFmb4ty+vCZ
6f0n1uVsKh1cCxrcI3U7y+SKH/05M+Qud2mPIdjbLwSq2MgeoDRUxmuLUx24kEz4hkAEWik6z6Xi
hZ1Y8atiQo3OT8TEbPArGtv5gCYj8z1fDc1jEdHjpNg88lyaXsHuIIHLqBYM9MLa0WBaP87gvQM7
APcehmpF1EEaJ6e2U5s0Ek1Cy3EmKBUfuDzuC3JRkUN2mIeRQ+ZiBjlJhMv5e1CzB0aQS2wogyWG
jwVRWq5v1NjxU1fE/P8NC2CEuQ+0fcJdbPxWn6i35DdK4gTadPkD1BYn6X8+edKDt8DR7Ear9NG/
/BFvvBJ5EBEIJZNNviiGMRRAmO9M/a1hHdLDMWGCv2mHagelrtP6YR0ghb1ukMPmAcNvYxMojv2l
i3tubXF9mebLCvjIYTiBrelLTwyy6ZnbuFg/cZ8j8VBzwoDpi2dnhjysiVw02QjRjXYlDetwJM4N
8vGA0zyqD2xq78Zu13YJpnGRgFUxbCVc2/Aw6RwfxQS2SbflxLipkx0V0co9pilfbr+Koat4zMfo
/jBUILcuTuLStil0yT9FLEjOkjHQ68zcuuEer6NIxU/+zo19cIrsgQgGk2at3s9TKMHgYKMY5lin
Rd04bp8U7A90jFjruXMTmYoRGRlWy9AKYeSiF4QuX3MQjgJt1kFQBDKR2iaYqeWlq9bKIASECG//
SJhHgliwoUeYUC42CkoR7uAYFAvwBYE8hCGezto0olvlBe25oyorkJ+aUZ+URq1YcYiT8wJRSNqG
Ot2uC21hXa4IleeEXo5a7O/kVHEhgpho2N0i3k5kT7N1xjn8tB5IyUphBqP8DjYJCJGvWsnNjTPZ
mw18kHxi/RbftaA0RyPbY5L259zDABAcUya4MrRas3EIuPmjODJxpODoM6wGjcKomSeoms6Hq3mM
fHMIi6Tmbri9uDPfR0sDC0KXk+c0f1Gaz6T2uGjMuR/5eIERbJx65ZfQgm0dR9xEWdAt8UORI1hX
UwnpsnYLjWVJW798wo4PCbU/vsAconOUzb4BaU2+Loa/iDzIHhSbJRKHUajNJtyvqaI8akpu4sb1
mzEgA3Gfjzo/ANAsg1KHU3JoAeoHp8eXYokISTZdeyoHZycvK44PEz8wy3/SzDZop2FyBBKtHgVw
FXTOR/wXqjo0Z081QrEz9/Tr5v1m/q27wfW83RUcridyRke6exNuOw4nUfvRaOMfoC+6asypsxgb
cu1iUbnuQ2KWFZ2qkQsFxir7f2JYor2CdkR9F48Xk94/VprpeU9bJs+AclR8fiZC3hsFE7+KAOBg
6aFRG01tX9Uz8yAimkvG0KQpp2GAKv/No0hrwmI56eTS8XKyRsYlJllagXmjPI33D7EDUXTXga27
XgsLIJSM8S7ZoLlTesLaqa63KlgV5YCpx0VzFUB6jETslEZwoQGAcEMMmwu3/VQeIHLp/7NR36P3
p0g4TdRzqyEq9Gy2L4S6LJ9DHZqBh36FcCU12qn/otWT4OtEfCQonEUWIRdzN8eG8KZriU3OxrjU
FlAtsE6vnY6fHI1BachdSXtVmoSBK1MR0YG9MV3VjbHH2m0pKqI/7gtVk71ownlZ2T1o+8OYuB9k
v0qxGwBQKaqCq2DyU0C5lzkXG68QMekCotUe4f+PmQBdRfqJgFMNmNCXsG9m9s3ZjvEvhJaXr7hN
1VzgpH8LebNYB0wrmjhweemRbb8kF/AVtzeUhgFq9L2VjlMMJbMt8RGARo9XRpmeX7m6UCkodKoE
pT3uQm6RMPdAcNKAM1flT27wB6nV3d3OMD8wiaAGv7VtS6GZn7fELlDtHX8/2kwkzyif39tV/KGV
RjcXk/N/hWZLpjNatwL3tY8R3kglElolghMAAb08j+fm8MTUhvnY90RRQN3QzTYaZYy7dWw0SQ0T
Q+qnoIzDszueUF6wASAT0ope/1Sg55RQC2a6Dq0ICCHbmKMbS+wAxVJHYLz0Yuh06/bCFCCPb0i0
DHFEaxJUSE6GMsgPNOrs3funnngYqNh4h1NzcniZc1xTeNBiP6RmyFjIpNXKs2BbpdXwy9FfmPV8
tFj16lFbGfASPVEaQesKmFZBkEtsdNoSWvWU+KtwjHRG8QlPBww2FFGYBga+7sSVdAgyt0fCVdH3
j74B4OaGIwmNR8LtNMsJVxnjRqB5KeIDsUn8S1G0JWQ5rTFvUJZQnt8APRet9P5KEoxgBDgLnua8
v59/eMZzd6MAtwqqWMHukqTpFo8XhzU+rfL8FB/BD0quonFAXvQCUzNGtTPlmP3ijvhhZc0uvmxP
NyDIA81/tcInnBgWhQVz5MdzJsJysp40wz0z7RYvo0DYlP7xCJsGufcYHWzuyHHMZ0xFTNngwfT+
fhVdEnXa04DtWr/d8+2Z3iH6KA/kFdIN0TmQXgVQ+uhi5MadeH1KAA/vbtN53YdIxOe0dssll8Wb
jTzDHZvYFeeifrIf0UvzVPUoT2YZokVH8vSOkZofWks+i9DQY0ixSWFqj1nGznAcnqRTbepf6REy
GkINZ5BZC3PdBlFqBtjfA7hL+uch7hQMmRIkVg5DQO0SVSwnVKUUAjhb/ZLsEptWh0a+fsKEco97
b2w7V1RCnH0BcKiYOsF3gSrWze6Ie4NsIGIS5T2VzQQnnA/ki0q5iKZbTWxfC7ZxOuhxYkFBgTGR
aZif6s9q19UQnxG8AkmrjK71YEwgTF44mjD++IJlcWddg6kCMMpw3BiyCawWGnqZ8VIZ4kwMAKFj
Vmns2RO4O4A/9iT1uPoP1uL8tqSSyzgEknYamW3Tquw2/M/oeU1eUV7KE/C5Xsd9F2F/Wrzp/Mg7
Mg6FFNuwdFS8ngYq56xPZud9gLpE9vFvqM3JzHZ7Mjkr93G+yzDbK/Ye4HHTJpnbVvg77qkmaUBY
6ZDtCkjymRdTiA+oZHPO58Mm/AH9MQD5tjG/66qrzkKk+PVguqJ4r4Kzkbswa908zggJixEGpILs
vQtZIanTSf53w/L7V56fYv3J1ETqtT6H8fVqAN4qLTYU9a3fL0mCN+RNg5xVKr77Jmit9grBI2Vg
gvbX1u9O4lHyl4CK0z+lB21roMNQ2UaVgD/GnY4RMiypqVp3c1XDO/tCXWG6lXw43pMJGVn8r8ha
IxmPKdt6JgfMti+LQO/HBDXullkKoWDTwGLXtdrzl5/QeBkQW/BLUYzHdlikA+iISO6F1jzaIq/K
02pZSZOhfL/zCGz3rCFoNI3Lse1FgzErmZfNzM+Re0Cecryczdy36tYchoYQirLMJZFs1HnfErd+
Y+QaGLIr677B7NlWeact1RADRbQ/43bQjd4OdgWGZugoRqWj88htH6qPdJu0g2y5el7H1hBA0frx
BDBoFO3rDgGvwJ6sxNsYlaPDQd+tvP7bL2uGOHvn7yw6wxLBaBvTgumDNNzK6Qy5fHICSR4DPbPq
/RAr/CYn4newefpyqEhLcwQn/vJ5WujxIiu5JcfsdO3EzQsV6Zme+02CNqoFIFik0uif32XMDzaC
wBFbpV6mCYxSu/EvaLB/IP94/WKOZyUUEyJlAfcj46unC4LG36LUCryK5lciaSWvFZwMM/9ThIuU
lwDYMqHYTvLRPyi4sYIHsjcKuhS8D5FBsoI8oc8iroR6uF4U/QkkuH2RVOT+SZ07dp6hcjyWZQ8K
yIv/BBYOEKOcZ426RFAsoLGsOU/Le0bvktSD5wToMpupB8qiqo6n4rLMIhpysczi0MeRmqv44RfF
z3Km3M60Cjch2gvbVdF+UMMLgOvvi9HvFZEv7+x7ORf93DHGOK4pjAxv5zHgbGIOvn6t4ZJE7MO2
p6WqvXvxz75Lp7Ib8bi4HZCggYcXmYwDQRO8ujbwc4KwrKK2D8poKadVTaosinB5W+BZO3tMe9fS
bigenUeEOzoHwIZL+T9bKMa2N3a/YPv0tTCD5fKcGCrbi2w2l2M2+7B1XC3BKXJ/EDj9OJL1S+/2
LbhwR94FoIEJiOK2+JqYyGFlhn41rduTJNdc06qpjjj4oYS0wkLndUiWBZIUDke/i6Ql1mG2yEQQ
hLc0YNom1Fy4sjRWsBEklExTLrFoQBisEcUmF4MMDGqITK0dv7Q0z15EFhOA/L7/f66Rh214pl9j
tGJSQkG4VxE99uWKshV6kYrHAAZRsciKUdVdN19a5cTpJ3FXQjcwiHJfv+oJqDp06Ci1qtAKw0Up
LSatv2rPGQU+ntFvq+8qwxSaTUGzGktEUDJAxnNlkC05OQI92UsJ5mWBGFvCHud2O/P/it0TBh2p
31L5DRd/0D47HPTSUF4V5vvMUXalxRxCIgkgQ1xvahxPIjxE/DIVQ6dm4AuUzoUQ4Jik7Jiqs+OT
oPWtzPkln1Q9HPE1hBPXGLrDvQB+OCssWbrpQMgv+gRK5i77t3/tXO/8lHN8km/Byzbr+Me0p7LU
wKzv1klq68OAdB42VW9Iedeu+PVRri9g5oqBupWHgtXcI2YeAg0+0ywjmX/0ORQA21kdOCsCpCG0
tRJBgTxpiEmiLtv2YA7gd86t+MtOQsqAvP0vQUxW3gk0WINWTSKAxHN0YLzwepe6VLComMQgxv19
ubdmeLCaWoO1p86+IlXK/e3RkK0wZLyrUrhIOb9NFi+vsOhQ122FdEAjYwXLZSwxxfbj77SQ/rY+
fuOmaYzLam70a9pmNB/ntD+G4n31X3a2kRhv0WTZU9pbW5ZXLJ7HN/uYxsB6JqzW7daIUlXzF3e8
6BLnSG4yI9dvBOKpFv9CmiZigwXRFLp0NfD2fcv3qJtf/1Cp2AO9MiTneS73WJ4ucEhQ9Mk9e7jI
kpLAmkXN61LeydQq5O4Xgcv/dG3bbgYRcoAWfHJM3sV+s9/DErUpmG1qEUR+yuDxQKX6lo+4zIFV
xkccL6rYg19thI9DHccsoCD6yVGcs6xNDHerG22IB8fePMX6wKsrvfXDwE2ecZdqVzyAre3I/nfA
2J5+DFigFcgVfmn29l6k4i7j9KL2Ro3UK7ny031n13aC9Jw3IxhFwXlJ+wTSuwghdp9uMPhX6gyg
hArp/ZUsJqQwkYG0asnP2LWTPYTWuNBgENdETSLjV8hym0sZdOVrVNCinUvYgmH9BCuYVc/d8Ryl
Uvg+Uwq5ZtDTzzoPdMlN8EoBpI49zApXKZi7lJ9YgATLaPSvURBTZhoZeSPHpiYjLgr35Y16Uihq
y+EeE5JmkkyDbi0tBsS5I2PsnYW15Xoo8oSho2MKDb71+tURtbl2DLnG3bulzqiO5JXJX+Dj8tOC
lqprIZgT2YlO2r6XH6GDvNNECDzCNKJz78bCJnYiPNQc1pI1No7CJ1xpnxNqaJ9+MlFq2nH3Z/YS
+f8r0wBT/ARBxsZlsyKumnafxhqNHFgY/EexCRljXa4nNFE+eu+OYWhtV6i2UZ532BEGtcWcSl9j
zBI3rlp9bmLvGstQMY9xdmkA4E3kqn8xC5aeCLX+mtEJyt2nOZb9Poph9jgoU1/ZalK57dFyDECt
5R3Z1EtxLX6ioqqwRiLN3up5bjwVfAXCjeoDICZwdWmBlP0OwazHE1vsFlasd+KhfDJZy6VuSwwq
T0p9I8nD+LDSz1aFKUbhqF/GJ4H3Yn+uSqOOCFJ5pFpgRSfMQbVQLG86XC1k+mmPpVac7ievQmjT
7l4Gvq0/xiG32mLomswkkYIiTK5z9CkoKCGANyT8kUAhLVDpPPZMve9hjr36zGsW7fbBVAfHk/zC
+vHLrpJ8eO90JPDWLpdIwVKwOi40hExIw/dHqAgYvzHl5240zpRuhL7FRe7VwzSGal9tx3OC4SFQ
SLjzeI6TOjsQ6bCZXc6xqiWAiBEjAhoVCHXwII78BiyADbAvbwofQuwMCus8P78Gj4ZB2ZKsp5ce
i83YVIMOhX4NcmcT9gJlRWLI4WmeOPCVchQVZLzwqDrFF6V9R2oSwwev7+mz1kwinYb3nWrQfgXq
i17eblV9y/JwWkFApNfezh/yzKoKD9cAGqO2P4g/elot2vSQt5zFhJARDR7noQYeFNUQzpOcmmsu
dWhH3Rx1l4rsipIs8GTS/4yUUOF5+jC6/r74fMIhqmmjeVmhxLBSBJmTY7ItxhfYcW/tV0Zrewu9
B4gCWm37ybuDXZFjSRu3+08HtND7ExuiexlFovJSwaOhgM6ax2pcEvk7Jt7G/bpn/yYkAZY4qkNa
Na2pKlm15oI/W9RS8up8ieIWkpyA/qUK2FFwHsQ/ttgpsLB/3Bkrk8ZW7bNDiDwiNaiYJwP3EAvh
e4wcebq0mdBCNqChvN+x2HPgTcEW6Ae0fT3hpQCQVfTQgC9vL/OPQT5Wfrmyi7vzu8PreoM40DBg
D+Ucp3L53hJHL2xspYW/pYrxEEk/245Nqrlgmb2BT8YqAnGnnhuBMd/CJNmcey+3HsbO9kLAfAr4
keFLeVCh/aX4pn0k29Q8q6bp0nLM2+9aKMp5+aYwDmjoBKMrNOtMJgtJZ7UslIEywJbU1EIWJu2R
XsMNBGFd1pMwzPNJLMl+MgRT3l78gbdAa67/FrmXgdNVRQCJc+U13V31po5H1J51Wpwb8sJDaMuH
36xWd68btNn2qRUBS2sCibvFlaUW+OpWyWw7lkQeMGSzAz/TRjdZQOTPD8zNIf4dUonZL64+VteN
jXMlHjJ+zqwpg+TalH7IPZ4PFnlNBQoy9KMDenm7rpEZVrVaZi5yTwtqhiNAT8AGDZar6ljEi/xY
2CbgMgi91C5KkdYUgmGPjOxTrPOr3x5X53FZ/0dvjobTIBCy58hCHqAIKEGnkDaBGVIdss/wlhKp
q7nKIYKsbhbdJ4R997N8n4Xp9GSYz2twxI73s+OziuJRdUgkqagz0bKcrLdSHnwekjXtwRebk2HK
eLlcofEdDvKn6w6bd8jlkBseLWLbPp74vwtApHPVbu5OSeZFS2I+4jX4lgISW5Iuenw20Uh9TwO9
28ZpFwUzbyalaUMli9HevuJNM+i53UmvNV58WNH8oviY9nnWNnwYUGz6dU0ZFtvBH+b4dT2ntuAa
eprhU3fGodOt7VkHFG3R8293+KCj6qeXTAM9eYaiAaAwo7BG9ZSoXe74Bs+UtacG2H3vAi2QgtZ9
htEKcgH8dyMcpDMU1jQF93DXP7glSc3PvwiunaPjoYB84udincDV0a8+Z3pl+wnHqHkQraDhQ8P0
jmnJDk9J9nwZnMIZH9FwylEHRjbl0Tr6BwbkhYNMrCTpBzcRFZe2RMfd/KTQgapZwMK7H96d1X2x
Oa18xv9cVUGt2mYKh59El0Mjf19m3IGwb5PJaZTue3FgKRCnHpQQSgK16f1JDFFnZe9jIkOhojlG
5w+FhuHR2gPn7eS8lrd37tOQyo4q0+4uzWH8omdR7KkS+kdthx8GHb8hMhxCaGcxCXrcmLjGgaSa
PnhP05wNXAvvNsTTQJPF3MrAAVEsX9mEV2lGX5pV6BcmkhmxBDXcX8btu7hj/mfEPLeA0Q1TE0p+
voKl9akbzEXmk8kQlwgcX3/VGR8qqjwd70ebePQKMoJgyENQtzaEICd7aiKqGVgB2P5w2nODwzY+
2ugGmr2/UmOuz91J/3N9H1CI50N+Q2gxSSxRo2bzfprznDY2ugyT9D5vj78zGH1ILpel+oYcQthh
99Z7HtR9KQP2/EgjY44yVqVz6dBS1JoslNLMLCQI+TU4/gDdhcuXo9eFVLFGD/lwIrW1dmSoIiBh
6DXACurBuTZEYnPl2l+2fCEZzUtB3AwuV0f22oxvGBbzwLnMjbi/cApxBs7GM5VKxq1KOV7DBzQz
pugRW3cbtSMIv5Y0c+uOR8gS/f8WThoqoe0zUJ69msrd3OazGSydfghWb26zyUZuU3X200Kp2ft/
t0yaJ19bBDWfh/aFjUZU+bmxIb3OAhy4k+O+gh8qTexLQBrqg+gXYKMYVnXI91msDoFDP3m4TmqR
u2mtXXNptooab5kAKySI3xiPXs+vQTuD52l7VWPOJnmFLdoM8N3EOfgJrxP59ivquJ3IM9OpUaXF
UHP1azWz5mE+BvK22CbYK2tcB+4YaNSCTnYegy35aVK43r0Cv06TCgzL1XDEtVBUAVY43nyMlNui
uor0bDQPDptMvIjYqVFgn5P6RzIJlC8D0XUxLJII9EBZ5j9YmAC9sUc0G/e8gOq8li0rmJHEgigf
ZMzvSl8QDxBRgoAF1Q7ov4u66IZ2bn4WLSK7D/TfGvAX8XewPjSgvLOetgyIB0X3F9QqAbAbGRrq
nxd1uCgpeyfOsfLSLLMcZsUA03sw8QYzDmtIWxNAa3to9CVMjdB9lTCCoRmxSWtMdTXBeS2NftYe
b5gG0kwcW+sXDjy7ij+7M2hKqKhn6vUCgISsTEJiV7iqrMVlojQ2sipGfA9RsZTHTDus8n80UHAv
FgpO8Z26ikRrp3dsPQYy9JkYNlIViTED4/Fkp1n1oWfEy4TNH6adsh6vJ2N2ZB+bNx4Ir6Wt9RuG
jqcUk+WjCm5CX5YJvrkFLE9oXIZbGxSD+7AvHMC/fbR9JXjRJpJoo3/oSEURHYraz47gU/mIV3Jt
22/7Exu1fz1DQF2Quc6kGyKaSW4x/NL821cHIq9wuWdc/6exW6L9uL3MlbM7yLMhkimR5UyAX+Sd
ldYLR7jVFCp7S5mjl7WfOG9HiKsA1/TNjP09rhriRqUPqXQFBNnBiigLrP4TWcpFNzNccfP4zTbV
Xpbk/J1jFIfFQwgqDE89FZxgRwCIR/fwbpEY3qKalLee65lBQwnsVerj1/E4VArM92T6djX55Hkg
jiybectNOG5PscnZzqurDx0nh6+AM9w16MSQLn5oC+naZSXMc15X+zltFLiT5MjVwdgvH02xqSXa
13j2zfz+F6eY8ggMekggQ7UFiCcrrEMyQdfJ+IcOcuN4Tu36N1MxWJtUP7EDRz7X+6yW1Ihquish
aIlLz0vz42MsQUf3XacYl0EIkYKXZkQXnviFpRKM76f4MBPr8EZnXuaH0MBo6aU0AIOrWvn+Ln4E
598XA7Kecqw+KaCVT5XNLdByRQrNokpbOPCz4V0yJsTDmSGdzpPentnijUw/wJhWzh5pLbgLEVpb
defgPYvmkA5C/8OFEHucBDuoHQWncb0ZbeZrJ2fACrMZ3qU7iQHF1c5t89TdqwmHX6lF1N+St4gC
VV3ZvJw/W/+Vt+IwkLFn41ylLz2+wgCA/5gOnvF3zWc6diMEj14YGC42syWQ63b+QEJQgTbQz0i4
D19Ks8L+RIz1hfp2NOoxVyCGu33DLnek3uk8M3ZbtZ42p4jcQ3eDWbhvof3CP5stpJt0MbWr9/CP
ikggEkcK2C2KbJwuQFkLvuEkZeH7s+eaokkECdcQWnxySMaSYrgIbVLg9hZ6bF+2uvz7ROHRn2mn
UQ9oqVG2ibcg44NQeMLu8ZAVIyXEBr6xY6YWSQsy9sRZAeh6oVQcWTNhuiF4ypUAYmGTwMR8NVYa
v0/SP6prCaZYPxX0D6kzzjT13c2LAUhtCZLbPhZ1CI1dIt/mJ6tLz4ri5390D71bQzBkfGEWdAIS
7cdkFEaNI9uz4WPN5EZfgio5nKWBPoJYiIL8ux5SuG08rB9zn2YnVLAWuXk7E6/t3il8yCJceWzV
16YK0ViNsXA8Y/zgj8Vt7QQQHOv5nCvc+Svsq6FakfWXXirJDoN8r2q0cnlA9CS5ZGzwBbtuj4iH
j1ubMP9x96cfLaKPh/c+klJAzKyXIzM5JpmWFhWMGdgbq7RiTnT9/JhUif+tmT5vajYGttGWOXUy
tvgkb2bd20P8op8IjfSfXHaDERCHNyiGqCvPflS6b5/Bv76f5vlmg65S59AHoqMHqHwBlpEST3c1
8uECgTEnqFU6Rq97ynnZcKk/H0bFZ/nsr7k1+6NEMYo504H29G2n3oZoN76eA+SPjHevKQRLjddR
2lLou3qoJs3Izz4jmAw56WXCSG7YejQV8LwA+lehEWwapKX8GcrhHpk7xA8SjdZCqKRJwAY/zgA8
EG/m7LYBFUyKum6xjqvRwd9n6hEHO6M6UPLI2szQH/3EJ4bQ6nalthDkK28zZKtoqMr2XhoC9bDj
ZnRSbn1sAEDwqUM4XTgRsPeUDWC+cjnAGzqRegq3MRTW9C+ylHWHhmwqTgTuGltwxHXGOHErwwBc
TTHqECzor7QpYOLPc8tqQJ4OV7eb5feTKecFa6P58Si7YnX6x6QL/C+FNWHo8YR45PehYCD9l+0J
2r13ObwfXQcgdNYurPQ3s+WPxX+Qo3mXq6+WIc4jOQRCAS2Dqk8Kgm1e2aAN3AjXpt3GmQVbhDii
R4V1sFT7ZcX2Jxap5gQVDCedjV5lWGU2wtrxfNPqhahtlraSku9+s9vc+Fqxs/bzW0TGV6hDdHKV
Wenil+QtBx4MIgQftRCiAg790NjIJm8rnjezD4hsGkekRt2Se1PntQRQhXcfZA07DW2hhJO9wSE6
NTAjVBD9Sb6VqD27OPpMZYRZlJqlUBj9WBxgAv92zj0XD2P4jd4Z8jPx7GlSZacIptMJW/VS8R/w
zi96DnbkUAY1rsKjPLktU6dA8tWR4CUuQKFOO30UhTupY9/WtNlenvWnZoHg6UG5U+wdR4rT5peP
BuHBbeGEQQS5Pqw+saJT8dvFVRrw0VmbnbHWeyO6GQM1tOCuxuK7dYfJo4krBAHE5qJ2SWWQ+LsB
LPRwPmiyJbE4thi1BUj3BAir3T+rkoMffiq4TieEKpLuc6LS9sOwR0wWGTygtg6WMpd3Gyno32TG
TKZCqt/QK6pgW5IN2R6eadfO4D8FUKlkeAYHNjKiM6zN1xMp23CcyEhi3ki/NpNfke+mI0hmAQwO
+zkMScv12y20JHvuB7x7xWHg61W8srSDWJ1bRI74P+SIOi3oFhB3bG8w1Txy3z1wRmzQDsMcbsef
wLNXVJLDp3gZKbdyzZ33t5ZyNsA9hmuc2hk6tTYx6WR0YUCvGHyk/pOMrsBvqKPObcn/VPzoO708
5fdBYJ4AluFwNFWHty6bxA/gnZExkMCLy3fZks2x18jm6JaTe5v7TEzNDTEjwYljyraM7vHIp8UF
2AgaOjxVeBVC0xh4ERvsqO3QyOiHtMuT1BVHUBxKWlLywTJtO99qZBUukqUB+DsGfewExunULYJJ
+xRG2rkhAxIPTNNQnBnz2tGQGQVq25+mrDiF8KriQwu6j8jfF4pgr10qiFoolIDWl3DCa1nqeJ4u
7uMibKEbFa3b8fQKLAlIL399hZgVdotgjMCShMOSVEBUIFZYdqL/0iPdh/32nH/kgxyeaPPjtkyL
oKc7Yg7p5jWzbKs99eRhYLpzkAwaV26+Ued+9ipKNL2JQXXuFxybgW4k282FsQ3OTc9badfBNFeK
pvi6cu7SatjzQWvUvw8CDsj+W0aG8cQPK0DY+FPlFWslx1jppwjBrF9QbwKKXDkjdC7HzltFIeFz
Yy5sAMbcwnsbe3i6dh6jTQAp4RQ9HvMUNEf7DCSeFF/pBZFCLaoHeOXNwB7ETPYTn4dR+S1rdq2S
OHGv+uKph/vhqiIUHGAmh11yeZPhE7rxRQDfXnkA0DJz8f8EiCDeBg7HPaxkFf6DT2/KcXfE1qbL
ajZTBqNYRK/TbuRQYOEE/W6Ze+2DKtgzAavQvNaVy6zKkjyard7kq+9zN02e2VF+DZXJ2JkFWGH7
eyQYZj0HMQEPh/TlYJvLJT+nJSOo/Cl5+07NM1eKHOWXf0hw2k5fuEhmICfA54La9LREue0eZz3J
flJxGPcf0fPRbdgF3yjs1fU7a7meeTDylT3FywuumQkK/Bc8D+JlWzOcvAvdIHAg70jgnpFn8I3o
HdDYhZJdKo4HJtDQXW/Nox/Hy1LRU3hJA69PZ8h8CgtudTMFf7YSDM9pvWpmb36BPXIPKsEK6VUG
zFnImuKK9eXVyykPLuz6EuRTG/jV79JGXyS4LP+C3KhfWm9Ngfa8FFatF+jQ91G8WYMZzTzMXmGJ
TCx/Ka3N8Tjr7UtmwbxwE5QW7nr6Qx7tZLwl+Qfy1Mi9FPRgWHZ2xFjgZEJ42F+khGfAvQr2S64g
LphLRdETSvsFpf1wceDnkr2oeC0sJDnvQ1YGS5iz3YSC2GT3R8k1sjUj4t3T1O4+WTZcKoxGUdd7
D4KkuCOcuDqwSewyYb9sbJ/cJUvBbbkiUnsIP6PajGMgZE/RvghWDmXm6PT5T/0f6Wv9qzaMYG3+
QBufFwY7IbRuLzD9cVuSgLwZNqxaqiNHDqeOAWQYY0PL9DmGc/NqcssepXobPpBoJtDUUTofmj6F
e20jQ4RtsGGW1SVglJRyat2Oets7+wtytGsPJR/bHHr8fytBv221ffKRTkb3S3a5eK+sFYIvUsQF
BsHpnkz8EdNL72lzmqbhS13Ro/jszQWG6B8eE3Run1gyzhnav5+cZvL/iJKxawJ/QDAEBi4RDLrO
zMFo9yhDET3XGx6IyKprfg8ZMCoeiV/lq3ZKQ2ITLG90zI2gjKjezd1dqrfblioJ2XFWI0NuZWwl
Z2H8rnZvN5r3jEobzIvdgMlhJuR0PiZCbJ+0bmjMAOunRd3RtMKQTOqK/gb4CE8DPI95MNHr2+rr
h+Cu7smJbYE8YTaf7eGB3h4BPMzSy7II3rTAXeWY5ci7IyQ5+Gs2bb7GN0V3cyS4jMGDFOgeCPXY
IKpgkkEZ8YKTLJRtsreWg8U/ahrSJkyxtNIILaBzdn+qnId2vaMADUqwAe7Pm/8YW6GLPU9sk/Hg
I1tkh791QJMD3asD5kNfaOzbnNkHNRdBt62ZiOKI4IEjmicYbezafZNvYGd/b2NHsRI4tuidyVSG
djufedIt9mbDx4i3YhUTaA0BMdLqyhQMJ7eb5xLDZwk6lp/Bri+wag264yUS0tzdgGxwF0Xd30TI
92jqlqdNqzoGXpW13KnFdfoZqFeKmQYgAEXaYhIGJCWew985NaAcRUK7Vhec+9rkhUcO2CqL6jW1
OR+SmuBw4ADi8YCvR+VAxq29U3CKyMLU5DE6AhB+ihY+YsGzGxlFChOTtdFCsNmPnLJrQZ62/MDO
XRD/TXc+xQ6Jpgbjpt7QmAGggVZgMr4sEVhCQeJqSiX62GBN7Z8kCiFZV9sMZo0NKJR+mIlrW53j
iYfjSRwjaGCH2YUJiQAvxlhHkXBJx/KKlqzU96C+IN8eWG1pQoXIrHHciNcH7L/TH/qbttw1mM8d
ECpaHg6lKG06XIyyMq0i+45//26pkwwVPSiz+aglO8XRlb9ry1P7jzhDiFAn4oXmuK0yFUQ5zAJw
UWkNux47WB3op3a3dk9edhJfdWl2CW600xk7D5iHMH9skfGbKQ1zpTLQ+nugFrxobekwVPqtR00S
yzhq2IxXzqNKUppmrsAMIOVpoejI0hvf+LRYnnrlrERcT8OT0ULuYrCTzRkPDwLuLfuBgWBcf5n2
YpUmSk6bf3yOj3r/w6JLU2Qx84EUAgZU9qSYLpYWTPIbXUYqbozT5WvWNLzaxzGcpi367dLwHHEb
ig6TsctSA7A6sJfJHdOtAbbEgs79ugkBgqKJIdiZnhjVgHrKDEzaGoMvW+tdEDGcO97K/0SLfN1m
V99SvLGsx1SDLyWmu5pzTCbxsxkyZToVFWS4JZ651rqrnT4CpFyk8trvLpzb6JXMC+Qn5iEzIDU4
EHLUm2iMAnvaVJep/5X9GXfhvRM7dtY+zMHYpxb12qoHTbngJxRxKaA0PNH1RHCXGWTzkbxfLaPP
EBvrZWfmB1igFs4+6J9AB/0SXuFU9CZS1w+KGIBk8qWXfauaBUiEE6HBOGCrwbrropMr5JCX2Ayp
9BPHMCzxvHCWblg+1yXQzt+2FxLNJpI1kDVHt+llFJjWvk0Tr1BmYQjJjZ36LVdtAAzjsKNMYmUo
heUB67zOJVtld5GnvuO+MDuQG/n9o3CmSEwnctaQs54pH7bRxF/s4ydrnaM05qKD6Nmtemy61XdP
xsJ/AL2ARX+SMwa2bpxL3a2tdYVwec3ER8LEVjgavQKzc3G40wMlEruhJVKVJ7B5/Ay+hq+9JeA+
R+7h3yg0W44W1x6ZgRnKT+qnc4+H8SInUk/JkxQwkyxKWwBhi49zqM/a6Oje50VKFWzjn6aEtAOA
Z7QD5SBua7koKOip2LO6MgnH6ron/9gpy1YJZnzDE0X+zNIYf1KFqOlS0Guy5fqs1dWRKJNN5mjY
BkmyGgvlbQCyONoIj33ew4gTWVGt5Nv/x/gzvebpyEiigElnQUsQD6oVcQT8ij5KNEv73VdxkPsL
btTqKKAEp9XWTv5718izH1Hkw4hGtpeVb6a4l7FHSNGWUtsvAheGDBfSvrvKwxYsheHWtcfctmfu
Smj8PrzbNu878rbwSRY33E8ChluEdwEXcIHugVrUaq02Lg1L880SGtjEcejtfMJEa7F0qwQy6RhJ
1gC+ATc9DJD+w+uWth2VYK7Y+oZuipVWUr9FHl+lPyQcAjpH/QQieVciteilVO4BDQAREetzycVp
bfgVMs02gDOZC+P4ArlS4yGOe6t3DvFJdPjX6KBDSUk+UxgOPTEdJHFS4PSNKOmvzk/Z5BYKVCyY
XK5X2Slh9e7BxR7Lu0pVTP9tOJFDdQ4Kx0jfnLQcQpinlGZ4scCB7Jw6nSSUR/bTRRT8pfF0GjBQ
Rjxqg0uZAntB/9tYu/j2K1m55sMDcSUpHfycSGYxBjB/jnEjIrB+66fh+iOtStAxxXUV0llt9fLd
XgBjl/wTBZna0dmW1qoFosElIV8dlhkq3TMTc8zjsq5TFIcedFPazcjAzBmR8JzhbggAqRBvtMbU
hLoRzIf0Xx72wCMSyKFowoS1u91jHUgkP+KT03JZDYBHNoG7N1oQqX34zd5m2N45hms46vZzVaOR
KQBD3x+rNFeewK/EBLjdRnhcy3oMrKvsYH3iPKUhAFZOtNDfUohjMlQpMhzHs0NuD1KMB0w5gENe
II1fNVYvU14nKsR4Bc/LMJa7SxuVusOCHL2OS1wh4mo2cUuolyNmmF7R3UsLjRhOT2bWoGnD6xu/
p6dxAbTbgozv5mCeyR/Lu7ExSHmAJRvZRPwp0z/YYJoUcev45hGj8yz1nRgi2TOnsY22yEKy70Co
b4XN4iWDHV3nEXjwNRFSkZcnS9iiMyxaqRuAcFxbxT4tFamI4lq2mM7QcYkgdGNNAXxxsMq/k5hi
KKjHjqciscp0FjxsKPkSbHsCbbkWMhbXl2v4FZoyYjvMRNNiVKeNSideP57c8iIcR6llr6Ykkjm3
REkJ3PveYKSampDrrhxbroQWYrLmc7uxc3G5NXy6N45BzDKWcOJCS0LpXvE3XVSjwlnNd71Do9RI
M+shefB6Lm1qp6h3sTKJPtHbmGU0U6Cb6bgR9ZaklGh7aRTKVSzhGyRNGlT0xXn3qzM5rAClOUv0
9OGoUcCOv9Q52a8EeSJb4XpKoZRNOtzpRqHWlvSI1FfdxLstAId0kql4Xk55KwDZzUtoQ6HVwAwd
a5wZ0ZnesKgU/T68Vtuv9nHeEMKwB+6258MgZlm/mWEPyXDEnmqN65i9BPkGI+TbjC4Dif+IxOLm
H4jLVb7Nsgtfw9ieMDwyDOqWv0k4JcIeXFm56iZKIRA6Cb6KO1nOrmfbatliipEObHQHtduUIEaM
NuNbuZyEuZopuwzKaXDf3ZXAmOJnSmX3h2EzF0Q1bl9lWNrAz0ZEV/Ji/iamkwmbPA/ju35ksMe5
ehw9N1md6LmMecnueYRRBi+xfYGP8+CTl1G4HgpiAx1298TSeC8K77hEEfMsnhptrnMwRPY4ZdM1
NO8obxbh2TMwkqgwSFIUrhwSdQqOAPLB9y5CMGW5ahYm/VLYdBh8+V1vCAhRpxFKD4AJhiqM1eC2
aVUGMRKggYI8Wl3sr9jZJe2i7WZXrypdYuORrzE4aKl4rKtsmuTLcEyFtjKpuSxu0nE0WfU2ga8C
XaH0RBf98/eJkl3+4iivdO/rIMm6HFq10eMmcf2HTtf0HD01guxY6Zce4+MAmTzXp9P55kT5sb8+
WyQeX0cJRZ6kS08DzKuQO7+xB2bk8ZYdf1uPG4o5rUZg1j5RLYlJ5n3qj1YwqvkMm4MiKgNfrI9J
Ght8gk72C9f4blD4q8tA1IT2lhMRWzxZ8PIU3LU+o0TX/d2IKVYydp61BmyL+Gex3YFCgPQdCsEx
y19W6+np+aVJ0+h9XKpi64wvoPSRqXHliPmkdC720+tPvIWR87TP+eHVcmeHtKxW0ARqgSv+wg7Y
6u027DS9T9O69HBp76ANHHLNFT8lb51I2uIMspjww/MzVWdyWnamk+WOPEiNzOJclkbBr+Dap3mk
INHGG+CO+uLe3ZpAVHCuxCvyc21GaBoqza+f3092gCJl4sA0uMAaPV90Af9ffWbbotZa5/MRhMNl
Spne2kHYLny9tDSJcOfWJNtg3THg5anKo0W9MAerDvxmdhvALAbRutudm5JYK66OxrM5cdQYEsET
Kmr9pLOJ4bj6YRUBVLdL53sUkcNJEURJgGIGwC96stDprcUDcbqBX/CKUtj7Kv6pprHZa3F99SlV
ZytsNTN1sfY4mqHd6DPmRU28XJm/su1pwQOxe8lgLMgtwNuih8J4oISxuJPypIXvHagQVxeAZqzB
prBLZd1l1aYiiaMSHvCVYmY/xqdY+WQaa2m4VxKdxfBal/U3TFH+QnFb43P0PZ5BYu/R0rRTu1Z3
Pi1vCqP2K3EGuzZ6V0AYeo1dCH1aFjSbAkgCA4HMGLqlTC5KiDLWVpP6RK/WsmSZhpL9Blz7Jg2l
qWxnDaCRj/tbSMUX7giGkwFIPHlyyg6uTZkv6Wr0Sqmy7aj+ohVrx7bxB6oKFQMc5ghtBRl/u0Xw
t5NNk7DeyKJaQCK2QRaUqqHl/ObY9Dn5F3JQT7eZFuNBH/TVIWQohCAFXDGl3M70Hsbu9ivcMx1M
IjgsaeKDi/fR7xDU4J1eBPRpAjUSr/efR2XjqwAN7BIn2YbKVE8esVufvdT9vT0YENHuMSzBTYw9
YG4QjR0KTC/kl+Rp6njgnFDYY0Qho2Y1DXgfgImDDNzKpACbRMrACTV+p+BXqK2zjdsckGq6zaW1
0GTXKwYw066YPHBhoHbv6bLngtbLSog6g/dP8ot+z0zma/25/nogXZokOrXr8vT5LGoS5tObgUkO
wMJenGKFO28u3AOcUo7d+2L6q4PdR3cXGovHLzFpmXMyufsFP8Oaus0FTpZcXlmZDHR1v2il6Xg8
oFaj/x+HN8OQAmvBdvEc0qPyfS/WOTjlx94Py81Jr+WQuNpbtn9PqoK0nJXkikhFJxReC4pTco9z
yBTy1HxpwRZIacBQXyxyAT+hgGIH47uSXVsRl0B9Ke2TzqVw3yakykuAv+guRDYgITg6AaTdIVxM
scMAcLjQxOPeBknCzY4o/VYXPbisbSWs8FvyAhXdknsqHbG6dFT8Bb9lioEra+hSSFZQyYQfwJVA
0dDhBHRrPgelfw6W4As/6gnOhMjbYHo29EMD6dw7Aj+Z8XErVzuzAtNM56Pd1ETY/ee3CBiFllha
kSVO92gskm0wbCh8M29JTyWhFiN/h7btPVoYdYBQmCHBupmI9XGUjVwdV/24XYgpPcdqmuxzqguV
kYHAQKbRb7h5wv18NukfqlStG7fSykbcUXgcoJfqCRSjhQiELNxPdKMVOyjjwC6s+FIa94Q/n9SB
WyCMWoVTUCfOS2bTHdl63jCWk+0+A53BsX+ynK72zm8ySt4UUy8AoInMILiEVC0UMd9a+sHgWpuQ
peJKMfFSp8O9HK6AJbEc7iyFvUKPsJ43VeZHXZiMlkWPKilwnWTBfHrsX00JpqcWktYokBH8eO5r
Vwy9X2oPw5+4et+fxkvSi9FuivLe+AJ1lr06LZ8GadgjI8xbgMNil9plaFUo3unDAen2b0fg6b28
Q2zi3DTC1O54c0pHbWKg4OIpkAhqpCpafs6HLyMx0LgBWf9se5AtrWLDV8H2VUCf+GUEBkL6lRtW
Lj9LIvGCaQn3sp+mlP1vk6NT2d+aKdUWWsub/jK6xa/ylNNNTKnz+ykcOAOyHzPeDGIlggOHGZqh
NAvdAQBqPdG1VxMHb7p3IH6AjnrwSjqerLJUihCDIgztsAQz1U1QmNphRNZzkonI+9LBokN8mgIT
YdMwsz7C+6t/BRCWN8b54UfrBldAIX8kFAfIC8yh0DCJ65KdY1o4WQbkwSfO+wit7KkBDXpSPi0j
Cq25Uih6zfiEYswuNoouV2W9r4XIm9mkqFiWneusAakvE7qoPX+FbBfKSPWIrGnY+4D0dN7M9UhL
cj1a3RqNJZ6MHCu5fz+YfI/YTeeUmcs0tVrL0y5TOVFslx1o5ItSsY+yVStFIcNRnBq0ytZOQlL3
/iuWw843EshQ7hqEa+VfRs+UYbQgnwtyO6hRJlrm+/rp9tUe2/9Rn7PqUatQqIzPbENVgh+KCLYV
oORXVcbSOjdL+KmkANQM7ielV14sL8yQb2LoG/qBdEMkBZwd/M7y1xzF+/Z/aB+qCiQ9y9NsaVB8
J8DgNBJPjCGFcD172XFXGV3M4K1yNUN+bHNyM3cDPxmgo2ZN2cKD5b2//l+jUWOfk1Qz3OdgKXdp
s3ozRCtSRr48ptvmcKmhqpVp9PgOASE9I5kpF8vhbqqF1d9dsV7q7hXg3VDm2OYjMPs39TnbWd5i
LnkkailzhHxGoeqoloA3FIEuaCOE3QjyV56vrjHr0hribo2Q8lFNTwJncqAztQmLRyl94EAnHyu8
LtkqZSmtdoSURFemTAiaEFz+3Ka5Umzo3tdfe62nlHL2gj3l2heoGkRgDyIRiPzISU852WghIv8F
xNoxz6Q5xxsZuYPrFDCsI9WXBCLlv0Sdv20GfXRhBPBTO93YFj3hiVNDDGsdfO4DqwD3OZ6ri6l1
3Sl9wurBB8jRw8qglpSmdWZL9ypgclC0RVEzgjeBjdQesCkiJQpK6EXvy38Mn+pqFEhO/JFGeP/p
fYX9XGM8qu46LuP91zvAfrFqhfMukRGtxR8uS5qBm0rEoFG1UXff5Kqm24RCMOGnGMNSM+Wjuv9H
RQLEfKnnxybbFkebFNR3PdgBTMS3N5Clyn4Dk+w2IrfVSrqm2KYBATKG8Rd7G3xFVraeOx5vkmap
XiJIW2HOI0d9u00YsfDZlVSdR5olRvMKZxK4WNu2O8AKl+AvqeaXSVDw8/6ng8NsNh52DdV9o1uH
xbcMIDaIyKCuMP8JdYxhifIdPbl6le5IlaUr/BWwc1m5kXvHeenrgyUcDA9qY0shdrwSOEO9V3dl
0MNTblp9IGbVHJ5Eu0+d/8C3SG5CngeR8KsaZXple0qeEMk+eto+Cq/E3Zpm9OjzSGSCoKW+EEEH
D/AOC66ivVFBBbJley/I6wmjkEO4tg7DTqPjha0+fIfWaPI3x6jBhMJogpuaFxUaKnHDcXsCQrti
LkwH2i0eEYir8pnJjqA1xZLhGCIKPsXt40PlI6mTHijqHM+QeEKPCC1MVoYn+a1lOV7/Ubz1ZoFG
a7bzLvcSOj7h+0AuiW+p05BUdT5C2fd/IzKA5Jg80QMjLiveQ6rwEeNynNeGYxZzL5W79TltBNFt
2pHC77k3e8vf4brLdKQvSDGhcC0n/wTGEKwnqS4zNNQpE/ofugUIgTitPmMX2ubkBJZkKoIcyq7B
JPC1d7mW/rIPtW5RZ0hLBX1gpJUVa4c+iZx3byLWAkzVTe7eAZBAlS3xhXjI+FCwjKsqpNc/o4iu
ggfUw3YJyXHusL8ZXBE+BjieJLEc5H/MzW42tJyt0eNa44nvYvgvZR6FZKMRNwQBq7fHg13CsRJ6
IhqAbrI+DvNIWM65pIhPZcRJiwf2foy3Dh52Qv++T5KN1q20EV1jopEqgc5qn9g57NZWVirT+/ZI
z2MkS4ylnB/TjfPzERidTdbXrqlnKI43ALQDHtkcLFMp3wVMUafWYL7+fTZEYP75xtYo629RGFkk
3j8uhkbxZZIQ7Y+5ovofT2mfC9KmDjDluLNeOSRPpwzpxEuAya9bvCYxXWbS2U9ZeZ4WHxgXFPWv
qL5RGD+nOiS+A8SmmuKCU5KN/rJx9UCj5HQUdIa+hSPtryJZAg0L4ckeL1bnh/M3JtbhG+8BHdh2
ojX6cw44LYSw0mLWItnvLGCgogkPVsxN8EMlWQMgp9vDP7C8Q4uOxSwGBvyz/5FjZO2Ebfl6uA25
3XNWF73MfE0Vdd/bKw5jwEHBSUdToQzqZ65tMbACGRJIPCIyYJkoCuCdvZRGalB3Zvu8gG1n7Sg0
G5WnP761tgvZ/femgNnB43+dZLQAw6VRkSrRbda5USdaAahsDFCEAYkY3AXEWMbnMtiPoOT3S7w7
iU0KLYa8Z0/mTsIoz7IgKwWMY6WSh1BvWk9tb9TBcaoBYZnCzoeGbb0r4cBWYVOOXh+A6MUW57po
sIRG7qncd08QE1TZrSLhyPODH2AcpLw4UOyfkKGk/zS3h3ySdgxCl14Gg4GjzIwHd3qHu4EQ5fzr
YQmKvFnbbAh389dGmjzjCuA48ZOYqwvJtkwzQL+ehakporFTVIpDga+Kn/U8I8HxGSL1FjB7lPLP
ubSzwrOUWe1/w2BA0R7Fp2qZna3leqMDVMIc1YKfIkft2U28m7si+0bVA5Lwg6tzVeVvMw50xrJ0
KO9bTKZLgROuD5Et9LbgPu8D7Z2ko5tMB7jYD1LsZh+kB9QDFC8b3ilVOSLNpUbvNr7fyF1FWVWS
zg1jz4C1SPeSK3hvX827iiYVBT8VOrmllPrskFvX4xs+D8z1mEjmq3QYad65AFLdpgmem41U2En+
t0sUND1o6uDXUKtxdn3Zf72MebK/EGlAsReJIXYkGhyDgWGbM/8J2Oll3ghSb5eO3R/weoZGJWMZ
EalJMrHhCdGalBasP4wp4QeOah61/8BQExNw2b19UzRiFh2j0Pw7MLONj3o33YRLMuGoe/8Far9G
tqECQ3my69nblPsqWWMD6FyON6iLaXo/lb9MzSNt38rfNXKh7gQD1iOh1Ia5K3PC5Xb9hZgQlKIA
2Gd3ris6wmVSVC2VBMI+gRo0TQaFLiqdoK0WHRlrpHxukYR4z7VrxW8yN3o4yXGrelYPDv6iiaBG
v6FsN0skvuosR9wvK4b5J42KE5sZ1WhiaIj83L9EPFd4+qPnep+M1XqdZmoFbx6C9WEQYQBYcrrF
o2l49PF7IMN9/Hc1/I+fYsDhjSjvKuN/xm3A9IcR+FRkDouBH+F/8EivDwYCOn6w8fOpnhMm4O4G
12STbno2mm4VIAzOobKQCkNQBKANowoAb2YQugdFBbxCtBX9iyXIlAGhnmmjXTbnLoVPqyeQX1Xb
lr8PgYR2WNETxu6AxxgFBINrmZ443t3WD9QGnZckAMUJWA/FvMoBxk0jMbmUbOSANiDfyhAKz4fr
/ZOH7bDSIfspDHTxBOGOeNzVGYiiQp9guOO4d09vwOUC3Lo5M23SNnrASlEdVIe2vp2YXm3pvRXD
Gpj0dOj52lXpyXqy4OqGUvjAlbmzYhEH6BFTen2ZaxNVxED0HCzKfE8adOytycHPcENqtJICMNM1
PzEiEkZQ5yKg++ASuqx3hC7uyav8iA9soblzITria241GbDsBdxt+7gT+nnd5rDmJ8scdeToSHIP
kb5r8LDz0jRbFvw+/eEDP9eRPwVB0Fh8/Gh+ZGbFmnkDNgFmJI6FRIgGRwBDl3z8X+K6xT263+iQ
EFMnk5mpfqU68ZynmdQxCSJAgEkj86QwWxnGp6xQsheTLPwN3hamQUsXneDDvqD+PIamQ8OmVDp8
uZeYchenmihSkDchEKSDMThToFCaXMEPB/46+Hn+dktatFS70GOlE+RF1kPHOjz+vw6Dev7odAiE
39gtcTW/ju5w4oLnJKDlMmIfIEJRT9PZ3JViqFNO4+cJTlMNvPx/jGdooC1JQSCEmx/eRIpWVpE6
NAo3bOVs2awAX6wPs++g1jKT+IxtFsVmAkGjO8Ovt19hrVstzLprebjajVoYO7kiGV8jGWhNjiWi
fKSu9+QW558su/6DSX+0kNfRRwuaLMikpNna1kFwq2Ho7sVsSHV2qAZh2W48GF1qGA6k8MMG42Kr
GbHeae/0NF9N93BwNx7/VSqLlzdeaBXCLa4tjbV3iH6MiKcyOIQHo0MiHnUPn9micaIB6Qa2WqeT
4ALRuo7v6b74g6NlxilFHMBjv9VzU4CpSwMqXdeY43D5AIZ0ilmCDcdoqTLo8DqD7twiZfkw+thN
lX9+/MKuRgxEWrB9H9tm39MI4uuN51/oAVC+82ZIx2ICle4idCRZIf9pvN+82T1ejfaO9stgklrN
J01SGiA5As+tHdBaRfmH+KYPr2DkoZlv5qBaTGuI+fkA+mZU3ajExbZ4RE4im6I+/NQ2gXrQJXLA
EajOp9u7387pXU3uPhKcKUWgHANaFq3nKbksN2P7t4NAY4jAypFVbSy97ne1Min1Dn7Uf3ABOETT
fu/DYsz/+n1WPeLWawHw79sdKdmX0RI5JGlAa/cTF5ERF9zCXreBDEo6Os6clqcmaIeYNkBGs92y
pcEwQ8ZvscedTUMNVJ3TYETthUXn/tKwnZS24GrVhQigabSzELoyE9i+L6BghAzEuMVJCnf65efq
ls2X0938Rl+07fvb/YA7/pMeTwZotneSkNpo9dWu6R2G/qrDDxbsM1VbaUNsdJggxFuIXbi3XQMh
ShQ9E4fQcQdJJooQ44KSXSCB7ZXA9sBlHaekawKfUf7auxtXVCUbwnOZEwzkf5nDfsOCo2HKothK
vVyA0FoU8rGBten6BFobwmGXQ9PjYapHFaaSuO3rKhKJR3I88Pxk5N32I2qJ0dMPeU4dlo399Jfu
x915+hE84u23mQAniJt7oYyi0xGi+8a+vOljovZ7kaPSKD5mDWSPsJ2GXIQdUSSPkDJMNVRh0hwC
DA4nG95/d7OWngyD+2E//2PlS+WUJNOwkhTIP61vxyoscXw7dRnvtOGuVkvo2k/CNR25yOJXHhtC
pxSdSfxXfoq3XwZFcRKdKCvxPzOkO1G74qfxxX3F+wZXWgZNDURCZFeuWbCkexW9yYfo8tV4Ct/M
GCbqAM22ODX25j+7pIv3kI/5Pnm74TcJD2SisEPS/FVMXM0zSsvnNLqr+AxK48sRAbhSgdNKTy4H
QEI2keUCmuyfavxodJu3z0kLpuHXbMMn6HpG1XN64G66x09qK+RBs9clCPMgQD+N2pAkQgM1LTbP
CU1JFXV2KdIN86g8L+q26PhsLA+eTvxkqm6o4ZZQSS73DEJBO5QBFMIehDlc1YcNjFL1GqoXgs1L
UBCo/5TOiikw1Wvbe5zJsmsNPgei7kedYrubjuuA5Z746Y3NjydtuqPv+FILw/Ehhpjn+D4Ja7/6
2Nu8JicTi7n8crz3tOcLVmb4n9+oy4BqROlimwPOQH3UreX1hg8vraKt67FyzVPOFABMueYJFECb
BDl3nDLXQ0OVmnyIftKTW0Hmhem3MXTtAsVp9eRlIvp1X9DNMBs2d+shPoZghuC2tii0neoPEEnt
+jSC1Fba0Ij9WWVQ1ED6JYcAVorsjxKNk3cQkwprOcKaixtW91ZFw9y6BSV41yptBog4eqbK3uoH
pwHHvdU5pHS0eIwWkDeRysv9rKJjYGVly3xrrNyw2jKuAVZ9KbK+vYrjlzyJohkVgHB4bbqSoUA8
UjkDMdlb+YJOwvJE5O0YabpURp7WnYcXUEaPE1KaPnF6HfT1zWHtouRM69v8AZGKCUxTKcKyARc2
mbcKg5fK4tGMCE6YHqclos495ngyrvTGhGP+Ai6mc4I220nIjEh+bV1uM82ILprp0UhAXGO112PF
k+ou/54wDDNqlvYUHNB4yVht627K4Z55tDUo3H4OEIqm6JBJqcWHzs66ekAiaEGgFV/PCXf2jsys
hz1W+ZOhuS9VyJxvOnfk4CcKTqytjRAhJob9EOJNndPeF+Lhp4zf1udw8lo4VH9aqDL7K4nBcUAS
lWziXrYt1z582kTyxNDe/OnixStfb9xNaT4LtIjKp3HpppnpLjadmtqPDie34crjF2Q/wM9nN0mk
bfW636ME2WF4AkdUUGrENAk+WrjcvLhZIE4EaxHnvT1qb+/kVs3hxeWfJoccUjYOrLrzEClgIsSz
jFK2xs9HCyTBcTqLdHL+tgmqLmElpPk6C4r4l1WJDMYH5mx+rmDfoo3nTypcUhWt3RW3SmPQggNn
9Tkt65FWpWoTaYZfLdbPsuM4L8IskAADui+hcnamCaOxAiV1imL+T+RxlTj5IDSWHvGIKMvzMWBn
iG9E1+fuV5S6YeFykWld7NDZfIExiAVZ8fM9dzTUH0D0KW9OpP2zNo7aLmQfxnTEv15NjEmAj4Nk
oTShQoWfVB4SFcHlzQa5QFS5GTvyk+honpFnsbP2AnQmajSTtBv4mLT5B5zejdXgATiOJfqvitgP
eRHdNbqlavqqd85KL9+rs+ODpet/84iVKLqs/wXUHK18QQVczPwQ6Pd4DgNhhtdDQkd8RiooBNpr
zaYkY0v2cptM8oWK/HdzBjBO4F+pLB0Kx7OcjwuirSYUq5JVp3YHY4fWialsETfbrT5b7zM057wY
3ljuOG+W2ZCSyTpAocHeexJ4N8Bd1YHZkTc1Yqv98aD0jdcthGWj0PoEdaPEDjBZQvMX3fwygR63
J0CmmujwvTXXSAlv7pk0KPhlWM/WuK620b2tyuI+2UsoGocdwj3KeKOcrp8uPLNgU1nsevCjLA5k
jEkCDSjVmhT7UOL1zjzSHDIWTV/TBvfEtMmrjTo8MLfCRBvMYBbai2DeyjZXquspHUKGArAV36S0
a27wRqgFr3ZeOQ+vyfniHB8Z63zXpA0z2fTL425FpUlmLUnKhblCjccJG+6E2YO1v4nzL88ABqEu
bkwdluTZLyKGueByGpvRvCkfV8abRKHALsYMuQc3D6aw5lc5mqoWsGfKUsN5P/+/LHw4ZDSTYt67
8xisn0sHKJCw/uVw4LCGQPg5ZFYE2CwXFznyutvsHVf2/kgCiD5HKZS6gwmnxaJmGND7c/Aw+yWv
od0fYyu4NHurl+GbzyVJ83QDMWwpMxj6FaKcD5UpXfl1NVSB7lEcm37EA0Qdx3bukrlNCX00s8Oo
0XwDfyCqsVvFCqs88DLHfcaWkd30sVsyKZFLSdSMg6+EcS1Akwwd/EPxH7u0WdS52cBXOSS3ZT3P
loUkqGA1B0DWLyhY4K6L1QD86QC/6tgkxHT3ZaifXIL4BlbYlWtDqImGV+9S1AyLfp1MF0j/OaPk
2NBT+u36HNedJfuT0n+uM6wPU52t3MecOfB60QyBof43bBu7IPNzOE9qTL4cOR2xdKKqxWKtYuGj
8fJ/RUqsa8MvA20KbL8npftnAtljbPYzAx2RU51J30muWvUrUNmmI6OjU/2aSGWSC8VTJZiW8OLm
bcu8Z1U3BQL8QvpKkjVag6/ulBES8NMevBE2j/RhJ23YQg5pAAiikkTnJXNxk7rPG3Dy3CcL8cgi
JLYAipvMGC2TDw6WOZTLwlOa26iW0p9qzqusk32JlSrtHwKP25j+HbXkDaGW6TIlpzxAihACgAlm
2TzeylBFwON04KPWclWsKCAHwSbsaK3MJ0g5NyxiFGpTcYJq3roOGidpfJbBLYt+UWkJHcmcNuIt
w6h5o7ShAcswpfov0Y/zWMnlbMxzkLd0QQo3obNrte+GIPkM2dRGpGsWbFxz65rvvqVtSemf5qVW
6oWCqALRyFbheYHyT3p+kQ9TAXyHkZ0FT0o5OqayXE75Xgx0CAhmnz7RjEi9v0dPheRLoFZHuszx
GxUC5ZbcfYg8a3Jvr/HVr2JDHUjhZjjxhsElntANPBev8NnnprWyq9I0MIZSL9z4b1K79/3D/fxQ
HdN4rF9Kd3hg7vLsWttEw2AWbJH/eaLmJek+2mMpT+BhX4gS7W7HDiKJaWjSFf/N28enmMLkUukk
RFpTRHK0o+eFbfSrU2TK6nZR5FXbSuovhWmwcDT/pQqcuKwBAZ1BAO3claBGrft4TmuL0gj9ANBX
f0KSG50jAiZwZ2c9O5F0Ul5VrDemKcNxfni9suSAJTwN6fmcCQHSM+zpan4jvFv/x/9zvw3LajJ7
+bVaWs02UV11GRWR6gVB26YoJFG0OY/XSFEiH+iA0pDB8zoYCnPts8ZDLlSOP5wOenjfuZmmMx7o
i4YT+BA7TsogVxfxccRb/46Pa+zYFtNXsR9WC9WCRqI4uwzHWEzdiK6rkKtXUN0iX+G3chkTUyra
vF8ty9zAADjsaQ+dVLxLR2gosLrhj9vKiOx76mx6fFuke15cqOjNTg0Y7lqT8EcRvXl3TFqOn2CZ
UFwyw90d/ZFB9iNwtJeqdnYSK52gW8XlMIkY7cuD+jRAeEh90pkapxHoyIwmcvT53rKz2WZo33hi
PrHM6sOLaeM8Jngak0Z/3xUnUWvOH0URPbt3oZToR05ZlJ99VEZFMoLs8/zMNj3+0zZS3WK9aWXf
Vd8KMI/rzHQKj8snAByONoGHav4PuopHBD+BuYgpnE8oLF0a+ub+K3jXhTmzLLwafXNFHTpyUayx
VzoTWKAvDMgtGXOw9Cuzc1RixGuDLCMYZtziS/eEVjukU2sh3ThxZQ4b97ULQFLrwOXhtwbibtwm
FDmpge9QwEZ97+platN7YUNd/eqe3bVLR4MXfVWJgBrlBDoJ8KQwBXF6P+vLNbN808WI3bwEkczA
X+3FaDaAv21XQ1XIKEyY2KBCbjdg2zTC5VrFUkdA75RXoSKUgjfkx4e1jJzkKzLsHsyZ8sZ/kNPX
m2QzqcC4fXVaOPCcS1F+ei/AZ1vQi/w8gdM5kq8cviYQTKbZdltfmvrBWneqswfcOVPGikUcsHjp
GcIAqVTOhPcPT0obt7GwCsR4maL7vIQFVWasUqTzdOz1f+Mq99fiBVmAoaC3A9Aavq6FfGBBVwnT
jeGoSJ8Fc/Bw0It5QAITR4Y+cAgsx498+iwtgvhXvNk2K08gaT/RC/milDYKWo/zkGqlGDVIR9pW
ob/pCHvTJB1iprlkaZmbt8Novj0ZtwQBPFH0ZA0Nsdzl3JM1BYvY7Kjl3C/gNgQHNzz4ql7UGBtI
G86SrbyAyR0SYkMnjPXdh7eGW1KLpb3NBMwTzCjFo8FXr4AH/e9+eXE5yNHQaub4D6hY51fTEIru
20b5ZoEEcSnR1GsVh7bkRT+qQC0GOnICROt7RjRVpXxAobpxAsFH7nUSAFqF3FBL/eri2AHnC36j
107OHhgfnL04S/ajzSTU1HvKUaKuF3komT2ILj6uH89M0fuQiMIFkMfOR47U0V8h0gZBFMenIOra
v+Lj+bZpgKF4Lj+OhresClVaOMmIoq8tnplHtUDetcEtEkGLRIw1zha4pVMv2YnT/IYYwaaKDDDl
V+iekx4t2Ig85AEqbyZKpMt4l7VjejdoLr8Ny9mieDtx/0bUZ4F2hZ/q6bPEVdoSVvE+oHZe3jBP
oCF8YqE0ENowJ3nGiWHjbueESxKv4CF9G7DDmQjm2z5u9nem/RYnkAFNTrzZt5RYrC/5VaO1cTjr
W0T2YJKOAkG3CR6rcvk2jsnyDXgcMsPRZ8xC0RNdOa9v1qFk1lno/pLXGrtNbOQad4N1vRhm1TQp
GcNSh5ceREyps+i50anWwF5GjrbxnI4zuz1Vdo4cznQfVpSmDq5YGbVJL2uOf4vESXYx83dOlyJX
t5g1FoI1KV0ptvzTb6aZzYxlbw1OOlL+CkIzMGqSlI+hP6Ot6p/eor3Mp5/p91por3YmLjm0Khi+
dwWc35yvaTL1HTYjkYU1pQiCIxuFlApbPFOiZ1vVWF2HFHIfkW9e/VHj3U+LHGJOeLy3SXOm13jf
dgq4ybXlXOQTYDS/o779gykspqP7tG7wGbHlP0mTJJou84L46oSh1u09+gmWSuXzv4YiRPxu9wpR
i4uMjntY32Ri28+TZUVUN57L5NTzPufbnmITI0aj6J5hSN8md0Wp96ORI6twwuIxS+6Pe1yANJQa
nQHfhoryPsTH6VnkSr8rbzUHl6gEgbfDTPq5hbFYMGg52Yna5NLFfJibs79QIffk+CmNuPw+vm/w
r8cx8mfrIqIy8Ihl0x45OLy/6vfUt6/6VL0XpfA7kKwxlPIeVfyZvfGG/7Al3UneKGipzvBdB/3K
J2OBSQws12q9TRraVs//1Rm1Qq5Ce2DY2tg48PFqztal3367ANkpsjKfxPrcCDbqegqoNDx8lw27
jZ2+ME47EO4H/T99LgeUpFkVPQZOQwjA7xWqfWeM6FeJQ7GTsRo3gFG9J6xanjdluZJ0H2cvWH9o
Ktqv39bf7gM0r5Slx5SCXLpOwwX6GSXLj2inPKrbBkAnwyjBd3gzVtV/Zsc0oT9Kk2OngN+N7M0U
VzTk/tmqIzqnncSKpWY/cqtIchN/S5tlj9amypPs1VnH2+6VGOjOq+Zv377w6M6JjYolhiUaQHk6
LSNcjeKnSAjz0/78mTJkELj/qjf96PSvy242nyqUM9B7NCgbasvffLwA5TCQbnyKjEhZysdHrBo2
rkRZSoN86rCKvSDPI105uRO7MedxAetNUXS4LcCuFKHbKvCGtZnGTM77W/rVmsLZLi3wBwWxGM9p
9+mCrBDzcBCTnL+tq20hZ5aWOLwyDz70pcFbUzDuKnaM0PaOYP7JIegR4U5v4B1yhqiq1Rdf2aj0
ZUiUegCSHr0BA25JtIlpuNfSjYhRDIAw32B5KIu3JXoMmV4yJ3ZMMTo4gcXkLh0fQzCv89pL2bdf
iIqLOrNJEw0JARjv5CpSMimPELmcgbV6ZnnntVNqXL3IizlUkPGNpWWyAxXkWCRismcTeJdY1nUB
+giaNx0M9ErggaFlOInUKeAVnLqVZXJ/7TeZ1xO1hMzyFQlk4vIYSxuu2+bHF1LUCCM6/GUtFsXa
N7nLJITMLiCm+lxS5b6I8VPZIz51oGwVwU5DaIzcHbh5YmXK3HN7EAaOH18VoLEGc3YlRiEgydRN
x9v1MaX+qH40LtDL6/AsYowt1Sx09YXdBTZ2QE6vKcAfN6rr+8L0wcEZXKeTCouwTtMmqMPzknCj
KeOH4kk+ovLYIbdJ1gpo77sEcEem4uqPmDZrF9OKw0xSkNKsNk8+8lG0l3GpgNlYVUHk2KF3w7Wr
o4iry3pWQfbYGFX6EWWGs6KGpCo/Wzs3F2q5Ij4LFf9rSZPEVeAWypOFMRpeKzCQ1bcmes3O8vso
VL5BoIbhEYiMpwPCsdXUnv1Yn0cuYK87S4Hpv6IEukTKO/TojNGmt0T6DHYVwtx2oBQgCOmdrEGZ
4/QRNx+DQbbPoz+b3yWcnPpmFxiYx0/8dJ+hwT6GEapLJblFLL24S68yoQsZnjWavGySYLyCAiAI
ELfdqaS2glkS8rOS80SoIY1W07gXcV9KAYBypboulLQPpcFkvZreoGObgPnXJqyv8od0Ev0EwP+m
1gJ5lNlVGCu2W+rJb2Y0Waz7EeFKKcpTtumNSsuUKR3p3JBqiKO9Nr2jrkbJmea1vd046CqPWb1I
8+6BmxoM3mxY0r8YMfAXGOMzsKEq8f8L1Lwv1c4c4kz3fcjtsK6GMAbubWUnw3Ej5IoH20ph7qOE
hrIS5sjod3Td2TJSluttYkIsnqldTfc8JfwMGXm4Jlz7aOzyvnB4/T3ls0lBTm4TtNzMG/8ijZXU
T98sHqMzrcQKScxf0ZFROVne5zCOlcK1wjfcl8LocTPPiBR43cQufvpeG1ZgyPRZkTdI6UASHVFt
b6PsxL54b3u8NKCLsND/Zf/xSxAVqFjDdtGPe41zIyVas1cOEHZ82bEa7y9ZNKHchKoyuyBS9qr7
Zzid88GFgblL4lWDsAYQ/BSsK9BH7bGqj/EqtIpfbLuuZCiNgB8N626my2R7n8YPSCRy7JiefKRf
/fCWKUFoc42HXA4PeMJ2XqqgKp+5gKnT9Rwn0HLjdW/1j2lITHQpXK7XI/J0SckTSBccGDahJb4S
xzg8x9uxboCB2OSduN+bF/FC4rh40q2H5GseL0PW+Wt4GuPh2X4dQ8wV8Nm7cGG2hKNAF0M/Bpte
RcX4sCml5kBSmyZbh+rlIRXfra+YocSd4tfKucBbEW7mH7f7YTEnazXMy29QLwk23JhULO1+r+Gl
HUX4hKlP3ohbYWRaftuvZJ5doHwW/zqUc46o4oK2ilc0hKyhlSMFMSFhIP/2h9KbJwHsMlUjKr4i
LrckpKT48kkeGYaJcZRH60lIV7zLasczptqdr7wwcZvw6R757J19+8IyztsAUxgzVVZbLI+8SICB
tBaSy4qB3iWb9DBw5JkObd3un/kBvaSkuuBWGyPSyjLl6gzqrM8B4jHVwMNYoXEahSh/0o1ZEDZu
odZwNiAoOp+xqDeOQztLbzOx6JWUMZQE07jKeD3pvWK14rEu4ui/rqxsGYUgVJ9XapKPT7Y16AJn
Qu5QQb2Mnm5wd3Iz9vNZbUvdsj1be0MoZi11p1GM0K3qUSX7FcD9UHdfaD7YpwnhkawIHD2AIs5D
9Fd/SZ0hf7kJ9dAENdjLvGHKYulmxZDOHFFeSifpvbUs0L8XqSvBQ2jxl6lOjMCvmDcoiv8JlCma
GGJFLVyzxlWS4a8iYDKGwkm7D4sznIDWTx08JXqw/9L4cj8p1M2UQ/kKpjo0S9AQGoJoRlBmLYJw
KHiXh5FicpF/RDqrsryaVW2MHiuvMWwg2xssto7OGyPZTTysDUYDhjrp9zT66KDHCq7P6MhEvgcW
wEc7zWmQ90iKoB9J7RbfC4h27+nLW55BaplkCo98die9THJ3/pDragLlbceR+Mam3C//rYOPoApA
+HrkN91WGmNOrUv6FL+zzZGFIPvhq8cbhUTX6R7hnxfwmnbk7hJBB/LXnRe5TYLwgK8qlwBJgbQW
MtX5Dy9CoHKG1E7lwGzFxvELGz5yQa9TGSm0+VDmz3BtXYieCK1ElxjF742OFIXWvQlowHn2yqgu
d0xhscrhummg/wzOQnR7kHde8iYQNTwsmVMc7iSlkrdUmfroJMqq6km1U+AvDjigWIvkyFnQAGiv
MnlQk8dmjokYnKyI0gRhltGXj8PHcJsZMBeeLQki0e0oHo5gcvjZSnzGKp+1NWhVp209KOfdveXU
J8CJwkPZEfBaV0WEge9dH40QTCWUcC2+0IiwUurZ5NMuyN8BLRDBJ93czYf2W45evCU99BqUUxuF
b9X0aFtpWM6ruhaVPXD0ogdg9SaEf7y7Ms7aHWJU1l/2lpEFWThCIWHgz8WYOjuwIDduvno7NSHF
447uLkYPeMGVr+IDlj25KWnXDbCGLY6ZtrWAEJxozr7cBcAAZ92SR1OZf3L6LqvgDtY6gvdIAgvT
pasZRVGcT+i0Skh35HbXNsHRDFv65BngiQBbBpfco9U5Slvhv7516HbbG+/8y77KJHp828dhVvCt
2OjlLlJUlkSp4/E2P2mFqq8gfYVqPGEgFZ5ewjaZ34vcOIRNGnsQtyp50gI1/DsjPhXKE9aQXP6C
dFXYFziNl1QBEN+RUXgzkDe+sbH58q4yEsl0/u5mjVlPjVSy999BqH3UvVyh6WrmZAejUp9RC3++
PHApBIDXK1pbIXDK9Fv4zCwVFd3Hk/vdih9YWwCOwCGwXuenSPmp8sH10j0CKeu4Qww5G7T8F89d
nwsyvk0mcDYzUJQGY89QXZUg3K5MV5jaKv5HPi+312AHjeqmGCes0g9ulSbU/gprVovnolaNI9cs
mxafooiFDtPesUyIsd7nsnNYHPLUTR9di0/pBkaaXH3ste+qV6OIe/RtoHKhVAuxbxJy/fBiwV0c
KU/7h9CFNWnAYDQ4wY3F5f4NYQsO/Hh1Jb0G6JXSkj+DAqnch4hNHdJQUT9yOamM6rLT3n3XG1X2
dcJztlWrcpOzRwOkY7nP4KJjxneNkLbRe29BqfhRrUrnUrQxuxB3yc+hOjEQO9rcletuCpqYkUDg
no8nzltS1yuMuBpuIEL/ybx1xqXsEKvlgVaEZSZl3xWwB4sAukGFsNT1QVYsc49jtnrpwAAfJZ9L
bxMjq9YkB9IQclAEbnoWZf+rq5DlFWRYvKjLQcfxQy07AXoxAA9EkCW7wTAufB+tpXLm2vqZy+71
BUxn75Wm92zZsYrRCEISHGH84UIAC2krBj6zseA75XL6IKUxsASe3wr0GnY8qv8UoSlFyX83ohkp
PdvX5xh8qvwkkibOxJhvcFGIhqq5eo3jRrn+V/A7ucx/7HcYyTMWh64Ny2XD6Pr7Ji7mkjQvPDpY
3grZJKWVqWHTwmApozR+yIQ8C0kja8GZNpHKhA7OF+IFt/lNMNFxIRAk0vcXywQogRvMhnaNvrC+
TXbJ73OzO1Lx8pcJgf0/4QrtsK2Tg8FWaIKJnPqAA9KRMNy9I9AlKNsIqwCXyUthJ/XYqLg41nfa
EpvuAPZP8TZuK3OoTFkVZGlXnLdRCFcKuwzTj93v4u1dO7C3SzggDs6igccpTmJOcpeGpoS7lnDO
bGtC1lU579F4Y4ypIqxkJdGHSQZwUEHStuTsoe7lPlW4+jCe8MPe3lg5mwmoESvf84urM+X7FyMH
kcajR3bfEWhgQvOO8luxvMiwm7r5cEEUmLFveocyjpfO+T28BN97idSLi7Eyzzko6oJ1pr/T5PZ6
6VLKnUDVo/nPPvyow5HwY7jNXYyBOvf9h9XmkkUpgEuh+3v/HZY9m1DTUcLSO1av5ZmEhuRYHS+M
1Hlz3Havimz2QoxYw8V7Vb+TfpB0FM9K4mIV85xrAl1CBeftLtzinAOTcs4ntq/U5spOSvka+eAH
5qyK3bw3cbzApKCGHKP8QynwzZ7NV5Wtk7UGHV+Qr1R5aHKmsRwC7X/k0XNUjdZ4BR5DKD/V39DI
p/OUVGxAR6BiUCC2ehclGNP4c2tsITnuYlu/pUH4Rr+PKogyyMUeEQ7QUrxoSvBO4OhbSnovOwzi
7waPXj69mp7AWLt+6gJulXQdnxvHFP3XK/hH/AmQRzOvgVEMQwJHtdMzN4EzybioRwdPVKLZp5xb
xRfJfNHG6PWkgSP2Z2+22akk+iHO17Y4YeeIPD73NGyr+zWN4m0YtLVShy7z/oMUpDM0SoTVN+8g
Fw7C/nfIt8Vt30GZauZpmJiEZaKYHsVcqJRrDqFAEeB4V1IvkGhi2dHj0hR6VCbQwFcU3qMBRSqW
JD/powTCyCrEDwTE4v1FaqYrOSO85HpabDWQQvlVxqx7pSDFn9kVQbONXDT7IuXY+YnO8+dPljFE
dMyPzTIESFNZJY193+iddBF28RK4YRijLs4nHKzmBFJrMLylP/TLOSlR5N7jNH6qAcNh/Q+bd/9B
eCL7PKp51aLpYod/bhNz3GkQpo5AnkHPTCOgYDbQoX7HjD8QJNcHzQ/x6IbYt2tjY6DwamkfrpfA
LxM1TcMO5kMuqFj0K4KwP01FwnSWSJw4vI5Z7LO6XaKisC+5ecvceppo1GJ2cJ0UbeLe1XrFqtrm
xtkCyAAjvGJOKp3fRYGqe7XmPwnAheNkwQ6R3vOG+IAHTwXSmnN2HbBC5KfsMoXh/yuj91dGoHuF
kSEQJmPq88RgPwl/YRYLDioUvGY2KaSdEL6ZgQx6yqtgvYR84bTuax9o1RLvpisfRnKTEkYLy0DH
XC4wQE0+3W7w6nqmIvDNKQt4vT0pYQ5stG8zFdPba2/rGxmmIbLcXkvE6lfRrV06TU3uH5ICTT2+
QzakOMWSgK5g6J/2VVh21aK5H6aRmRqF5AYnllwZUO6FzvDOzIOMmozTIc0HRoRktY00cV/yREuB
W6xOdbsntrqUiegkJYzbgJCjaIFSSId4YWtuhLixvn5Dk9fkLleG7TVlFfRI7UVprKAwqKLcgeWv
cdfDXDs/ZjZlw9TN826UJOHwULTzsl19YQ4P5y/989QPrvsIHwRroOPU04BdFR/WUWVd+HyU9Fxh
kJN0NX83OJOOYtVG8ZBSfW+Ftq6wNZEM6lJnBpnnj5sDw4CBQW87wXA+cyjDRLWLH2DptfLQFwGD
RrD/zOzXzZl5Zo1081EWkF2b9tIphF2sEJNzQSqcd28k6b0vgyDwL4sv5E4wbesMnsihCsgUSlBG
9RuqKaUNzooTFUQDJlBnC89VZIxvaWwoP3rzzfMgoS+Y9zGetdx5o+nfNYqx6sJ02qmZh0E2ATqw
RQStmKVpjevmavjchYIKhQ5UxpN950HGXjJTVZZCgxu4DDbwsmUh4BD0+4DYALjbCIcLJxX2CE2v
mZaY/+vLwxWnChMOaOIz5XXlzip+Q45ppJzMegwmaagype7HIMU5tda4Lu+ZgGBgzZKqXNla5hRs
z/oFoYLhubVclk9VyusinT8H31H1g04SlV4eDPITwEvnsRGpbj/0SE1ldM4Uuv7Xn9BdxUU3Go+w
THhSG/z5XpXKPgwo9ti8oOHqFr8gw1Cj5yv9Xm2bPPl1w8GMFlYGc+q1RBjBvULijlki8xIWfXza
u8ShUkC4u6MArddj87IGfaiH5dU0R3XDBLnwKBP0GpMlCE/K4Wm4AV4xg8ZkAqb/pSP3Mel7GGNz
ACtdcoMijknFlh4a0GiWJou7j4MFyHnHEb6N55zOCiOTi3qCLYGFuVlkYT7LT2G1yfMpy0RetmAJ
85di4mWYWZDZ55lWTD1aqiOySwKfn8WMW5FhtndONbk/026MEOoMdH/b/y3Ri7pDkcU2MgW/P5r6
Y4lvii1Q1HHqAlL69VcG4yuJW4+JDfwn+VTjfhIt3PHi/YxgSUTQxD7mTl4aKw7ZBuQK7cYDMMun
an0EQ/4/cjP1CeL2pNtIkHih1yLFT7h8YhRQKxyt40pgGY59NDHNqmJs0hl0+gHYjb8Mr+SYa0Ar
B2JiqoQ3LMntXIjrQCEFggn5dwh1xVSzkMTu/D/7APG+za/W+AVftcUHnfmEAcEt9e4+m4xnvmgw
/WnF/Xq6kZc7JPFyOnTEgbVthx1pROZDkEscWoORE/TxzpwYrbggNLakKFc+JQy0cYdssACbUWCO
WOzhrfJCsdIDsEg3v0D/dXhRfTEDsCQrw+b8O2+JyFFk0FkFdbBFBCq8h1a6gvkmxF3siIGQaCWZ
/2QqoBGSbsMRbGaylQqgpK36s4Zy/Uaa2pz34oVeXTnmf+DRDY15eniiTI3KwZCZLNyMr9y3A033
9hlNc6UuY/DKFgLZ/jU80rqNxVhA5Svl199T12J7ymbxv3ch3xU0WlruqQhYap3l2MqEIoCuYymA
XvqaklADqrgM79NWclW/VsiaDDBc4SWlNifMctSJ4y6hC1bGOCGWPjakRerNYzVyTm6Ge0x24d6w
gGY7Jk9Cdwnm9hp+3uPEQAn7+qQWsjRC2draMav1wnV1fBMaThcqIFFx8WxjKATZMPFOKCPHKuIf
OvSmGW4YV+f3GofN+POEvvxGGiSeF+FdAJ7aA5927+se8ZpQO5ZfjfOauYfyUb70DIbXnrRvqpIR
KxX51nsgDmVcQ+ThoLx0E+kNhLRYnSYCgiY37Oc/qN6jtDNTh5VfWcP5bZ0wKfqkcdBwEmJakgk9
HyiwMCgjlTrRozd6sSWh7ZhKSOf/+GqMSvHu9ZNLIx/Xv7UAEjwqYKxaUJdcLuEIcj+Hhl25fa5h
YA+Obz0gketwAL5sXh2qYzs6eGoN/t+p+wcVB8odn8n2fXJv82UFQgvVpDZDiky4yrXQOzqcC3a/
80t28KCwFxc5dIPWMtPZBRnL9psn+Cuu9E55yC990cxXlwVdRKy8JlBV7PCj3VKJ7CSWUwsvsy/A
Xco3cRJq2I9K6ryNO1I0aby7fDz/FTOp+DGKFAZ6mpVVU86yvV26nbyI2NFnCYqH3eRyXs45ZP1w
/rU6/lZVvcKVg3Ph/9GaCbaavZL7ExMQKFrn4oRKqxDWu/sX3Onb+hEKvABQMokbvZhnzRykFBuZ
HqLJNNB4Zv5DgwJL0hNzQZ2OrdKkZmmRdVUAlZRo8nJjKLWH7wnQl6kfVr+v8tb2lotto2kpYdSx
AxFoEEw2czrM0I1QoOAOiQituL1oSTa3c4Sp31GzZOE8pNjO9m9d0KLZjux0y1wzA8P0ebfxgmAk
pYK5kl8Jz4WDwLBTUG3NLEflB2CUZ1+sPmNe7QE0CPQtlIOsQryRGdfWSNrfzMleMbY5p/lGg4UE
3Y0WxnXxXQ9R6iPYM758gYB6na6idkIbiz4ZyUjiS42BsloS4AEWBkOoqCHyQGX59wlIVkwnm5rF
Q4CU1V5axBaegHnbRTMlgm6AnYKgT8LkjwneTZ0T7a630aaEXTzd5vcYLgpbu+fN8sdjdMjbX0Tg
NkO0TWHTJz6jRaqHcwMkxNKTCT/oIaOikgHF2thb+zyF6OJmG0UyDhPplexpqZa9Ij0hrh6Xw+1G
Bv38bXdUGqVv9KIcEY4IYRMh0cciFe4pKm9avcul5i9iEiuR5GYO0DHABgW254d/OOlwcJp/xMXr
oKH/HY/g6FXQDNqtkB3Kymz3qqtZIhUdDy09i5yg6DCWFY0jDREJZZDLSZ0m1T0zWTHRiE2QgxE3
R2xWkIi3ipat5HEMzQn25GPEax1g0ZArPwP0yiY29ZRSPP4I3F/7hbIE1ZeLRvyK7d5FEoMQ2rEJ
ku6o2sJgCIrc+dOstJmvGih3Mtj1FzkBX+swxdbt2vg4ODcZyyNBD+iEXTnWIZY8AWTeNbjbZjSO
zmpsqv3MAkBiym/7NyAzUhgqshsL//FhJiC+2aPNsssTMgcz/t4EpUtBL3Bkm6JBK8sYsnGQJS0P
H9sLp75XTXobu6ACTjL3yzlbrzgMP3wQZiEwYneCfgBo/TgNdJUZp3d6TdtDSbXP12WUrL+Jzh9Y
tnNfLurC0JzyVoW5JjLYEk9/ijAQM6BrCVx7edjrqX+ntcFAcA5hzGHq6g87z62IbqmGK6dM7w5k
YFBKyor0yH4sk4KdJqW0O26K+/sNibJHkwS7VnegZTHgTn9VledJqE/ArmzB6FFQ9hfWfo4c7z4z
G0m78vT58X8CnY0ij/Ph2VhtZFiYnBK5gB4YDY14kcMt2nrhy0hhcLfueY9i636HG9oHbwWfCLDk
z+V6gzTGlPNSx7/oZG6ao68JNLWeF/Nc3WscGNVOS8p1LRvTDhKBdYQo6VqDKfCb87S1ziNlpmO2
gNH0cL75T4Pkw3NKKeAoHKrO6kd7x2wcRYJlsM+a+VODRWu4uCapHVvEu0JyWuIsUozzvJSI9026
ob+T+ySupd4EHCIm1D5V3ENwoh+T7KxvZdBV+KLFvyvHFPzkikLxTXmpaYt0V+J5/Y+KrOyAs1BU
//ALwULSv2lKohgd4IuD34r3O5GDADGEA0YVXdT2OmEoCAuuyiVWJXIgf+bTxFgDfgi0clb5SMWU
SIHCAYOXIr3xG1uwGBZ24nMTJg91iOtcxdvuDoQVExrLFXj8J9/040FyEPmq4t0sqfjidCpxxrnK
UMTaBocBcm2vpabdkK6dvSCeAEfRp5ZTewfP28e21LM8VLdV2lePAIHUdM/k6LaryevCOkO/+xNH
APAt4ji5iBwupK6pXiJO2g7MN2+0ozzggIVXhJL00Cs4OkZWc3cLQJIE1TS+RfZIrGT3S9cg6vsT
oB5eRedwe+qICqrAjhkrDp3ihB6GoWhaNW+Z6pgHuhtC66qvhQIMFg36zlnxppAWDN9HBbp6NfqH
2sVZaIZCt3uAy+dkLPi4UVLc8FKA+OVoBsfsMw5fNf7g8r/kwJwZ2tyxgMNTTh+INkRmm+wtQ/gz
Cd9clVQq7arTB2eh6fogY37iDbgMDEHPiTyQlc2GbUuM71/WC4fV3MrZyAFu47KUbPV5Q1FWjHha
iwAy7HYcRIK1HwMzqcF6LChyNiPKFNCXvRBeNbiPnluEZ3LckB7esyS1tiqj/zGo//MKfukyvvK8
AXLOglA5YEuiqo1N5jKIS2VQJ0cNGGqSX4H5MSk2YhapegKM1+y5kNuC6H1hp7O0diOIgHpLdtem
h4cUALntVxMMdyhQWIChlV+/djakT9uFlcVaE+zhVTvPOxHexbiJm5rIS8fi2RxYSul5qngzSnG6
Hb1r8n17Ez5xiX7d/J2rZZ7JUF/Fjgx9uiBLFSp6XLuE7mf/+9i7GIB+7vqLFpS+tyL1qV7vH/lG
dKyq+fZrv6ssX7GPRQx1PBYLIYh17YeQDFu1feiOTW/lhz8towzpsVl1mc1OCtx+cMj/KS6vhHmO
9vFx44J7IF9gL8v4fRbFW+cDepEF7Ji3VcEKs9AYEMgtU95eIKuIsssNOmgDTQIG4MWU2viQ3ZX2
M3VI38pOhimbR+DS1c2NzpTNvynRmblmZC2A1+20mGf1kuNAFQ6XwM38vvha5Am+YxQPWi9O4wXO
5LEiXtGDEekEVngX+9zu1a/B/DtHyGVEdB73P4O9qTk6yatltnYM8zKDm6nTcG0vRoMI8+2p7Rww
TSajqL+D+VTdAjErm3UlJACPfj266ljgqBcVOvff7KG926RiyCQcyXmUSFQhZkUlY8LwBeuqk4xl
h2rHBu2JpxeKl5Rc5iKvZsimqUVDqQ4j0N+lvZ1BCWrLQ/Ah0mNcdYiRzGeu3I//qyqtbOw2KX1P
DOykNGvcQKcxiDDgSU3df+5eSs8sEPNkVHY3inER9GCRO0/kpYzpmwQwhByIXJU7wuxSOqIdH+gz
LvLBBp+IMdXV4wWsNFaGoObXMS4Hgk1USEmgEGK8I9LFFWysK22wHJf50TGe/209Miyc0kLDdc2j
GScGF/jUTj5pAkZPapMnu8wiM5v2rDSqjb0FdRg0trZ2Vsc/cKHiLepZvqAMdCbwQS+Anwxo0ixw
V2njATbk3kflCvf9I5HjYVYh7SI2IaZTbhmbBIFWs4gMQrYTy5EmeeMgoEY9EDmHZ3r+6m2NqddJ
a+6mmh8vflOMfmtuzChwgT3G2fjLB6VtMr9ialCB0Lj8zac6LeX4wfahZ2BoIDftEDEr8d5loQdD
/y4TfzOe2DO+utNtjveFCbXxJOvmjhncVdrf1eAM5pBR3VrHUgMqke3c4iSJUJBizs2zSl+Jf5bQ
hkI8720H9/wEZofblZ2+oV+GsUsiqH0ZfRVOKjacYO4ugBgdH/Pr17Xzj1rftN25vWonnxLPMRlf
f4ewTd2YDDrmpC8pDL1xdu4owHSSceyuVwe9mEMFTSmLvsqwJzMWeohgiM3lpnmxomuF07fDVTvt
Lp5OycY0ESFYIlJXbLAwXKtZRlxPWSsn3CQyAAxJA+LBO1xeq0AyuuPst6zh0IyJwZqx0n9ls7J9
/tgoVXgHn6kTB8ja82W1X+MV+X2mAn6oQrfllXgnYeXWzZT/5ALDdIX4q0k3qI8KFm5QbZZkC+C8
ABjgCxsLsFhbEP+rlj6BZjzg94wgvLZ6We9hNGmaoO7KINrbYCVKtkrZ38QjlFcKPeUUo7ouffFd
wE9JdopGejY1bSqa08agpvAUfYmfav1fC/vQUFMk09l1ORwIZ7fukKggkcMn4oKVSoqTC45rUF+1
HuG5L5Et7TuILpyYHuSfoIYrRzPMinsHxuW2psWTwC5MBR77+7C86mR6tw34PhK5DGQCrD91/ZhW
XQwRXNMCIRj0tVoYYIkbcFkbjf89twc22L6JiJyCizQaoVta3LwD1DZGH9WUkEboBt75KdzXuRFv
9b8f2LMy5hX3zixnYDX3TGfohzl9sfhe6K9mCD2kVAg9qUOpDW+JY9oMASkx9dsUSUXGyYe02tkD
efxNgnKY08vFnPW8F3TGx8+eBUWkGOycOhR6LD3l1PdHO3ncOqR+kT1A//91qCSWMNEsJOq9WTkq
LPk0coM4X01y8Sx0bwMyDMXO9mMuwNklqappEAwYIZE06uqAvwBApElGOdrEcwF1xIFCOStWSa/v
+EdVIxgLSf4MeuA4fTZGCTCfudyzYZP7ZJ9ix+HJ14ZCr8vmo/vsGJlvgyqJ5FuRQvRMKeRa3+2I
WNNKHmZz6QYoRTD5Ezd5jM9fp1pLydyjDZJx0JsgrFNQQiswfUPh68i4BcGhZ6ZgwaURLKZosxnA
9GtiZ6wN84Kes1pMWzIOJKOm/+NhqsIa7aM8Lj4tQc8AB4ENWjikPdpatozNDslcM8Kbga+drE0o
kwHgxTEnwn2TGxZBMkw0EQ+s5TUzLNytC4hWFYomtT4TEZZ7pemZNjGJlyPSpXRW1d9Uxo0xbIuC
Q3L8JVtM0tgPvpGO3zP9KfCi/iHBd3PvHRE0Ll2kuVa+M9an2za3S/mFMpUQe6lz5FfCbRAg8An5
sgavX9WHKgfA+xV9hQGkWTmKmToDN2gCu2OJtVMlD8UkE0YHHMu/RVwUsUSQiTDmghGM57dxkjoV
QJe48z3gMZVZr2JONjQysFVstp8r5CHDwaGekijdgeI+wzeQab/01uE9FuMRlqlhu5v3ZdQhqLY5
Kfn7zGjRVMNg8YpvmnDz0KuXi1k7PqcwZosVGWMACzLBMvhFmuhCamSxpDHOcm1qs8H2tUEdXW+7
04MU5Jm9YyISmOIt9g1mDGq5B4CyrS7bqLPajTLm92rg1uTl7YYIEAx0gjS0JD86Y2Pw0hV7RCIC
Fg1vzRFbofyOR/Oe9/XlEsV0T8ONWExq1UoFEpyHYxZp5a0PxS9+2PCbtK0dBth1dQ+O+uySwSBM
5w7JqLxIiwwxwHOwsEaDTRlJ4CmZtbPgLAm8Bu7i4sLLH38wOsC3l1rII7Eo5bvPB4kPHZmutTwG
LIffBg3kQooLLmbVu1k4YaficpH0GaZkgEzAK0T/TTUT7jFtoB+mk5JfHaL3XV2NpOxAG1rA1XxM
/UAiRa1YAH+HFQdLE096dbnJZ+pEfIqBii6/4VyuoKB8MYx9+Mz9jM4QfTKmjQWfyZ5jjc0x9Wcj
q8ira7dyGTtNsjzDipmcDpuqenBrj3VwAADErjzi5IVmGkfdfUousrCSx5E5lnP6E9DYUkhdUtyJ
53Dd5Fn4jE2jFroRaEQ2jFAnaFus/QyxFyH4zDmT/92YYlYrmoiDuloAYi5aQo7AWbXkJmwVN2mM
GmHmYGIHBC7isvxIWfVUONl+hl+5ib5UKoirY3LwgwC+OME33xCyvjmmesaHX5OdERSeH582mMPn
nVHjJ64F01OL5pzq7jL0jPTDGCbf1+8w7KhzBsj7PYxFyLUvjhVR8Q6Y5MnNWokRfxYZHI78W64Y
IB+oNUJqL9SuUzzUgbmboQcbmJ0Mrh3vKJWZb2cbkh4JBWTJQmw7YC6X3zUnGUEzxIAFgPjOl1is
PDHww9PJDE3aTcEIzmq7BwOA4s3rYqhHmeBqM8WyA2guFCVzkiRgencSsUd6Mvn6GH5jlDTmsTbm
3fE89/eJX2c10a69QpzmGTeZM3rhvyqjIJ3gwi+uOqgw7zciop5Vkx/FRb9w+H2aAwx9XH/2KLP6
W1BZvyCXjSHLc/mMjN+3H2s3TRJQ89MKRS3vQURGL7RwKbascsysJsKHYwI2RpZC/kkBGq0gxrsq
SSaxM7PG8J1sMUgg6Ab59czLvUldmh8BurSmaqLUvwn/Y8ZZzKXYRAjNiaDZbXuRFAB8Hufz5sv+
TkW5KIYBrd/ePN2ccCP4AIfdAH22nsYPcIUez28tmoDQQEB/5xbJyG1OMz4YZRXYhUlZ4AIoBspJ
eiD0eSc0YktJBX35qWEDxNS5vjWNrFDhZnvvr2xs83IzNNCFiTFtbziOe0ki51P5GVYxdMxiKmFo
q2OtkE3R9XjguLCJ0CRlePBFSm9ogZ5SD25Doe/HR5Uh6M9kuVe8WXChnZGV95K1Vx7ZubvXkdHt
AeJ8IBStcEUg0Igx2DbB5F9wFv6Mvb9Fcw2pZYkji50LPsM6xCo+J5SC3XBn1m3a/qLLJ9ZP48Cl
+LC+ebpcqYeZL9tSAn2Aqm7t6hC+rhkJfVGXaiDqpQ5kS7Gsk3hGBnaqXx8vGi53xraKoAKYKEXH
Kl3s+Ui/uy1/5B2/Fq/T5M7SlW5c4FxbcokJiEIH26KOXzqQCqAuno8n3sk0o104oy5y3aTkR4mJ
cVZvrXc2dKegdZxQZ9j/hE6rjqkYA0iFVJItm2E8AELLbWFInk2/bFNbaGj0M8616kcXs3bBEI59
gmfGysZLARToDCgJjVuEpvZta3iNG+HYoP+BiAdBEIAJt+Di3ofZgBynS1IZRkU6t0kLHsl/alsP
dlGv3VQwj6GmxHL3DDLYE5zNp61x3w8Jo7Kb5Ya937akJsBJx57XG2sqciqRDXgTMxLT7Maauc3i
ZQlH8b4l0gcuNdTiHhzrveniO+5ANxZIt/qJ5mPeVbZPgWN5YWCaDcmZCv511PTmSO0Gwbx+7CpQ
51TCCda0trtI7wVFYa+L3mnLdHq/6+aYA5RvB8oW35MzX3wdU7AhIQgTMqZ099WIczU0KBZ6X1F7
pOhq0eO/yg6FIWfgPNgwpsZbIaRtA4Mo/GEE3B1MmxdffkVdbVg3MCK6dul2RZGVEzAdsP8cZTmb
+ib8yrvqjz6cabRQ68wgGoF7KOlpuwfUHzSMtQH3qJyR5JjbtAfwkCkqTiOSoImkyCnzh2KQMPbG
uycsHUMVuHHXUh9CfAwRxGbqou5CTOOIXmMjb67rASGC9gFJD6RaWrqktVLdRgtUg/R9gs0aCvmz
Y/fLFH2vgBM9A5OHhsTxv6j+hMr+lqf6rO8v2WSsOA8rEjsMBU/wfT/0bBE4pulfWxLFH2ThoZcI
T6NJIoONBxo6GN44fRRlIFKINSmrdqCGh/KMQnPIZi7EiRDpgblQFKzBJzSpvmnC9lnLlARET9it
+kgxEFZqlCJvX6bs1kFuMRMkOjJb5f0PV7tqruRlYU+vf/Olz0SaD84Dty9WEyJkoVNaihBig+dl
zSxtCrDaIKa4QQfjC2LFvLbrphvVQ/b8xOzjMrwGxVJnLGOlO5DaExGySsO4inDwRt/uX72SLVkr
C4oJ02YdXUwPOGymqbf19vODtLWC00lkgZvqj9f2YCIRHF5jZiqHUkOKN43rvM4HJFE3UCDO0FX/
zQSB97JKm3LCQ1dhLmxR1EWKAX/eeGvDE9wmr7AkfLlqot506Tk1kxQyYlN7xjaQrnTFzPOUqUJy
LDATLkrxGRTIQK5faDcVOXePFLy7iWr5Qo+QGWHUGfARdMGjk3G16QYHsvSAu2VvnMK3G4fD9cZE
rio2IG+c+fR/ZA/NyIuJZNXCffnE22/h5k6ISl6g9vLBA7HG5TRiijNL8LaoxCFMxhDvJet2Hu1H
PRKWVz5dI5Cd+/QZl98fmmbRug2LiB98ipqOob95krYh5iwlQ58HyJnMhhUDgdzAhscCuaf14Fkh
CfUcPM4KLUHVjOddbyz9WcxvNAL1BvJQI66GHrzwzVhTENqlDaLgiN1bX/Z5P1E/0pOLIHrSz1L+
MlmSr1f4PfBdtFsqt7R8jtbK4vArpSK18CahVVMQp3ZLAxsNj1VUgbzQOsSsbBCbldMEB/J6jfB9
v9XNY4VKXFSry5KnKoE+upkeyjS6ue3mKzV8Vc6J1etpyki8uCqJGNqSEus3ZpzCKWXTp0uyKPDo
xEjKqwnuJoYwCO2DJWy4XaxdFkDQpRfOTd/CLeFC1lUT9Kkd8Ab+9gT7fjwMpRB6KL5BDBca897J
e0PnM8FhadDjO5Q2FFcOIWKOSUD7SKHgpIBAH5xPNmA3oqr9ST+XMKR9qjQpxc5ycfCImKELvee1
WgR0YlnSRspGqJ19CYWgTnrz1t66t9DyK0qUl0GrYBII15EiYRipGNe7Ev9Smpa5rydHUH7SBkTi
mi1qMw7UafA5SKNR5bsv9ZnkqIZuZ3xQXhPg9VMavqbghTGOLXE9tQX8MLWBLc66KfNZWLFwmEdd
GXTNEJRS1Xak+TeIkN6j0YX6qk9HowijNX27Hi+2PzkfNNsshlqc+BkkXIFVK6T+V1uitxuEKSK6
ZZuzDcaxcfvo2EqCK7zKa2mvV3xl1gbMLJCTM//hKoZ0vpi5321jiPLDHGgXLETKFz/2l3SCf/XH
dXlLFiqeT8Xhm0Xqsecg2qC8ALw9QaYC6UF3fXKdVdzSYoONNsmAc5wmJVmiuQpyL2ySyBqnA5Zs
N9S2xQNK9v+536+6VOOk4nUC+GQQwSM8nnQu14C2OvfI9R+vzY55s1ET2quT0aQgU1QfvucDhn2V
ITuQy1pm2nzFGwy9e5W7QD+mq8YdNIXZ/73sUX/fMq6nQK1FiQQyoR2oHyNo34tyuYc5tHEJ7Gh0
/cB4X80PBvZn/aQ4I6wC6Hr9ZsIfaCti15lmoxq+Da9b2e+DYbFNE9mJoIcbl42jmVeunw1L+idM
IP3ZIEsuyBG5Tkm1wHjsUil7EFH3Dci+z48e03SiKDrD+XvKMLavSgjOp86BkdAsp9WuEEmZlphC
QMvO/KvqTCiXSirZ1lu9ECGx6KjTNJ7vBZp3s3KFqQEiwqdJhR8Z5gwxIwJlfJwFw3KVIzl4Ajoo
lumtovBZdEKkejMIrTADWeYemXifWjP6wEwbJAD97M1+6Wu9CiOJ/CR0KJOLpnhmwaGhxP6nx1QF
c0Fc+WGkPt1vjsftcK4MiRbRPlyGyYiXJ0Bjf7z+MsO53t814SEmOgS54lZQpowxn2bIIJcF/kae
YAVMzqhlpAUMLn7wXG0hyJk6PPNg3Cv85AGPcvQzXxYEsOUsF20etKc/iqBusUWSnB2Wlts6wieo
BMd3HeBtI7UB0kRUZiVz0QEtJzpTIra8L4EPP/CWoLdw6rf3sjQ1z/KGQhnhk5fpnzqmEj/I3nfO
4ko8gO9J5oV6IN0dFjOPMisf1OWavjA9cL8lOU4AlMR0xx450r9EDUxi0QROSZRvry4lBwux5AKv
AE7nNyLrjGLXb5dvKiM14GN8YmDum7FY6xu80An9/qdCSq1IJ16C2DEw4zTQusGlCOisXRE1maka
7oyvcZEp98X9KKpUxR2ZQb+AoT0u8mV70pBrYLdseP33NSvPmTCYNRgF4+e8DWLoxVWOXLSBAMlP
NtoNLWrR7jrdG6s0F3aYz6yCECDJGc0Z2rzxdSMe4733cy7xlxX08hvjwb+H12RzLM/k/qJ+q9Y+
ETt/iiyENJvdXp3tmN2NFoXdbHaL3/dwK9nsYuHB7YcVn8MBlz6t1fmO1lEqdgSffG6CLbpa8w54
OlQyRd7M0LJWs6931xYAfsKbbkPISkWKbCZ0lI9mvfKEfzuhdL2lT1J1TauGzghyCr4eUqA1u04S
9MOwWCXMkKV9dX6hu8rQuKpw6esi5BdngDPXxYh0aTSuiIH8XRIidpEW4uigE8rlXGW/NiLIBzdx
8Oc+mVAsV39vwOvXX10fufkedj2y25r2mH/vDPoFAxJqo8LbTi2+tMx3W5mdfn/2wQPeBnnfq2ai
MIm+vrYX9U13++A9zqfHs5J7qMxnujJNOSmnebTxI+sAiu9uFSmXW3am4Jqea85JhAOYqJWLix5U
ghSAg6d7BAnMg9nvMv/FT5Wbw9mrXorT/i+0DauKfELF9KI8TXxFAz8wKYKIUIsV49d52NAfhLYh
427Gd0stxf3w0bUa77Q7H+YtFxYEJ01WyJRS7oRVJZaB6YxPnvNFxD8Upndd6Mu57yTQ0+N0LUlM
AzZugE2Dwx6AzWs6+ObdRlIRA7w9U/TfEZ4ZB7HDfasR2xaXkgs6JSrO6TBnUaHmgIJsoehyeX4R
nds8Q5f9LTTmM4lhNUkKVt2aP9myF/VKvmQqni9BVkWaRLMvG2OWsxRqIP8rsQBWFqlJOtBPB9Qx
IaNpCbJ1l7oYfnF7FaRt9fLEDidjW/NFkwu9xgsi8b02LNOodK6h4Booxrc2snyb5PBBNze92At/
Ea9ZJonnLVX+6OiVcu+dIaFdO+2LgVUVg3QdJtEYFDq4Su/GadOU9JM3TXXeGxc66IaG2vY59Nd5
fxDpF2Tbo5QWGcmVvd3vt6e85mAI7dJ6v4AkYC5qJcB6/uRbifsook0R/eTOmU8jACK5dMDWqxkf
sNACYMgoji2ylGCB2LxoFfkYmxgWT1FMfEKRVii53943SKe45NMF/NuZ6bALuzAGtaN5m43XG1Y2
9QNVGLK6nyA99qUWrcw/WZru6h1xihr41etfaubtxRA4QepDnvMASIdfr3pA+KtJOgTfaDpxZIDp
80ZYlqcDyGc3Pbc6cwL8V2yV4gS25CntZfxRnhT9ReVEiBvLaASRl86nETgZ+D4UOS3Fde5L6hhX
mBnq0JewPA+MNIW9+uNvBlGBuckX7L0PA0y9pXjD1TwYwaMqGn61HoyAhp6cRJxvrSYvRe1ae2j7
f0V/L0fNSvLTGDwa/O8Y0H9ESgX/TmLrOH/gTatF5UtpB261KQMmKbMy0Toy8o34udUi0s5oVvol
o20ajGRL3RAYtsdpYU5QdUJaeQl6P/5KfMrREjGtCOd/GrUYgMdxLUAcnqLcHX8/nmrnghqtXupm
7kNwWFNY/fIcxDIoOq0m43USMKLLgM2th50e9s3emD5xUBEd7Ee4CS32z6s3JPOoTzBcBFIxiYHj
UMmhYOCh9saseLBsszK6k5bmodpyGT5XTFry/WOoaeS4IkgQdrIWMgjDLB5kATQUP4O9rsFGCNGj
MknHLxY0aPpNlpkNrgdzCwUWDiayP7gRrwQKjAOJxDKxaF4IjKlY8ZefbkqgscGuUjLSWI59J3os
ZzLXVTXLml/M2XgettScim5iR+F+b9xLxR6mOZYgogClQlKUoIhQtZdZigakyUvU0inqNiMyhYuW
NoDhhmFyB5g+8gWxszgPDMIMD5Bqwm0vKCCl/zJ1W2TRO7gQ1R0ACpHUKW+efKTviXetjmDxIhjg
8weFFD3A/3F59f8EdHKlGX8dlQASQmmkXooa3tg373heYhzRbjWxQ/DB7YAtYgUPqM0cyUpQeeQv
bcZIlyp4gEbTNV9QqLg6X0XI7OrmPe8UFGZEghX/xZ/BH2sap1E2zot/TUQv/3lWMfrhU3LaRLQL
nmFXu5B/Zr10h/tsbxd7R9g3JjRkUtF6DfyriPih5hWoASUqWFpzs3y+9pV0hz/UrmGGM/hzexwq
9wkwpnNNN8l320gzbVxAtD0KRZtOyEdwc+4et6RePSViu1YOAkmfnBFIxu2L8wUrT3680NtdlqeZ
8qwo/nr5t9NlogKp0sPjBP2DmzRoCa2KG/EzdLbvOgzGMaeAohunRKuEl2BUHVJxHz8zxT0UZrnf
EU2QedX1o63Xc7slxGfJCHiVdWPfvZo7GsBd7odYB33gjWe2TgD6Z5VZD5HUBZ/83NcYtkp3NLxu
HUuWOaxLwadZGTnMQeDLetLBeHnIjyXfjZRZkIlpqzYbOqwe7OXB6hfCE06WXexQN/+vkzSSsPjm
YwIYExpT2Gj9drFzOY/fW4Ski+TnMwdWzYHAcRKSD49kOvh9mVXkqzErR24TfktwRC4svdR8ZjvF
3ynjcRLaJrNeRXZpOR6wthwNMxtwXd0fCI5Y34w8WGcfLj+8M9Ekt5Tj0XEmVo+BJG1NV83IR0PK
hf3ExcKeZvpWrFYVh0P+x3LmMD/+m0lF7PdJuWoTR7SQ03B0k+hCccf856ksGyqZT2xg+XIORmTt
hvIb8sXLhLx/jqYFVc93s5dCzBCYAy6XYnm0plTLMIhhoeRCRnlY4WphK4Yn8JJqyCQIY2y4FdoD
RFJ3MjR7T9Kt/Q4aT4NGRNTfIdYMnm7klFm5MakgCS2aBf0IMn+wS5hlz6gDqp7X7qdQ9rpEaAcz
QLHgoStRGqJ6YS4FO0TORELODeUnCFl4dn4NXNuWKmtWS+ME4CyP0LNw93CH4EkjOmB8ed2Q979E
kzs8cPoqLC//y6wWQUW4uM+cUoZgCVQvMji/jMVMU5Eqz/FZEUVurpwvHsyXYGA+yU5sW0H7CcIR
r69b2xAAtXMXITgr9RAiTNOIHvPtDH/G0lZ9WvLB6ssbv9b2GlKrcTNdQ1RiH1hXjU5B3LaUIpBg
DCpd6a6RPawlKCdgd9s2qYfP1BteA+4Vh2WsbpFTC358UfauWv4a0N3yBYkSv9qxIdkUDeJlDIvb
Es9gn2bIHb7d+RnASG3FhebY1UfYh0Gxd6T3r+X/RMyzqxoY4Mv6Oe2HtVmu4MPzfkcbPhLZznkG
31zvXhnxWM4lDMg9tcGw5g7AuIbgEnm41TXIOm9lW8Wn0gUm9Wx2+qYvqZe0UHotraytyeqFEPEF
rjlfqm5ik8aMolCKCucj2BGRVY4A7dEjM5aOv38Dy6itoMqg8CRF8qTx7J7p0V3QaZY0sXd2m64x
Wi7LOEurdCHjo60eEb2JR0KDPZBdy4lg/pJa0obrx+EaMqL45/kERvy/iJQI5BJBkOR3+xoJmEkg
LLWiwgEZMYXpkUT5RwX7CQaImPk5Vok6Uj5iCLJskoNbutUxpuPixCuqTweL51gjmuRuXsPvb0kw
OFXu9H/l/op29P+T4wmLm11p0zHqg9lvHgnJdwQpnDMcjGMBH6QUGbGIC045JEqctTK3v9ue7Ljg
PnI3wTO2MLgcTPGFwOqCW/eIFy5xBzpczm1wNJSlIzHPcbKhZst458ogAq//+/9Xd9B5DM7RTtw8
i5H2A2OyumFNSawhJ5YYN1S1s+Q1PN4PMIMxKcBw7AHUwpjPkmD00ZsfwNG/XMrnfHv9wfePjeNR
pO9VJ27yyncBXiGD2PXNhvtdWm10Eug123orP14Eba0s0LqhpaytiajDS4V7NIu4W8ioUpJs3zZI
hMHizUOXEXZFLCECehMybBSgTX5rTXMqF2zmaxpReQsDyFxxmLuwNDq95+sKL9/NuNpeNoFPecgZ
ViWoMNNFkbSXGTM0LhxVBKcvh4cO6/zzZqkwLcGzmCJkCjZBEr8fcX7EIT1dnLG3liOZg4d1tECb
AwjBwjGycR+6BQgqGQgdJeOYUkR0DYInk6ykshun5rSKgl7B5wVtlOxj3/IuE3i9U7yheK6upS7b
y2zBbybp/Gm8HnoQr0blyNx6LymrFREaWRIBIlGukchlDojBHKFIq6Jnv/Ov/R8v1Um/Z0Z8JjjR
iES0Q0Y+YbzHikokaZjfT3zrfJscLHQ3RJI0r0hf/Sa1Ho9v6Qn8PRxb+zRz/Jl2gB4FrtlrAUY2
TIN3IxqyjFJuGiY9eNyppEnSARoDchfwHmNLNpcZ08ZLwvs05Au6es4PJMNFVyt6oog/NBtvyXIW
QzGapyFE7GOZh6UXDFoVps4H2Iz/GpKJCSbDoexJeZmazJ0bd1oCHuVgiRwtc5yytPeWmDKESjpZ
Ca97rCwKPkS1LVGukUI2iZDcH6/abbz7HQ9nT2l8svRYwlRIUVNVSLx44ntKANKTEGGDBVNQUCAh
W9GxMq13DLr0B98eAvH558cLP6TR1sqvJrvFD+UmS4aIGqWsDz4ALeOlmSkrl6C9du9A48fm+JA4
f4yGzJuUy1l3MXOyZlRdlWSJPJdQouyvznEs0kikGd5BYwKOSuV8G7WHwkG9tdc0p2pDXlmcBcEb
Z1Cy43XE3gJoO7W9mopmkWK7ACtzsoxawzuqYinenhKdP7dBdNE92kY/7L3FrCMsB8Z1RXYbBbnb
xLCBnTBnDW1UPL6Bkfokem+CySdlYu4RA4HGHqNyk8Tpd+S6jfboGsUp7mpmfsAlX9w7X8blZWAH
OaCo9VbGLhpmQd9cxoIkXh0EoJ0ZlbYZRPszWWyPO/7IkHgt4uVeZ0kPBl5o6WUfBCWiTVtufpAi
ZPV4y6GAlK4MJ3YoLOt95GlPio03GQz1z1d/IG0NUDmSfZP+yIhDLs/lhx03yNwNNDammEu7yT7H
4huTiZdpvZ5EOfi6ZW9NWA9JeacnDYwy/b4uX4yMeJDQwRlvh1qAJ2WJwY5Q4lDjPNedv3s9EEzc
cv4StEACLUc5fIoLAjNG+HEUQm1LCVEf/KrpxnScOfE1lM1unbqrglEqP8UTQCSDAZ6K218S1XVl
bjgAXRuHqRl6CZrpNuHE849Uxmd9JCPg0485kJAfi56dNjhNj17gZhlAZeDBvyrMjBxqG9F+iJD0
yMBNuLjaj/69//OQBGc8wpoOt8+3bDMHOAcdMUAt/+mqgV05xXrfeZ9g41y9NObN5L5G9XWPE001
Yr12S03nbMLbQ7NuzZDUNY2lcuThs1D6SFAvNf9nrKbgkhtFYDBYIyqTFn06WC+qBcausSSMyR60
8fw9MjjVk/6wLhhWAygWlDdNIpNZpbNdIWTFy8v7I/nFfJ1JMgrSjhgWwonaLNn1gvk90g+OUpPa
MzZTYqmP6Gf/3nFEl3crLDxJDmWRqtAUNL8KSNCxYp795ubXd3JbWRAvX23uT4WEXc63nVd+yMMM
OapJy/M6SNJQ4yreI81aPTu2O5zc8qLI84zQpM5PvPBWk0Y4gvJI5EbSE3oHSHcAWDW6Lg8Izd0p
Z+ty+basp5H0UNm5Mjs+NisxGcGTbZNbBXRBUASNKjTayrHXt5kayWJ0ATWdmj/AjHpXhDOQUN1w
ELB80GbUXCTTrReSUI/1FbZBTns47Qtc98RCl3Zj4DHO+taXPk2FIrm9u/s+uAX7OExxDv8HdfQt
ijOGgoyPGRATtBcA1963Z+GM/u/TAilo7wC5EhIM+9wNJNA+VN1eZbO6firFnJ6JbgFZavDp1Ngc
T3bQoOxsEYwtGqqD9W3tA82bCkHim5TpET7sxabV18bdK8EWWgewiKkc+/vE8TQrkFogMupQprIs
vPT7nIqtWhSHp5W6/9rHvQoSRJRzPR4k8vxxUdLdEKSONUNQ6ES9E8nvb24cg2riJtUjh9G+cmvV
hRfv2z7Zw9zDuj9bZj83l7ruDiODxmnhNPWoeeL4GHi2PbNlTUhWueeAyrut2SJFK6QS3QW2BR/1
6JBHRkpkNF5VOypDo5+AkNW3WeHyM/pWlPuG8dWOqa/z1dNYLJRi911yuFvgOGUkVcWJ9e6DYv8+
wPUOWJCiRoN2TYddFZDKX/mZkCcxqJNVIRxXddTsUhbTgEIit7YT+ztvVJqGrbfY8uolGF9R49Pw
bE7oQ83JrPjRoDAKNccHFl8tMraEcL0tqhO1CdxKsmxzz69gCAowjNPRid7rNdxQ+yr63JQvskFc
YDySPNKvRd6fSWky2yceLct/GbWSLDbsTuwASZWOPOgHNgB1s+rygTv8Fh2LmgW/RXdXWU8c7vYa
GhfKAYdQASaXUoZcTqwDXyH0ny4smSTsTLTHa+Dcjg/vt7FF6jgOlh5lzfb/jO9fe5102F9vOiFL
o1wHTIYRbKiqKqotOgJJIDdQWsb4ToTWgAwkgHadkj1OshIRfV038WwooMPM46cEY3p9Sd7mLHYE
TUEissEC9bvHMxUc1U5jqJPl4iic6LZsgJ2hDrLq8UdYv8mymJlzvYfQSfRfF3s1+xOUxagMlIaw
66Js14E+pb72OyFwRgZDJorkdIBiXVIiwitblHKiJlmPiBECAs7QYlrfKDGZGEJJWbLoYY2hTE8h
F4npD4DK4v/+b2mif7g1m5sYbFcSNCgGcYu0KkAXIQ1FMosUNUS7C+hpdzbQd7GwubxNF4X40aJu
GXBf9bODA6BtyQyaU3M0qIRHahT7pLdSLboaz5SZDHi4+PNMba5BOYH4nYZGoBaawWqk2Aipris2
dhjkPgspkrg8Pd2f0VpTBO958KV5Qz6s/m15NnELpMLFRikyXHJnC6ht5sZCSM/ZMHhrwlOEKSrK
VhBIqliidvDYwRMkGGdJajjn4hYmtBrQG7mkydgJJpPY0+eQm8hoh3NoKHleHM2GzqmuNUTuWefS
jmapZrTF2c0v3D1V4uRxoxmQ5aDnWRl6mvRt06s9RmfqXOnDhoWKnPLDweuJgKe4DP5uc39gi005
5hPpqvnlz9xAlNAKXHLlsC5/mACseFUuPRXIZWAHiErXzUCnrY1U5bYAiLp2cCz711AZaNKlkgXm
FQP9h2FULy1xlOwxj98lKlWw6IYY5lS7MfopxhgVTJHkAJhiGwgjDvjHXqmKxVvRgeTFU6N/BnL4
uRUNZJu5oLe04QBFEF9acfU2kbfocQjHHJltZaoE87FOCN9y+VHVMt+KJvPUnX9t8m2w/QzjGnpp
owPE06qryvmE4t/H9uYzjGb1fy1cLjTL7+dTJ2FAbr4vFZ+nCyGaKmPIYUUw8m5YF17FwSE8pM3s
Y/Tkerm5Rq0RD3FmaGPXM6jR1/lUn71bFjDEhQoptFR9j9DfZK06C+penum4TNdbg4gBpFkPbJUS
Q45eg0HkhA7DMPyk9wxTx/ntYO3zTDm4vzPThnFu4fo9O1lQ+LQtQydTBtx8ZGd7K6bFHK5XX0iw
7pAWv9lebqKBFoM4WWkh53xJlhxZXEuKDf9v8RWauXpi/XkWDElZVvNs7mHOkUP7JqXvz/0s0OC9
XYK9DrT8brzKqs3VcrW3mEUVCyaEsHzSDSbKNvaoWGhdRYpfYVLtTmrZoMtOP5xgdR+4oqm3XUwX
C4P0BaMPx3UZdvqDzdlb82o+nnyU1GagB7I4tYcuPspOow5Tdv+oEuGyJzOr9Mz6F4Nsy36Abr8f
xLCNvIsimLu4P3yaCuIcn4zPIIbXKldA9OojfNT6kVRgLfYVk6b/VyLFTnebnKFprW0fhdzfI6PP
bwUNoPrhk3xzQx7fYHrfibdFfU4g29cEUfN4kvXEgcksmr8TEgwBpKArPm0MCOXqdwR9G/ZIvjF9
YPulWmNpRHU6rb71vyi2eVm8lzjKEUlIwIFcL2DEb1bSDkCuaPAXx+gjs2wGyI/C8yQmsapMAcn6
DhFf0YHJhkhe30oDgmBy7Zpl7Uf/8Qak/iekfIB02vI4LyeVkdsw9YVXX0jZVxbIXsyfqoVau5AI
lhJdrAHMXqi8Cu+CCS66SxGU4ZHsyhcs4ksrNRKCUTFWxkFtrutarl0jh8NAQTYZ3vVKExnUm6ux
O2BkyeeByvuddV5JdVDeNx+ds2v488Y9y907rrHOeXPnGXQliNYeU09ObQX1ma/58GR+51JkxLHB
wgNbSVVry1xQZITrCVCTZYD4a7A0flldAO3acE/dyI1xsLDSyZtwqmziU4EWnT35Xu9m2VpxrdmU
sT5mC4fhd2FQPNj5Y0KKV/c9MwXgZ3ceOG9PN7UyyavMV2mAHT/JSK8hzApMRbD00GgIS0eQYslc
6r+MCzgkZpZO9PP9Aqr5Pua3fUmM6dOu7Fk7mqU/NtJ16sIgecHkYAGRbSAFKHyrCd+hTQZV4d9t
mi0SsVEuKPe0LqBBrKBKQ6qrxOSBB/idC8xHRqC8brOIz5sUs6IgJeXqgZACafl0hAJOgXJgcWix
jznFs/HYnyOeGBft2jpFlTRyQDYpRw1hac3AxHP3Ft9lfxZkVqek+SUldI6LQ8sEsLrRvuEKPrPq
Io4/Pv0xNSyt1chTUsyT6cG2N+/gTRiOuxmjnEOyFc8og8JqL/p4onvgnb0RrYf0AFkgT42MhGLs
D2V/ssHnli1BLjjIvNoYECUkh8bWNEkelunz68fmhKBrCJLaZ0kEIAiLs68mI9RXN0gjTvQxpd4V
0sCDKPjKkUUrnsz/O3pVTHDhEofhSro38bxbWDqP7gGSHdKA1GwCVU8m4ovqZ+Gecm3PsPc8SOyb
r0mIeJt9FnkrsyiHrrwnifK5JtRYli83HJaqWbTF6NJG/PFkRoLeWUQKyu/A47q62d9P1yMXyEqU
sz+j/Yt8OHz+/VaOLSgy/0+H+/QpiO8Fn9pmr4GIszDdrzBsvMFzO7qVlpIoKE4rVTO1I7wm5SsI
mjhI6Nhh4543/G5utnz7V3W8J+oEgfUF5Pr2XDXxbf6pdwBIP1HFV5EeqsokzTtduOB7KpSJMMtc
pjeL2+yieQdYnn0V7QjWOA5E+hgxKIkt5Y9mYO9NzKReHrHk3sGeSlq28/nCd6I2xvqVo+MxpApe
BOP+4HRXwwQkXpTu5QueCoLJQ02qMV2kdAnIIDzbG7jTJBhF87X5pnMmK1vk4HZ3G7Ht7eo5jcL6
1Dqn8E+6pQYB5rAyH26CaVEhaFtKVqxMlxmjWsgZC6G2IROyeIgILuK663/1ucb49JFEwwcsEDB0
lZ3qT7D6ouJ18mRUKYc4FJf/ga559wApehKm5K0CFBFy67aHE/h7UKHMpsRyMJ49ZLCjPn/Yj7SX
6Tk5gcj/3pe/WkLb2skRot1+HBmeFiRbRIIYU59eQWL9vfgnplBlUHOlqDzy/rJGCfqcIRLjYvwt
jwEUIBw7anPFHOEEeRYE2Jg3mu7jmbccMwe+0vsJ/gFMCKvk42cliKYo60JQBJBVumkw9tDVzYb9
Up0r3pKlcZrJN10rRmzBnnYG4P+1rm+8Ags4QOYqoRtt2B/mVI3JS7Xoec6VnXC3K0bW4bkn/+yT
9jpKdjfcYCkcnhApeBxFESuVCvA+mPDgndj2k3N+8xxEaLH6dikM/gDPy39PLuuV3QoJCyEzuBD6
ajIbk+skenbpOn/XBbYVO7UTk/vE3CnXFt4ZJpXqdBLeqZT3FlZ+xoDe3W3qfprlM3KC4q3swlRf
AhbxEms55gAV9gQGg1n95wiNx9FtV3HnXJWsK7s1AX3zE2neVMRU3KdZ9uRUBBLkD+Sx7KCB1/yU
lmBQ0+2YPpq/M+/tywWy2x65UXbOQizMCD9xVoDqIq/PfnFI7XWFjCsvuf4sxXNU86uddCmOFcT1
POhxyNWnXZHMpXY7+Srbw4zsX/PEZTfQyphOKW+DCuPwP2Kz60Ksc9ZYfndMM7TybUbAdoe5QWPu
8MXeCWNfOATcqX5PNl69pghobkbun1ldjRMnyho2cu28YkfNGiRyj0pB6i8lfq9niMmg9D5NhFXX
vVmWPckFK3oArGAB15YbXBQq8h+KvgKAUJKrBy4PwPNctx1S4nvCsUlcjGNk9QhHD0wxbmRbhVzt
SsOytj1QKJ+aEFXt9RUhoURUJx0yi34bPVyT3hTBobHreW4FuUYaYHU3YOGz4/xno+fD8WvJ2Orq
+0BR3l9QSGUm9lNM3upL+pRscXoitRpU3Af5ZduxlUOaiRR+OxJuIInd1E5e9DNjzpPDNtd/inq8
1sKsy6TVPV5XkMTLAfWnTbOn0obxPPyTC7du/MZX8EjF+D0DbOOC5prhZSBwWkgJ7iv4uuDbZ+Sq
ZXqRZnDz1VFpVkzj89wuKt+qf+QAVAcsJh8YqkickBzrHgwK7RO2oBvHuYDQLY6icOCO+9jMuTAo
wLpB0ds3pBIEXEDrfoVb62s30KL6LcHCGlFQ4E2AUYJYKWxqoQvvSM7D8YUIueTBqK5BVhbg4JXv
a9fu1vD4y5maE+fVvJTuDODa6kK+s7MVqj8WqA7hnNobpFvw4LuZSCix7pEiKWMT5RxAjyRcM+3r
OPQWrqHoX07z619ggU12bRmpnGoWsZtpMeoXYZyOlTDqemRa+govbz3XI2OP2QN3YKgOgNTR8TR5
5ka3ZCUz259ZsXJuh03K9W7mUAj+MSmSaWsaIyYya21qQIAVvSpGAWpxFFp8cm3xxnlJccnRI4vM
9iebOYFzFMHPbU5C0afOIPGwZI9A4z/f+zLzWaPMSqgzKu6HeoF53vysKmwEn5eitZ1VKwwmLvga
jcq6PXZS2mz3tjWuc2ECC987HPzyGnXltDkdnpIqMQYU0gmJ8Kx7NBIqTC+dhCniLSlKGJNNuUaH
Zi/T2Z6pYo3J/LGjeVzt+cSucsAUwufz4nJAMat624S6l3ZFAab1qztS27Z+08o31btNP3n8hgi0
/hVzIhbkRpaNA0JD7uZlvkTXJaj4vFqzcvqXyjAtd6j7wou0cyMrdB66AX/LV79RhPewjmTgE4Th
4KQ7/9ku5Jx+IAZl5/NH5CKmQ+yUdqvYfKuTLSt/cUyBWpp9QDtwvaprBWR4cJZyVn+MptLtHkjT
Fqu291I+qq28RA59seVljoEiYFxDE7kzXxJEaFfz7bYv6EKpm7CodFWUfuBRX9odKyJn8I7aeoXv
AuYdmxu0l8RWySyi9KrTdtG2/kM3jCgE+aYGY6sID5IrEJtcR3ujenuALgM1ifurwX487ICaIOBf
uIYiXH+1CiK3chZI7gbY7wGSX2qMAfVh14rl3v9q02lnlfqi7hcblftj4/znnTlfqNMiGefvbFpD
IzQlG8aEmlp4XIkmVzherE6ckv4jrUuxiNAl2ubqf6lgeCIOt9efIZthMCB5A3BHYb+8veKwgPHl
2QHmVCQInGUE4sdlmatWwH42u07Q9hhClRds6UA30QDRfpX6kRRqW4LpkrGLJj/o9hjnqB17IBzA
6x5bcRlBy7Wy8sBTZpGekOm6aq75uwUpnffUf4g58Zf33S5wUsTjZ5aTjVkyYfPAjdxuH6tYehWU
01kcwWfovNcKfu8P1rFCz0dtB1/sMo6vMMNFHCJbiMGOCmIYYDMkK8oRf6AtjogpGLTI57y4O0RN
mC17wV6AhTEPO9B/ygTJvr+H5RobvvlKyZsrSxWQndlay1EmZm+HqlGrxzTsHc7p9WN9Al5Jw3lZ
KIXsXKUuz0iUMxz8hMm14htagZ75pU4aoYxxrF3kZgnN5+5+KOhcFJkN7IfFD13/W37WptIi05g1
P/JMvDGPi1YX42vCLFr3dfsizmjXXtM8kJKF9fi8MUI79ufOKsgsg/71roO+Gl+kd/qoizdEdAY0
KKhgwLT/GfgFOMA51WuHYaMzHOUGVRjocrklFewCOlxsDlLiQagjkpMQvkpUnbfrSYAVkDjlfhuK
bEEuc3t4h+al0wBakvrw58RGkF9Jax/XyRJOG14bPNYLQZv3kMuzJtzfuqfT6eg1pYb8RafxrV4V
uoiUJwAfReNKHk9ZRr8pIhGBkXrrhR86CB1B/yaJ3Vhgop3bhcb28rmpROESBWJH2Dpze4e2KCSp
eFJQABOdrQ+sv7bQug1U1gpw8L4GLK6F6LSNln+WBa468qWf3GdS9QrLh4vhttKqVyQJOsmausH8
LYv4t+himnRC2pWr7M7CA3XHXQDGRxn95Gd8zlY+iiq1fs5L957iw28BSZU0G68V/yk4+kmz9jMh
Ws2wToCwI9MIDUtRS9rfrySi77WyjTbYU33k7OvaBFUI9iRCyvDPlKb9PR0OBKDL0v3XjxUUq2D8
5sNx7XHBQwioHYmbfmA3By+O7urQ04T/c+36m2HJuQqkTRNYsSTKd1ggLwOsBZzP8PxOqjCSTXl5
RUlZVr5uYSLWANahAiJ9PO8/VvX4jTo9GMJEQ9UNULuuy6zbWjfrugDBiqYvq4MokQxjThV+rVFb
djkELXBadK9aO06b6/nyggk8afve54ZfQaiQO470h9NmaNJD6USbwyr1/VDUACGZTwLVlQNLE70Z
0i/awa6Ainav6xp78xc+U8qwTqEmFjwzhQuHSCUQnP1uF6jTUT7NWmBGh1xuZG8LiEbPD94mSgTL
OOsS1De1YqS0YhqtKJg8nYoFOoT5PlMBbYiLQiBbujpa37Vbm62gRVAXhGWVcGHShlr1d3I7ZFqp
GsAIxdrHF5qDJdZnGwRq5AGG4hIfbIoBBsh01HagmGOI1TGiGxs5p8mIsL7Pr+/hLL7A+KzMdeq5
JzzqA13z2JV0V3zMbIBHG4Gj89NG90zB4UbNGvc1BLeS9i20m6yjrjJKPrv49xEmJvo1lLFYkIWk
Xz0SJNCFmvVj6beKPuqYz4QLOx/a+BLlBVPlePXtRlthCtqRhuBad3mmB78v/h6HYfyCIFifs++a
VnsCw58pwOgdSNprMOj5Pxyxn/tZAfpm14ikbnnqZBf2Qm2xnTFXNOc0QK2ou3ywHO/3MDK3S927
XtKUjXOstfcNWoRFy7ziQCkHwBFawHWUEtciXgE/BxQijh+ELX9+gEpuE/hTmEHCFKZ3U2xs2Eus
pnnbQKMV1EUcgUwf7luiGJ/rM4uyHRxGVW46f9+X2ZJ64bPvNmijqYAABHIEXLQTsWoyNNsKehlu
FUZQEVssRzLoe8jgwu5a75BBzdJPMwSAb9LkMJlj/MwzxFwjwfC1YCaj4BArtD9iMPnMS7c3szUr
N19KmU1qKu/4cf4f8MdstL9fgwQfEQLCOOYUKwbxfAXjcfLeXmxRZSKjbaj/lTHERvBCeoi9/h72
Tbb9L0hS3v1vaFfdfCmN3HdlYY0BymJZkYrmVOFEcm9sU3x8IiP5eQ+V+jHwUhB/B1H0cn58CHN6
AvBVqm2ULVKSsjeb064jbopBOM3TevScPaHl8Ja39WRJD59q5TNGfiJor5qL2kl1oph4WWp+Tfpd
pzCqCeMyLgdWCUMxoTklflUHofgDmTXwAfstOkZrcLNeV9i5KrgyT3PSBPh9JaOUZik5RGzflMg4
f7wQ2ukQ56wkL7u9PTAsuglYJjHBYylg2eP0eCJhT0rqB0K9sa6LWz0FTo2eBGYn1QSLOdLgqhgr
4RlILtF5a34SQIw1pvYWIPPiNZAZiJVdX1/uWlZqBc/8K65pl0lMJlZLx48xRtBjeT9ViF+KNJgF
CQ3HIerAg1httW/jtFPAwugJlmJAbf2wFyZXhdpOc6PE3zSE8lYtS1HbGycEfbtG0jd/JXLJcmJ/
vWeFITiJ4GLOrjRdGi2AyP+y2DWEs6YKW63nMey5tPaeXLhBwbyflPGVZz9DShKMB/fneKSdeRld
DGtf4kYOQvJ9Usr5Qxt6olJtOlYVMp/Zg/nZbh2pTjWK0tFvevD6OBZQOn/UE1oaoNv0+q42ax2o
QG2K+umJ0Akg/0gUbCdJNlgcSgnHTipq0Uj6ezGIAxOiP9YHKvHBhDicswi5G/Zs4Q0Ks9miAS7x
c/CEFxSH+nUNQJeQKfiJ7hXOlcE1YIBfbY4rACBM7Lkmahd4FChRliKClkzChc+Lws8onD7wP83a
LNLUsH/eIYiHaAeNdIgt4ay08OQfoYWyXzgwOPf5C8SWP4GbsHXBJY4oGvqO9gVax+kFMPZLvYHK
ze5IWsu3VO8VBN49GEykkDdSO5CicljjNqgB8tbY2U3rXq8YdKy6l2apTVh30i8SMO4djuZ3NqtR
eWP6PcdmsHRVTbrRGH50n5GMJLwABS1FYJj3fTZFah+RZJEeZ5fLTFxmOoWMH/enSVnHMTmbr4HJ
E5qAFRYKDGauT6pOq23lRAKEALqskITfPhduYKAMGMGp235bgBZ4fpZ1MTKGlKebBeHiw6l+X+uk
hBO+EWC7NSCSPIqR3QEPet8dt0z7LzPNJoD8qDv3YkUS9GNqo4naBHoGsL2F/CJ+fAfEE3xSAoFu
MaYBDJbsCkc4PaFgd5RMwhhuTleVO7FIf/jpv5jL+jmoGWeR4vQezfgDugKZ0EvpM8SFQB/qCV2V
T+Y7EzlkAbNbu5cLSV/Ldv67c/rAfwWtvYdi6024guQKvckePVJQaWOEsFZPdP9PTRH8wl9ltVHX
fbwFk+UvcUpttdY/QngaOB4zmhC86YN7V1jsJhtLKZnVMhY4LSHY4IbVAg7YVRajlBY2ygmGGEpk
6gAYjNYeZB9lrltgLMeq5nJ8PgkNJWWPWZcvKPpUIf3402YTPujT9eLEH0H2gCIPQhlv0Ificntn
OUuS1Pg2gG6pgyFcU4VxZ2Ngp4m9EDTI3a1pbrs9FNlDHsd5LtOXfPiW1njvz6IYaFcKxqXDyPRZ
m+BgQtFSbNL3cW+9SpcuoNG3ExPOpA5UhtiookVXxBRNpgbfr0+GAs8o59sGu0dc0vAo2UDCxjsX
Zhj1nq0wL2NVO6DQa53OVtuL4LfiVn7sNW9ecBK5EEaQISPoi5mmBXivUkhYbCmAkPda8aaQpxUE
YB4EHty/tGcqHlPwHlDHfk9nkLrixpyhdu5PyuMCptcVFf3VNMseickA6Z0JTLN3+OuBxaTvv/5J
p2GgFZXXriW+zf9NFdg2uzxiFKrxhCRi+3ocNQRcAIMZlzAM87G71K0Ni9WrO6mjWiyPk2q5uX48
9p1mG/rVjT8IH4ylcwQI7Nflvsn3EbnEKptmodDZ+afyn5Z6Hb/Xur/HsGb00e4zuy8WU/vpcwkk
G5/fGUeYxR6WiS5zI/BsGLX8UiyOPfNQdSgeXo3msxHIE7ypHhz/lMdVwpqYJFP3Uf48Iy9XajlU
35FRMIhsT9plPqPQ7Yxzi33uUGabPt3QH1caHcjpo5wtYssfYz91d+Gk1pKSiXNJA/8GJC3zYaYZ
iJmAb4Rn4QCxOsNBBP6yMllc3fltjQ2tQUzSl7Hlw9kh/5XHM6u2MG5yAasDBwE0njvARyaRhG+s
DXMN434YOq4Tl6qrJAKwMN7KM+5c3tsLfUNFDmtLe+pPdGosAuEfLlJaJt16UDSWhbmDJA09ZoYc
SvRc2YgGQoS3tLM9ip6AQE0/BY205D5djn51v8rJ5X6nFxkV6C5Im8gzB5C2tTaKp46v3BnSS93H
6tXD9EEKmrnwB3cvu6bqSROnux2AkywOl31C6eZ+4s6V5/MmIQBIyCoOPLT/x1cp7AghD+hC/beW
m4QF9ncPL9emXh+BTYyXBLPRMmn1527f70X+66ksp2s5bST9y+tG82BfMKtMHWJjM4Vf+y69DSVo
Kr2QidKrfUyZXb/kFcXdVEh/nn36OY0d9No1w35lEul+hsT2i8FZ6CkgKxkBa7V0qS7wMlRztqAq
+MDF0y+HssSMqz9cySremXSNxkwj2uu181fkZHeVoR/tO2HIffE5yPJOlhI6qWBkGed3XDZSHhXx
/g+1rhYMPjRMmmrBGjdy+Cnis1rrjdpVpROXcGkw1WZ1eLuKlSdzb8yVbuoXO8aM9tO/tusS/RCP
iYd+vaYNwDlIix8ps3hv3Yi+KuSXUDJNgbvoHKm4lKF/LEWHQx5CuUitaYBScHlMqOj+k3KVMB9U
KhlGkID681iVN0/rTpIAvtRFKWX2SSmmf38GFBcQ+oUXpdz5FqStVYiSEXfjfBSQtqAzULrZSQeJ
ai/Qj6o36Zas6w17YloHsYVlXU5sxVHpYACCGLWHm5WZzhuVdJPJR1nmsbHIw8J/4oxptfXwB4Pv
FfdVLbKX9UyHSUf0heHCKlCbBg8thmiJr3HKfuLFE05+M+Af5EvAGPWXlO9v4Jezs0ZUZou0AkZH
ICQdTL1zUPlaa7RFBdXFYYmMwrsE4TSwKfFWncLT0ZDvg64xjSR/L8bW0Ubgu96+lsoy5IenSWEZ
99bL1wiG4bE/D+mptdapL0lrEnlh6AzHZ3mIj77qiUaFtS9YLgBiBrO9T5dOzcQtNnGh/+N6E8An
ElWKXT9l4oXQQUsJ2IYRywZtkGTS+dnU6EhgetmO0F8yjh6H3L7wPbirzBmHI+lZ82D6kjTtxMR1
nfAwjaME6sY1ky71yVCoch5ytxEQcxRCsCsFx6vCUAUGfsybr22Hkrv8SbjUghtfuGC5PgIv+eyX
SfmRq7mF+69Ns7IJaDlgW1eMJywamzPXJYmurwr/VXmOUGXIKv4V9vVCGI0CjoGEx1mO+8aQ1BEw
OEIrerkFRZHgU9nxffjDUHVHlNv0vQB5VYCqQEuC9QnDXtV9rrn8YE0th+/14AT+m6Xo6gCxLyu+
9APsnaQGZnxFZn5x+oOlcNObISayNbGq0s7QyUVO6rn9XlN0tLhbRoaTF2dg5+9M2z1SY2uNrayU
N2My+1ilJyMp6kduybeX8q9sYc3NnF9RxjaV1FsAs7XjyDZQv4sdOLv9P++inarXRZ5UwPsYWaGA
EwK/CdkK5phVGnjDdwj9zdKuFhXlQuNGYXl8IYCMTy0pDaO9gS9sLmhg7yEsCCKHzX2yFsG83Rz2
IBkLTb8zMvp+dkNu9JbP4UKEeKyX5ruCdYeSzMOKT9cZ0bHrU0a1InkM75NmvRxl2OeMlpD1dOqL
iVxjiJlP++RnJiOurJxmWuOerkQ7iQe5NFCWjvGU85k3sUbE5MlkKo/9MqiWWEYNk/VlLUUlnjCL
9wYaoyY5dB4RWvTa9GL8qoNQECLUMkExgsatwM2E5BgNS1dc0hMPk/6bwniv5njB/95txq4rT6Mc
G3FkV8dBZXDp2qUfppmtCO+Pxz16LMRrUR39k5oPFm5pb5TSkrR7/9YbxhaCArsWqmj4h38DYq7N
JIiN6bzJE+6BV83hjZTjDceciojHttDwHp20YSJCJWyK9WpPDn1gaTgGzA48pEOvTn4V9gh0trcO
nANtfSYl7WuaNwJ48dZTUPzgWfkAFffAI6f3Of1KhHlKuuPY/8Gl1hhqGQJQxO1YD8tMk009DuLe
Gv12VkBKIVaqRX2GCRk+HOliKtM5XXCUBe3N0AITQq7JGfUJSu90pQVc76nUylh72AgSF0cbP7CK
9loyHQtByO+baBbQ4WgOURDQfqGYhXagCDd2EeXtuS/PsW5RRGUowtAIEOI9NgnSlp9HGVBGKI8d
sLbutD5tiY9c0CJHre3sxVauiqRRLKxQMfVN7+4OWdTC4PEF6gFiRCCvqCommMfUZiKhmtVHohAF
TR62v/vj3VyYarQjYv7UKgbkvgsGI/2Eco4Lp4Mk0cUwDeJR2tUxHe83oSEfy6QtL2LG3bQxYZW4
warjRAsFGy/unS5Ga/fO7qRk7K4iwLIrTy4S1J1Aqi+OvgHrfI923SOZR1qM853EyhdHkNo5B3ig
9Y0LGh3EBemeugDqrFjz3Ou1I2zDZduuaKGgYFife0NqLKz6suQkVw0EWX8PQAKLRjvvEIneFseq
cUc+JvnDxfgI5KMt19qM3cKlZT19aPLzVbc6Io9T4zkzhSOlXZKc94SoeMS5jHWyJzEhYyQEOcyR
uhd4AoUcBHXS8JbsSbKJi562juoN1rE6C46xN4+dwESMY08jZn/7jRCNJqeiO7zmRjKZPZF8d8aU
LSR9ikV0i0a5UbtBQGteRbXrPCoYMYKVY4a2b7QqlDyDddZVQfrgCKLTdY6ULb6ZKBjks6Cp3O7Z
Gsh9TasVNQ1cJLEI3Z6ppxCo5TK3M45Cml6ASyKlIReELoP4zlQ0k7pSa8EUj2L0WsTGeyvXVBcQ
GlAEoHCqEUFIDdxI2udFVSXlngTEPJ3KU3fZlw92FDQAHNsXT9ekqr+CD1ww8+OePxJKOjBAZdqu
HAV2ir0mp5QkUeoEiEzkXr0Wl4X2cmIDplyZWeKMMLSS9GQTG5T1vpUpmq7mQARPDxzhF6AkG0zG
JdIXZr9vujAbGIaj/awV6yP42GWwn8BUQrT9B0+vS7+1cP4Ae9btkCpseqzuqApvcM4q9h2O/CFt
VrgK+WsXzA0axpFC1ScUpuHiDlG534uw1vaEDXljG90HJMC3XVCznzTPZB7J5CbnBYi9mlxFZ/b7
v93GhAvYzCtpeuQ0ZdQZXhmQrk7xhPB3R7SnfZLGpyP54748QoZP0sWD08OZiTMQz7l/nceNHPMf
RunL+hHs12w5dt8uie+/k7MXOuhqpBWZyOV6LyvZxg/4IFcirMECE8N8kZugWCx8L9It0YFUG00I
vVjSzSSoIGiCVE2JGdP+qOhJq3vQvYtffIA2LOVeBbtVAvD2wGcPjsfhBfThHJMIH0jyk5h9xz2i
q6emLQKWIyxbHazZyQ7iuTMTBat0x1XjFUkAbGtjjwjeuEKGobEIT+GD42KutkVYzuiwzS/7+rWQ
eNT2+vG/ILrE2ADeXILsxZGoQNdCXz6a3XamrEkyoBGgAH21Hh05dzINFPGrIVrQSlULmUum7GXW
jbdvhtmrzMD04APkmMnoglB+Y24ctoCSZ1lRQYVzAvIE5ZLW4uxeqAEXqOyrjQCbL6s98gGCq+oy
kvY9e83JnSnb4m1DQ8AmpD/nB+6buuaSzmnLvabrpow6unkj2foE00NnUSg6uV/SevHLw2SrwUtm
1Yf8ZC0JrDpYL8osvhzXSt0x2++6MbX9+LNX3Zf/aFzcwmZ8Fe4eZmms6yw+0bxPKtkseOcN2Sis
Qhrwv/roR9nKT5YhGheQcOsI13tHQt4VBk0cO+weWse9QF1NJNWBJf181B/XejNAYS8s1b7jRSlH
CIjZgLQDhgH9NA1tRKyvL+SbSPNz0afH10M0JX5w8KwVopiha7LEA5/Ezu2bo1XkdDJKsNNiY94i
YFpnkEZ7077xDsgc0kWobSvxR/d39W+Ge+FBy8YI9yjynsTPY/cJjpz5OD4wW7LUEjtJP5K69+gw
sX/e98dFcMZKZX5gd58y05yzuZTlCsRP/u87NhO7eX9S9MLh9PdcfZCLU3GTgznbuJsI8mAintRQ
MUoSlLCo35GtCiEQTXiLweLqrnKlf1AM0AKAoPY2KIPE5KgPE01TXBER+w34QNHo6dZnGBIpAbGB
9/ZGMR6gwGMjXXNVih4aQSEFTp2jxK5MG2BpDaSzzpd+y+9qGGOutl3QAeli+J6DzlnuoMGG4x0/
4WH1lfr0iwGia47e70CU/DV2PUCjUbdRv8YTzrxmAvyBd6a3DXRSG+ahwlnePwlh+qf9N7rV42S9
TYXibFOyIy/mDwA5zj3F3+rr3FaP275IbZ0/KFeR7bCRu3cFvE1pbGPZXMdOuByADNUJ8N9YbVFO
e7Crvl5iIwYguiCMEJL+KHl0eHaJlyp85TYSjtXM7M4qEV29G0V5pYrygx5ilJc2pl0ywc33KiYy
5DMhDEVn0TNUAGMeYdyaGJDylkJbTh4c7Pl77e3Yo8Fuk7W1MyhthjhFoDM3G61A3MbfALuL72M1
NVC9yDgZ3v4vn4BslmA39zdhVB6Ixq9L27uY/lFxSLcwpO6v7N1tMs46H0gW5n7S31WXNRApS8Rw
0K9+xN/b5uQQ7SCXqzpsaPltiHZw+squa1T1tKElezL7axEd6tuhUaJKs8Ink6xqJ+NV9pD5PFU2
3QpNXmfAUCopLepPOpbyL59vc0kCQGNQrA2iGNsC8fxHIOMq53Pvq3JkgIKK/TZJ58gsY9BNKyQB
Ipi48LxwRETIsONNIPD4cGibf0h3ABAPASTdiDNiE+duJA/Ne2nI6UdtmhELcQSKecv+Dc/RpIAl
/bBFmm6WLQYd1TdBqP6sUUA5DzADSMqk960P2U6xp2fQyQY+TAPjzhDbf9PUC1mDXoKCKdafwazV
t1q/r77PycOc6F9E3Dac5mCzUOQwRdD/xOpNR7doPjWYC+f7glnMDU9CEVuNUuqVHebRyMGDMUTw
0DF607vnUDA0mNw+mEIJSyQ2Q6LrUfS3rGBQ2RZFnnD99m41CLX1iiFp7vDpsHtI5YR7JLla3WHX
4BCpuvC+FDMKsYuD2j7C/JEWWiH1r0RuTUz7G+FKN9nUQ4T9yVj9CNk7P24NvlyMIVNHKZLaO6ED
xkMKADyEunlULm+8KSewk5FiFKCW0b8CxArVQb6gkwEWEte+o4jRLlkHP5xh+3Oph1NNw18viQcj
WCZ2BTTFbBmVtv4mHwRM3n51EC5R54wlXMO8dPmXGyh+5lZgxyhTiDR5r1mvRKZwroZOgxcUhH+Q
ZelUWo46JMEvA6lDY6NZqLhv6L9W0teGLMM5Vyx8Bzy88aglXEHjdr4JP/C/KrVw3DE+YgMIGHZP
QR6zRqNpOGA1xD9iuUkT3HOx5h4sjaAenena90AT3PwB9dGDFEosiT4aPrz612UtZI0/6ICdtWRF
6HLKudv03/xAIkXlR2psYstDQfBXiQeK4JApjwU65FFhHRAuo47wAvdTUhc8rNilCIneKDaNNIfb
mBtkUjhEZ5F9qRCle8Ux8Efvihwjp0KrJdywMGEVwTv68n3Nk21BgSNMYMwKQIOU8Eb9b3XW0rV5
kxPmvc2BGyyXKL3SRoZ3MgaartJw4lir1M8+i171B+tM/H1WRtdwhhRbrHWoUn+YuqqBwhdFyLtc
chAYGQ6Qe8UcnZ80IPJFj10isENlD45eXM6aIf+MFEGI/3gWUbEBkUpe7PMX4UKjNyZtY+x1YgDE
4zC/qbx0wTvYpuHiBLXRnpcsyHPtFYjhlCCnIiW0ImOdaO9PDopCDCWay9RRwpgp9/AQB6gvvzBb
HlsumUXX0YPM0CfY76//xX3UOK2RldOB6tU96ie79UQZZSRTB5IN5iHFV7Z3MUNYIC2/8ue+MSvE
g12YXh0EPmElZstC+Q1vBi5JgwLsWkZXBpNiX3vBuRFKW9NzVVLA3bOk0o7+1kN2O6TbrBUb1MCR
ZdCrIOppK0TRHDJ2uWj+IRcblaSzhWZPP0YXOK8OJ3avVRiyyUiROxRi2HwkU91pBgTgBMIP6gf+
9mQKZPWnLzOr729Px6Tvdf8lc3vToJmeJS+PBab61FV24fDKWIFE2S4saenmwi1noCSAeOdEmmTi
G1azLsSCE02RupHw4yZ2vnIBfXdSdi3k9EEaavO1iPWlTkQXPb1xfIz7n8wi1y3uA3nMwlL2QWK0
MUJx/N7ni3qVON59FThpGcbpYdGs92EMqCvL47OIyEBt4Kkr4WUfY3Iv9l2x4vS3VXTb8+3f7SXl
8vXlHJjyguz1wugFx0jk2Zvry56UV1Q0egZEE2EneET2O1LxgVO7MrJnGwUeWDiniEq6btDlujPp
Ck2h4j51N0PUzqdRuNOAjvF81Shi8G0n7wio2og3ng5mwekAL7TA7BtvsF4wvwLGFdp78EtfqoZD
E3CxPCWHueCB9Ul2TjIkSGXndhURMY1I3BcbAT+bErRRckTFFJ/5rDxMVKukNGYDxQjLaqhmLWrV
PoLezELiD61aj0Pz/RCU/SP/EfDtLeJGGNjoxVGgNVdPd3B2YTP4fYTzNVuaaSEvAqSDjxVzEGeS
j7FcdLZ4N0YVaPLKqVxjGjNzpfRPp5AW5B95nSWkDCAMsKYOHAn0/Rj2yAlZ8JLksC8gMTryG5M2
74ozprmSp/T8zo1XbT5NyHUCAxg3Qn8l72Q8lnxQk9uZVbHKIyQm6YznVOSrxcrpwyjcPodkP60e
NvPpPpvhtyhjI3ALCcdEandf+rXgJ5NdIqXKCPwmAVmXN9Hp3E7rLAv8zsy5aH+D7OOG5g8MC/Jd
jxgTv/8/9oEQz1TsPb3OgwayN6l9XNPcoGM8fwTIWINYEfGPuSAAzd4FOMr7pBQhK0d5qPfbh9zI
JjtOP8PPCdwOopZk74JZGGZL0VDoVXnslFPMklEAlsusbtu62BvLGKKkmz6Fxl49/JfFfz1gou4o
qcEyhls06VByBV+qz9A7AoKFr0WaAyLZvfhib5HmVpX8+e+wd62UkaZ6SajYdV1XUgcgBPtuVUvO
0lfxGY3yOdlU28kuj+fJEed+WSMyB59OikwI6HK1rsnVlkYjs21sfdcfhHdqV9Kkyai/uKId+Qfo
q69qWg2cpyzpxcv18R4HfOHRQUOG+3g+J1tfBIORTL5yKm4W84JnD//sT7Hv/oqVB++0gI8krA5b
7KNhysTLHbp9mA5WIcNIuSG1ea3714kyrvZwqmzmrXNHGeoKnf5C7tPNC0nxjHlc4Za9Hw6sW/Wj
g5bMHahdFNzVPvabK/BHVF3hBEI3NTtNjgaMq96z9TH2OTFzo7jy+Nfs1/A1EBS3btQroq7294mV
kbyGuq7/0acCl01KQ4rUhWqFA9o75DUVqNZ9PTKpbkmCg1WjooAP0TRLOdgZPYSyvKfngv3J9Lnz
onlEyM6I2PRAmev8yTTilkKVpFj733OWAf9hKXddIjzTDRMr2/ukdUg75QAPaEeucridj9pr1N12
/owWGU0WGVLE7oVvGbSkwQACa/mB2DVpf6Y3pUyNe5D/0MrSLIKEA4/+m3lp10de+EZr5+QN8xY3
TF0dy+kSVKi7WjL+DMfq3b1NP6jN+j3yS1nMi/QlOW66m1Mlfqlj6Io47nPiTFqDlSHRPxaCzsmY
oWXHxuf8yXtPYy3zOXcLnIecF50nFV6yHLc8y6FGl+3EInRSYva5t0k4f6jAZ2xHxOCWNX4Fm66H
AA+xjLO3obYlrURmu7Y0I7Rs0SKuKBtaC8kcpI4uyVzmgTqaDKn/JcwCbA9n442RzH7QNkw+ZvD5
fvDZZeRE1Urqr+SWY+0npMN0NZB1RKhyGqhqatHdxhxi/lbar6i6qx/V2y6FNIoQVFZ/fC3m3Wqq
MFawWmRXlUa9qAaT2+uGemLIxasdiL6twIY2hfjogdGqPuJet0MJZEeV6ohO2f5TDm1U3XyHq2fU
0A/J4lqFTv/5hQZrgbQEFyrfLfwzLe4D446QNcbHq+HmHxJ78fge5dr+LtpGrnU75ZpewsFCJRrz
6w7t+IQm0LX0/Qytv/eLCCWGgOTaaKGfEyIZc7J0+fZaC39NqMq59n1z8CIH5IlV/MJ06xqPLLRA
Uv6Kz4IT1ynHpZfiUaGOQalbIw2yfTdIVhuMTWGrz4gAQbEILUeuRZOBmxJT0SA4YqseTqsMvEt0
42So2zFHHyIJTU4RK9q8985ElCExy4vf6zHo/X5AB/WEu9zxkrGKwVBy/DoqxyO4YnsQx13Q+Pa5
vA+eVPayXKCs4XlFLAwzdCQoPJTJ/LeVN1uOIVVTNtBBuQBi5V3ZakSx3NdxbZrSBJNRkrL6Jo2k
8aJGJAqiVQXDIA+ygl/XkV7o2YTy3KAYXVYDJ0E9gDFQX6rBmT2n4GIDl/vRx/HT/U/Bwv7YpZCa
FRGVs3AxhltbdYdyFgGoelXVksPckfLStrl1UBnT9kWKHUNRHn60x/LyZFZVb7Diy3NpPZZmlRKF
KB3mn40zZB2IqtfCdCqk9KtejhnI9PEdRKdlGwolbcOOGNCKHEnvGvoarypmQW5+u0G9Q/Cg9901
khsCU+YXgFzhkWX06yaD/xnW4HG/VDFDsOwG+Hpcz7anL2lcXe3ickeSx4oP7ftDcMyQTNWHxEK2
LE2EsJ/BoOf+ACr7HWRB5BEF2GGzygGcwMoG0gviUijKusa7ghurxLRlF0v7TiTfn06wMFo6S763
NQoNzPFe7terkNz7Row0WLeLQBdz3aqh9gyf8lel/7WXgjTGAUd7fLWHuaD3gPDrzy2w6XnkCWQD
cSsJbZ7r4ckBNFK4Dqf52WIBZuzKYh3jGjjxkZf2nnPc67qDRizkW2znPz4TnSt6YqG7VCWWK8Rq
umuYIylDZjUCCxRc1HbvkrTaWeqB99QQSgiay9eoI0dSu25d0AWHf8LT5wZpW4YdEj7CVAusurlO
SlrOBur6BrLMm7LWZNZCKzkcJBS+mIcaayQdGFiV0s8d4ik/GU+Esfa9FORn3lEIkBMLtgjjdSZ/
uSjjSZgqdAyiUvzhsghbDy/xV+GDPGH6tM+KO0qBp7/Livhn16U2ZTyP+lRdDZiqY5Ux1ooEaH71
T0WGScpfY1t4LEIraCx7z6pyCaXlFB8mQmsjY896ywjKGkPGuYnJF+lJu1VG7eAJgFzbsvPGbX81
wJ9g2ybJ847mVRFL+a7sV2N1/HlN4N71Zv2jjdGiIxa//i8tlBiV6Igxj9RW1UoxzbIfhx8nzNND
5PUTMULyePPNEMZp+nWG6efu8oqdXTPXXON/T0XdWqH1KjRQm59BmU71cIa0m4Hc7KPnUKkN3/es
0ZRIq0PcQKYGB+AvrqMmdhboiEbbnLUHXSC5oWnvHrcM/BiSfihGFd631ZvgHK0jti0PJ/EvGUgz
QpGvoPmnfnabudUvWoJ1XymflwX9wfvkwKZ5f60/1f3fBYs+P+kZFdLpg52vOyi90bjk8RSOqDma
NT1T+JsJXM6lbDPx7RAL5lyDLBjR0/WABotDeUlx634OlWc0xT1dvT7YwkMOYTHGmZTkUUvSeZAP
/uzK8KgGouk6hK08O9CZVXQDAL1lBUMlGJwsVDkkYeCj++iBIGK7k8w/cll2pJYV+46POPxaQN7j
Qfp7LySJAyjD0alXAuGQ4jw69Qvbf2RMeQAZ4aCpo/mbDIh0uWNxm1FXlj5bf5N+H/IFlWBzn7sM
KnZ0eeRGxS9Qw7Vk4jeK4+BkNzJ9TPh/z8YZwQwfyiJHXOdaFmvgB0SLeUo+wdn7gYKBdEA0rXBQ
vQma35qc0WC0/QVN/D+UZHN/11BovRJWT6fdKUSHM5QSLsbqfSdO665tzHJ1rWny82VysW5Mq1Af
SikBpO9uCXzpFHmSX2X5aK5BAtQjVjl/hhHiVtiCPhQagNLNNPFv1jGiAFicdQV2fx3kiQZz4rEE
hK9wanvDxf66UxeTU/WYBztAhlcOeciH7D5SEy24AAUPtBV3xJ0OWQ+PIpeLzkAAg2/ljwFcnAQO
gdi79zFwZNFGhv4rpeN6weQVnZPy6KIMAoZ0ZIeCKKUi3y7PHfpW6jO1Rl0Ux7ngfPWnu+2qLPJD
irIoJHmMkjMsBHLHeq0C5KDuyeA+7rR0Mjen8bcfVkFI5ad+tbukTCJ+livAp3yStppMp9+p0mJD
GnmHAxqMmJI/wNJOsAzLTNdFhXQcJjViUViWuDzseJHe8VUYKApf7GrL8GCo7oyOtgtRmXJRb/e0
47P4evKNTDJtQko1KRSAq+encbxMIxYsn3uR2TOaqbz38gwJyGVoCRdhNf+JgceXqO3FBUV1mhGJ
qurAo1bPhWA64W+j9cE1aGzH7Ind2HqEmuf1E38NfZTV0EfXIMcJtwT3olQB0Zju1ttDNVRVBrRe
/W8Begda0Mydymd6SI+x6XLDCT3QJIz3a8kw3PlwHEHK3XT2vqbnKlllVJoG8tKCjilUzkPrvS/7
D1/rfHpa6h7pC5oZNg3cTppOg5UECpn1x07djMdjKptHIbbWrbvzxb6tn5ow1ZxzVHllO8lBQqqk
117E47r/S6C+j+aveDjJqXmMPwgZ5Mz4Vu0Uu//GvrQN72R8UoAVTjtJY9XJgsjQeULjtKSpTiZL
QWT5Scl5nY9oPXXt7z8SqoQ3beSg6hIkZ5BB/0IqClf3jHKsbew7tn06hafY1YDGDXP2N2IAot3Z
4RahXj6kuMQhPOBpADPO4mNhZ/OHBNkOWROr362OotT0TdrIEPSjlSZ4ho+ujWIN3BXLdx/cKTYV
afzBcJ4yR5VnnXf77iGYu7QgYpE/EzXa1bWusqpbHTOAHNxqMmwc0dXn+k4pS8+mSH48Fa3FbCgg
eXXGz8a429dOKJdHs4Op1Hjy+UX9kQWQtm4uqmEWPRL7mL+JOcUCN7v1IWL+ms7vFf5NQ+U31BqG
6pugtkNHHNjhB+guIYOlY0RsWh284tzAXDGkyniJ9kWQ3fr6uqc4+uSwkiFqLJRrdWr1YkL4ny9X
wNoHQz7waif93Qm8qSGTOVr1V6KJ3VesTj3Gjs3SyJBCPb/k8Tf2du79ZqvHXqnz/DDkaiotMsmR
PX+NjqiF4WHesAiTlYXp387OdnrY1vGX0cvlhAOd6LcKh+t3pSbhcrAt7FUWJ6oIFBXRrxd1rjeQ
hR0Okga4gcgVGhda64G/G606P6+CZNr2rM8Rdaqfm7LG+pzbSZsQzNoQ73D4CgjSBKc1of3PNzXr
NFRLN4bM2rLiibWo13lnfPNssAn8XSyDpuEwpRcVbFfc0K7U0BjRjWGP1mnFA4W5uPDhjF/VO7iC
kDiJxnu3uGojOL3gl+oJLvKHxwygDJaNgK6bNp/6Al0r6lQs/2VMNadE7d/llnbhb9n9eKZbbywL
x6xlLvYSnrBC8+88SUta2DxCJT725GzozY3BlnEnbnFQ0UuCYOAVR24WYon81iN8UpTDJU3pssft
9Ndu/oXB7hU4RvpZgY4vIK9UMba11L6G9GZiGdk+XAjRuU5c3ePy6SK05MAw3vgjQG+oG7HBQnBJ
brBvw//aL4OK2+MVgvKm+hPtp3YVeuKefJV2br1+tA+QpAa3N74dmEzQnpHJi3mOZu8JuiVUjl5T
aeyTdxcxgOVMYFa2GCZbvAbZc3jESQwCKjen5GUmrfKnGF/lHiLZSTbIZV+GtDEFCnTrKXgvv0jv
+8iIovBzloSPRVqsoLK1cUbu3wYXYZVNjlOO3Jx/RseihRQu/ZlvhytQ3UeDhCv6XW4s0nHafxxG
24pg0zXuzQfrK8ZFYmO8Fk6fNXfKchp9C/bjL3NVxTonc5QTa8aDRtQo+cj3rBYSzD4HPnPYYiux
b6z0BOpK8Hly4pezlO7vU99gobyoXsWFBo4KJNZ2cjenQcBEGyyVnop1iHd7oq8jzuA17J6p8Xbh
O3w4qPHEERrny+uNBw/5vtGBYO7QmlNqf7/rYLwQBf8Orc2di6q4kwMD45MbXz1wPjjHnaRqr9pL
e2yIiwayma/VrJ7yK7sxNdym3ce6HaxcFLGOhcEUuX7K3yg0fjDqQwV/iwiIBBZdNKL2DtoIlSfX
Up1mT4ho4ONkv1h2pmUhaefWb4cqsGTVwPss/Ptofx03X1AfWjny6qRsAhnycC/5163P43iS+mxG
vj0qiGUDprlvOV2JqdZgezj7yfHEkzAWf1kiRN0PNJOOATF7Gzk9ODPY387uv5juNU3L2QUCuIr5
pzZfK7ExXvM9TVizJ7AFFrzzDznpCKxeV5OOgqwIth30kGbqUZfC3XKPq2Y8QAilWQnZYOSfhNmB
hSW1/dOmm8nlPcEfamqgyMDbE/PnUB414YkX92hRVNEka8DHUBkv689dtBdFzTzLrCvi0SalgDmS
53MwHHrJ/WD5zdc1WtnsXhlXPxreEDKYPNAnVi3eTXyRQddrY0wzJE8iLY/g/q7hsedL4H7lvYRA
GNifULFxhGhnuOdDsS2irxxcKbhU4KyqxKW5249WzPCh4wPPfxNVLKjcP/Ua/E264acIUKeYoEHm
+ThxuP3ksG9pDyeGN3/hBsumuVTO7P2131T3Jaw42FQ9BGZct1WioYN2Uy/LhK5DQ+DkEKXMBNIw
Puexz6LNp+H9OlH5e9EqujrR1pRkO1myQIS4icQJZirCfB+fCfkrl+Z6V/P1Rb4TQsUpKjvc8uyq
FYYwqJDt0udZVyledKwpWv4bulqe4TOcieMYqXVB2epvEKN9SeSxOYtNODy1oz+osT1xzPBFEi7B
wFIR+FC5IVLoQykj96VhIBvEwQ3dxvkLa8y0+jJ0lE5dYXVbL6I6bhSjCM01iAjSF+A0XEHbH58d
ehXreNKG2jIg/vb1b/jRbegSRfd1KSwMMzNnrv2csEZBuHK78WTSni8bbTRnogJnN/FmDbGCiywL
IJhSSOMS1l8fkPC/r/yCNPX+qMYsB5zp9pDx/v24pGwUjVkL8CpU9aIDLLqp2m8Xm/yvq+LNScoy
FgvpVFN9fFHhoi3+BjkDBN17YrGcDnwaL6+Lr7E/z3fuiMDo7rerajIvDD5R51e2UE7aNJw70wAm
0WbbjuqGU5e21dKVqctD1nh7no/wi/lx/Pfalc3KtKudwd1A5EFeQCIVZcWy92NhYYjbxg4tDroE
q3xzT92hSjPlZC/RpdCakRaD0KRVpcx9WImS7fq7woGUzT0/lulAB0xn5WSnq4P8wQWZT3UlAJ51
jsFT+ODUUEfgdH3wpUlwy+xCvC/1KiMnoM0igBtG+q7qmLJIXT1wIqtsyAxM5UfABYEqjFsKlfv1
ADrlvl87KEUOL9Tpd/L5OACJMCombBSisj/Ayx+iFJ4crOjMS5RJdDRz2rYP4fa8l+0dHv1lSUPz
2RnTAx+Ue2crLED/jOCMfOVBKhYo0h9PG+0+AwOLk6BtPTA9R631WXkMHQhSgz6GsQxfrc2zsRQP
GpwPXURZapcXi4xyyXXPmqbvTyhzParm88cJ4yoklqn1SN9AgioXhi+CaVmXy1nQKNCL2L7Vl8tc
DoF8LYStNp/EwS0p4ZsehksKtG49kCFDhhkocr6ADV4wPQLo0QlAhgyaEwXgw49ub7/ylRuGEB+P
LFTjTPNI7b2AVjgJLbiavcS45LZeVAX0Ru+sdkYMzhpZm3ANet2t7KCjZ1SskH3W0JFJ6zcTsDSR
sG+G+QhA4t8YwlJJ8qLkFzVxYZC1NSPyJjushACpIyJ1EgHDOn91uNtOpmYswNtjuBIHwzvVJ0Mj
e1KfyHr2ALz+N3x2uLjd133biyQEQJtzq1J7IY8duYjiIko10+6fj5FO+C6nb7ZfY5mGZFelHB+1
wW9Drp4woN6E2baIjDJfbCFAQ8mPeAPlgnBpI8SALw++iRPNktQC6ulBwQoY0JFBvfXTL1lZ9dGW
/sWP/yr0RdXsrkAOr/knxU3vAwZDsIiE6drtFIGt76saDgyRQxrhERbDqmFdHKAexlFeDxsNapw2
WOLfMVtUq5z4AqhijhJohklombhhZ/DvG7mqQThwJJdE6ALEVAL2QiJI0uplxdsh6IqwfQVG8uhf
uOz3G9Sot4FDTBrMLhRFKaeKX2NDPHE8y4sg9OGAS+zt/IUc89AjRTIVAvRIYzqcBaPthi6BdGr+
KhjT7oWPuJr8xYEWPeh9zWVF65xuiVhhNuOliv9qzrzzNwM546hhC/vT68A5zovPSYs2pI1Xs6bS
gfImFSJKTNpyjmH+9axy6t1bJtLyMSZlt9P04dT3kZUG0dG7liveN6PSl4OaIQKyVtzc2PXouU7z
aODUwlbzb4lss+qQkBk6ttLbFKFjbP95D5ASygOqmUvc/hIFpbs0k18McLIBFwl9Vj/3Z+yc+/kq
nDVeiu/B+ZIj1aPIigvUbth6jW29FRcpOugbI91xv8sWeKn7M1JOIsTpnSNKUvDaBziIVcwTry+7
Frc9xuxwroxe4XxvIo+b1Cpj9gDHq/HQeHV3/rfe7BSPXKNq2jbxnj+iayGBY9uIzFyZN98MkGvg
hUcVlcHzAEQ3tVEVohLW3mjN5QIkNQeZvXvH36hB/N5UGavt8XL7QOAjTwm42u6J6CC1K+/AyXsY
d+D9g3iTqrVp3TQM0U1ti/qTRrGG0Qk78MNzlsjySiwfNtj7016D59imnEQiALDtLivxMKFWp/ZB
DGpAXBY4XpHDVK7OhxfxkuDjssMENGFVlC/5XyKxmptKwZAFkOYjyEl5T51/rKyzxW66k3jjScYm
tC25KPv2ZhGHsr1egRkwt9UCHUIlx6qN67Y3qNsE3N3b8lw9KZPrK4hAtRCNmjsf2J/5Nj1TBohf
DWrRvjCO3cJXAQ+mD9QpXZGBNkIQ8WLlMp3brBd6CH6FSA6/rU1enXztSRuGIRH0OiQ/xQAz9NvF
Rybqmn+EKeo9+KE92RdjxDH7kqAryu0xqNttIlyuWR3Ozcw3quQEZ8OYKUKjChpgpaiXllP9BIuo
8GjHlVw63lQZTeH0EALRcTQKUGkt5YHWbNNKaHWA6ctMwlFiLqkpvBUbwqEnJmQF18nuM1hn6USN
YSeY7bK/SNrzFZv5oKKS1/xBq1dgi2t//vt1WjrQVBh9HvEL1unez2fMpTJ1HoA2oi01JNZwBFQ9
a9tKfvj492rhGZtmSJiKC3zh/zClrKuz3eiim4jNVbAJBZgq10P939bOBwPtrzE9MbtKo11CTFRD
NlBaV0NF5WfU+pZQs1MZinO5PSu9bh2IbbkH++vZIuZfrc9OdM1kMrM6gLk6o2n0PidHc6+FI2VQ
slGqwqx8eFopCZ3FkUkmBCAGMsCClRQ3xighDm7LZ30oECoyWnvm5BaQhj/pjv/v76wVXVTCBUpx
96lgF0vTZbFH3Z9jlw==
`protect end_protected

