

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
p7OtZBpltt/h9CD5IsJBmAQ+bQJxazkQVbRBjNJ7LWO+cgudo/XA7alKhPL+qAE8nYmt8n/nhFV7
1FHJnU9EmQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o0V8lbvMs2u7Pr48iEK+soyjigqgrrzx5HsGK4k7Ph8gI81XWNRtIljFPpaeGwucYu/H+gPVGgh4
LxNZUBJhgeC8kZr5P0UJ497gR4WHGLQSo0hvtVYHYDlrxnVk2S/+il/2gMAwvI5YF/lKiRUCJMb0
2mL6cpx+2git922rE9I=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hIqrLT0Q92Qul/GeORaSvJHHAIqLk6EmPwtSD3Sw8K7TFMN/pzvjFhA6g78oxGwtYju17YRUOAPP
BxWjMZac0YPGSx1A1AySaj/jWf8/sND51mJS4hxixMPKgd+iJln4gROFDpToYNAZ0eBhqGsKoRPf
Exo4YtwLGOksTW6jkb5XyScrMy9eg1uc2W3HXgQfQg9hr9gpWWe4xqhKUCFXFb9eiIDe3eaUQ22t
Qgz9S0YooH+uhgkKhXgOsKoG8s8RO9q+oyyLd0ANkoAdDySOy1H2+qKDhuJHoo8oHgkWp+t8x1nO
sbVK5ZibMfLbKeRbGwFkFsj+EKfWfOy4ck2AmA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
O+omGGx7WVLIBeJijOGvFCJZ1IO2vxCm1x3fAW3H6+gw883MkRTmRZO0ddVzk3pvzQaBPeJUDRsY
1XbF7OM1C/khYSkVv9TjyhihrgNNT2rgkTkWtfQNoOMnsmtYkK2fHBBMyNXzHPZRBh+2VgTZHxjv
olfJ+wvlLAdf8BqZKWo1gutmRCut9sBqwVpKtMbEKFGRBnt2pETIJcWkewW45hEmUxoPlXpgWrRg
sESpeoKuutTTWJor2paEV2RoktNIWs/+x82raY47L1AIZ3uy3vEVemolA7/fyBhQXHdXuWEXntN5
bzesBXIrWmoZpCMSf+IISz8dywoKgC/dpdCKGQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pc9IPtPXrLLm2VmqSrmdhsB2/sqloTepqxhS9rXzXINDRuCWOADiBYd/5aw6fJ/PtHP6hvfQmgPM
pe5Rbb9vXhfZlTdZe6IYAV6ajOneMnpE0SRKlyLpgkbpQbwWF8Ta9x699vjybNfWF62AYBS3D7DQ
b0t7dD7uNK3C2oBkpBFbB3y/rTrUlQxN4AZtlp8BUDmTdKIOwvLfH64R9omltAgRoa9eT5fKR+NB
hJulrR0XnMdnz4MTDv9F/TNStcRrNIf5MM0b3o9Lm2heOPvkpoBOr22fj5c2jTQHuYFT3gyiU8GP
rFykj34Hi9/EcnhfJs9E3mtp1Tszf4e89AyXHw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Rp2qWT1ngiwszVInFfAgNDsqirvFBRH0fhGMVLdTcJjuZF6cagj0r5deSp/lHSGQXbQ6hn2NE/pT
sVS4xwCY2B03TkdpZqI4G+dZXB8686b5iwRUQ7S4WwcHb3WXRb4Df1OHJ6dgH8h0dIOxvwXXNlqh
PKzd3cQ77q4ZzFc8bvI=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JmHrUUSZT8PLNYfmwBtqUH6qJ1p97BdaA2q40RVMw79ZG2/5JMAd6P3xNNzdIISzZU+jzu0NYPxL
Z/zfPbolJrCwAck6UGljZ/OOpPHLUDGkBAu8BIP536kFNfmsl2/w8PHTByudSnwDI/YKiNqfsxGP
M6Sq3+TkXml3dJEoLhHWDNi1mL1f4wADZ5vEh09j4ryxXNWZ0T1vCwLDq6JQfC0fF5S+fWguWeoy
y4GDwuB3WNo6v4nkxnIBm5jk34GhklMVorbQQ90znGRfAejdTRlBiH1jH/CASbqnXiNzj4+1wJ6K
83Kv1+Hi6TU2vQtu3O5wYTXjTMpJrASuG6iNvA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
e9asiFlPlMhHebvyhrXodkSb+NOW1z3GfRmx+mGmNkvzC26DFe0MNgsYsbYULzPnFNt2Jph5a/qQ
la4+MGYuu6kPTujJHRAMXjPbrQy3NuEI+bFALotLuYulCGeYXOHECHkCQDzwE7cOgWofB6M9nMDI
MrLhlrFd4RIgHL47h6tXTX625M4FWH/nJM1zOgV4FtdkDNqrfdMVvfKsGlHhYjjtp1SRu8Hspgqu
l3IIfXh7PB8k7mC0mT+l7qcJgo2DarCHHeprDgNdO1zGCmntW6VIiHesLxPgNuzqP+AZ4J47uWLl
7QcIfX4fFpKHciTrZd/pRl5sAuSX4o+7XQp5wRlXj2huCXK1zmK2I0r75nQc8rZh5sOggF0lD7rk
1tqYUAbYuMwkJxroFYiYKGXPZcObY3yMRJTQgZGWKFDJVA6/yDnvjJTnNRHjdbVVJ/VuleBivEgf
vf9X2/VBBdXbJ/f3PMrMNxSh2HXOYj/gRRaVOYJ4/WOolrt5gy1/myf+UNSQupA5BQXOqw0xr72b
rJ9fHAAG4CyKkFS/yoM0wlLVvlcNJFf3Zkc5cClW50NoXjnTSeOyyGjqV6l/UylClVQ6YSKxv4Cb
2ElyCpM95qxOI6oOtQU5ASOMp3QNsOD4kElgSRew6/oD95KLnhgzI4Lme/RqnsgVjRKTzYC/pmp1
bFBmpSnb7OqWPZe2Vr2quCiLG4CdvxTAUv6ZktbMi1E1VkePKX35RMXAvj/xTOWPfbLz1TzJ0pDK
RQzrohpLOt8JeIXgw9Al1BONObYrLkdLo3zD8Ocop/hGa5+l41O2bib2mUjU8PZmeJIEtD7mQaNc
GjKql7W1Tww1ZOKKKtvqP2K9Qs8iRGnnCXfdWkwGxzKky2SKA/TQ/Ctb6gfg/VLRhfBt4sjGukXu
2+PgXrnzs9mw0/12Xu7+h7eFAybv1YVXZ4pAp+zNAMBE3+MTbVReii7yCtQjVitt3D+I0REmIFK2
jE2MgGAr8KPpCJeR0t7tMy+BzOMdpdt6cvPrTwRdp+amiqwdfM4azn9trtyMbbXK+eR2mnP8ulLi
Qj4ztPX3dUPVzCTahW4Aig2nVxImQXBfreoQHatEkPRxhgf+frdEQaBJ35Oc/wvfOfq823ipS6nX
cbCeSkWwl9cm6yr0Kx1eoGPpIFs8qcOI8FPYFTfhjEKfLWcXrG+39tK5zXKKbj6k6YXketMMU7JP
D7kUFHfnAOBZpvnpcdVWu6S2rKmq0QJfxFBOx4mXphb3es4pOse02X2knQxx17/eafnyh+3seFaw
4/IDeWKf0yLGxtfSOijOesKYXwSrUgTnZhpzMKGuDww08HTt8ENr/f5lPYw/jSdIeKDgx2eILHR4
iEJUkZdAKaDKCMLM2gSYhhk+q3/JFXZMi3gm2rLQ8XJZSluMjUAB2EN8XeDmUGp4aaM9WaQ/3KRH
Iq1VtCI98MCsezoPumRGynJEznqBMaUgc8uEW+N5v3MrP+S6SdM8kZ3kDahxRIKThC9Jvzlulgn5
t2rTPEp/Pb5UrCpV+3Q3GcEHcEkoJE1KFwNOez6UrW+lzv1pLt5BESz/SsF+cDdpFhYwI+JON76x
MlLBvU13TR7Vp+EOud8s9TS9nye6/fYSXOuejZJd54bee3dZFVkf4txv9PUfFrmI07Sk4Cy7ebhg
pBUQOB+KheYCo5SC2EwhBxd6GfTdfYPesg2E9Gn+tBMi2A2togC8bENMuNpjumkyR3gvyWj73Trw
HaxQAYx5MDzMWBVAB1rKcxRcQYF+qpU1/VwF+tE2ujU956bQl5EY9djjjUJQpWr38DduRuUSzKdf
D5cSbX/aXKROURYZSGiOzE1a+nPAfwg5HZlPJMLnGxjmeDFw0K1npNmHxmIrsSDLjSX6+8I2tRpT
eF1t8XJd0UT2apHSTfdckfKQHSCn5v22ZeHDEhGKPe8TrFWJFvn/XWeUU7Bia4rWt2negHN0HQ5T
z5CldeIaEAke3Fztb6m8HhegeVhd8/VjXkYvertNN/aJ6ocPq0yOZZDZCy2pmV9nTpSjnLsXydHl
XRtTnLqhCtk+o/TL+ndZ1FTIPa/WgWOI13Fii134DTm9VQ4k0lCIrbb8W7dLnoIquJphLDxd4Hpg
ZG3GHlWDA1zQB6bQWb8nUQ1KQ27y4GEYcdMxJbzXOF5TH3Hrw1yn+67OKmyo4/yrk5FHJERkYjM6
4332ykbPdim0NR4l4hxn4MlR8RZ3ICRsHJgSFfAIfrVQRRjGSkAUZcumxBMNPMhRl7gkfw7PqqM2
C2EeKBG4uPjDdrU6qtPwYK9ehRV8DmrJzZqZz8Y86zoVJC5fhPI/+cjv6Jcc0cvqxN5nQMwZvC/h
bzfr3ytb+5cVMga8YJ53S3YkvZzpzPKhVdtezisq9ociWuFeKPuNVBQp9eXCbna0Q3f+UYxHrplf
YJcrCU8RqHo2IEglv5xiQn6jlBUmUiqL+mbZNrZz5jQsicJH8JbCzGAqdFNARm8FQh1hfAZGeo/y
iL7t3/PuFDFvolI9OtTf52wtZjBgnPcvxOYhLrwbiceXHQocj/8JwuGPZSyocE1I6PhUX4btQ13G
Vz2skdiKcQOvm/W9kV+9bnuHO3Rl1/fiTg04fWO1aVPQOUrIOIFg3UMlJJAkvY3PsFWgTlW3ha19
8n6TDdvgV4VOAKJT3VcQuqYhLQpJWieusE4HB5EsiKMjgnorl19gI3v/WkiqCeMxV64eHtyCrwKR
If+sLPn0K9b3ESiZbWXk7UnumnErXagQ6uLOTc4ffyZu8ONcO0V4JTnmTLWAd2QaYl+zD01+HfMU
hvawqn1CGdS+saFdnoW+3zXWQQ2bB57kuCnYXMG+PnJkgyNkECNTMxnExtyXMlu7nUarmaN16/Yk
IIYY8zhOJ3puQRZaodq+7gf6XRBpvaIUUwzEZvTln77gqGKuI07vfxKseO63ST7X5AD1ph3MZ1e1
uo7/YBA4EGcz/+eUDyraI2TzNtkv7iN8zqtMY9QvxTAmig1L9gsT6lepmXCy73Ta+0F9h4SH7B+i
BfTsn7n/jvhugJ2ayWTCgG8byJLSAJR1Mzy94NQejwc35e9ScNT0hns/T9sAGs11WXtql0jLMmZO
g/JzfxwaG0zpdbaxEbNGulmrpuzMppO6lfJLFkeqAOamgt+8t02jp6agE+3AaFZAobTQy26up2lH
TbnHA3wQsrd7ZxtwvxtNkeYsaS7t90f/gqQj0Sv6aH87137JoBXe9ibZHzXt2BcHKycr+fm6igpC
BmhNbbzYWpZBJ7lqlm9Nb/scHbkN4qrou7c2urd2uogqd/LV4WPMJOoVgl/CnL3eqZNG1EQlkO/9
T6rlBvVvWg9iG4X0S0V1+0F08fqqHpnf8umnKsMxqXskWN7ojvNWr8WoiP9uST/KL30woEzEQFop
4Kh+ZEjcJ+L4UWvLhir/Y4JrxyceLTpoIucvPqNyVZ3yTjyWC/shxAqVhfmafbFrIlIOT0p2xxvw
6zs+PvHm20DpQhAXPm7qmyeRQwbRXpIxDOVoP4W4h0Vx5HnwU7TTygj9z1qhSkmbkanC14I35K3t
wlCEgMwaStXlqnhyfuIk8NFYwf/awdmR7ycHXvzXF6mK/qEnhLjzHdKLkrNF5BuGWf7f1omMMaML
qNLiAuf5sXX+KX5k+FLlsCjIAOGesqs8j6AAEw9ItMi7EUIUWPyxEdDZ/rT4JK/A0CA95UmixxLT
r7xckw8/KHPLytbA4603IM4hWd1CydI4Y/ANgL6yp63oXllPRdkxfCW64dk4hFQczse3Q3CviM32
fHNdM1dddyqkrK9RjYuNdcHF/MRjmqZTo3PZ7slMWn7E3svr55prcpX24SBuezHawOWbxfQ11ciS
fjiLx5eqrRaQRbseFFSkCkRqSAgxOKrC58Dzzon4nLaESypXliSuW8NtkfJBNVLcgUulZBGYHZUp
XSzqOjgW0at91DDRwbc6JvYqQTRXgCIJjo1hhsbPxmcZj9R7FtzgQS2relZ2EyUCvFlSOtAYdM9a
BqJ9XIg+x+nQmS+lYjmY7CbL5cVsZQFjc+zjoefIgKD8I4wz7ojEhYGY1kUgc51VO97slsPZgf17
DmEeZ4DG0yalw00+x1oHIrdPPTYuO3ADWocrPKTsfGR4aNzzXZ2Q79sDkjogisHaXknTeYol9VO6
EY52YmzxUduLPLYKjj1lByh4NxhfskGdpVuANoVURnbVFW8uoLBj++j5zE2B68emztGxgSldG5V8
sV428D2bfev1I8JA8tACnf+GlLXKfKndWyV1K0ADjOHVMa5EBcXAg+f0LR8rgawRtUQpN4MghQNG
KQNzJm8P2uKjKB7O6Q5/2Ec4XOwfHxgGZ+0Ya6qhr00cqkoZZpAXcoQm5evOpZY/Y7SYeMPhZFbC
ynsmPrU2QbxVxO4NaB3dCDAsnozsy3moJKNhNLfnP5+NiYSoXelyPGsS5wdmv7RbLMie8U3z6GWq
fycJMIag4hzy7YW8LprBxbd15/tyDJ0M1fQYIgHqGlcNdDm96bro/63SK7Zy+GTd8ePAXZJsJv47
uuuovE1pBofv1cgWdyvWI90Dsl4Nf5RldLWwuau0UW43qU+qnZoz/+mf/Jwh3EsQXcP/+xmP03LU
/2FDbLtmDjaVU6gKqLX1GvgA9sF11N++x0t7FQe656/g7xBUKH9W7bx8LTTE2yajapkC+EsGTNWj
viqDwzOUaRxwgDdEefwSSIoYBOSgvSBQrHWecTu/G2u2DkpDdjwWafl4fJTrEbflZUpitRrkW/QZ
6aI1QLGWMtVAmgnSC8qAt+ihd8TVBCjCpuAbtDubcWoCedptOXMc8rWSBjc1fhALqsj1f93c7DQn
/60G9rqhiwfFKGNUvEELkdVFYQfJD54HunSZDRAYHQsSHeBYLkF0xGdSV4Qtd7ljuINX/JJCElWV
Ytz5/IExZBqY8712cFu8ob1RPCoD0GDjscitiZVWVCHfeNxkXNkuBrjInFOrdUmHvD/w+1zIFwRX
hPHyYUqKE/D4Zh1FS+J6HFQUStyPK1qc9OrjpO9z49lAUJT5dHiyE5B0J86DJsUIGPncM8QsZpB0
Lx+UOSEDZquNzPcT4R1P3O4TcLtPeTsmrQvazSaauOeTPj9x2LwSf2vYBpVw4HuihF3ozE9OEkbx
8fe7qqqefxI4p6FNpF5vjAjA12hR/LujEq6De9RP176pVyGyvK/pepf+NyBufluEpBHNufVo/lru
Lbvfbxxfrx+mFV+t5uBBJ964PCHZHsh3UwSGRS1iRLvuBF/ULSUNPF7uygIOXxIGgnWkVOQGrHwJ
qw2frFL77JcUy7TLhxynb/z4ow1AtRKQw7VxrS3JTck0dxT0MSYIc/XYg+P5ZzSOcbsemy2GhBQs
FlE2P+KC5sPmtzD+yJVhmlcvviVLiUv+xMFyLV4mUU6FAHL3aVy914oUR/ccPwY9XcdJslmqfZbk
b09O2xQ3qIzPn9e88oCzjv930LPY9GiXxoKyRvHVN4PLcR88Bcw21iN96hfZ5HHtYTih9Pvab50H
G1MoYdWXv6L4Bi0v2j3ndt7MtbzGJrMHmBMlsJ3/iuCSjtRevtBxoh4BB8/CBjkb/iv1oLAS4XUl
lfxiEbXqkJIWOkX3Ooo0H6wHtDA+l0gfGP4kHUyab9y02w2iaiEO5PUpz/VdD1J0BHnBvpvXtG3D
hm3IPDj9ROZ/loOwqLwG22Bo7NngcD9efqo5uKnhTwC7vot5I6Jv0xJdUhQUWELvjVa7BFKfxApl
qXsiStiXjVVs2Dv73NQwCKe7GYSn0wDINzhgNOMqmn+tSdp6uuPblfucc5C9KFoTo+3HJmklICnL
5HGJF6UASJW/BQiluMgJA+mY1vbTA9VGZmSCmD6J1xN5D6DkHfpOC7HBdwKjDHoIOuyHgdjqiIdX
fuyyjfFBIvbXxRVL+TUfPGSz1Tdzpuiw2sjp7z64o3NkD2MRvs8SwGPBr7CGmb7Z5zzv+hmVQ63H
zc+KsW4VElOxiWkUA149eXAlLYQibsGa0S6I2SjZUF1WlbgrSgMnYcEh1OPX3mwHpwT4Nt4eXgKJ
6Yb3oEMJ5ZsdcwBQ34GumqFm3LAQEP+fFngyD8m729/RtLdFifm6dA1NpcC3VZyk8ntrBGmiVjwt
qnaQsEEZdqZUSDLQiHrFxMUDQnCfW5DTBz5rT+vGBkh+Vr4gaIoL8LkJzUB5thiu7zbghaaKY1ck
1tQ6Gsq/kNMInVJqSxR0XG4mpDzzGx6kZNg9boHfO32VgH5Hs9i3sDLulSLn3tU8eBGhXcD+ti3y
xFjFqS6p/1XgKe1tcKs+/va8XZwGVlQXm67am8DT6Wcszx6zZjY2meX+4Gt+ABsM4pfmZAQ/5vRY
IsKQ3ZCkCEyug9GVUscH2P6GgQ47z+xUVctc8HrQXAdEA4mOhW9iJckgfLs+TTpFm8ooa+0NLjOt
f0WweDl2XwtlWOQHEfGXTi3bX8iiYQnbeOAe3QGUMODk463Pvp0RcwUL9IN3c17tN5WhUstPS8Ur
Qprdo2+Klr3nXxNBy8i3uJ+2uEsOZzS9U+02zrHlnvrYSGHWvtRcCfhTOhC9DL4lo+1yfxrJjikk
1Guhhvt+otvzPgOi2NM1oA4PuY4dQ88PyFXg3/nGD3TqKzQfFMXvW3mcGj1Ja5Fio8ROVi7C8jzg
ukbSci36SPyiaG7gb+5LB6KUSgmKv3xhS9BLSBOwdXX1OUsMVkccmBJAF/CKbAjwlvZwEN26hTh6
6qvn73+yrNf4c0mzc64mmInuyjAgT+bKK23/cuKlwhbR+9bbaAq3/d1xILzxNzXnZvA+Kh4Cyu9A
gREJYZdiPMxPJMEYBok5YQjwDNao4zl6eTxKdNnvdk8Xf16GE+ji0wYRLxNQe6hMui6NClPsWzMc
QtIJ3hFmAystX+CgKEIdmuApkwri0AazL8+BZjdIqY/IRzx+EW+RjjHJUODcVT0NkultD+uGENr5
5wE7IZvZWd/zy1eXipU14rTvr+5Nl3z2NRXpXKjZ47Xb9xCW221PISR9UaYpnTxwllk4SfpCEjQZ
dEtrFdHATCcvQOxjiXgIlCpGhqMF0VhnqVlRAx8QlG65WlpG96qqIdszs1thsprBFV25ZFi/cztZ
ABXPDTukBTL62iJ3cIZiJXIYhRyuMPJSh4IN3drwzolMVvORbvVczWTv/BX49lRNICZtXPA2PKQp
6YSP8TlzDSl8zXkGzHEWk5UqW+IjuaZEikeK97xMc2y359uvt0Q0S9Xh2nKPX7cVC3JXEMp3/3N1
23My3+7UPHYgpKfK8fv9onfrdH0J0me/xUj0yQ6EvCqGOKq9AmceatS8P7/THLND1BkDcBztA85x
BroAc5u1LpzbhRCDj6PYXHOUE1QxeN0kjBSk0FcKdm3FDXxzcS4OKISAEnjwbEuTLPmYki+Ks8tG
3kyKfMHvU2stTcLvSuJGVFPwIW5rmUl8WVRJNC01wdI7XnaknOQJy1NLPLkZmBzXq+HmES5cb9F3
ywDzsabi5h5uHmGhhLMSmS9ryigVsDb7YIw95x/gAfjDV+Dg6w0Cd7GcaWPFO4vRW8+zu9jd4Lse
c8DCBvmg70qTLnsVshFRt6CVuqfgpmY8ZTLtCkZAm2S7Ea1alRAkvt8HpTMax75rlcpQRA8+y4RA
zdR8ZgChbLwPMZ1Gz4ykOY9lrjd/pa0OtII5oPt8OhsEbb4vBD4BxdcJi12YRjLO2dMfG+EBZBgx
Pk6yHW9+aQV7g9CzM8sunlkG7VTc1CcPgLNN7uOmdabpLIGFkU5sblNuRb9tRMXiSoYReSPgQe2X
zHjv9pnEDGY9wvY/t/4AZ17Sb/PdAS2+4z6RpuHP/ifnfPoBP1xgDfj5D7uruRLAjP5OcvU/+fj8
qwAEYn8VK80GGLWlFdSj5py4kfdVEkPDt6QbeapoYnVIKr1ttLjx3ZPe5bPRBOG+EBMgENeT3yFv
pT+dw0542TGJN91Jc6V3Cs2Tjt/li/5N+Bs2wWgOu6H98bJQqmpEQC8kMkalSiJrmll5JSB4q/CH
kM9cesabnGHVrXBrvuYKZSEFyOOM+H51ykcNyJbQlMtzgjSmcgQnKxKGZCO2nl+CceObH8502d/W
07jnYMTGisXri0a6dLyGw3+wKLLrJ6wqWtVYmPjxiAZATWqA3RwTknTlcvgGH4OowlVBwLjAL0G/
TYpV/DKangydzS/KApSfVQQ2ViOD5CqKqJWLigtsO7239uEkck84yGcRkJX4r8Q5g4lj91VadjfI
VzVh25kVM0TG/1Qx/yRF66tLCcAoUyWLbzciz02MhVaqc5aXobYn2SBw8FGlSzu3MGb7W3QRkTJ9
T695Otsb+fSDzfeVqwGh1sRYa2miwo2P7X+5EfdD37Sq2ZZRjySPoMwqzt/81ZiyPJ3ZCRhb9P7i
DYj9409NKZDvR836aYcUXpAbFNwLeLC168gPFjoKGkGsE8zhEqfRbulIxb3xy0gGR9/o8sgHCt0l
cZ6Kv60pZuelonVUGU4FPnyId6fYnfYewG/JhBwOA4c0KXkvvSrGaWIP06iNPHwE+jUVThROMs+7
lTYykmm+OuUNLKcd0o+FTybFby7j4zwbDEcYdJDkTtsEJsIWkoucWzgVxq6woBwnoLf5q9DZMbbS
0T8Qnx2MZx9I4zxmvSdm+5TrKlWMpew6ibwZ13TBikN1S5ARIb7cR/XVhJL/jyUI2s+nqb0GKhtP
oW/nLfmWcJddGyhFlp299YkPOwPV84IiP8hSZ3G7RC+v6dBByh+V4mHUNBUjFF+37SLYnwloYuV+
Q7k/MIkoWbpjBPlKZx0XmLqvatqqbyDYwuvQ+NewkhjUMKZm5hu8QNdfht9NoA7EZ5cOnyj46FLT
1k+YqMdLcIuEopGVM349CQW3D+LTgQcCnNG5Au6jJsfbcQTW2P/jf94kL81sNeF8n/pfiPzr2Rtn
iXoVjkSQqjRAeF8fYP8cIRvVdd1uhOcbdXaTn+DYpArvm3GXWQ2hpP9NIPODhAIg+r4Mo5K+7lio
mN8LrTYTBSvGE5qRUyfL5MkE0mlawKLGFwDa3RhqI+tlyA9i2u3vqM+iqQf11kJDZFOphDqY/Q6G
/TjvitQu1yXFe6uxaJXcVhrNXAre4rPd3XQVF0sGj3JUhZmvbcZYSf8t2VK97R123ype7GuvVWaa
ryJTjdSxQsV54GMgBgy/Atow5d+qKzNDCTkVdwBkPrss1ZQqndXFWK2myBbsIlPxmJk87UThFrqM
zOC+tb8seoqO/RC21t49ayr6Tb41Hj7xbpi/4t8/GfBOj25Nf1f3jJq2jMgU26QV6vcg/17gn5xP
jL2kLiKzD7mtKVcG1btKM3dRMXMVzlreA1t5l2n57De6HHKZMGBCrkR+N4rDjUAmw/WT7cVLpS1M
CN7mDJGDq+/P55ZK+kDMKkITn1Laos+9AowH5U1zR7mTbxwrQsuq3riPncV8625je2hil9gYxUcZ
QQ1Xu4fjPqv/gS0zKRhLyiU8UUcm+5Oxw8DSDnXHBqJpAtJyjuLpmLOpcZYbJJdVYNsUjgBHMbJY
wFOjPJ9J3o3NM6oVi8hLSrxjUadSmr8PQ9tbt4cX41LuwtwQAIa2ZT38LIe1dsPMAlGHDqc6mn01
Vd8OBEov/b0g1/d3FAwNaJMINPzbgwm9ABQDM0355i6TPrvCho7GzRquiOncp5gqH0zgRqQpRTTN
36S/i1FfcXpx/kvMenPO+eoVG68/VERoH5cOyO79t4vHV0fDbwVKHmWo9WoVyRLaVwVVZ5rdb/y2
L9FkaUqeOJUe+WgjYfSNrJSxi3DWGGn7+WcQv5ldd03kQTfgYpdIdZx870jN+nzl6S5SWFuSnfPL
CvNfWzR+p2j30xMdrn2NXjMZRm1HX8fkxPq4P1TXgP/dzrHBgHi4gybQGENmLxko+k6OE4xp7Wt1
4ZbESU5LQLamPa/Dg2e+ddmJ4w8wyZ61yxQzUAH5W+1wUCBgSBdoRN0gES32wcrcDmvmLP620KjN
c9ZPksOMEP4xL/f+t+P/U2ER0YcNjQcwukvHb3B0NmOGnQcngAs3ZQ0LvAfrrhFHMIbsoFX/VIYd
7z/p+x8MvDTtC2BBiiYvsrKku49BX1gBWlEPqfOaTtlU5SV8d7d3hLgmVO1azOADYK5e44dUJK+l
iDQlI/qIPGNHY9lozzpXMXPPFknqb5cUbtU2XGxlpwIO8IpHQuPEp4BwBdxVePUXs7G9abPsDKoj
1dqdHwOdc30bTAkOQhmValC19pfeCI9ocTtWq22c7GbcK/h5Liof47HralP4SuVlLLPBX7816DQM
i1/EImD0tz9YpHWmJBj02iHwzel1RefQlV58DfImI4UKuTY3SG1u9m9/xXk27M67XZwN6pK/HXq2
iEnpb8eNGMxRNgxGWOe1zECmuyrVevQg48oDtYmBnU6kZUCjEKsxfkZKE+hNNM2LqGWegRb0Nsgo
tQTVF07a6gBKyQj84HQ0fjf8lPVfIK8wYFH735paW6MIlCbM3mMQaLCvz8Hj9wzinJO+m7wfOAbH
bHYncpC32zaFMHHkOLpMlIaGsoHC+TKQbvbEKP4ZF6GxF9IA0xM7HJfqhLJbcEGPTND+rIMgjOwY
9LnRwJShUJhRkss2HTRIH1j8pzRp1wF0Kg+M0iElolmeLwfQvqEcGWHGnPWwLKrgqFAI9AxWQ9nH
4VlSOmlQ+UGVSQENKe5YPMYP+uZw1CeLDTjC2wXoMMCgv3jjPWCOrRrY4+CV+FPUywJYsKZEufZD
xxJ5IL1/Hj51QJke7kHjeoYP9hZAr2kf0LAyoUKMO1LhnRpV9mvWLlO6Tb1UZBMbOeWd2VGm/zIq
ciGBdO9t50DY/lyRwS9S2HYC4S8yX15fVFGidpcM8+SgUjY5ccyIdNbINW6ZjZJxP6tfX00Nuv7G
l6jL79aGg2zeLzS+sV5f3cd8thbcaSqSHvp84/5+wYqPc4Ho88CETXaiuqcrzpQgtzkteAHApmNH
9BPRP5sLb7Z3e8nNwL7qwlUT1DKPDLb+55lZzgZKC0o8XY9QAPfehGIFF8N+v7lfUiAbxpGB2flh
pXT6XDOPIBfy7EzbkknXo7+LJGRxld2A3O8AY5oNh36HsIGzTz0e0iIjUey65JB1MNsyaSu8co4D
01UDK98j/MxC1vGRFKaOkEO/WCH+awACQNIVt0g46s26kTHGDBRnYz2PFP9sbIAaPGGtfyHuh/jr
WxOvUWXP4rB/6rxZsGvTlyaHtuotRvF2e1RZO0FwXB4BSfUGgyWkmbDBJ+AIQrYlY9Uvusury3TN
WCeIp4xR101PZoqt1UR66RVikMqeIxxPhrp5KX3LgwKOFN2loxdwJ6HCUaBl2GwQW3NKTw7EU/vj
gn/xymGldbipaNNG0tF6tfTYh0YR2UFjpBWa6QrHRfeklXihxHfoKGXcUSl3uj3/YY6Pb1olI1xt
5S3ae+RBHzMXsQxHtsBpwJDR5RrEsLSrsRUGuCf2PFmDF/3H1G9D7ThCeth5ENjkAOtTe6IEo5EM
QyAJiVjyjvjAbIfgmXp6eCjFv/8MtFJk/Uei9fZGklFYT9p5rzP6gON+emptEkuZQl5uDw3Rn5MP
1yUGNz1h8BK/C/KLXX2x6Bs8LVt9QTcm3d117UiKNF118kTiVDgfDZVl0NXYmAItiIJoRFWE3f7r
id7BIstH4iazypeQ0HkfdmHf1ExJAJbjk0jOhxNosKm+TfIJjO0bmyl11PYv8OJKC5ciMIJabTF9
OOrUIrxIVHVSXMo17zbHuVeaHLUl5J3jtpDozu8tha/mCkHpzgTALTR4xhL5attdodlx9iuAKpA5
qB7n0RVfyceI8efGckbui+0ELdsHQ3K3pyv/+cU0vMjHntoaC2y1esZRZ/MWIBClPfoBXaQMiJK1
wylx2F98mjoqDQ3krmhhcVQ5vXd87FTMznmmTr9MmoGixt5J/OLoiB3VAIfNF7u01edHrj81j5Dr
oWwL6eQ0cSbeFaQBO3hJdhK2iDjOZt4bG1l9M7+eRyIBSfszFKcF1lY8KCCEJK2gIhA3UL18BOvE
jqBVviUFhkB6G8TrGQst+QAcWORHI5HEm4ptGVdfIdtcNia7LFR7LvjyMAoosgpBq06GzopDHzTM
Ch0anB0W/5uOhiNZ8vSeo68Y4VPlosJndDQTayis9mNqp/Gb0ba2hY1rZXwqKnlk+dNRKSsIE75E
xTiJ7ilH3S8rsquqvyEzkAq8sCTDHmtc36/s1y1yeNSgGN8YZyu8q3T3QvO10/+gVkdtK36zmiKx
Etc3zxmLikoGgUuhrtMRAmNaGqa3FSVLMFbK+cANgJhRZfrykyq8DEuBYseqHfR1IBRoTPgQF2jc
/hjfPUrPpqeSAOrcFHLNgNGRs2BXEwamakmjMhevxgrgMHsBxRjrT62XJCHFSvUd6FdLeNMn96dq
3GpiYn8te62UVkViqYIsw/urYr5KX1vbHMgPDyXUnrN6Ek24mQro2ZiJuXWGbxCDzK4hBdtPAnbd
Bq8PT39jc5qyqHHWWR7gSIGa7fiq2X7PgIoOgOQ0OjMI37RmdAXGOP9g1iIsPpXfs2XXCG4DAUil
/OhHnM4TiUy/hfruyQRiGz6bL9R95WbPnhh1Gabes056ZTSc9mNh5DhfC7SGKt6Hb4xsp9Cisz5n
Xccg0LaDv6Zv6eVae5UsO2dvgVH/REJNJe7Tnmmkz+rjMzm8pubFvNwaRFbSz0HBM58MWR8ZwWxa
FUdKSmauJxen3jdrSbS216TR8+kykuciOOJtPDwcKulq1tSLJFuzkeQDreZgCSB1ovhGrUWO9mop
Q7d69Zs4wd01zgJheyMxspIPUV5dWvNiwYzXITY3zIu9pocWpcPMsHc/OMepAoWaHknELMAs57T5
/ZDxu09G86J2fQk29gjfo0LmuIdO3BG9V6dHtwutb6dnuQiw0SuxflBtB4S/sg/IH8MoTGlSt6c9
ulvBohWcyVrOYAUaFRaEfslHCYnTxu/NyEqeJ/v+xngd5PHnq+KHUMCcH/m5naSntTVLE1put5z1
3W6fHzImlI6Ok9BimRHxZYnpfz9qgltgYnCLYMoUWNmZ8JAXr6iv3EN441g0TYodlg6QvyWpfzl9
mkLQem2L5J2tpXQ/9C6CnEzU/nvgUXI4YTlbm7rmhKu/h1SuOmgOwSOngQKFIIufwLhd2jRHiua2
zLlkh18SHHTjBTkTQocn1EjlJ7quKQ3pykqow81OWwc4F1NxTn0FFKoK9r2rm+kCckAthyOIqWfB
j4hqUtRUt7TDMZp9s1r/OrReINHfmyAekrB7Civc3UOSnbDHMFkymjMcJ36IvAoCfZq3uKjQCF+T
Yuoe/eTSRQbY1E30cNgqbPspfBVrhvWemoy+ywZ6NYrKWwDUfsZdCoMsNy5oq9J5iNTxMl2IITSf
ApsLlLBSxkbCc6gpqwe30GWNI96wfxiC1vjxBW469P/XNZVZE7JqnpizWxvOP7ZdKQ3l8dRFNo/H
6bmJ9iEujWTCU41bQSQS1fE/n8BZf8ZLGmevZ5tPl5GXdVfcJxG/MPs1/1t+GU/oiphyX1hW/F1C
gOJKqB/9cHHw0tz7KrehwdAwBSInHSD/7uhyCqYbZj/66NdBpQ+hBSHRnK82qaLIOWrq0EROmraj
rQ2V+sDUimYRk0dEEebgv5A1M0eaFWJLzYgHHXPsyLAYGgZMuAejd3NXzgWgaoGvn4s+tfOtepjr
5hm2qnK83hW4dYP8nqfn4BaOpNlG+D0mJdOT/TQc2Z47q10n2Sp3A3HiqLBGSF8LF0OS85i+523E
quckaoLm8FGVHKz9dMrTEC/OzPHu5yW0nvxhP7bFf41mUTEHpddWU38jlg9icESMAnUuBqyd+DXK
DOQLsyvFKzwRf+Uvf+9YmKQBwfuOZB1BVWJjcA5KiuoY4ZFhYVsRbLTNePd+KuOlEdSeYYgdwLjI
4nr7h3zRuIRtrDa+VRRJH4Lhu4H+klwUzQ3Rh+kpVPPeRz07ClkFUCM9sEqizgg7Fai5vHVU2wlr
+4uHwg+L1yVoirX7xjGOS9nxH+/AHjegBl+fmknn3i6xqdF3cCZ8fzxE9f6L3x/eIdIveebSND4t
vdRjgsclORnKZcbnPwW1bcNj4RjvW0Yvj8sol8qZ1iR8ECDoFRU39Oj+SpNVixp/TcVwuwyYGtjF
v57JN2WT15oTiKXyU0Zf0n6ifqZUUyHVWI2uThrWhEIHHSN+/ig/7RCdIOrv9CaFmNSvcoloJmH5
SDRi1ngvR60fTR06DHtdPUdJIWTRYK7SkskF4tJNwZSk7vxcIazCgN+qOt1RJ25+rMOH+/bKeZVQ
DEdBAuudRoI1sYEotj5aMfhRB9Gh8S4pmSd8tg7hc5xv/+w6Tqk0UCFMOTEKFFUscrF5r7wq64NV
nkavpW6mIv8XErJZNviN1hblzN1WY0ccNJ7u3PPyLtsx6ctxDziLDOrlkyDABrWqScyiTZnosr8W
tYpQidVMZRqkvUOy/+gfldyuqFLwf9VuUDWQnSyK1SKyjTuMCdlKEOO2dS0oz5LsqhK2uEHzAj4l
Hrv8dKBKIoxAsmIx2MbaHiW4TFNXEgmzugw8j4tCnG/AiNnY9K7D+W7rpPHFFDqMfWeV7e3eM5Qx
tFVgK6rF4+RiRYXPDg6ibcD4KGx4XKNycayWkJmQGD5nZ6Yx9/KdIzN8dNjAq46pE9jkVQf1g0YX
8tSnR2LnLJA8DAi7+EKBDd/SNRttZYhMOjPrSCa/IsPfUXwfxWJfFB6fWBVKnCs+/vpdky7tWRZW
lDLTAvoUA8raHrEGh5XfHO0j6LOLQ5BY9W4+XjrIQB5RDCN7e8E1yJodsb9Cc+InOYviptBstpjQ
V5SrAZuHI0sKor4nz60ta2AQGoVSZ+nDhlNtUglL4iIgC4ikq/DAe5q/XE3hi/SGfGpwIF2GwrX0
lnDZqfO1F67Cg23T2C4nH9wf6ZW/bjglBrGst/61NI49njmeKKCPMyBXYdNXiGxf7qHIqeDmmHoy
5Pk7AOUXplcjMLLQeMUFNIKI/+XISuxPiEQdR6MBJXN6ng8/mpXye6NvWU/HYT4j1J1GfhBgRUqp
xvJ8Ow6F4gSvro0k8Ex+mm1s+fPUbRlhvD2fReDDE7pJHcf+lD7gEJpmCvRrxPU3iQsIA/RGrqZu
E2C0iwgoz29I2xoG43fvi5wJ7sP/cAZ8umHFIisP5SXvyqR8ojZ7GzI2hugy2cqDoAGaji4Fd6QB
gpEdlQwRKsbAwOChElAfA0q1H29NOSNtNXcbbGbiiROA8GJRGgkNzHLtgDcQI3y4hTfA6VHHhceM
iNXQ67296iveYHXTPTkgSPu8SsRNpnIYliPQ43MZyjMXY1v2EhdWZ5yAgtySyN23QAOnQ1fEL90Z
8kKSy4P8cBDRnUIU1DoRE2JrzxKvunEl9/H0tzmwAGsfCtyh10jIgnVgeyRKLmbG8Wc0jGgWk6vv
2CIeY4+LRVAXpv3FxPsb+fYaBkXbBU5mHwS+GSXfqdesoPB/ZfjUsQmTqm4DA2kOmOdhQhmCxYpB
Ns4Npl/5e8ajKcE5I8WWgUYliXjZeZgf9wZQkz0mgU5+pZqBxxiPqY0atD7Mj9L0IooZIncXlaUD
IsNPlb5RCBO0aPwfuXUrURcpZU6Fi5ykCBEu5w0lqv0nPc1eCIbnZIvUrJ+fgph774OmLDwSR6s2
V/2EtxHpQbfp8aaBIdXoI2x3826io8hfursXAA6lH4Zy6fy4KcEZttlocvQVofmUy+/pG0vzdlhI
n2krPSMrZ+R6QblUx7QlYlRTje+Cn4VHf/NZXOjONwCCHfO9NyyG0VHKwLdUTvZAiqefxQq8dOC2
c57HHh+3ak5M4Ytn5Gv1dcVYFb/x2gUVnasRneHTJu9WfH8SfGNUOi+iK0LZrS1CQvr4fXiy844I
I1il0J4AleeKRjLVCSPJsyGyxBKaJh10C8laMgj8xxFGT9JvGHzfwBbJaJHxBIHdei9lUli12wh5
S5q4HglzULPryx6c/nPlN7f5iq3k99qh2Hn4vidKv8faY1CMhVa11tgfZ7EJBa3rRjCNl06KUQ1/
ufa8BJdIfemyeWy39TC50qR/9kYSC2tyz4rKdhlPtQgO1W3rG1r1HysZzk2hajNHh2N8WVV5+9o0
b97s8vn4k8jl3s70YUR26UpilvPgn5gExrlufBxA87ZFyAPRxR3Qpku1B35u0dL4+DHe3+wOpKid
qLzup3l1993yT1iRn8HHW3X3rlgkXtoWuS8vbd1Kc7acm2WuvimdA89OTGuGpq/oWzCBR5g+wMzd
YhVKr/nspa+WwAFKiFSxuJg+12bVeLvKzoMM/M4o5PYEUCGX9UY1mc12xDPMyGtYhbixxucMuRtF
UR11HJDhLTzybw2BEeOCCjWOAWWni+imMf6MN57IyI8KxdxJ9RnHcH7WV1OIuuANckukOwqNO9ik
vgOk/xU4B2xiJOCyWkw3PyeuzWaaoWevbsrfUg9sSQl/6khyu9cqHF8R8/yka1A4VUvUGfA3f3vb
Nw67zHbwovfX8vFLdCPkONzCx0zSTiFICNptAzqIARmcqSl4C9ot3Jyix9hEgFU56ri2WS+t9Ytc
6SV9XX1p8ALI6nqlwgtboba8fSks+GgQfXQ7VACvMVI3/fCbcBGptKQB7aFJYhDimGt5dyeKGfsk
3EB0Kzu6Dg6H4OcxuJHpw6YyusQSK+Q2TwlNYIVHbPFQt0WOeu88qvtkRQYtDdp7EJrqCi9mi/j+
oX44KxuiwtY5WyRKBroBCpb/y1QzsqVP4L2A6GhsGxckpsLX4DO/cHnyIxyYlOfooXlaif2VhVgT
mlQF4UbdrLw17Hn82vGCd9wxzEDSA/mZoymGulf5FJ/TCsV8ioOQDHko6B2DMLoSbkawJZu9Cb/d
hMjAp6DNlE//mcEI+cKcfRGWO977vZMgF5e258cVZWYCi9vZm0/cfdpolzGkUyO9vXEimbyIPXU9
Xe6Z1vCg9biTFk3S2K1im5hxOeDWEjMh3pqKY0uxBR6PlqDthkmlxoEXVfaY3TRtUhYeGZBd700G
QfWOvpZus46qwh5T03a7zPXjaKVYF0nbBIjxRlfHqtrXNkDFAeFzWY1X2oZ3nJ/JN/GVtAO94Rdr
h3YrELam2VoLMICGzLN73KRtW7thY9dLsqh4R0oVBcxLi/rF1zhYi+9CkamV/jaHv13WwnjaaeB6
rl0T6D/BeALDZ7JyESIgwYc6nPyOky/FMPwlLZfvsLJ3uYOyXRsXCflTfc2F/Mko4uax1Nq02g3T
zoWUWAnOaDGjngygkakjF/BuJH5fmpffthKDSAdsb/42ZeQjmsA5b6VFQPb6ts1+/CqVE5ItGJjE
VkCzAwtsEgN7jiSVHTZXtUKPdFP7vBGxFx3UOdNcv+bMERfBlfIVnVr9cKYQh+INEQ33kbaLResG
GuG2CJsUz6G55IQLJIbpTfKC77AkF2vu8+JBEoFNEFpOr7X9xVdr51Qj28Vn26rCB4cH5afZCyDL
0aTaEaxmCn/YpD3wXwQ+5I+h/gmoy3cghN5G2UocnWRdI/WVVpcQu57VNQTh6J78wcu05t0zFHLy
s0CThWT7mg7P4lDFd+LbqTE0ddfh90mWE1dEJJP5XmCSuVQw3SSYJNO7pD39pX1F2fKhToSGNs40
xlLojbYegqCidM8sn3tVcog8QC93ifZTehiv4nK2hfn4UuVEd37mkyZ6IlrMngmACaPYGhhErPnF
tth7t2UtFzJ6qbR8vAi0fDjFasyOxhyk4gHWXuZdksAFHSnxMQ1Mj+h6wr+QU2eFowzF5e7o+lYV
2QztcQyY//FxQmvkrSfMTjKvuewg5XSPr1wWmtCNKUznq1Zr7vJhC5AyQAXkg9H377oGAx4/9V4l
Z+P4Qe5Dugla3414g9T9/xXHH+kn4fKpYhSDupTMnXPObJ8ck4/VSQj7BXElflTnHL5tN6uf4aHI
v+VN0FdIDh2PM6tOZnV+FdtUnK6bHAQOhFCWEWAoRjZkwvtnjifryZHuxgYfJ/TzwUxQ3GNMhblv
J3kKtujaSavI0Sn/2qQt5n79UioZJFVubEhR5WCn3/30zHlzVnJ3M/HOPIEwpq9ManvbiTUObTaW
Ox9Z4asXxXdMSPJ7cRaqEpXBuEtZ64a4+T7NrcwZt+geBvZf5bAA24J+m0/ys+5B3LpF6oU9gs7S
GXwvVAoxRZ3jKomaLBPVWS/+Nxr53vLA6xN+K3D3hB0X7UpFEeMIbr+Ixpd4jN7+/tuEIhxh0Dpw
zjqdrmc3SnhnarA4XGcVFlWds9sIj4PDtDc9FFsgO+BOyKm/Vjene9xND3kXvqLlSKjQPlKpOYD6
SOtSPqF0/k5sd7el52PE1sybFa7X0KTPotLzAPpmzepF9ksHIs+DZLeDEpRgRR2tfMuB2YZp81od
Oq5Nz3NYVbFYg7//YrDtHjhvI/Tg5hUTkVzX2oXzv1kJj9GDUcXzrazjL+LYbmVHdhv662RYCKZW
2MF+PsRMNxXW0t/83e+899eigWXGWhS94CWYqMxWfPEt6DnSwptYJECPmYvk7/3xGEYx8i8LSyS2
+NtN4R9+nlyAElmrQyzSgJhlqiHN4awz+zqCs3rhNAh4x1kNU079mDg52aNMgcL7uZ2wdcqFwmt/
eVcxgA1EzYcvVC7RS/5nBcJz1eR06rRFA4uKidTeeV929z3ZgXBIUl53WTzxIdkdIXzFXmZ8nMS4
W4kMxl1Ugtd0g4B+P4exxpiODtnvVvv2bczab5Bju3zqZTtfC8DJWt0BEo8Ep2sjzKhTH452P1Y+
DJEfiKchOB/Bnch/FqwZ+VbQ1b3uzttWlHk+OISjgJ40vqdj2Zol+PX+FMn7gnrLJJpK0fUeRm4c
5fR1PHkMV6tyBytOEp8aHdsoZr+WH2i5wNEziVd3bnj4MTKMd0W1fl6q7d/8rTns/7gxCCT/F2x6
83Lrl3SxuJwpzCElf4zwYpAeRZMmZTq/SH70UB0JrAYqzdsxN9d092JRqhKyzrVLdouRBWWpJu38
OEkIM6njRk9fmvioK0VWlCirN6DFiuOK7aftaLra/dGBSBrwhjFjLWH88c+16ZjBMy4bulP3AKab
cl3THCiRBYFgiRSbVQSakWouirqCW4WApxKAeTvjdQ9sdZIzp/5BFmOwpCAQHnWUlEXz90AzYCVW
KKUGQPeiOuCIHB5mU3Fis9uKGIKAHulzrfv4SoFbctDkqiXlKppQcc1xZWnEjlwVEszxQqugpNKc
QaMhGOOs6cnE4Xw14rUmnbk6J4RQXmU5rAfMeDuXnfOlYhizkwhrOxtOcNi+f21NK5lLTxOdh6wB
eUT+EzXAsNb+YiZmGXAgSQI6hr190PMjpDWCV7eETNl0mujfYdKZY+mxtOioVmzzUs/WVvGzp3Ng
HNdN9ukS+8t7Wpny+XciBh9PinWZ5wz9Jq4h5hsp5bHEq9Ou5rc7NmLXAvZf934cEuTgKkXpE2xh
HWFcLzqoglLdBnCY1yZJ59dJfgDg2Zm7mfr/SZ0HNka4ZG+HgEfxlAtxuEEQdA+bzklKUQHdChRP
xY8+HRFlXlwMVpRN3M/Xo0tiq4DkCGHurynC/4sPGX4c6sJgQc8Rh1JADbPW+3gw3P5HOELZ41mk
xKPAVY10eLWwNH8FwLCQz6xF6UjVCGeFKlStZIoZ2NESXC0pp3nY2UJkWRczTF1VAvJ7BpqgQrSU
V3swQuRTwFdBZK7+SmVJxFOmL3Oyj7UtwMgnCsFRHfdIMhUw+6e2IJ5hqwb3h0L99YqU+Ym2MQs9
wQu583lj99I/xxRbN8Vlmf9G5SE2HuJti6VlfNQq2XoTf8xaJ3BNFY9hi0xj4naJm13Ps9ZVGfDa
OJzRag1wPujTGzmIG4aQ7V5/J0y8kgmmAjHW2pUyDAGbkASRiar46NVJ2iFuAEWWp6Aa6rKrN1ps
XqCpR8aH0ExP0daZ/U+fvdDevvO9KJAqCyj/fXRrGbCS+0Fo3hNCYQlVuSpJzl0oia68f/ZbhnTy
C+KNJeIv351JDNe2OoZdSuliKQsMUa9jDBz3tQgptRFtJ2dSjqw1tE5mOzprb5u5fSrd26+gW2/m
BoqvLb2m43uzqnK6wFTMFdxF8vmcHMAnbHhGwgss+/Ked8uQZC6orddJof7SFgPqcBA/Pb0Pe/sH
Eijqi1MTGKSQiloVOV0epK+Z+R6wzs8iN82NrCnQKmRil4Wv8x0DliZI8+jySAj/apO8cTlC6rCF
aQRro4LWqEXJAlx64vdXL5n80p1dxjfcAoG2awRKJBqGnBRCwUTdyKPMoe8gMmGkyEPyqR6gADo1
SeMk1sXMt/M47egx1zT+uXPjzNNB53/3IpCjoTwfth3VrAD9lSJGWiXWIb3xwWPXIyMNsHp/XmD7
VB7UYKOb+cXj/Z745wmFWBJFJQuL25ajkXTCYNF+eQDCBcZsqnjQEwsJANEZhV22f6P+TV0saaqr
Aic+HcE6ngbvEswV0f8dqzM/oVRD/3XJ8Pro2myz/trpCi9qzeXQOF+7216QSzpTUy40meYK7y6Q
ZhkFHyQr79A42yKBSx4W82NiZbqXasG/e1ZKj3zKZoEwYvPql6puivHpUDmesl69ZFpGpG4wyoNR
NqOrJqH8HQ3ANQF6lFblOB8uMlbIjbGW7obd7s7L3OqBV3tzrC6rudOpXLDQwcpTKsyuH9bQD9RL
clesZafJWIaWe10pppbnMapII8cNSMcii5mM/1/0E2HL7RZT0MkUWeCzvjYBTo7mgXDHkkWJTCE0
S0NsRRZPLhcQuVp45GBXMDwnC1ZKjlsp14lakgpn90MPXEGxF8G/zBYY+dYyYCMA7YrNRuKZNRl+
M6AOKmtwNu9olcTxlRimngcBJPKdEy+6Pe5QXA21l/5PbCQE6F1w0OR4HeBltFBI+SJTnO3pt4lJ
7YcXw9VC7M1H8eJ5hud/5hGcBze6sC364xuyvREeHerVFq3oMeFJgcklwj6CUSznpgiF3Ai60bMn
ADgEj3cpdyLO5PqA6bmJ8rGJDcLAy7wNlkRK5zqrhIVy2bnYxeI3WEyWRKx9UcKMUfRwd22gDQNW
1EVfIs8gzMfDbhDu0DvyJZNjJyo3IoJd9AD8T3So6W/kgVDqr3goU9bxT2aKyyhS4XgeC1/iGeoy
PUIRjKbE4ahUsI1FPWJkK1lfk+ALEfmdEorqWW83ctb/3FONil5MZS2RP7cqKeFze7+V4orIatSz
pnUiOt5NhIOy5C0UITMG3mY2u1fO6pPJLZg+IkkmpRBMFKqL4G8KhA/hKY6SBKGEmQcsbVUsh/8H
BCKJm3F11hnZF6nnzTs8mbv8i5MI/Qx1gnydURgI4keuVOEtXp7lZcpLHCelbtYPrikjT+02H/kk
Fw0IXm/0eu3Rvixg/Keq8uymWxtKkLQo2UUSC/60dBB6KhBp7geLhm3e7PoqZg0QY1RExObsWLPP
kR1l/wqzfwj/XRnm5xgO+jjXnx35hJ2pSBGzSzgZ/z1ZMYW5llxYM46FdazTRItglK2sYQ/V/+ww
bpse0rgh10QWjfUnA2uI0xnNxfU+szn/vzN3TGelcX+M9aZTW6boCq2PR1HmdlkLmpNVPSQvDMPc
3wInlMjdEwdHDaakUIOieLLdD6wvbnZf1RPfY85zsK9yWh+8PFTQunPhpzAzIlfZQpWt/ka2cUue
FjV/RYkzsxmTJTIKyT/eghEXOVSE5OZU5vm9CXYnfWubjkC4E0iP8akDdLAsQaBvVQG2a874yv58
CZHqUuuYEb50ovFYkP+ZHbQDEgw4ZGzm5NGwZwYtz79b/K5tcvhJ9yQzRAmEBuU49HEMscTO81FZ
sPxKKx7e0vSmtF96GZoPHbZahAQHYPoX0ZKBstzz8M0hldfMkbeXegMn3fMrNryTbGSCm/gZxmOD
WsUcxsmgv/tVJvVFQqSgMApbjxqdhwh29x7Kjg2vj+Mmq6d4B5/+28rCusSPYVzRohSbGf4B0ZEd
vVNgZY7ThgrxGy1PBnseUO8oCClyePLQC8dE8iGq1rXi2mpMBMLQ0z7Fx8Zvx6gGC9yAfThh9t05
+CQ7UPF0BNGQUxpOJ8fiuOLNEUr2YrZKGb5uUKf1sLxNfwNRitPzi6ihfse4dQps4S2SoGM5i1gd
ceQ/uNmB5Zyodz459pwXA7o1pTiVaIPNDqdGMhZpKA/67VqXXH4AFWRhmM8CxnH9K5yXlf/vGAyR
amjgEd4cGGuA+wNBZ2AgxQJ45saU/jwQ6DPXdDfjtyIwsVAxUlRkCE+GaT2CUz/aCe5Dt3jIoauF
Fm0qcVuXMYxwjgUIwFvtWTS5DA0TFEWCCv1L1Q+9FMZxheg6G5LrczHbCDlCc7n64+1VGNmHBb8Z
+R4SJcekhUKnf5zR02i5pcX795D3OC1HRWVhTrSQMIVp97sTka/Fb7SutvYZ6/nRr5Jc0UoX64WS
Cg5eSIf1jpSCvQD7y88Z8GZesmtoAfug//kOlthEO9b4vNI00jATRJph+Xbg1IMV6MQNVDfF8dtK
+2Zlxa4WfPSMCzjUMNoygvBWXI2jL8q9W6xCeIIC4kzRZHEPWTxLQ0iCLO337INPX9YDANgq6bPh
92JW7V48MQZS0hFici7APNFZjgsrTfcqXg9xKFDjQxBX1cehCI5JdB5RIEbeyEm6aHGEzl1V1cB6
hWq7/oTvdlJLRKQYqfY85ei0SIQF00j/Zyi1UVwdJ80CknNrqTGp5yB6Es3K3ZukDk3FR7uva3qv
+0NgyxnhjYUp+Oi9Du4V6K06ak6saT7+vb7scstaknF6SsHBKUZlYfq1ZER7aZ2e+c1dsck4b3ss
3fLjw1cjEGsS+zGKx2RsYKz3eVSOJPfb18a7iSs6SFcseFUCRGa+tnlXhUxj+TkuYAyALFyBFyVo
jxynXC2TXsGfHucYtWSuO0Mky0sGmMpIaYzA42DFwiCuGk+UJjkIArDr8lG6dqIgoGExIo6rhVWj
YYh2Ard6UI4CIFE0JrwLXzrZvyjY8ZoNF/AFgsLpuixlyP2GgziMKMsqvRcNotN5ikXQevvnlwN3
0+dEKxjvqnfODM65F1edHj8iwFIIFyiA5tfYdKrP+Nk02YPX34WFaKvS5rTELiW6xLo/KTrw4BvG
YcVVcNOSeDUE2dqlpoGiE8zjADsy03ZVmC/F8PYIJZBZ6iYUX4WYaTiKEcNYi6eVs+/wOH+b0hDX
gXtSWL/IehFwc3z5YFEn9h9HdTz9vusHmx8Q+eLIMDH1KBWhw2hy8OfHRt8SSV6vtT107ecSxW+5
d/QvLutRO7lAVh46RnZJT49mVx64nHSeVNAajVKp0ec/J8MzMdx8mFr+ZFJ+RSLyBUVNX7ARAkZ4
O8IjpYv3bSacFaCmB9R4egaX2KaFFHrBc+5a3YN2Rv7EPw+ak2Trx1wu1irxLOjlD1Cd0H3uE4s5
AgYjs4jIB0jhK1YmQiwxVUQd8id9myT0Cx7nc6PpCyWWYVWkugRtYbLWvMxij3nEo/iPvQjFktX8
KKYQka1tQIiHnLuJyLgL4dqjBUFgXqor4odVwY3QU6nl8SlvjzxkVgfzTjms+ZWHs+ed+ogFzseu
qcuWv8RPkCV4RN8Vp9woblBD5pyPMJI/qIE++0CfhywvtckwPVOVS+lDdZEAD+u5nYu+h9IzMRCz
0kwuQtCj0WdfoJcz0sq9mFuDKzGzli3DICpydO29DSy5JgL8stLh6zFxDUNiFqTdgpSjszx+sUIW
SqS9gCoS18AbT/XUvtEduKQRhxKl0VDczzo1azyDN20ELw/83KEleKx5x/cbQ4UihS1vzHoimnea
Q70y19CzXXUK8tfp//hua4GWffnjR1qGXPjQSpx6bYDyKJRESYWVMHb53t5TUY9UHzAbMonqx/jf
QReGPwlX0dIJDV/Fui7dMTfO3q0QXkfoDmbll6slevqp4kmmQ8qlUjsvXOBNZPg4qARCki4gtMPi
l10TR7wyjcCxUfobJakBFgMIBAoceDVrv64uVff7AJkEuJ9EOBI3YvNCwctez+Ft18i30/RFsHlb
TZgklPnJtOZJi4KiO1epr7sSlm8rITpdBavhT+xhCrUhz9Z3pptzk3p/89+00Gu5m5jpWsBrX8RA
qxqQnhkYfMJe+NDMN0qYDXnP8/jIo96Vp6K+KWms7hwyW9F6EuHD4PRvl/Nk1rj8jrHFLzH83d/d
TePf9t8detWzJDVyeL8SDsDokFfSGBPi7eaowLzkIk0/hE+QeEgfw5rJObVzmmudl7C7d849UpYU
AOeGNlPMYsVunQxM03dKMFKQOHSw53TcMZ24L+RYb9uo+yKUE/sugnBkT5/Y9/Ege7IAm8jfN7bK
EJyVAp+wYzygxV/xwh6zRv6uLKyOoc6e7yuzHZeSQwLjppMGGXEzWoEDuhE+1hEBGYmJmEi1+QJe
a4UbtOHJppZjJ7RmaY8g83zuPwzp8LJ/LTi7BN85OtJGc1uBhJnbtDmytHjJgLJ3q5Ja/GScil/1
NPVTp+ZKT6e2V9Pts8L8eqgnQuAqm0iYMRKRsYBT4Rreoo3LyybYksLwpyN1bBIgFCq8QV7zfOez
PGOqzuQHSYw7ARL655qcRWdqf78/R2hwzjJf5iUIC8XxknP1WesRoqhb+L3SSoxc8+r/OwP+SeLb
DSLk54EPVXKXGw+HMx/WEylgXS9wijnnfs5DNRXoTgwUTB/+CSlRPK4wZhR4SoTBw4bnLLvu59oQ
579ptVIN9sK3x8xqRIERmBOa4JoQG2HP89mvSs3zFVM96mNyB4v7iidsSBL+WqKvqlcEKo8BHCjK
/RdEEqhz6FN4kTmJkUQUNMTE24WvZ5nrsu13suRnsx1gVTHgJLrJQZEa657Ptwsd67wYKm2yJR+r
ZySohEoSM4HLsvOKuspSqNIKYOpNYN+v9I8Ei6ycmrDPYqS0Jcd3nveeHCiGbqrMUfNvQsHgo/EE
U3AfpoDG2ZOrnAaxMTjCvc+kG+0XabXOZ1TenC12dMXvO7XHVWzkWP9TH/8zGMh7WxBn2wMXplHA
bNFb6YhhKU0zxMT9wATX/G5rpbcVeaS2dCY+IljOT9+kvRdB7fLvATy4I1ebJ0TLqb23cqPra68E
TcY3XiyuDuuIqiPPn9NufQ4jJulF/M9p8iI/wtBAvslT2+PmajUb2lKbg6jI8MTOs09h7JB0wS5t
8cHwR37QD74VZ692LHgj6sdLy2gQkWcv4q/sDSpPWh/mXATUgmbw3P9enhsgrnZonGDEv4KIxSP8
uAjJk+7/2GxUZ81mQtesfjSOj23IalHN4+CCY7Es3OHOqFpEfk6DUHYrKM9TSl9JxNN81dLuUH8P
gOiVLrYmbJMLAZeTTT2lL9NVn4Srd7DLZ8QzTD+RjOZDB6qgD/0OewzU+il6hcaA8kvfGijoilP/
Cg29Fggf8MvAGoBOwCdNnmHENakXnandccOVZjcTB4n5RBC4HK8y4Z9Ajsu6Zzvi07QJVcO7rP+C
6Ia1QBWyWD/qTgr8RuUKwaLnZqFSP2rfqq2ePzWPMF1y6wMiLFr+AV6v76O+6vG/5vDZX5+psVf8
Nmvof6HE8oG7FmaGJjtzkcZCF+IapZZETV/ecZgyz1t9JJ4D6eigSlwsVZPlF+LfR9oRHgKYFnxl
HuU0Ssl0P01FPYKMCtf0f4PPCrvjJSvnB3AaH9tIaCRL27/KvMQByZWZKz4ABTyqrA6UXqGLOcps
WMELqn2WkR+6JGtenuOwxj8VWUE58dhg5cH0wFX6bqA3xbMdMXkwveL9u68djwEFPbLvOIBUxJ7M
lzQAkDRgi0hXNEDU4r7HGk3ouLQdTNqKT7Fh6Sa8F+DdZISOQpuSMPrAEbrIGvS2pG0fGTpyoIlQ
9NXRHOo3meiwWKOvIxzh2xP6P4QSyWwaL6OGPDjQDBpmZn9a5M2b6xHEb5VNB3djHIcwMRkB7jXX
n69W5qx7JsMbaWb1gRn2u8u0h4FBbYwpE6z73XX5/fUlPnipM2isbDRbW27DetgEQwRTpQAZQqVT
QWztKBpXNTUmNQPpF+duJh5Rfaxsvidc/5ZHX+wUQV6Pa6bhf5xl2ATXsb+SGk0+ZaxHu6Oejaa2
x+qJ18ogTb7YaiTX4zuASDlvvDkiwpedQP8Whszj5ZwJ1ddSRfID2fJRbYunyGlWyu9gT6zaTIOx
xeqpScscYBvuWxNT/83uAoUp12gvuEwLJ+GGwuiCslvbldRrOKktrVPEIhqB0pGLN+XYIk0TaNUf
QHqqL72q2XimGErQko7VO53bKdaofLxBb1a4yIcT1d/WJzS0M6yd9AP4StN/Z+X+aopddNpD/dLq
iHxYDOZshU+cI6PSy9Rm3cXxfQGOCSdmYkLr4SwndAvq0oIF0gr+56npUykMUxWFGZGUnA8818YF
SLkoHJz1OQxjuH8g3jbq2LAobSQfZeFc24GE0scRpYPw6FNWeKFfsYuXWmZiRCtP0dKnxGfziimG
JKukxL/BFuej9GrI1rItJAvX+yG2CQ+eh6H2OoGbKlrlHczdKJKEVmzTWU9/FMqHfT0PZR27RtIn
4tkL6jwA6TPsJ7F7DZ+sF0FN5awh2Jpn8xFTw/LND83YB47Ki7yyTDu5KwXtz0HrTcvrPqxyL2wZ
UuxNrye4y4YA3BTK7PWXopOm5IOWT9gXs2DSKH1VgPHcXIdjI+VruL2uideLTyTYMT6HOnJp6RwF
Ymq3eYgxrMRw/QKSMq3VWSN8YNOTpMO2QvBJt7tDA5ZTQPUW6ZDTcX7894fxzSPJ6JrBTz/9b2jM
+HTErBuDQA==
`protect end_protected

