

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YWwSN+9l5ahBqN8tuQHA+pe+2Q7Fh9//dR3H5K2w3KRc2pla5S5ifvTi8Ak4V+dzPFwrZE+Uv4ZM
WqK4mWAaDw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WcjiphsvP4YifX33L+r4vrauIXRkGno8B+olsJNjoqAxagaZzNDAFnvGiJsIWLTLoEkntxsgRnIo
WVce53gFCvnJJkmdaYhg6W308/4ThcXkZ2dT7Q+TUTpvKAEe2vDwO0foHspYl4iLWX2KqDyY9jge
moxvN6KH420mg96l6zY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wvng0RPku5m5MHpJv9WwJDWJ8F5PUKDSPU7V99zR5erdP7PcyDhypTKxqOMHkizg+gEusr/QYxdH
b3OK1yRKUZ44xzg4dZxpsvitjqx51I8wGaS5oiuyKX8hGtgTVrbfoHo6u9pcLQZn9XK2J/iSrjf5
dyOg2xTIXw233HzwIrCKg5RT8dfxa+iICMhoGVZIGJ68DJPwrJbT6Swg5gWMje7MS+Ppwgv0Jxqb
7HSKZuEIyqOKVjWI9mOWG9o9+LBatVHO9cQqYlFkeCwc3YeZbVHELaty1PZ3GYbJhCtr7obXWCNH
f42iQcUXnPWhD7j92uOOj9mnGCfQwEtmFpOg0A==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mnRNLVCxq+sgQJhai+B5fZRsJzZ93rdvyaCrmwTY5fIgoqSgRC5N+TQCYgevu6oU/nSzurf6krRP
lHQ0Ztrjgg2Tj4+uhFcaWXWp3gef6Qsz8XcVJ4aB4xMaBhgkUeweDC7vzOKD05WXxyBd0/qZdLtt
lS8j7xW/2WXeJFqpGaMZ30TpyNYKEPbTG0s7zfxCOI79Vadm9yVGLdGkntvGV8guzxeaRo2Qkmsm
e1+jXsDbdOr2euBE7JiOnNqartejTWUhtjRbkQnS4YCtUcNrW9+ObOoPjivEDKhArV2d5T5dFhZd
vZIU/RR6j3BExhd071LKzolsdnCqR62C9tEZ5A==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
E6549NUXinEnqZcngO+xA/zs1xe2Bus1VEuxweH9iD+10PgNtRJtsG9EF7ZdZas4DjOhgJh7DHf8
ndbSlKTeJx/4QdIH6iyjSx9xrJbjCC8TeQlSsBzTcSKNDMh3HuElLUknuM+x5+UC+hkdrw0waGjh
tjj70YkP+K8Te1Nhfp5PHo+OirttOLZY7Bnhq7x3KDxVSyWnLuCBlLcRqRosb6oaQVAF5dnEKVG3
DDqNFX/V0KONWbfs5QSo5gM8f237iV+nwxPmst+L5casdH0vfnMagphcYI2Gs12f9zJ/qipttgTQ
46Pj/rGC5IRv5Z5f3c9wnJBWRVPQ0uHojBicwg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ogp/UkagRFxN6D0Tvatf3PJ+RNRc6aGWLVAuekDtCdp1urxgWDpgdUpLAqv4gVFTloxR/WYTIPAy
tqnoQwfvxF8+1H1sANWUqIMweNpcUZzEYS0M2VRPa5yH9GDRSd+LmMbbrq6RbwvXiR0tPlJ+qF//
xXzjGxQQlbn5MtTPwO8=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WS3NnUM3tGvHLrK1+gyTpPfI4oWwTOYDJPYfQBcc9ol/GaO7Z5AyMRqRkk+WEY00WrbCfviFYMzU
pGl2IHT4VRRzqqLR91kr2OFbN6OGXGirK/a2SoQqoRH7NbdhMzwc2r2DD8mzssXGs2HnjNYorDiE
Vs1axIRZ0Xwgll0Xql9UnW3+H+bZdCSjNWd63t2LxcoNPpatkn50Aa0uZrOTFNGicGTTryERIIjE
tD/W23CkHq3rM2LwJimtfOkZfT6H17TZIlmdf4GzYYEZqzxs/jkYFtiD89KMP+/WhCVPGWSzHT/R
ZumbUYGnUPG9wSLIU2c4b/c9CXNngT5yj0uIjA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74224)
`protect data_block
ejA+3/GyNSF5c2mG4a+IOhurK6tqajaZSjTyZ1QUDyW7d7y55UO1EWwYkeZ4F5ePNMk7J9GCPl1y
jVpvgnPV8QsYzKp62R7yLxM5XdNBzaKp+G6UwIM40+txgZmJV2V4RqZxJpKnEHDz7sAmj+QtG0JN
PTDWwF+2/Ch1xDTbfTOKhtvQBm/3/mgRBLWoB6tgRENW54Ar+iyWdZuKUHWHml3S5uZD+6+kXwdc
u4sJDqoGTF7dB1Sy1d5Rztz6d3TnFnU6wRZ8w5t7X3gOUjrPkekF4b7UvjXiFCm7Oo3wwqE+FXJR
dHfzrX43O17uNLRZHBsrVUKMczt0L3tXGkeqSuODHYOPgJ4ts123u4BYnvGYf8iEmdS7hHYkmJ7/
JWGwi76g906Q2Wu6I9LdSLreBPOg7QYJVtiRRfg+jqTKhMxk/97RSy8qyJ1ul2VkyK9urfwc8wpX
Vv4INZGNaAcgzXjq++51/72wvmOTTsvss/VMRvg1aO7tm7V6urAFLUWMhUiF4GtQfauXj94fRf5W
m/oKJRwfip++WlJmK14XnefPsUyg0moi0S2vDc7HM27YfOn+bxeDZdMviy88p6ahsbpqmT2WP9Nb
2n3eDfkvXVgyNmpXwmxEBYohU4jcZVxPc8u+Zg6RjomDLKGKKWA17tTpICMGMjxbfHwVJ+5YHcMo
dqCSbqio6BJ7B8FLaa8rbfLOSNYg0mhiMf95GxtSjXNw6Cypu/HQqan7nx6RqfwSARlh5U5Kr4gd
LOv1Ul9gxD/dkhM1sqzUpJwsPit0SCX3sz0IurVyHM9ZxTAwaE9qGqLQQBoktDT4l5SO3awNGIhJ
wmHbjGN5HHRug82KLtbFfuL4O+aGWaMHz/Dg5B77TDMdJrS4fSpwYLPDDaQoBgI3zyDYqE3txX5r
hhA+gp8sHkVVQu0uMUE8BU6ZlWfhhydDGpiB1/zmEGB2tsNOyyh19g+hU3k+kS2/2BUnQwlnn497
NIcLsVozOIckioM4X+qRDtiSTeLxTIcTYlZoa8D9xSXZEV/EoJ8lksqf1EzGaHYFpi2tEHL8muhI
8yoIg1dB0463GHjfNZLCNrAjGFDVyqQmGqqFrDyb5WQAzrei7LJOlpIoJt5AfIF7xGlS9EgSbNhi
HhyBO1gJkY+mSn2E5+BkJnsxyLjtNb+O9EjWI3IelNGeOH9/ZfAzhnY731Mi4PsvUl90ZTTt3uzI
IH0+38UAOmNDUV/9CnIvS/oiT9AZbUGSaBR2hkSHwP+yso6XOcb7SeN2CjI8wTIaJlrl2FGDSXx8
gSLJxUBSEHXMUcqWk95OEHv51hau796PKKQReAVypkvtPLpqZD/+NVMNIBkHLE9LWA5FHa8mGUVd
qDgS7PiA6ZdEH6qkVUAPCO2exbsVyMqwHZ5H/1tm9eYXx3RP8oIySAbGoJ7eOdJLlW8qEBreRNEP
60UfkjG1gZxfdka0ilC675blk8pequ6xqY7XppxpAW5SHMxa06fUna3doXk9ziGaT6NxOqCZopPJ
Rw8NToofMmM0BphVj9JF/Vo0VHMrw0ApX7Vekuvs4huXN9U00dBqnJ6XWCleP6VGs2rLzqR9RHYr
4NJ/TCVAyP3bvESRjrB3ZRgoMOxGbEzy9waa49pp8eZ/qHVmHKsm02owpjCfzv7CFArfHdjrKYNE
AAH0a3cAchkZCKVn2VmhslKODe5T3htoETLd59W8cZyHSodvLg2p6eps22m3rgZLcbEFQwd90Ed6
fXiqXyYI6l7jSp5XtcBh6Y6wG6CMYN3aOnvVze0fMDJUv8cJuEoro9I6EPRWnfXFFaPGTp+q3yLC
xpUWYaYc/B0YbOHjNlGhDyiLErWEkZvaibEIfZeEknNPQ0Hf/X2m7U71R98KCEnEYeyCtb4OLaSX
QNniYZXTRjtXQruuxdcTKvQp5nsGxLbPi5Od0+rpL1sE8H6SGptsOAU2WtCnoOnTYxNX5wp5N1N+
lo21hnJX5v0fQ6vpE9cfLC9YvtRFsZ7fE3llZ1AKgQDfe8BrU8q82wWpewpm5ErVqqGyC9AXU4xp
DmEp63+CaJPcC4XpxgkB+k9cvEdqDZfRdeeyvMTfDJ8DN0ByLczID/BDcB0offAHvVg/enhKEnXn
edeLN88dj7WIrOxmKJPKNViVxAS6p4H4mwMpmJtcDvYHlgq5wEguOdjBqJIHPKqscRVHKpB3nv7D
6dgq2vTWww7jag92EyY98NIXV3K7PMwREZ0Kc1tkv+jtTyXclqrDv0EqWidpzGveZsMhm8C/HZc/
K8SY/w480J7AMEyj/uCzT3TyY6VmZKTlYbTYWQRXWf3C6OmWebOajhHYdvVvo9IqdmnGQZSp87DS
h5MzUddQQ4pt8s4FWtDr79gdrEgrvPhToyGNJvlV2tI5cJ+SOJGbfVE/RbiZJCdlL0jTDF/6UibK
J2K+GExHa/n1h9Y0aaSR5q+jb9zjcXLQXr0CgyK2ysa3AyAWVeOzTZ/XnyTZ8D4hCQlZjwTYzff8
38uele5g3HKvmWoZBKbKKsbQQPj8DY+H2nPigNftlEpMkQqXZbxLQy1p0y/0RVdeRF+Wc1DJcjYu
aEz1Ks1afEbeloxUwf3kfj1G6CimqI9DaD57NAie1saKREoahR/rs7ZIXhiKOBztrehV6AjMxQ9U
cRE226CBnp1eiISXE5KoBDcqFeuIK+f9dqlQZKSBo0WkRyAXu64En1WjDUCfPsPvDD03bOSFQXgs
ty8qqQyHxpGLnVqkktqe40VS7+WzW+u/+8UaWl1VZpbO/xrlpZAIiXwZu/ybl8sTKwkRVOKSAsJy
DcPEufZePKHn4SE4GldWTN02pKVNeqhRNYnQbYxLH5o8tjXOFr5BFIyz1W97EafsaMurgw35kxcM
0orsLQkBcz9Pz/8a1epxsJcUHG9uQReBS2J/dFiHfHsq7z6DiPUkl3kBc04Xqt1UVCzthyoxEmGj
WfRBZ7bknEA3PdNvuY8zbnRCnvfn2sN8zrteIAFTydNLIJ5b3ZLg67Q+u8dCq8CyUUuNy8Wm79zP
itNaBeAJSdudtorQTn7vILlYBaqC/jEEZHqDgrccQaA6RW6k7W3Zypiq3KdBXdGL9zCuzoZZQ15f
Wa/xVqjz4C+snt3P5QSkPvTYyme3HrSjQm4XJVmfEztUyWbxtR6fqtUkP1imq4YKLmMn/eZ5NcpW
MGr9UFAEgWsGwF8ep1aXYm9hdqaN5K+1aPqlEJjEhpouJVYTQ8xQzy8uYA9TbL0hV192M2oKU+Fi
XjQPERXBOIC/wUm3FyS5GETPrlaVxmfpDaEtmQsqWxtqX9ICAF4xVy4qPuSrcErf+Dy/tjdDvYKa
PXS/9PootEgwrMuXVNvQp8H2IG7MSw7ttmkk/fMqUL/j9bzu76Co9NGd4fOMtHPTiUZVGnx0YsVg
vhTIV49mloIpN7cIV+oIzqxgVLF96m7UMFMvmAEB+rg9NkLV/mCkBc2dQUUwJL1tgjBXimHQ26pQ
KzRzQuxx9jkPKyykeYYKBJdqG53nXmXb0m7anIFmtn+uKk6qcKS6OoeeAaJIUp/eT72d3H/VeC2D
YB3sYRqy8yHb/qa9fPbqQhbFweXbtJZWOOde5+rYnLFk6HvBe+WeYXWPekyZTmWe+JvIJwcDZa/2
Hc/d68crXMQDDaeNHtGdkSwdZW9AL1F54Hgera2uqkH9freXs+6u5JWD9cV8PtZuCkoxANPleipk
fP7xYgm/lSKEpbu6/IW8ihs6fuLc6DfUUAlF/NLySh/Zys1GqyyaC8BZsp4d7xKdME80UQv0xCuj
AReEk7UoGq7kVDVTMKCzfw4ZrXNxSKA5HN1a8sFg3o4VkbX2Ar36XUlRywR48ndEBtIq41LeFCjm
1xG73h/96s6gTxjR/Zl+6AIb10GU+V8ps9aRCL6g/NGn+rjGTFv7tvk2V+l2OAFDPzlBWQC+mB+K
pHNww2yd3/sO4TsO1IcsBUVaYF7x5IMHLii90l6po2EcVtKoNdeGS7Lz4UpIddm8JvPef4d6SP1z
unjOgFBRupOyRrShf4TMvFmvCKlbWWL25J81bIHolgUDdnsfebU97zXfKBiDcoIsb+w0+31kJYQ6
1W4i+cAT6IxGenRVt+/5dcgXqQKvCElajCarxf8pbskCwtwJN3e8KjqnQBZ/0oPLncDxKB7ZbExb
FCEguDi3nSHWZzGRSrN3QTjxr93PVmCrEf+rG8Q3F5KyozgMhAZPrLLyCRZKi5BVErdfelzRHptA
gxS1lcmSK+92as+/mWxnDSQk5BfnJX+fK3sX/DHoqfYsXNTXT9woD9cCoeKGFU2wDX9kC1M6k+ac
qyViW33n5misJA6+DDabQeEJNHsSQ37leZ0H8h+3VfxGlt92gGsldpChE0w9Bm5AHbv6R5u2dVt5
W8wbn27Z5O/Xmiv49C3mdpERO8addnv49cE9c2Kn7ghOksA8d53fIW4xBPBtaVxewU1OArIovuUK
CFn7K8GRL0iCXKBgEgT9bEnqV/bGgA1o7wegifNliB5aohYAjxnAXd+q8WYxrGz4NF5DZQDexJOc
fOmIow3hj+0hJenqgu+8J4fYqkt7Ys9yng+iQEhgWR9gbLmUoVaAZ85B9poljVNatKJgKcjhYWA3
B9OWdcW4Aa7c7tYmTeQtKMtv10R9K3X/DfKCm38RudLZjjAM52RdwREeiTko8YH77AXOw5jkS/JY
TxCjEEQxAynU8GmlxwaleNvIAbEPeb8MvnGj62U/78wQBe/ovBMuJj7BbR8/bWUwY9YjeUMZMVjI
AqfD9CE1YKQPZ8f1qm1TlNZupuUyvVyiPD/dfNvo0U3UjIoO57TvsGSMkagTFI3gQADB7SaN8fII
qraqbvF2Gwp67fz8IJlGfCTIrlLFxGEX9aEJHBhK6rUXYAt7Ki4DG+mk4OFeFJObaibl/3x24fYM
eE/ng2+c3EK9YwP+nG4MP6O0ZjmEt2XA0/4UPQY/wd80xgTqugUx8ODuckqg38Fj6AH5WDSP54pz
jEL50cP1VWh37vWPprDL3bxa/+UE8T5oX0rZ208ZIEHORIA3WdkKF8io7sEavoYlXikrOxSSrq62
YHY7ZG/cFlCIADGYaer9zaUju0NvmcYykuZqL7jlVkrBmyXJCBD6u9jEpjDACUt25SqgJGRAG6aV
1akVxs3F1RnItTT3TX3F3w3xLr/HLIfs6uoLIOZynTo/XCni2KoqosOwhdgh4i5ubxO8n/bIzqbi
BBRWgM9Po4wERwY1O8nXKplFqRAIXHM2lHFyWnsP708KJN7ekgr9QxK+Gr6Mutza7k5zbx/upRlL
yV5pCW6Y6rFpXbgz+oRukHv6gV+oUaGjWg5ElBsofL0Wx7pz5NkBDbr17BUYNhnTMLu+IXfLBJbk
/bkYq/vL9HxfCF4M3abl3GOhFwXRem6ixX+dGfmex3s8ddit3Fm4aBb/JmZ1sehKJCkXvy5lipKQ
hbNFNvsIC8SiyJb0qUcM1lZ/XxZ1gjW9x37t1S5xT4VcMfjEBFs4LsvpqkfxolRw9fhsoSDjVs5o
qKNWJAKjXaBc3/ORpMyIe2OqZcIEaHohTg4URtONEL0/i4LkxT2C8is9s4Ko8bAl4p1/xQQKsoZE
TD9DY06Yv+Ic6AWqDYjlyplsO65MtYKu5nm1CRAfqSAxBHWBVd8s39qDXuMf4c3AbBEIddkvzcCd
7lnL3Sr180faChIFPqkRbvb5A5HTuoxfAtXHkM1nsuefEQHLffjIwpZCZxe9u4LJsz+0Tnp2dUXE
q9dTHE4J0WZ6hpB4A2HNEWEs1naKNwBAeP++tTKw7lVACI1eVzR1i4IaAX6znNGdGlDL4ep1/i3d
Ral0F6ywV8sHala+sHudEEvyRch7PQ5Qiq4Wqm/z6g/jrm+7fmFalheFQbrH76037kmiyKM1MzZs
o5wrAVEYYKWU8bCaeKzkXfiLdHErhMfWokToJnY2STA2DVjWdOLz6eCaqyswvn1qqIWqaGBWBROq
7ItEqgc9l/FhnPXe7Y8Vh2V1i4/S63xu7ZgkptCR2qBSfq7OOsf6B3ObK2mhdqxVjX3+CzksaTSw
QJLKHfHRu2C8KZXlFUwL2CSpIUOEy3qGhP9J2z8honiBuQQ45+n/G/EanAMCl8g/A6GNshgdj++9
godCZPqwN4hCwBDHjIGIaPQbHFfN50dzyrDOwU3uB/uyUz4g2yxIiCuN4f6emMgxz4okEENhvga7
+REXBf1u/7mPaUN9v4KURdpCEg101Q8JDPU6TmA9amgPcYdtc3Ab9kgr7PJ+G5oEWRQ+dtD3SDRj
CzYaLMtZPZu236uhFRuOa3P0d+U0Up0OiZztQ4aBzG677Np5/t1VpCrYAsuFl1R30PLyQwSA/459
vsAs51yQaqboSkU6aYAHi4Uv+hT3a+8XMbzWpMvjv3gxlSj6z1kXH0qGiOCGCRiWuXsma2Z9F2fP
IOuxwCIb25zJOLLZia38GDth+M5tpnsbut8/QZr8eRE0mjedHjZ89E3pMJO1QQXrWsloeSXw18B+
ORbIIfG/bAo+zwKVpJWYdT6NtCk4HbbTlGSe7lu5y3l1TahEOETdwrm65AMOwKoaZc4gu+sIKR76
s4k2KotFX016UBCfvzfi75y0wqebJGA+qEfQNGr+VJDLDPoZCoQzg/1wlOofWQr6Tm7dwkvUIH7G
KGj36TAsQ33ZkOi/Ahls62UghW3GIbDK5Cg+hX7/H4KBprBSh/c1aDcNuDGiwuFeR38w8H083E1B
PYrpB3S/wuoEvnXzDUeQwC23n/D0RdYCqul+tVEH7bGUW97iB0GOGux9GlC4jbLcFicSQAtxJpVQ
xGqCOP1pcmX1xHikeaaeyqPHWMBtYfcidgMt9d+PrdaH3AV1qo+jNlKFZxFD83vwq8am9Unr4dNF
Uz5BmtCzzK0/SUh8Rqz8bFhn0VrCohxeFOZ7xLP/53j5u4zeepXtN6GqkSjQtAsxL6VtXtd2lYwk
SH/HxPSa6hoTmzYwORNBpQ8aOVNQQ20EKkamwdtMy6IxXWo11ot5KXOa9pdx0W+2fQ8sx88PXzX3
9AZfIJ2KKLldKkvYU2winslm4VDdblXJ3Dfb44DZQZMXn9Z4Ss7wCE24Y7y9yI3Fa9R0GF0z3dJT
Ub9SkSuO3+ihz9hjgrT1t3xEJF7yvLB07wn8/krdKmazEoD2/V1uCZ+3cv0GHJKbKVkbzI5ZTK9L
aeVVOQBtA5UZ7RoaBRnheM9Kwk73azvKwKdGLcfgm8LnQgO4CnCoU/tAPi0BDEj2Ph1BQsg20R5h
HN28wKiXLsdbkTJ7q2NdgOyyWXWrU+/AUj+fGSxUuFrvHxNkXo2a15Dl1VLs3LYs8NTtAtb+FQL/
NoiB0k9wfrf2qSm9ESzzKS6oTCc0MMTngUV6Nh+suCeNMo4q+ap2iTNW9CoufJ6zVjRy0Vy+Ps7e
bPEV4DEWd0rMspbZ6sX6rkHCg+hlkzZCm4SAveyoeOpHDMvDlAREvtbJC8YutgErLlYAKDYJno7V
UsHgyT1gz9RZjfgQZykkN04wJrnxQW0V1Eg/lbCCfHp5KP8WfdJRUKcIM65a0f1ihVYVzRpGgrNH
HaD9M3HrbkE/XiLAo7n5FukE2EqLRNaySs2qBkn3ujqUDBXMDpHXFDSBhefJ549DnB4OGZX/luvj
tvownV/hUjcsCmx3OE/C4DQXn3ZmxSerEbbESc5zL/WY79geU/m3t3ltAA3HJrP4/2MRGR4Uj6zn
1mFRILlrBHvxgk6IuqwwC56UH0LiwfXFj8OIfcOi9XMEDel6yaluMpvNv2wI3MUFSW0Y3Brodxtr
htoR0AS0WvLJZc5ks6ODNHdkbJfymQel6zGfA9dhHuNbypV4EHaeADNI5vCM4aMxP4qqBObWQjOt
v7snT0PbfoD5fV8lab5NT7IiPekjMRUS49vbButdBAf6A8pDn46JY4mZK5xboq3GY0XNlxvujgEI
7Udoqnm4L0MhXGK2ORCyHvTxPzTJuceg/vc2snO+/OXxiOP7geXAR35mdIoUgMwiCjEycWCcoxiA
/tGU4fqaW7c5B3TAi75QheMidHgHUTb5/bbspH7SLpqf2IhIcbDxlW/kw2c5G/H0z4OaNFgeLCHi
nacX0qWOZslAgRID0m6mI6eagjr23Vro867gr2III0duAmv7l2RXPC3WA45pStJekUVVyFYIlYx0
c8Gq7iVT8KuzECpS8qI/lzu8XD4JSUiPd2MRgZTRHSbAHGzlovRb7TzZbWFRTe8fgVI9V/VB2wEj
e0cX8pExUBFCVxlHJw+Pux3DSVbNmdkTRtDEDOkYCNtd+w7RjEoGPYjLd7nxUkUJkx0a/8rqFk/8
VtD9O/GybwPmJ3aUS83jC5BeEHgkAxQA3pkUzk9N8uy12mOMRRPc549+H+4fXyhiO8hM/OQXJH/9
2FZLf0yb61gnNh5DgWHhcbshTQvWSs9TnQP6mUoOaX0E4vYgcJA2we+UIvD3ISA3EQJbDsQ1JLgG
tTw3gjT0k+f2vzmn74CJdtAJHxuhRcwJ5k+rUxX8RrbZHSKNnP3mbecIlC6a0fNmyagIC1lC2DxY
1CbsccFxqJqmen5FbCrJrRjInQjjQuvjXldyvc1Hhp+vNtoDt3lGoTIrEb3chpCyhk+sHOcsb1Yj
d95Hmcl68f3kU2po3Emu7nIhoVceYJ5BbRHiVqjaNR69aseLFCTpF0fX2APC2troRTyWr0c5P5Zg
mp4BLFlDmctBBcv5zUnhvcYoELEubueF8fnQLmbDOoM8Jf+HnCebSBlWwKdrYEObmQZMV9b1d8Fx
n8dKsF+zyZ6fk3vUpaW3EYGd8abYW+/ZQJ7bPaz2g40dMFtReHM2VWRvOtzR4l6h0jWLRlMzxJ0r
FAThY8SZO5hr+s2mfP6rGL9djAVMdl7cXONUH2X+9gkKUGlothk2DhEcYnmlTbZrbESygWt4mHTQ
GzXEY3Xg6psQCPxk8PZsAEUq4setN3kfyrrFX3vUkZ8wTDIL28aLViduLmlKGkrV1H0C7+5sXLdO
8i7IhJfqV/T4dGjZt8QZ7SPQaM6rl9EMAZWROrIIF5VAeebXtD28HaQPwXc1BJ7VumjhEDGpjtEi
YlLx/VAI/ZcSXQGzhp4onXmeHS0sLYqsW92qRE/w7O7+Ir3hlqMtiSUro2DJVvn1b0hOtK5hDREW
cD7lc4GY4T46ydNcfMvW8UCS+tN37c1DeCLV2a9x7UwtFtyFAmGj7YysKeoB2+qzgHLJl6TrOS+2
Xd6qxNucUzZmWNgsC7u0owM1skS1Z61dL4VAwdWt8j69FHEI4F3hbOEnznsYH2cS/gwnAB6BJGWc
NCuwcC8fJ3PGVnegEMvMeYBEWetXUj3p/AE4K5XWkSzpyY3kzjik9SIf1j8jr7EOhEaH/LP1KC0t
A56ZWyCCZVMEHvZRHSR+jlpG/VDKbodTbT3G4L+DuMULxcDYOxRYQ+FAjn9tsdcsBoBaniYoKdz9
BaM8n65vMuzXSymMV9HHlSfTGMIZjnTFKhHW2tdkraCT66C6Sg9hZz0Ol8LVlp/+i0IGU4KUE4hm
71lr9JIQDxoC4p3U7n++Xz6eJTBn1Lt7GsnIgPB0YbtLuutR1sM3lJZD5vcLT5z0L16E9TtoK89R
2oT56Q779/KnfLnttDJNMqmLMhvZlXF8UXbtLoktwMFwA/3dccIwL/Bpd/gXZnfRId3w9Kcbb6ai
ZdEuUJdD68uFMRg9s5JIhaRYhfqrfNRXcyrx9fqEtYk7RZQhhT1YPEv/UZYbwABSzcu+3/JlReS7
dX0Tl+kQOgdFT50XA/+OaS6W3eccGowog4MLYd6ZQw4NR6+fAtzkxdw99T5gHgEYj7p5QiotO4a4
P8NUwEunldEipKB9YAO13LD9vvc9XMjixC2qVmwoac3Cqxsrrk+NCHRmvpoC/ee3CJpx0vc7gCbU
MO+h4Cnl7oSwD/n7mqJbSkOnnmdnz1aUpVi7RODLAkFhmauo37/0lFlU2weRBdYEKsK5IKQR6DuM
lJ81roQuqxcTJ3ayJ02vzjxALqe/FF7QWmzHrvULp39YtWLD/GKv3twzxvPJ49M8LaIcKw4fAsCp
y/GN9R53ztLVb3u4nnfrIgRC32OAqnd6/J0ZZ19aLJVW0/OwUpFsBS+norxD/PqrH4UKcaCFIaul
KixEY+nQGeqEjYCW31p+xUL85dq6LFRo8IaAQ3cTImklCU6YKTYEs92uNiOPpBxCnoCLHR99NH9X
83Er7hVcacQFDA2Etkbmt1FeG8f1EyNt13GoeecQqXJoMG7wA0+cw91GNhnq3+qap/01XAC+qO3b
MCsUWp0kkDV6O7q0yLLQaWcDFlIiou3eNroizSyjJpUd1XajblYalaz5mS+tV5GEBVleUC5jGGHp
dEr2j2Gc4yV1TywTavMNiRfr3GrU19XxSq7HYg25yR++c53YvTyLnCAh+31977yQDzLNZ+B+dCk7
Bq7I2GQDbeM+FkkUosDjqTHxqbvqG9N7mBBSAe0r3UCjV/a5A33CJ/eT6CDjwd6ZU8wLrs7A7jtm
MS56kfdtdGLgSaBdAnJq0/H78vmGnuQTvt2O3cB8BmmjbKg6Mjbf5M9gBIV0tMwCz4iLScb7CyvG
avFYNhnU418WBqyaRUC2ZiQaG5LUbGVNWTU21MA+M96IeKZKf+wAg9/gRgdo4FLjxUkXTM+mx6JO
+OmqfpOI1dTbxKBxHiAknc0o2x219G2JT+TjiRT4RPhHrtVv3p2kWVIRkgx7ETrmIOq7pvtDZUpT
0iNIAo81xmhRR6peAP6nBxoftT4qkXFd6Th4UJLmO53qbNJfc4otkpe3Il97HONd+ZFCUZ7xZxOV
uIOeM4h1NTKRK3IMOpNWUdcUv1bER0qGl6/VSNYkpFGNfFZZup8k2wCcbpc807TvTU+AZ3DA3DVx
J2ajbwRbxYyDyO0tmCNk6I4uyhMpqkr6GK27Ae+HjN1wXvv1T7MaCOfyTrAZKW1yLClE7oX9WoC7
MflWzHSafd9Oix7u6DqTBLm+YYQS6rpydPQJmqHmQisLFJ4uKR+ePzyYXbib+QQrVP/p9n9mQJod
ekVBJaKDrrwvT4WYGRGBtHrgowqkQpLVOw3gXEeU0dRfVeKPaTDJOVzzCI/G0rL9/LG2dKbda5bW
qYgJ66k7GW2NUviTE8J2rJSWyNHscH4sIf3c7RpIDI4pf3inlD3gmsnI17p0dxOWuTHLbx8rAenT
XnqED4ICYj+eu797gIccJK0rGvQNeQa070yltKUpGc190lJQslgFt49iIew2lDdV79pxvK6VL7YF
JV6nRuqLZZ8PBE/KZtnH3VchqWZ+WciNQ8SjmWZaxiwGWkjJPWMBG4+wSVnu2chl6RNKuRUO+xOX
VADjwJj1nOOrwC49Aol6/98cZqg0yaq9mYvfuh3aG27ER5sAfjInkxDPaxGnMUKH4cB/d33L57/t
mbea6T2hnpF7L5TaK/IpDB5bHefubfseHTZBV+a8E0ekT0oEIFsiyXvUAmQaha0m+VO/IY3TPlUK
kLh13tUfXjbK1t03l+KhgPuaqwYyPj2tNo9526a3gH5+Odg14UvQUhW9QumNx/Ykp4n6K2ek3M2S
GYx88hR1YWvErZzVBJ1NgPserSuJTsKeFk5QBNcr0JJNkUJf0q1v1tuddaRr0fp/9KA6rDAlgF4O
61fi9mX9ZpDZYx3EAftfebV4P6PK//g30Br+WzNVsEr+GLYOwT3rWHaqFv9q6ol1w9t4lHIrC3DE
W0kEtrfCxkSPyR3++nP7/+pdqUNxtKer0O2i8rZ9ToCNgnzxQoCr7aPGNuaGaKRLEaadPjjipRSW
Km8dJN0N41rD86wSjz/mx4RVBS/ZIaLmgaiE65QoiOg4Ekr1Ic1r3IvBBcCsn8YJ9V/d9XpungS4
uTN2aaHGou7HTFFS5Ydt19N1YIMrRDJrAnL8hwEv1MF+ss3/WUTtBBXAX9Ev5CR1M3cotGwSGH3a
ous8dKft1BHTtU9D5dw44eytEGZXOIxbgvLxb1hp/2EPk9X0RzEL/Ug9A/C0WcfJ7yeV93ge8Y3W
+FejGcynQA/7aIJJjI3prXYBdQ0g/zXXG4hkadsz2GODX5CctxzG5AWwL9BUaMSZzKm8TrMgMGZD
LshtIzDfWDnvZcEK1nvJq1LxmwLhwPfT8x2OP8MGW/iKynnU1kA2AjEt80DXxQL/63XNOLBtlkBa
2SExZe69/3azSyOtUJre1RxRopX4aeuj3KwxRRMI4xvalQXdKproSeX49r1S8jcXI9EXsVDNMIXB
sBLDOI3bkTl1TZe64/w70TePIK5gh8uUihzNiQYdT4aAtkRtxGB7BVTq7xSy5sPw+WwrE2HOrKde
Bf3+CvCPANiNxIf+YKW4G/Yc3uK19mrRwXNgzZltYZQBqUsQUbSJ7+paLBjuO8I4csp6MlifVT0A
Bxn3h9DZppotfcaM7Zy/6JiGkYQOQ6OipLFiT1wmHQs6PxmRypRvZmUFbCkcmKaEXQC/xh6zV9Nt
vfTdo8azMHFUSWnKKNRLvPBKgoURAFq3L3Nl3QaxX9NapvuPm0M2ZvjSpskqHCAjljUurqPC2pt0
0L2W9vLK+4q5XInfiAJxSmRDbZmVPExldDjcpjUYbftX+if9H/uO/IyWRaey0D7tVmjzvSuhXWoO
EIgg860zajGxMX30Adj64EVmR/6/AXM42ZNARJttHRHarHbTovmu6i5gtUBnTZncsEA6I0fe0ueI
5hbcQMdDdkYoEaJPK/6dhoP2nGWPgfIUaNFmdWhMYcDrfcRdPtfpI2f4ltKNVgbmW1qfJ2e0HXlE
w17whYsNxkmgUAMgiDznLub6PasGTp0s+SH43ccPZDWBJ8kdZVWrC+DMqSvn6gBS+AN4ZkBPR5KY
T4Ry67tn42cLWVD1eGLU1D0tA8qGB7S/IFExnZkhibWkclyYr69lwPig15w3TVUHAugIxYpiUUrL
21E06pSszIZpOkRK7R/g0EPuk9Bp23beru4fa6njTLaRDSA6bBEAoQNX91v0GJGHIwZukvxLxbsE
muWn9neO1miUWCiO5MgIhJfnjhvdULxQYFi9h7FzN51vk1I/UBEaZqi8FXMjqK/AngOh9zIqgSSe
QjRNot/k5JGd/tQZHcvtdwsob5aQ8DIICDfMu7SRHHPcgtypjuup9c15wzIQfQJut8YkWZkIl3h/
Nvigjn/b/qT2cQVk7cZae2rRoNJD7lXOIygTmZnnONJY21DWWjCeEHJE3rUgw8hc2hsO4HqxJZbX
Fo4bAXrd5xMJwqVB002mYok6puynI73mZb8tt36S7070vlA3yYCk18MXY7jUcc9Ve1CAsWPSkSfx
kWaecZfSnB5vVNjRRMfaw6Vn+tnoNII258NxxaPrf4r/0IiNoXwtGUqHMO5CYpSvdVkLquHda0Bt
AjSvgDkUg2REqvNfBKGu0CSRqSVtb9Ef/H11yEvVLTXafzLRekVqwaeUnJtdv0OHCtyVHPIao5jg
x0Obk/OXofndf0l5DybHH+NSyuB8LAXL70eXjH4+dMLvXPGR1I8FcZmkTfqSNc7lx0GzMB7MXe7J
klcBPTtxMHST6cfR2m6aoVuI26GQ0ukzN1N/1ye/611BecZON2NBX1HoUIBjB0lgOWCXjTSl+eLZ
HQYhpTlcUZy3VfY33GqT/7nZ+XyQOvMxUCanNft4ouSrZ1DJYyueiZUR3mV6A30rd6iVOIZcOCOI
CpRPFid6e7kbqitUxrbjsGJMPaeNCf8WqhFAbia4UhQxcYKF6ittIuuv64udFyQen5pzM8pHTurg
YI/jvOE3rCvqNi7qVweTRf9RMDHqFuBaNazAZ1ETDK5h/nXaIB5Y63TKwkKuovVBoEMXAW1UCxHs
nIfVjtxGv8IO1q77frFzigZnnrADJwIuAfhqScNthi+/8DKetghy3kchO0SN9GscK+LxSq3Onca0
M+fEvcESkBjpJboWIKpF86rrC0iGllCZKbGRZf7xJShKj+waGQbIJfAUWo4rluZ+OAlHWvebW0TY
ZeRzn0f0t/hfNugfftbuXX/47aVwQXlDvShVgq39Ek0FRliUv+yiuybnLOwyizWLFUyUxQbpSQl3
U+YtQY8TdqdMV+Q7JEakAwT2CQQ2jii35LvgQAzjQEexrPiuHM8diclGgZBDMamQ2WDdcU9jO+R/
ntKl0ovWAlqh3zjsohLPvTiZ8h0/Metd723jHfxAPM+uJLYPncO+3e59ibMMsqPTIsbtSabdE7He
YLZJVyXUxewkZEgDQTippmJUNfaTkhSfMCmg0/mrFABSIJhjthSq4skbYIPXkuQ8Pcnl2QttQtYG
empnPL6Qz228mqjunWNg67RZBw1BStlzSNIdLL+Yxco4weorIa0CMbIXI7jccOFFxVRDnKT26xuX
zp4rP0sFiuTwT6Qbn01245D8wt0FebN53VJ4YAqmH46TctcExYghXJcXE3tz1Q2LgDC9NCZILTu2
fDpWFe/DykTp8B2A5DYY+bjGs7vIu2LMcHEBPSUtVctgRk0lqBJQtDYwlyoO6z/a4EyCbUOJ0o+5
l1dyrAGB1UvT9ofxggFvhzvVJ2JoPmdoyfqYajrl7P6kyjtKN/mti/+W7OfaY8I/EgS+bd8L0Tif
nFz01Mj/O/pmIxL+tqOdT8BOz4MkfynZJrWM416wMrHIlhqMYmvqJiZjvwyS0ZNyS7yNxnizCow0
PaHr8NKqCuPLS9+3pyr70+Rko7vuYlibHWfT/3yD8UyNgnhoH/Ra27G9tLIWz/tZMaLVsb3uYsP5
0MyOLqHdfESuC/KhUBRJfhCeC0EhSsqyEEXB+iT9FEfubuGhhU0ejnIDoteg1KiaNAfk3dwyUaI+
ayIoTxD1nWouw1rNwt6nqXBzA9oeDPr/ocHe7341WbqQPPfBE5ILtFpdeT+dkNx2q+3yysFtyl6W
mHSOmjHP+r0iNOjRvny5WIbn+CkqokayjHDw9DiC5XLrxFIqJPk51zQCzpR9+6B/vCW+EB/kg6Qu
qYnPKTKafYk4XV1bTRcNC/SFIcdZfnNoYzRL+BT6GS7hRpb+3k1o3wUGA39raSI9KUW/IVALM5wd
1C0snYfBk3NQpB6zj0oeMyPIEy8uy8GuCky3f4ux1l+TnxtPMgR8xk0UvKb4+6MzKYXG9vpdeczn
2A1+y6kD/hbn57sMD4TK4YmZnvD4kOIaQhoqQac0EwhsgTDRf6sNySS/M3CyADRlH7Rlts++JvSJ
Sqk28RoDQYpzYirkpYaU3pXvPyOQ+ke2UupE2ioe4s2QL0NlrIjc+ZdB/Xq6UgZTPKvbJDJlZFtK
MQuFVNy4IL9mrMAM6lbkyypcJSb1lR92MAb+dTEzyHb53rqoWWnRLrDGnfGJGEPx0ZOj7mbqY/K0
Gw6UOz6CuJC3tjiIwvalyhY7gUyKai3HK8Y4Gn5moTxrQ8/MmgSiHk9IMQVOG8D4W1WYCkDA6oOc
L70pgJFjcmU9VJcmdxyBmyoGRHdTscvLYCSCBlcP2lTCsnnyXCGxvugajMFKAofNTnrdZs5gp5FX
3JzT/0Tyb3OuRL8HjU8F3AUW+HgjJS4Jq7JmNxFlKM9XKL52nMx5g5WwZeit+z+2xEuFEz7vwBty
zbzexTqZSOIROwAHqfxtLtwMr371yTthEae7Lf8zW91yYNSrqqD9oCVKthh5w/ecEgAQhCy6iHgv
nuQyBnZ9g9g+9DWuxbd7gpNZVxcGmPkEsDC2dBBnPMUFgMo3FQkXzCbXTXKtiY8hULUcia5Xdy6p
BTA1l+GVGMdXLYNXjX+XcSqkScU0vy42m3QNbOGi2LTr+KuQAslRGH1mLGpsj4YP6cW5oMg4H7FK
FD+hqZJogBhroEl0Ht/hTPByShRgrFjgHJXKoqXtdorXEtZpZRtFxrndqfb+HQNwGYPeeCvdZP6b
UfuuP3s03JwzpDqjMz70QS3RnlqvEbu39uxDTq23GrMGKFDWPi+UBngmCHjdERsd14e8UptBRGNW
YJYgzFMQGWeLu4m8k8X3v9xEUjiX4Qdd4H+ko44BjMincCE55ii0ZshZt+g/JV30k62mSkgcgCqV
GJaIBq0bDXZE7wG84hWKNiI8ZvMOBqZQErUEeIIz+MdWFEvp+qZdxvnWlZ8+uJwTZMB8YM+X7DLo
r0zwSuFL+nasrnQY7xzo/YqOtsj5QfVJk4NXmzMZgS5jjo2uMYofPvQC5xMGMqqoQItVBGs070LX
eNKDKDqhCLnFS4kHmEp4o8KrBVTuf5UmtA7xQtg3Esm9ub7atTssz9Xc5y1iverbcbiIiSdgHFha
ZhBx2toMBGlcXN1FlhtaYVDzOYmHeMkbI8K5BvPY4OGCesbVfoS3kMxweIdGD1vfI4RhHiixI9I7
2KbZjZYqqzlYA92reU2SSDeLZvRGEG1MkAXUDwSpPsofcs2uF4jxz0ykai9ZM0czugFwWXi8/nBu
fhm22sBk6vbPQFQfoAZho+vAYyAliBBp3zcH1Rb3rivjp5eZ6B0NOVBmayOXy4ye8mMiWw5KYqU8
o7lZgXQejQSyxy2YpF8qrxI85pSS9d3ZcpJf1atSa/QAfhb6oUSLfoz3Dmg8c9HtIg1e/udDWxi9
czwnLUnUtxtlgMmbIgs63kIdVOm488aNepiYulFGZ64uU1gPsY7/M8ydkoEv1NBnvOT+QujKPt87
iUkMEJTp7jx/dux2hPuKBA8t5OpMXBkfsaQ92RqVzbbBIsFzwtio2laWBf1ORae7k1u1Qig3ek7e
4vV4hv18Jrk7f0dipp5R7Wh/ttw0mhbSuWWFRnluu91RbpModNgRQi6Y9P3r3f90SOl7uaWQpGJo
joQJXMMlThGhwqCfqYU2YSUlQ+Wja4No1+HWbCz/RKFVFTkge2KA3NZdXjSJR3Ze0sYyHPRj/mEU
4pCvLFHcJSivf7LU0ftMC4Gin51LlnnjSa4qgGODv7xZYvSirEA9xZYR27xur16wl1Eb3Ic+OsKL
rHg9+u0rvrjFNtMFRVmmvkINmj1Bg+uXAOISOv5+VCar2gl9tbJVce06r4a33kBGtGDwy+y/OjI9
IvieLnZcahn78Txvs3DScfWNzpWNE8Kn6MrNWxbzFeSa1LVRsDl38SBLU09YOFs2/5xS27GWODIC
gPfvgm7z6YIL+anCcXThZ0xS3MmWJObDijhcRAoejaYc19RD3oPQTcP2sodScUG/X2jz8kFTbsOE
2iat+LRjU3CZ4g+gRWw/PvD2zJ8HDI7+yFVzGGFG6nAXL65eQfX+x8IJ8IVCq43F7tbwEgeeil67
AsqMRaULXqIZ/yQaWhWZwCKL+aNoF9DrOCiD9Iyx6Ffr/KPTinASDNq4fLXVAyIS6WoDN0LvMkpw
a2EIho6C8dT3uiirY/PNQUVUEQsqPWjhMZIXQ36/gR2pvAVBszuiDguYMsaOuWuWRjR9w+139vYI
vqA60gF4INa6fk/uvb5Ty8f6sRMhr+TWRNDD+JshYE5qc22tjwnwQxVAOVlyYl0yinnPjSeLO/U7
1d/1FkBPJREez3VdhnjpzJ3Y0oF/qxcOfbrm7BaG1fta2Q58oUh/v6kCe8OJWkFw0pWYSmhUaVGd
QNiNVQrjrgLy9Yin0wRcq9QNPK8oHqAjvS34T4Ui8zNDHHJcTS8Qte+nkKLTmC5CMYTGSPIUrrEb
CsAuHppT5NUzHUlTM9ylicl18LbnfCeRkOw0sYzwL13iQdjjZ5+JGn8MeBpd2yySR/psRfePop+n
AS8lhkyfhe3nnVMaM4hCxIzOBUnZhiUntvUfNtFm5cpUmkL0aKNmX9vi5YgFvWBOC61kSZEQ8nwO
LqdEDZ5k2b5bEKKstHhWQPaa8/ZG1s9CNX/Jv7ndB7vFq3tsXXtwkcVmAgX8jWoceZfYq5MCgtxN
1f8klwc5oT7MwPF+pE2HaRujFs02b5xPFRYDZelVfU68ve8MUHt8cKER+j2GSNgz2FRxyLv45fQT
BIyjme+qLdt5F0apZ24KsJvtQmK6ub9KV5lDlCtW3BM3H+kKckmt6f5LbdSC7OATyMNkYcijQ0KT
HRcZzJ1WuBOTZ8syrIQagvhIj85lZAm3y3S4oKTRSj8/QyDJmI8oVP4a2ptrwDBG9GjsEvpi7xc7
8oKzHTFZWu13DpS7l4Gce31inh7n934dAnuReG82Wz/jOVyfBQSuz8o84rRIUu8RVXbbKbuG+UKM
Kb02W3suZ9PSjvtxCMp278gRhFYdsXmgBMO8PfPyMeVL6RGZ8xRuQYJn0pp+7bV180i3xNDLOg66
JHXfg49ujEt8JE0n7k9gr8Red1NDbhHOj7EAwG8gmIK4B1beUucg911Kn43XCs1YU2kfBRIXgZ0N
0vV5KKeDUX+76vLHZfJxwbqDr68duQB3zzjwocq2dtgBsUuzV2b+iFxiibdJXf+fSjsezO0a4Tdk
PzNyIpX0NJc9sGfdea5+RYIpvZAdsC6rt8ztKs6daMTwfaYME4Bxb9uOfyotTlw1hU2it7U/OVBQ
6QL/6VPwzEppBXL3K/yBQwlks8oA6YyfMmklOQ6pYAECW14CPNh7Vc2Ngfr6WMdVh1UEEuTb4nVR
l+hp+kXBcplWN2s30C6pIc7S3PqpiUOhaoRbBJ8k3nwBXwicxljeav1g/hsBqMqQGL8poycn8qm/
cAPAf8x/v4tZeg0si+DilIK3sg2YN8iIW8tx6RX8HgAjfqn4WU6HbLgIZj9us+5Z+CnJ0/6A+P/I
+vzo4VqZyAyU8YSI1l0A08nptYJfBLLl/oRL8NlQFAPngvKLaUXAjA8jXdo3GRj0pnLird2D3wFw
cBaZF8LuHADJpteIFwH6xH81DCReasffhtvZLUz8gK/k9bD4m9mnvfIZ2ZMmqdGXIxbQ0ESdhZjp
KivV6pph1ere+fwlqqweiP/kfqPXdpabCLzmJuuilZ9tSncxUrTRuafPq45b9Adzqb7LebdHlvbR
8ELAoe63bexCNMA8h43BkSxo6Gypw7ZWJnx8r08Wnpr1ZMlyN7uNmBWUbyeafdKt/s2D1bexwu2V
JXX9dK3zanFadPYe2RLA9pXacnrDOKm512dZqog9e/1a0w9wh1nKX5Jk4oNONadVAgyhAeWF9/yv
/rjXFWfrQMVa0WQcCbipRvucF54U5PnEYEFeGrMJFeDuG1mEzy1VUV9Jki1d04IV3Pcj/kKSsxZA
GpO3hxYvp9TVhNbhyRy0Z/zreBUvI1znwlNvb92gmj/bPTZe+HaAsMurOAwpUJq2IY1GG6fuuB8L
46Rh2ID8TClbzNxqXtcfXtjWROxe4nV2e2UoQMO105u1g6RFgqq5G+328d7733eqQOyclMRRE8W1
7OgFBq75S1G+ACXzd646IUFhWni0LW2jMlDtGG4QUW4pkBb56g8fx+N+oSS3fVSC2roVZNYWTUKU
cVXsRGupBiCOMujC1yfsTU7Ssp7YK56JkoQ17qB5zzdeWBBmX/Wsm8+syLue/KqnkmFYX2P8VSMa
cLceqwrv3hn9TDZ2A6csJPJPNJak3wICfiXhplN1mqYH+MTssqWN9hry/S4XGN7EhA+d+fVNu539
r4stfw0R/JfF2zHn/+RrQ2tl+3j+YmAtdDWz453CvTYteHszRCDJKHph/gM4M/ZCIFaCv8Zw3zze
Y/acxCALm2bFY3m6F8aXxg8ZfG1uW2JlLteqF08zYcCxa4uNZAPgT8ETjUnn9sngzKBUrShsKXy5
9srz7qsKpWM2Cj/FZndY6sWWuV55tigC97evrjpaobI6YE8e4WNeuvKZt9YwUAeQWJfNxXDjVH8H
ck/tbgJ6kPVB+BKhblsiIjh7H34TCB5I1sAOVkyerIJRnXYCwfpiHvKZHQ0/JfMKjycau/zU4s1m
IWf77WqLx86uX1DRisOFxG4W1VFmt2T1rifWn8klGrKuoLENiku7nm6Qw8xmJvaWZp+3c7L1CbEd
0TJ0/n/BVWtWkeWVx2g3EQrUAAl6jF9gZedfyqRvT4q11DgNBBmYe2FM4/AEhvGG61838fNx72Vo
FpfRD7qOdu6Uopp+JK13pBns415DWOSj2aHa+J9zCfhrw+FvgN2U8qoAFJEviO8Uo1g4NOJew4cp
oC2l87sZY7oWXOUS4OQsXO3MdePfbiJe9vnCEQS3McPeDQRNY2QA0fZE+eYgwgR3zUR4N3qKd/H1
YTYZRtVRhW/exVKEWLOLZHGA5pdMcCKukoYqvMNsBBAuhLzYUzdy5s9ZkZ6hRKOwZUgbOyOjHPB8
pT5aS5hZRpZxnurpMUJiWHfdasIvIqdOpa56AzLCTBSrzo8TL38Hl8Z0R/6hHan5xt9ViPLYdtI1
U8FmeiOG1BLTs0YMsVKRKC8JAW+4CCIPhVgcR4ugRlLLjFuualh6Oz2VdlKzS1Syu5jsJe7eaxoZ
JbXrhpYVsEpIfaZyhBf4olBfKXepaBQN5CA6QWp99zr15MESRjN7BG99jxLum8fPU/dP2GyL0Zaf
P/57j5TFCJU4Q9oI9pw462KM90xNZjYIUWhDNGQo9Tq0bdptIgGJBiGJlVWEjEIveRFslvLwF3d1
Tb7Eea7Ykwukm4EC6Gs4tz4q24h/CjjSqI0BK3RPfEjyPYqkxoUcSL6BfXrF/LdgysERUlr/gFiL
SRCQCGwMH+fvJ+5SJnzfoI+Gt40EyWJKvpYoeQwwTzq3lG+70QSoDu4xm4x5bYZMg1F8Wz5LzElS
/G9Pd8+9uqhV9RFsXsEq3rBqDZ4kV1EM7uAWTpgN6CzdeGrrGOC+rTRuBAQmCoFgzZzxrIiClldz
AAUeDR3ldKVLTPizcktY64cSFDQZYvYZ4z08oAur0fXYbPcATMpY8+G2xhZ9H1cTtg35j+693fSb
9BKPdxfVH8wLHPEtFT1uqzy531D1eIHce0bhLXEsEXAEJxh0cBbaYvL6WQJCOpYFsGAmy+p3PUqY
Uo1S7IbMzKs/hhA74xAMe76g3tRcstzPoN63YXDWlLUVffKsJDB1PPWxMsoEivGBjSKs8s7pNOIc
DnX1xxYTdKk1Tx2vxBrb+QLOxsUs3h93rsXxOYT07VzA6X7ZIUNhH+eIJIKKiixHiVv5tP/3N8QM
gNPJ1U/ELjh6d7zx1Sz2S4e4qBXmG6RzSjecSsCjyccymGGBQQ3oAX+SBLjQbZt9qfQJNebCClYj
uOrGVpIzCOpdqOfC8ZQh6ysA9HlhEZu4kXfmbXXpuy91/0duZ8+iuON/VM7/YiXkOLL2WXxUuIN0
N5/KPBoTHKKoi/9zYsEkeoC+htCZyQx4sG1Y9kYIZjLJeFSIcQFgo+KDuRuYA7/tuMLbhDiTO8UW
QGl9xNo9LKyFUCl7/4z5houZArINH7OyFWsRAabwQloHf3SrsLBfQbesOQjomTKbrLMF10Y3jArG
bBKzp38Fm6ySdV08hODQ0XWwf2ywGjRrd6mMfaIglc31hAYf4ntJyiQUqfWZwhT+q8m8IZBq0eme
Yr3TABFMr6jH+QQJgLNIZnYwOg4n/8YG72J4aHpnQoXLVaw5YtkcAyPH4My9j4/fMYyHC7weutnl
iSNbeO5LKCh5o7ubZzy6BgoUE1LWEinvtve9isnP4h0Nq1p6/9JShXm9ng2OeOBnayjzraHyfffb
P0H+lZ8fpsSuqmZlyMBxUGiQ/W7oS7GQwmWnT8eN6VPBnLP5eXe6NkURTFZTm+0e/qL3oQXoRJGY
VsNMPtlZnbCghqQPvNsLRbfLVEcnAnsyy7GzH4+z55FKF+TFo3LQd4oQYuGDhpQkWBNXdAkiGZWt
67HADQZqfhSx+/lxY2ikOKzJRjHTbcrHmH2/Vx0YrkiDBICmjBNcKOpNjEEmIQ56mca2EpZG4GQK
y/EGuyOppfXJU2Ge56u1Qe1P88/X0UdEXNlKnjD5SH/+6mSDQXTRnNx83eTlpahfDl+Cm2pxd0g2
syTMIJXeP7qTZdgZDa1la1x7fpNzbwiZPGmfq/Duq7XchnqIq3AA5z+Z8y/rrDTQjNzwso0MKfcv
b5GBdT16A9latx/pirVmHwb/Ood8aOeRUBcpWMl3nmsaaYE+84nRDBE1mggUs+pHWzClYn7XBtUi
M0ui+BOEVpLQpYUoMVidLMsnyPIbuYIh1PfRxhrQ3sHrZAMM1Zmi8bo4u3lvYJZD3NOghryB5Kvq
0sQh7s0zTn8g7l8S3Y3WAh6N8EFTYEvMbQMw/0Yit9kep+4adhSMsz6e+H6pYpkjk1foqaRv9EEn
uASce2xtaBnhvD6S53T1z2s39V9918K8sa1BirCLN5NfAJW9KW/cv2dew9y2B/fKOBOTX2jfdAhW
OMdOmfEe0jNvPMaJIr9t7c+ZZH1tm64EcnK71EuVAe9RZwU+Cc+oGWW/hEZxmK0667l2f8K3Y7m0
iPGv9NRkV/3bvytOJAlcv8wpLg5ulR+VQkjOcE2LHjGaWAMZpCmwPVcsAE4ztuZmtsuTgzvYJmg8
BxuRgn9J8udPZBCkahRhu2CwjxkYyBoE/x5LzGhdTcY4BXGnoWaBlQkCj3dGsIneHrtLW9L2WcsK
bnhLr022zMcXWNViQaGxVCbRazAPIz338kBhsodBogTG40G9U11gKLroiqXXc+0Oy3xy0gTAjBBb
E5FAK41JvuDxfYkDFaPn+dQjGRXIhC7I15QhJZvarK/QNeWfYqFTi3i2Pexh0aknTa/WMe1erdew
aNs3cUYPOaKzt2pPy38+KczitOiDUJwTY0qZfOIbo0y3RHlbAQKyhfOivveq5ZN19ObaS3d8ejoa
nToc6GTZKQ4QWyQK1cnY+trZcETeqeBEOHSrJBAclZTZBgaLRNaGNWRUs5oP4Okm8tdnpj9Ij8H7
lIyOdnfeCg/oElwj1z2/JggWOt3rkq1EDZ9lshATebUObhrMo5JHz9mS4Y4cq9l+S4fPmTuHESB2
SYhX/LATs3h7XQW+zzo5RAKyW99DbLPCO7ltn4sNg4WLf8ljNY5FAyrCIcUju4cN19OmnEkAhis6
uQOEsVjppGRY5boLs0l/vmRyh4R/ymo6Vem8uYuJZJRx8RhOHMgH39TT6DEfSc+jraZiOfvNNb1R
Z6MG41l54KV0MaqLsk1FdWHKH+5d3+T+/SOESJa/po82uj0tCWT+gh2FW399Q4kPKXzqbzI44hts
jSo+sSHEEMQLEQRF+gk8XfgAXbANt4v8lt/nlJyrkp7NT0j6wNBuySfRB7X22DQCHxykroQoeIJC
bRhe41e14wqkzg8kO4qaTj7zqqq+u7PJg3JyofkCCSLSwuIVlr4m8NvQ/cw2g4hbdSePhgzTsbO4
GUUweobfvF25VtQi/uBMhqH/tp3VxOsbDtQFPjo+9SDYGQ8sVLVhdujti0itfydDvSGwjChD5lNU
a6CHIICJu0CerrlawbUMfKx47lGdqS8DKKJ8WaXNouZnNFknU0Lwz/pkdylFvDk+3CZ4QlA9vLwU
kxsW2sxl95THF7j6BOjx3Al7YLkOEg7Ba8oZpipwIqDPHREXnVtM1zUlPZA3YeEYYNhIyYjpb8rf
jQSwgcpDKp5GRu71vILpriXjE2qbO5LL+OjSXSDj33pl/mMJ2iHCoVnRKn0DQyjsxUxmi5bUtvys
s/gC7oAByMa4yYBhLuac7z1I+0mExyFPRatbS44bYlU9ytU9UkhjFQeiqLp2QI+DwT3aP3RYWRSW
FT0pr5LacmNMpLIE5a4+JcAb4Tgc9eSo7P1bi2YgMZh+1Ues9S8b3gjNbETWuDFOk3gvqNKn8JFd
gK+PbBQgbPQWz+eB7xOv9S0hEZk6//HuUj7NqQjRuXCS6I9dd9sPmlc/Fim0ueokua8zgTI/Ca2T
JVp/t7Fzan/ULZJ0hPimD7HJO2x/syEBrIU05pyP2/l2WHS5iXXid+bH7aS9/s2+Tv7LGizfZtAC
BRNXntYQ0f6ZH0oQk9hHp7cCT8J5iQyShb7F5pePX3L2vUFP0/A3jDl8AWu0i6BAnyw0JHmnyAJJ
a54rzTjVIQy5qIydyVQtPvSFf21RmVACTuL9LJpdkWnztoe2gj6VgUvHqsfkeI1IuLbodyH3/PER
EpOybSzNWIdXU0+K4pt8jTkokWbspEPQNIh6DlLpydHxc3RM4GI5egIhiQeadfaR6jp6WmDyevs2
q8HS+J0FfDU7W/8xC0aVUKBmDiE+YYOfev7+Emrl9kMft4qSRvEk4ZLHtzfJMJLzeojBopPvG+1i
NiiW/Px2v013HpzHZoEG1MUvjZDV831uObRxbbNYKoigECYu8c9MiHaXbmQ42vBgVU3ZzQ6TNmDF
zPczfNBN5bTOo77hMoKKwBjmFJVyYAQTxQ4JPWvVaOD3FWxeQ0iLeOogSl1eAo1k5otIxkuvBoZq
M2dpgsOoKsCj3zYK5aDr9XXu7VQeO9v6Rwa3UjWiI/u1DA9tSKDuxmzqo1TMw55GPr8psKvR3VNA
gHBMLKwdYVtiwz0QaL7qqbKdBTi7qaRaubt03GhjOmyYOg8zqugw30ziYPCnQxt/pDfuDX3f6hrN
O9U0RelaZKq5eJJKbnEl0qSNJ5lTgMjQAYxCsWWx6DNlY4onOYL0islU9fjIukrmC+byYQvn2jFo
GqNmY4awyjZmEkujx352yTnUNub2/olPF2mO5UuDMZtHKsvJ4YESYpXB5SNfzDROt3Pjj8tp2A+F
Wm9vywo8WmfzGQ9TOsKZfuHlD4ciGYoeyeFQJ4HKu/AkVmBA2qbCr7Uxg0L7o+tDnUjrqkVzUfdl
Ob396ioqMmsRiDZffgo6WEhOkOfYV1cElxtprqzd1er0XMVV9XYVZSIh+XZTG5bLS6QTICJoTG3e
mXko3XewbsYyV4y/wBVYfejBqALKIbSOKPd/J4JUYnSSPAZvXuhfYWYf7hdCxtM55ms/9BKltUhi
FDg0igmMdTGj5+o7SqE+dbZPoaxn9ZrXt9r3jPXITLIO3bU/0FCf9Jz+EFqiiTQYM2xbzwin9gXK
0IpwuRlO2CjTxKLAsKYMOjPZ7OpKOGBz8ybhVtEWrnAEvGtyijHKRS/FbvaMI8qP33AZnosXQhX+
PcX8AhLb/Lccnx/OfoXtmZMfTFBq9vjIQ4zks8zb+5zknO+Op6nf2++kLTsRe7u4TfvCA+t6t+6P
2bKV90TlyhYJOAWvmITDUIufpFu0a6DGjfrslyQYmQHmeQMQYEMc8AN3xQMviyLuule1yBQ/Stmo
WBpxf2FvlBc4WdMGnOeyYWU8401dnDu0dYChbz3DJf28RBKPU0F0t6vZew7VYpHZ6fSYWBXM2G06
ZsqcrRAHZnfw1uajdIIwBm6ZXB+0NIhivZppeFIQrSnQnIvd0zLW4BVw8WQc37HHmIrSrPbtNi7w
zJ8tTvaBGNNzw0yEVkvCKEF9c9vsy8VgCyyJWqLft4Jt314TFmW1ks9c+k0UApjTKsxRiIKZUzAz
l3NJdnrZL44YkPbLmjvlh4RP2ZxkftY2MydumLDsX08ZLX9cHBFzHsmR2MjIrP0yJpxBL05djYtc
SgKkSHbiCpPGYRbSzI3q0f+vvkk+p2RwTN6q6luZg0AFdoa3XLoXPD2D9fMH0dQkbchWZWLOlO9g
l3B1IOFfu4R4jCTuD8LlWlZVOmzktyGtmXtfgZ9M5r72XnicrAfwgGmaWTOUByj8LUxlBuPloLg2
RLLm+Mgbsmbd2BpftJ3I3MpD8SkiSNEc+k8xorXmqityWLezV5hpA1CZ1/GdxC6nkDNwT8ChXABv
3jt+f5CO1qFXf9Mez/t9z/8hW4wQN82/bFBPBwy8Taqe9Tg1mdrTnYakIQvNm8hXqWivrwu0rs0V
0d/u5BdJ3LtPIK4SeCT4qdE1lrxMfcIreSL0KKqrC1R1sJ6bo4TH8Ni1aycXyge4AhE2cdrFP702
32YU2SutxYeoEzD3MrNfOhixDM9e2YHQ2R6olPzupCSE1axhX2X3uDUbyicCOdbjRBRiOzf5eSS6
/KAIJXOf7wSPiRtIDMYFKlrnp+Qd5UvrRNPji9zmrI0OQHV9jgUN9xNpVLhQg+SzdssAy0P3w6N4
x0b/7+4dHvIJqDRW6xv7zxqzT/XldhHHMVOGbmDe922TPKLtYp766vchKgZJKcemh8so/gEl0r2j
fku6xbWeYdpDxR8UyiTNLxYQkWrovK7B4xJpxSzTRZdF7OClyTvYwJr53a//BPYTCIaEkkE7U2x3
GmIy2QOgc5rfjh6CLLlLa2hL0U3e4wsgSszrNoz9z5sevftNtRr4ggIBdMYqstg+UpDhdMDcKa4A
uNcnSy8A0EWqwW5qLJN6E8BSo82CM3gNEqsg/4zgAchxcXh/LCxSZq8X9hInCWhyADpzfuhVTb8y
wTiz0+tkFIsVPgC3lb70nGJnE3ES6cq/Up9rM4tTOs9lQdx9zjaW20Gp9fGUwRVY4I2xWQLbIoUZ
VmvSsqw4X4B5PuONbOyljw8QW5waHMyU1tOHdOXvaqziir5HDv5N9YHDMidorqFp8cH+M7MpWJyh
ViTj8G5TzDnj55ookv05lzSfgPhR+ApPec61v3J2cc8KnNqSC5zTvYMvjAEcbP96SlkF92sjxSy2
CyyMLg4ilVfO5z60Cx+XPYflrX9rVr56d7r7RILieXR1vQ2U53TH17xZI5JfU2WUNnDqRpinCqEM
hJHMBNZ0MKuVVWlO/Bp+4RYKludypG82qN2r52+6ob7JQ9+3eA1nRyHCTC+VNZGtlB+RrqIGzOcv
hW/MY1ZBBDwQLY0vXkch/UCLHRI61LZvbUaSkreyVoS3UVQI9M4j7+LeuSFCOasTg6M0Op3QevfH
vQGNzAmy9mFsQ/71TxPGd9ze2Cb7hg4Rm8U1xdWvbUaoLokPtfe8vo6A9cVC3HbliKTRJb1ff3pC
xo0WkTfJyQEp7L113ongGMpfFCrAuSyTTArk9TfDran3OX6+5F8zyFepzHBJOXnqyshX6vf761PO
S/OUcWdl554UTMMG3hpjo62okAITm3mNZSWaysqkSnvNF9zJd3jB1SgOLWIog8mPqYfXmLIVX4o8
0PT3pmIdG1aWaNkjoEvzS65hEX9DndHEfxeMUa5aaoXV+yg4apAq87cv9mEhuvmN9+1FnzZdCQMw
epp7JfUNwyaBpXiMA5kwR1aVgDxJw+uBz4CX7DDg+ufJlqteayAA7Fs4L76AfNCt/bm8hvQ8SLpk
Ewd3Do7g6wgirBX3lTwD9IM4QvwBu598wMR9f6gRPzHYWAFwWnHPsZAY7HPMUanWAnTjGkdIljA5
uASk3NXzeEV8l3w21/ao6Yf+HZzm0G3TkXQ03pwREVr/DC9z4gJDlHmc822N9nfkcECHCCjRwyGF
UB8qt4v2wbT5G8lmc2fpcLJVyvsxxk4hEYG0ZtCf1M0OI+itdz/Mb6vn3miyLeC86O+XbPTlun8g
WC7wg7/x9uKEmQZ4reqOmVXJGE7KGRrCnYKDsYafXZimU0p5FQ65Lz+k8kxtf8mJqWBr/xFvGp5Q
aQ2otomUmTIUxybeuKHp9BHJC93qMr3Mtc6VJY3EDXWC07bhnivrBEaTaJJQbF2Q4SRCFPLEWne8
DNwV7mFFGM92IrSGJ4y5zumrf1bjcCZ47NAYyI/wUG3QyCX0YnXB9JCt0fhk8jENtVsV3xfmkcrn
xaESBiAAIBzbnUf7NTgFN0MNTyd0Fl/bGngr6U1H2Js8+vshvKnUCSNtrvyprDJ7dYHBa4txfuhP
IvtDlkWmzvaDfcr5c/9GNWjtT+REVtS6AnqODBhVJac7l5Ze74/qxfSxU54iY/sc2oJtHMJ+lwQp
JXP8irsKzNyt2A1xIO+B3J1xTbcx4QnM2nlhTRzz+AIkVuWfTb5/6pZ7xseU1pSZypoEPETfMvih
ph5kYrszXL/xMFTcTEgpYtUoodaMeGYDlcsUj+Nlh6BM1oEWoUqyKd0Dixc7C4u3sEMErMX8qSnU
2MGAXOdBJPTJsqkisFIR8uyODZzslInYAi5su2CQtP/ZzDlLhD4ak4uHwDsY7KjcUsgAwo2bJglG
FYAMl5oNIuh2lwjcgbmgavoyS/MQ3i6/Lg/70CkNqASTV016K3Tz7PTulGfhWWmCYR2BNzzfzsOJ
r55Uu74vTXbDiQo5KaI+dlu55IgK6nidKYL6jzjDut8BeGgHAZzX9CiRHLySPqRz+cFD+A+LPhdU
uIkcU4m78ACswUKFJn15j1fc2PRayh5foe8wX/dv7xY4vcI2Ss3vJOqlV9n/GpDVLjdSV05Sc3w8
lT9M/SefCgcD1FWGA6C29fPfQghasGhD6mv3FT4ozaBCV4cYa+uwWiW+w+5btcCcSj2rIkYQXXfz
EM4Wp4PopJbZhR/JryADw+SIUAEDZiLYfw2LHmOQ8IT749aPyLQyuzA8aYvb0C84A46scqFIDvj1
1zmjXFRrYtQeWzEYQNQoZFTMeswtRw/nyOS8xvbwSL8knHglDBMZrxbwRVAp3g5lr4gfTchIS1m1
kEpvWtOQKvpezr0dqbWe0yZMUxoDN4hXCjQSVT4a9HBK8fAtwTGOsc67pQC0rQrs/rMq5Cuy6XVl
ab9Pj8CHlk+uzZBCLmOuCkyHWF7IrvzXEo1IHkqW5KrUq0wEMMe1gtn2BxXGiaDvLJhPwIh6hP/G
LDq+ZmsqB5FTHz3muIl+NmZ/k3zsDPcic1+xQbEQVo00Dhb9gcrPPk4bCV4EvsZZn8TZko4CPE7n
LCZuiLfopgRKAHvuwlEhNsdDnFvyu5ZA9YbZ/e9DIZGBDzIfNMOKj0SRrsXsjMeokRQQ0VfJhisl
rwPjZQlDI1GvPkcMr0CuR+51tyIscmxSMkkReZhZ0v0S7TxWe510KklLsCX8LuTa1ENvNNa1A1Kz
ry9T28kIaPPDHTTp6A50xmv0TQoDdEak0q9UPNiia7SKjSWsUlZV63Od12UG7C3pLY4OPWsrGEZs
bx3hhAEwrsq2cRG02HtVz0teS/WRNq3I6t2GKTfoLkKYBMVPv0kqK08eDVlQZuBOc3RbD5E9zIAW
Bc3odYaQYDVoxhLnI56adv+f4K3Q6R01UXRLlcXZqPMM9fzjmd4H8cEyBQ9N/v5J/JQrXvE3ByK5
pvGlpPo+taMsD5kVfu4Izk1mVvbqEEVP6whQTIYHQpiUgm5RP4eWJgk0IKxpvB8YiPA3JPU+Vjni
ly+ysn9LI8UAmIcI4c38NDuofGQlmWWcwDnh1zdFTHodlMSuM3DAV3Kv9XJq/skDYMUMzdkJEcTE
7zPHHCXAkjpJG9b9QpBPD4n3LCOF5louF+p518k5qj7jFBQj9pEK3nkwl2wyhTp18XmVQkS3VMWb
fj+rVK0SbBJets6q9oTfYjCRfSOoft6clB9ay/S5sguD2dDiQ9tj2fOcBwkXVqWgU5RpnC0yHAIz
CCgyo0J/Pn7+Z9qzOGWo6xF8GtHA9JwpOzQFnCMepxtV9oMcp/7y1DW1g7F7Y/gTegkCBsegqfpL
0G87RflMNvy8h44kOMYCg7k6pyk94fw8m5jgsHOrgvGvwRvlul40FPnICEG4sqi7k9UZveoZ0eTE
1Es4i/srywXzSOUw853APEL2Va59Ox1w+IkGWZHXTtnY8n5eKyusnSmrcKr3L+6veszYignNk0sL
Hfxcl3ALuz2KiiYJhMzevsuy/uHeZH4ZYXyZtOIv/G2FmtnUwkxzi8wNEwT3e5mh7jnr9JqxQUR6
jdYTZs638IbF2KMkqFB5OKNV8kmss2CQ98wU/ajVk7b3BOKHAPsLMPeQyvY4R/pBpAZepFLGYI7M
5R8qFRkhzBPU743P+vpOdPD4dJO54uPJ5dynQAiQWJg5g2O6PvPjR+bhSsqz7jSJwOXrF3bzhWk2
wW3dWtNlbO7fAK0HmaULoTmfHYHuxHbt9kjJ9wtc+T1SJs9ywdrp7Pk2xc+LeDa1Su97+xCEsSbt
rFJD8AoH8f1aak9/vuLW3yIhYVjtgFvIo0LakMj2zgQ7oNfiQYZYrhVEMLiTHan/5j3fgdav7di+
fdBH2HZjVpVWspnjqG43aai4oFhdOp4mLaJpc0967PYHRtxYGpcUw4abqN+K4BiBOQUeTywMaTBd
E/3T7E1TgobDYfNwOG85UMOgYe0HG2yE0Wntz0O7SlT47Z+H5leyI5lleXbq+Ype/5Bvmn9Zhz1p
cuAIet98YwWG6FocaPWi4dKwtm8DWeNp3Hv4LPlmSWbFywzKjHrt3YCZEVeTc2+RZqnx5i1wBNQS
lxS06RaYlyvXWemAMQx0TQ3tMH36fAaIYPBkMZtgSlylJrYuGwwvaEDQCucGkK7bE0l4x32c9i+s
ljFHfgYg2RnwGMdewlBvB6H94V8ONo9lGdr6Zrr4x0p9JVcAt/rBrURuEQ4mVNLzXX9i3yhaAuLV
MxKtSVV3SFmOQqBGlCVCYMbnMjQfLFjNeUNdJTbz2K5JIgHiNbJMOJMYbIRqEecuFSE2croDJt2+
E8LzREC/JmFvxycHbejKHkk0Hjtfx6ByYuQLDlDqNt3DvOzqfwNDu/7h3gf+cN7r+9UHMpMzeCqe
0HdR/8lE2JiSg9pZj83SYziD+oRJxOPoiYcQ/I2snkSmP57EfFjDmlHd3QntiX72I6NwNjnZYrsc
KNXsf6Nyw+OHG5u8hX3NbMuuwKqHTmMkaPxL8AWumBX+qWI4oDTEJPRU1B77rsXhG2xJk84fG8DK
DeZZO4hupTGn2/i4Ptqu2DKqAH70IF8sDF0Nh65bespk75EiZcraf0YNOJ0+n9szzyIASv9xe806
e7kmhlpbhQRnZ67Tl3GMVN9BjFFSVNFHzJYyhhDlUQQuM/CwGpulXkb5+238uQI3daErIxAIU1/5
RC9L7MPEP0SNQ2hPxrJbVQoIhUEdOYYS+ovGuMF4WOHGdwvasywt0k7WfGcDtyFIv2AR6JhMNU7c
A32VfCxTJtW0sWf5uazLBrOuRQxar+Uf70YHW8awtIx0m+D2dYzcGsrS5z+pbzaA8tY6xVPlwAVp
S+tYaXmYUhQj7uLnGLIKclvioUjOY+TMd/rs4upaut/AoLsiHEszR+CoCa3RXKqeb48qfSbFZMNs
Gz1YyO6wica05DNjOeLZHrpIQ9wSyG7uK/i7TzDpJ4FylAsxtbjHA0/MRUkx6oZzgmbdX8f2QaBc
JT0jd7+4veRC7TDO4SrNn8Qgq5te70R4DP/SX9JerEylAat9x+KociReWF9Z47cqHWQ9zpSZeuba
62U+lg7UruiQZgVRuyd+uKNFuokptlE44s3V/kCgbpNPo4ay3vZ4J20WIQi+tGMjY/nWeBQ8oIxA
TSRB43aimkAh1LTUB7LUbWKzmZQ/QrMQyxjzfbAZtYqJ9UiUiPiXyDFHWpuhVG0YiYNgNi67drPl
NlNwC+MPRnVma5MQaQ/6ia7o64oh4aG6fl1xp0mqkXrUYiXgSU2jkivmsYgWrfro0NQBcV9oWyOu
ALcQWaM0llOiM719etQ46wXN5gmjgQY4lE15t4vKKI+omU6Q/XVVodF9/SCO0KuCgQ//dqqlhY0W
mlijmCQZ/dGQzOBGQhzzi8BgXWIunff6PSfKewKoQvbEUWV21wq+fBj5d5cSTQJ9gXVjcfxbTFjX
3Scv7MQ2qcVBQUhGZwFj6joP3Mh4u7VjQXD9pBwvy5gmAegZqe7RqfjRlluZngwcxIzYYhbqgInD
hm4fSWXDrW2kFZzfC3UFAdJjulcU3XDarR4TVvVz03dks7g3vOoDoGsn0+/n6mu5UTu+GJsvlYdx
9veKOBqdgvPHxmtbfNuB2fRtRcCy0olVb5GYAcb9jr1SeHUuV1TTm6WcEhdV3POl0foF/PVjyDTY
pfOvy+DYwJUFnfB6r7e40JvvzupMnzu4T2AaQQQ12d5/ltAPcbQNBg4dwuNXS5g0Zv2DDA1W44Ht
QbfVLOpKMfpZtouZWS0HKa45NAkTI7aSBK1nBbHvHWGDYHmRL6YGn9WfjwMKUKMlb0sX5efOjoty
ZiClUSTZVpM9uqUg5IHSG3F4JLfJkiQ7Nnq9ljDv9n7HVvIBE5s8S6yI9GHaz8RMctF2iohlW6hN
MK/5GmIvKjACCM/hRLZoYB3HO8G13HFW3KbtYgcNez+I609dRMv6Lm2Yc0mn7SKoPL0tTdjjF4wu
XhuAswLLd8+Nhg/TSvX9LDoBCwIxpRF5+cTqIa9Fae4K2LzvnYv3q4wP/VkMk4NRGRJ9mBxCksju
jT1mguvlPQrATZBm8Kl9eQZxbb9krimZrdj9Npx+I+DRSEJRGp04y5Li+K9dDm0X74qyekhSCZ7m
w+IygaQGK+LVSnyDJjCZN3XWBPD2gdOkkVvjsZ92NAlOu1y2an5+RsCsTQ0UUTMVLPu9wEiBZDWN
m4ohKqvAMU0M2a1oThlePochUrABgqdsfXKnwER0hxJ6HwRnp7L1zeVaKejB3ao05G3X/rHGXe0E
JCgVK2JOqPdQWUPHJ33SsQoPoRdwoMYHVtlXy+6/dNna+YnMMcMZl1qEmxQxDs9LI6QKoxa4zZEY
9fhlfakxssJ+wtlbkzXILJslJj5QkdTetUzyEePerbpDPL1Im5uLtnL34h0X5H9XNFbfVAcmzPNn
3UD6X5o/NpWjCTK9mqrrezZiSQdCbJK7XR28WJuoKEe1Yiw9jPurNtJAthYuSbX5M8GljrQegpr6
BP6ABcS5I/QMWgOgYDUUvVfaOf6yLK2+8pz56VAAuwyDpMyUKU9/u6+BXXnuq+zxQi5EDhPP5BOi
Olw2gyTKp+/D78jIiWSWmuqwr9JQwOkBj70QWOXDy3LKSCVrKxzk6Quie5odyG9S1A/QjBRKETA/
YAt83wlNTDVei7CLSeon7Y/cao93SwsKwuKg6i3vodIZAviyPSgAM07gBxnntonixZ3CdfhoOJKS
WDQQSZfi64VnkiTAwYdMs8TfA3PtbJ2ue+Vu1RfKpSrDrdz7OuRzqS+s7/E6ocN9zd8S0T0PfXHp
58TcoDTEWihA0jOW7Ndw0bBiQi/GlUQjIFe9kfChiYBuULXjQzRNfToW0PrANvxMPvFEuxXhCy5s
0ZRn/vAxhhO694bg03wvhz24K1xjqia4pAADyYSU/+mxl4rgd4blaATuRdC1Vd9bqrwbbna/vboT
mPkhXp3a80jqZmihCVMk+UUzvzpvZk7jceKCA0ivowWVXZfV6Akvlz0nGEEr/rpO8yms7GO/1/DE
DgdfmJuM9tsUl+oKuYUytiWYz7ktSUha6UaZMZxJPnPTPLQ3NPnpDlPhgEZ2j35EQ3btMXZuCYdF
jWSesEZB+J54+RLxWOS6qYCuKatshHflOG23Js/At9shQ3vw3ZQV/cOlUMbVDKYw9+9hs0FrNO8p
s+nYRMy72Ml/uVA8bejOKEAhjE8I8gHIZshG9hTtwtsm4cxr1wWTzDURORLDv/uUNY0Z0sbjBzY2
Aq46qC3GQMb9AYvvxYD/8mjF1L4sV9Jmyjuc18cMY919CRMmVXw9CPRbeOSlX91AGcm2bSVj+jkD
VIWde43E7MH6WjNcQf5+69r45xhxM7GDimuhRAzcd/0EVf+hItqFt9co+ztLmpjm9W0OB8ho+uzr
FgB0/OofMC7AHMJjmYc1Pcz28uwLl7fkUq4459AAp+WfiTPocalJAnlGrf1nU95RKOLYHFfLVBKR
M27P2ereNc+TR4Eg1AOtr3dBoB4OjOsQNIpHXxMLFytCuBoIuIqfxvFHfQ2QWQjvOrtUHtINQzPb
N9XRPwxPW7n4y3s0vccEG0EdolP2P8kAZXybq8kw2VsyFKR9hzId8QA39Tq4EXpgQjtGm2jd4Tl5
a5hJ39Ww70imGDbWFFBqWiBFSHkVGimNFmZa1qwLN29Nu57Ycjct8VD4k0NqN2HMcFZkDPzWslb7
STz1vpPWEjs6lADx0Usw2Z0ja2rfAUQWN3OZf2Lebd4QTLEdxpQ0VBKVB7ZTZL/6vn8heMwitWMw
Yly6/5WtjzRhMDp/0AA2qjxtxoXI5hlEp/UiIg6JuRSrqYf4XDeLGVfKAMDr1NJR2OJQvY0a4Zc0
Fj3SRfIywVjbQtxmJO2wvyNSibPiBBfkTZr0rMsk+UXaKLts7Ife+YfvEbCeSk7xz0pZKD7CF251
Owwy+TFI+OBNrU6XNZhX3KhkrMELFYb1E84VHCYu+obiFa1kyNrkyFRs4juiU0jMaxzwuRUunU8V
S7euesq/8MwgTz5i3PmrAKISixuqHiiWsJ0AexhKe5bji0+eEmie01UI15me3kbmm+KAKi5xxGZW
vZAlzXBwUpNcnQb4esxB615s8c528Pfk6aXh6t6Jg7WJ3vMtOhlAHHWEFyIcqfsvL50SA13elSID
i9tE9lPl/DjVx5qrz7AQPEaqftIJxMFhgHVcRiEa9sx1TAGO6NlPw55wsx1yq7NG8WA+OzrllQxs
TpvSnrUg8MK1+KfRAPk39Fef+rJTe5uYbtnMR1ZuiFsmQuCE3TThr6feswJ7uj8wE+Lr9CLObS83
oTwv03eF+jGwk7eJpZgshTSEFgrVOwYpTAs7anoR3/ilAXYF8v2WNh9BAflboLOK/fu79wc2QBx2
5Nvoy2owlQPBL1pww/Pcyl0Pm01YOyYblwNKjjdKYJKNpDR+6QQeyZxVNWWZtEmH3dPXzHwAU3s7
uAKrVxf2IOx34Mo2jF9yFUmRPsjMt9C+hUnQMcptFcsLKYmtaaZpzVXrI+dNB4uBhXm4SuORNcg7
xKiaXCxU7GOS1SUqxDg/usrhvPhLoJFPQPCKxY1tR7WAAhDRoumCaJTk0B6Lu0w2TYPMA/sOE5tk
O6TJPq8cLzpHeOcPURC9anojOmHk1vcM8s2WtXMOwy128ST8h1L+4XComYOzxa+Z2FLaO+e5PaT6
F69AqFboZms41YsSJ4sxjsVxetttrBZbBIEpArRnIIeobJHPZz7+qetG1tZTlqFRtUU+VJREMWEa
e+ptI6zekCHY/wLe37BRG2K/jSk1m9rKeW6x+LvQvGHz7UxeHfByOgLNEalidKxWPFwQe49OhH8q
qlLbBJ01JsrIagwk3u3cRtY7rJZnBO0EQ62RfgiOy2ubJEqSB5xU2ILZ71guWroVuFKc0sdk3Xqi
LNcc08fGvmspLzv8uq5E/28joTPuW9a5c0ZFBnUZWJjGy1SxhbTOVnKwOuvAvoz6kJaI4jj7yKw+
Xvdh84/EY8w+C6DhJOaru6Y/o9kZznpnlq34RPZIvJJhFM9RE3XbfrMspZrZzhz/xgG0lIxFVqXW
BR2eZghRtxVzjXifbnieeZGDxjGoGnersgM9VB/0KjTf4/lICTm69Pg1s+bcBhfb/HmPqJ88gP8D
lbeIq3qYhqObFTi3OHdIyxnmKZH9RlVfILBc8SARvWguDXmnCikC3VKX+f93Raqf6B1NV0/PsG11
wCs0UW1YSahzAsKGqCQttQh/fsLRVtUZaGPOxZ44gG16IQVq+RZJ3FrkKBvU3p824jwHfCgmOmcE
fMrKi37sFchg7fxZTCX3pDqojTetVm2BecHaN+6OwDI0mfMxQ1Ur9JD1E8z+N5FaSg4NsPHE5SVj
baSp4mI8gllLwX38+sIq/eYQR+RN6q+D38YDSSVgCAeYZ50UTg3/Q+U8UTSnROy0iKrhAVfDcseu
KUdwlmPxc/6o+VUw3BBdMoSPskQm7QmP9IPPbKGVLAc8zx/7dXKogBK+0jZgHnP7BPZen/nGL1wW
YvX8efmjR9VZUKI4qNf7LSppsEkFuJ9SsAYOKCVJZAqQUadYWGF4h35nwUZTXw++Td0MhoDE0z7K
6fmIlfrTqlHDI/t77rISPUjXqH3rwIJU6rYxIlhrLjn1Sq1t0RiVuRAlfZQO3noqJar0qgMg5nm1
w/goeXdKEKfb4pFknFv/FI2sRA5R0rMTLfQ4Eo0j3eB53TAGv8LD6un5lp3m7xT3gBfx2lqW9a0k
o7J5Z/8819fxdpHGnl1UQAyw4RIQlNuaZya43JTuW5woRNY+r/fyBSvkemCCaZIyRooTFf8Km26+
81USXYl5AZbqRPVX7hNBhfYjtvjlzgKOYXCCgVwq9fQdfo73VQPreItTU+k3NpLyJqu1WKMbfMwY
IKJZgGIzcCm1fjJ1s8TizS4R02JebZkCZOWHzVPD1yMOp9+oQBHwktTMonVP/6NQMaJWnnEWoxc6
Cnum28l2q/cP+CGVMUrmptKXHmsRmFJNZAclP+MSq28jh6tQcSFaLN8pckpzh5vzSK+MH+bDqpV0
Tgg8zN5chd9UbI4/O0Odr/3FUB7/ulxGJVUoFKb++sCSx3OXtVTPZcN8U1OdfnSg5BJ1DHqA3DCa
eVZgTHpCyQicRsGXlRb2IYergM3n2ycsw2176Xx/xyqhhVMrsIR1ZlPYuvkMVaVbsNgGMvhv28ii
HuLN2oIzlbFJyo31G+N7NUyVVRCRlEw5e2jTT+AnWnl8iKuaJqpGS+sQEDi1g8SkadQRWgMt8P8y
5qw3ZOQEOB/e98NKAeKFwBMCNkUI+5XpxcbXCLA7126lOIjvW3ahVLYXwD6sQFG2NGZYI0qWr+nc
Hhp/VDdKf47PV6LUac+cJyUdJJT49oXY+K7HNe5FRPgVZQEU1I/fc4KjT2+w87neljbVxC/SYKde
/VtWZUt//Adg7MDQ/ON0sJ/b46kr+I/86ZUqIOPzmCYuZzUs5BbcZ++Kl4pyu3BCawjMlQtFKt5Z
Nn73dSwj7ugfKuu8l2AvLJ8iU22WFRWHz+hHZNjyC3U+lIFqdiDjLSO7OMaiyW7Vigi7tflSM77q
zltsiqxpw6ryZoaLF9rxOdnf8w1GVZX6Yadz2kNVJsWiYkioD7hYSBK6dzQPllmC83AAY+kofgoS
d21+hxjYVFZBR83HDaR6SaXdiNxzTiU52DRX9GaxT+OBkEgT5rQ+1cB7QbTx+/tdfzr3WoHoxNzb
M6xKnZ7Ku26PO3+Ux8H+Y3QUFkY3U3iH317y2yFKd3/BD2up4gZt8EfBsK1F8e1yEtrPRCXWMuXq
ObJnMWSTOeUlycxHK7F7AJbzHL89tQxt0KjaNr/SX+i3Y5TrVNNgpAKr84eY1VWsZsTln/TB98As
Y8WsPqNMqRFlsjPWigDh8Z8lo8rBpDIofKan/u2xL9GSIhYFYs7RHdDCAnG328uj3JjJI7byXtvB
eE2msCSv5tSdkvU+DGV/Vb62vZ4c2dkHaPLMdHhUzSLPlCw+oBWrPXmCH1Cj9yGplPUnPSnkZXBp
pJzbYIj3snXOPquLiekNI4GBtowDnpusAov9c5P0WfB5Z09wwBdMxGLGrbhkFR3tvhAGz2ldaDjG
zFJ4AgkNg7u0wqpMz5532TlMxpE4BEP+leW5LV9AEqDITqQYE8GBiMj/HycZ5+ZusE4RWgBWweaI
jR1V3cVZNrx8v5qao1miesm1fjj2uHp0URGr0cSaZyw8tN9PtVR/WbH7TnI83SsooxwJ95M/5VgB
MsmqOTxUQBHj5cbgDRh3TdB+ufJAuFwYTsytqaZnUg139jf29fnG6dKRA23xBQVcJBya76m+Lfnb
uBSqfBJTkRYMD/9+5sWt7l56/+H5J2jRqP+dXnavV+4pD00jw34l5qNgxVtSHukF7jJW75rvCk/S
dejATpCK5rbBjFtL/q4026I6LhBcmgiOdSISLe+Ga40Nwd6Wm6hIg7iDxCwygOg6hu4+J5Eag5/r
zPxWt5ckCiVijgYXiRFP2mZcj7apb0lViwgSrmqnnNvJSI9IYhUTRUxUxa8hr3QZQ1vYS+bkz7ug
/9QbSftSog/S9wPDMsTpvLdqdHsJAw6+GvI1KaPk1bAY4jKaQ3oecVE4Ic/buH/aoLP0FAvkBT0N
xUf1YnPI/rxO/hs7bG1nAdKsZCJ3w2Cco6FZkxkyA7kR1dXU9esD0r7LiAqT557Iwq3ZMLAgcAFB
lmOkb5SRAXDBJMQfIt3n2SLFLA2+l8Ydp39X88aeYsKtrGoX1hMRfibLj2f6I6L6DvcGBCagZ9v1
D30zhmZyBAhJKvsnfGGhH7t9cTMj5imtkzn4g747nLpTUegZ0LxgcaPqBtnh5iCIvwFTYHzeMiVT
8+JxRu4kgaFVoM9JmcEefXCI9JNoQG9JFEMrYxIPEd1XoAFKfSVYlQuh7vrnfmVEcaRG+HXPxAnQ
vszORzEIsqE7CF0QPXfPwJuTnfdBDrL2XCjZUZcYfHeE6eTQZTIGS6s8L6uTKFQKM1cU4brXZLF5
MER4gB/0WdVQcb4LZvxtxJ9/PmlPdmEbqzYWNhPIqNrvv4E6hv0QX9Ki8yceGCV5uswR91+pN/eC
iiSkNhnrYxkzQrpICR2/EthSCaoBzwzXbPuT7EpFvsHh5WQlxpvZTpwCj3WIjAT8us2d853qcu7G
MnP8kXsAA/jz+Gyq+wc/yLU6tXO648xCSQWa1PJBaLC4lrWk12Ol+jMoI3UQFdMEvXdg5jdh/FTE
cKfoohf/PppfMnqO75vTrGFkhKVMKyG9Yxn2ghcWfBMgxtAnm3ZrIou8R1+Bnk593aL5X13ikvAv
1rcWKccTJyVh6Udi1pPKVyfFm+0bixvDleyd7sOysOhKlkqHxvFj+ubuLMEbc9XVRO6QFjqI/Yfz
qOq5XRvCySljSN2yYV8vVG4l6qcLuzYgERPGctG1P9aj6UBud9KzMrOBPs1ZyqTgQlm3JKp3gha2
vrqaG8/8/fKQJJhsbKUsn10lD46/rLP0+JdSWY1LSFz7PA4wIJjbgmiVNIos1YyxoTjtj71EOxKp
45OiZyWrNoclZ2h4VfaN5xSxXVnpVqrrpT2NgGY9irlwFcIU5DLW1VDTIgZw3l/ebJ/FgZMRalAK
jIjLQMi0lX5QVoN7bmArrWKuj74ecxjuJh72wkYlRIEOISKsKBpoXcT6M0Y7ZSD05ImQFzO+YGEu
VQZyUM23NC6PpMYQR+WwXhCPnRdVA6mXJFCRDhcsg5Ns9ZzlJl5VGpBsLeW8FP/mNHJW7BigQluF
t4iigjOlJxGTTeBO+Oi6FOB4G7Xi5R/6qVVUC6CttqNZGY0TjmkvU9pvZC55bwCeohT8h+9E5NTL
lA8YxKOz219Sv35FqUl2UjK5KNI58sT+iJXiXyGaeYR/Ps0BfX+wto0YBnnPfGBcSH3uQQIJ5YZ3
zUhesUkTjOlS4ceknCWRvcTyi0aPaR2SGqHBPpjG9uo8e4bs9EtFS/Yuiws65nxK3lcqI8TurSsX
qgM6tgy6235xyutKbvnZTM7GxlX4tkGGsx8n/W/XGwLK96a6ilYY5ZEkPrvrjGDffHr0zP/Vjy6d
wuYX5O0Vs/o7Yfv/dN8Q/Cz5cRr87FF5G8hOzEDfwQAdrCnGgUMNaZxmnShHPzkZRjByYhWGlsiZ
eKo/smFbdjrXMchlqIrr5Jkw60aYuyZkro2uWy372NPg/Z6Z8fWG7Wtb7AC+EDFGFYwFl1Fcdpxg
a3LAuQeDpqFPsgv4tfooIs1H1HegmA119KUv9M/rIi62kwabHXPUyyP5ZubY4v5jw/qZR4orOUbe
y5Z3gnT/v2yXo8Rd9SZiFt6KKQGW5nsvSuoE3H0+tWmk+31SPfGWdL2tKlOJMQ6fW5af+7p6spAU
V2RlUcHqMQoN/XQMEe7MdZtb5/4sTynJVzdYL3Zbckivoi/rW8MNoXoEvyb8qit0Tz6jSJFc6tqF
BCMZQDFZmLrQspf4DKJCpZTuoYhboJ0INrxmGEnGit5oWLDdcel7Z39nz1kcdK0eLpblw5rPdCE+
OBqbdykao7PsT3rJwYrm+lHF2Z7h9v3QmxdJ+erXyiI61Cg7IDkxTIH3PrC9TSvrYy1a0swBlDpj
9O56C51Ioa6vmJX44E/issqY3xHiFBz0JCWPhz/CCwv/bmLvJ8FDbGxmQWUdpC16XUntj+naYWfn
JdjJ08eCzZWwkw5h+CkLtW1mmolS4hLEFg6wqYxe8aY4QyAQu5fWNmIAk84OxvVWbNond3W6GGXv
AdTN7Tcs2LnPhwYFhVBgmN6RXy1iwHLiHoyee7FG1ygI2Ykii1btDUnBAUT6nqqgJuSrjVOGVa+Y
CMZgQnW1Ysb8J1pnsZeu8dVjUuES78rF5E+xEHauGE8Z86dHobvX+CvFoDAY8huiht2ltb1Af/do
xj6P57BFBmIaJ16iLecQLwd/Mxo8d6uzm/msHVoMb4gysBLXJ4awh2IB07TNc8pgqipVa04RDIzR
yndWB//e8FbH17YptYB6AAfdYpsS10mxQAAG3pqvLmn9SB573mqm3xamTXa/MoOcjGlFL9yxciUV
vnJMYtdYQXOsqnF7gSSerT3Wf6fV37IBihQzNNAQXkqFbOAbzDRFhJa4FiKw+DkVz11GPQ765C2r
+1n39hVhpHbn00/bjG/7EzsDJ5lpwQHz+iUvyjhqHf+WjfU/H0UutNeVq2KiVxZnpttHIVCVWFix
9gZ91it4Ir8Hx8sr7r6Fm9TsVY0Zri7KrxkZngvfeZtnMJL0fzki/Er1nnJ4/SIRBOBM9Z6XUv8+
9HKHujG2lKY4ZAQa8CAkDpVng375YJJNGTAonfVp2B6IUGTjoqg443GH0fAcYEmwqbpNS5sClUBd
eUrxZal6p15QEX97Yk3y3mjNkxHRfx+EY+oxTrbeTYfvmakcCIKisgBQzlpS4u5jGxonE6hf3VeL
TGQqIL4R5b7a8P9t/n+rdYf+zVS5KvzyqNSQ/WQ9qSl+iaw6U5xd7lVih+L7mKZXBztj60ggIe70
83cDNCH9btK9N/m9f7Kx840heujDknzPKySaVu11KQ8jSh/3IBIQkdMbLpbkEDCDXr//S49b6zxt
uQEG4ou3UTNYLJ3u/khW2C5pW7UgcXpXLeGeyVXGttd+j8mo7eyi1MbN9CRtRA4qZ/A7HD0b6O5r
aBSONY4AOj1uAJuhu4HqriSrejcpeXXxnPRizhhwD7bR31jE4z0k64c5p0WTBaFSNVEmQ5EiqwaJ
JSqV5OgEETTL0qzBmk9SGhMxsh7UvZ56F+80KBUqPJn261aKzP+V56T5bqsACLc0hckjfVKQGk6q
08KB2T5rOB5U4OaoMOyxGjo6UvzuZLfp6N6HCXv88Fb9iAUL7MMJXenONVrMCBYofD6EHI+H1Kxs
SKEuI0jM43RbXa1nqzTVYrqmXIbFjxMrRsQjPuW3dEVnrZu48r4sFUnp1zJwMOyTaafkCcJIp63B
7k/iDCtGM25bsjFUt7yVeJI/X2T1BzL8WVBQTmij9ngJDg7viOSByWeCoVp67rov3VOsUvPpnFY9
64TwS059d+85SxOiILqvPukHJ+mK2lAPCmPmt02ZZ2EZyOPRxMZHklHqJiF0JcwiUC0KY/4AV+2+
O8oso+qdOyzavbWP9iJvf4AqXv42oQXBtW5AUWWIH2EHeY3mLW02ga9KIxq5OPDChhwX83oWpQGL
4Fj0f7O6s1GXCJeaNhMJrKkx6qOYKEg98lfMAwOUes2SsPjZSYwVNJInp0aDeeyu6XU6cdg5zchL
n4jzSkKxHsIqWkN24TjAKUNxp7leV29bkT47o+KcC+OXReztTnntdrq/8o6XDxZiMwwRxFNU+IiD
MtcoNbCFneMGizqLlf9RaBQtRJhjxoWf+XQrse76E0XNdzdzRCPz0PnrmqoDAcyaAiuhfgSckeoi
Oy/0PfZTyDLnrfxEnUn896pdAPNNRxVxE2u9fVrxYtpRnf4ZtQtSAODkdTnj+lo4wa72pmJ5WtoE
KBKM2P6dMnt1VIevlnVv1AqsaBo4x+G/guYMySiwOtwDdT2Qf9BdTwUG2u+SOou74N6d5SbYR3W4
pmcuTnS6BNFsyBQVJoL7AHWcSKU4GQcx728YZAYPvcYGJX+scpUb37cGeQD5CD48mwuHqZAAgOyw
OSdVpRwOr+DyUyVNEISEp3p7ONFl/xjeXNEkvd97mq8sGaj+dCQ9SaYKVDH781ow7sZOD91F/oj4
B+1Ybu5jU3xD8qh4RCBKV72rGUaxIiDAUO3tOq4+dYUWVht5vyUZ/94qnZV9iwP14z60z/UX2L5b
SS4Eb3YRB4xZQOZfFsLENU0qx6mVqs+Z1qPWfROwk7pgxDk6lyRTySNmBRPt04IfYbpxKhSpG6OR
4H7Fe7w8jHbU+iVqdM5HqSzYQtstWfcwGaQ2KUyq7y2mxIHrRqtKI4LLM3n1T3xGIZ2SmW7LwNGd
ZlvdIREgXBUMvIPx1CIjPMsaCox9Q5VYksYjSrxwmsYj4cbqQ+DPzTuN9358X1Ep474idij5LeVa
rwHoOiyyTX0dhopA1xcTIgvf7hz/q+IXpMNnmha2kKZO/A5aSTUra20CXC2GSXo3HGq5h0I5ph+3
K4carYwxek64b9chBucjvHmUSJazDk1tKUypJV4lezFvGchysow16AoD6NJmVKjUY6wwsy2NBLvj
PDDmuScib4e3H68wvgfeVQRZzVyTatlGn239r25m8YBg+TS0Tt1XqoIVII06qNyEpAJEUPWJiJl4
IrxDcsFa7CCu2J52DwB3r1q4J59n1XOxfMuTnG7qTCK0CDtwxfVaBEpIaDUC+avy4XS8ZvYDIsCg
djP8Nz3Ut9PyLbsALcfiX01YBT8dWieByS6vdezeQTGQqAzZYscSoiZXL6U2TmXWDebcI9lF34Hd
+hkofWPCll+Z3yxZ1TzFVDwQmRkT9g4y4oRDjLu+6FGjwIhsog0+ySkMzLVszE9sHHprcxII1KU0
jFoT+0vZk6nwIk9vzPGkWZ4Z9D0dgySoAtVPdPh6ye8OwreJcfxnZftyxksu39uuSMYmR/bSyMem
PV+/PQRJuqMAa4094S+w5G4Ip1Ztp68e4+lWtVTsl0+NmFw8wVdw6QieZQSnbx0+wLdSMGjFI24t
BEA63mN05enj6x2E7luft7MZcWz0ouvQoHc9FfQhg+r+xeMunRC36rYyUgrQaKO2HJtftLxiXajR
x8xXJTh+Fi/XZRTBL0fq5zrpNsl5HG7jxCew5hZCm5Z3lqFmJl97lblyxCF8Xt0r9HQxX/3LYBD/
yq8WwQ/ie0c85mOj4HFK/+DekPxdaBOGI5/8xMXguEcD0EwuCapHRtB7WJgvMwuar5XICxqebmwJ
FZyplPzU/d2npa0BMTzo8yskqj9SiICbpUKdIxwlBSk7YQYb0Zzllm0uNV2QLhW7opzv9+q9wO7Z
EEUFNCa2JtqfdGi8Vhxj1y5VDZi8XxgsMg9QPgq05YeWom8pGTnlScVOq/qki0vd/LfE2XQ8aNge
XV5wMneLLLUTPWjXuYkmJlTbWw4tMZVyVSnFoGQoP6o5BvGC9qPAmpuyqTgkgT51Q4km6YppluWg
wSXbF5ho0Li05LXaI3NaySs6eAWdhf0M146KVcLORlsF2kAh7xK4CfdZkXF+Wyhlw3p4P5URujey
96eCy3DN8xZK1RggIPMib7/Os90rFc00d4w6T3mkBuqjAF7134VNa7GyPrl0Ven5ygPfHvksMDHw
G57LPXP08a20HS9hNyuY85fNv+TUDXAX7pWHcRn+RHIWSmMaRcilpjWgF1fj/Qpw0oWK+IJ+EAWA
ST+YIwa2LP10ENiN6eV16ccx482XXTOdmZjywNwLPdaf7iJcCLJ44qOyAtgTQWHtp8Q6A4yIKDKo
QjR9XXolDSE+zmnJIs0XmWy7k04gwzzzQDeZEoA9ZBkWB4KGT918WirdDy2EHm7yPQQcfjoYqwUT
OoppE35DwY/xGB9wgZFBELWgdatuWHXYfVbl0ox7fZQtwdrDu1hu9CwOf4V2eUWkq2ukjWgwm6Zb
EptpeoXH8Wq2BLnepivrdMsCakMhC7H5qNlpXLz/nb511wkDIjw+CfI+c91Cx5q/yBFH5zu/kFAh
BKQPFxNFLl/IINPaJ0OETiCiqF18CB1Cd+Evvz/FxJw19k1Q8E6ZbvUOuzJhwAyETCWH3SgTLOte
zT2EgVPUotoRJPluR8PhCAM+eY4Xqwz/bPhRxdvk8mH7hCix58PwsNnzPsZfsFHm3NEZ4X7IVRLU
hDtzgJgO19NIiv6jejC0nuHTb3a7uiTovqOD64L8u8vrSMowZMWAafR7+94bEHGVenucBSvhR6LH
FFezf9JJpxY8Y09f+cnnV4FS41b3oOU8rHflkyMVv9ieo5JzFN5CmBiZrcjE9lTu+6gvkdbHWkFX
1A+rO6143Fg1CyAVDVAviaQAzX0Hc7OrPWf8exXWzp0zDNVpsA8oFoPP4CmzUYfUqwQYB95PXKhh
DUpQRdj8q2NO0k0KrOdtjWRWDoUFQqnaC/zbCHfe/wsFzlCN/sINtV5hiNIxGnWSqoNrdC8/Porv
zfx7pPWnbcnhvHEtHUPuYHwkM5YDbJfRVfg0gaQbiTN1n0yGLboSsrskPpQEnnANNN8qkMSGG0Ge
DoItj41ytaCsu6DxyrxvuumH6M/tmwQmYLvxGyzE4lDCvX6j8YUJze7A2R/Q1txaLDyH6Twmzlo4
icwXfSMz5kJGvvueSYzZWwhj+pJV3MYDM6QrwNkEmsgrWnLFq+1Q1qD6D9EFwuMuX7R6uwSbHsSI
hlc6Ve57yTef0g1k2I6J32FDEdFUOqF6pXSBLApoARFh7q/RfYq1+39/McOd1lyDCOJPsLheJQUU
7j508LWWNIWtbHwcF3uiAGzInNI50VAZg4vkvWgpub9CZnE2Dbd/Zf1KPX2J+0jGb9fcxODFvmeD
lx7jG9pthc8tqcs81mnIsdU+EWNl0ah38ZXEOXmHDi5kuYHlKhmBze5p29Y9DSD6UAL/pBrpApXe
BhY6KMAYL7bRZkdAcq5khxh6QHwp4aOXyFY2joGdNvS6Au8Pr/r+6N/8ZjQijHLwR2zCtSNFV+hj
eo9/2jlt1PBcPImn5Hqz1KUtblarLxHrlOZpDxev9CXvmUKRBqDhqNeKoi3pafLhLT0x6Oe6W9JM
kPV9K8npw3mdM0XdIoLr34WQ/UKrJQlbfC3R5Mi5ONyjhve3lgMfix1Tw0WaCrLWzZBMnv3umnXV
4nzjd416GzjildArS8RB+DBfFx3+z/iSDJSdyyTLOLgNHM1Yj8hyTFFxj+Ck+j7ep6+wuMPLPFpP
WtBz0N8oMi4rySVxq0U7/cuitJ+s3stJtSotbjdbUl/ZHcjDUV7jHdnZHqA/uJYE4Q2NCTaojsH2
9LQ9VA/wN3hr2vWRVmStdo9puKb6ezjlt14Lv76NSrSLZuP8XnFILfFXunl2uaEl0bvAGDMQrRBC
1uiUCxUyw/xdy3pf8S2Dhhh7GU2Ji3eUH1/3vedQ3N7F/wYcpCAZ/Vt3YShaFLRDWzOfuce10ZNP
G8HSkI1YDMGfKJmAP0XSlRou1z2lp1KMpL+qevSa4HlcO326gpvfi8zEv3f1ncLfloYFHEySlSke
z4JUKnhBd+PNdklzrNlU/4dcULzrFX756K+4B+tlYa0F9YlXw9c13SLn8R6Iyg9rj8YadVehOrtJ
ApG60COUx2DVCNuJiYIMZtbaftxrBLxELIiXec3b5eKgMyZpb5DAbV+9BiYI0jkh14VZVaCeNsvQ
3Xg17GDkBSIdnN1/+MX19/HBvfq0qQOeV5G9HFgJha/ecYkk7H4E6us0jsUaJ7TlCaEQvNG8nsbC
y0lgp0N26oWERDJzVOQpu7aErRCAL3rdmRpjWhzmRK4pwtFhlbXpD3E8TJ3gD7Fxmeu4/ZQjlwtJ
9PIx+vJ+dyKeAXIlVdWy2hXjbqY90K5FK6QK+X/uuvNaiE15i4/BzuiyojsT/M1wavyjUMZ3ATcd
covucAqB5EJ7bq3sEuDFWZk+2PZC5nfiaRK745QAn56aSa5hCQAOLMrICWBuZryVdPVW3Z0ZkUt+
WgL5LjAZBqR06qJXyebKIxirqMBfedx+QUx4ETt/ZfEh8lstfpihcX0GiYLCL2WRdBBAz0Y2CR4A
XY2lqI+7pH0TRaYtanb+jB0WRMIRQ+KhNT5cUTURYhGvAb5gRaJi40YC606KgTQuTi0dS6mWhijK
oOYGK1hCov8Z0x8tHGCPnXabeh45j6TQBQvYNLO4hybPQ99FKLR2XJXrpStORA/FJ+yz/NDf25MW
6yGPwEMl1o/TTmwCYcZso7ZTqX8cQN4L2wS+4bZoFw7fGQrx1N3Zx9RJioV3H3zuCbjGnA6jtudd
MGPooU/Gmj97twZ75q73aUD/wqORe0PWbHHAsQn+xFabQyJ9bkxrYrHPwGvXAXUF8tHhsOZnMSFO
+9jDIXjcnazYeDTlNPsf413a0jAn6OWkmesu2D+BX+f7KWOYmmFWNyIH7dykl9IACEkynFWkc23f
e28mLKeSZ2yKVdMMqKkBZBJQhDSIY97CO2OU7ggkyUjlwUuRJQp77+CwXzkV7acg9vick+3KefRI
qvfttCcQDS08+OjcCI9t2J8AyX/LlccAl3mHu1AFb8i0M5iG1kFLCv8lE71qEWsMcWTOv4plAn/H
5Ias/mk1rBWPuNRL3uzRx6RWCu4itVuX0vW1hgnzOb5I37OaDxaNak7nDBVcjKZdMtI6FwId0UIK
rbA7tT5dxZI3JUA1fyBlhZ6SBlW3GMk8qRrM4RO5EF/Rhn1g/aPaEqL5SSXkTfbcfAtLRN1vnD/U
Hvz6CU16yD6fwYTPbQMQJeTmgAL1I8n18VA7a4FrnEptbdsKezCbmL5XL2AI/EIsA5LI7QcQVsKU
30b6NwpxNGHlpgT57eNp3E/7soOgUMrDfp1cVHvabumT8+59IPGfckGZ1K60u221CS+0XxWq1nym
+tL+GXNWXzctAsYboW1gXITwnicCjHWk0ERlzuuH5NTCNyX4mF9ukSvriMNe/eAEafdptdJ2gGWr
aLkv2maMDZt6NMnfeDa+/mW/5MxwbccrMvC01u71xqIhX+oJQjPiM/x6yvy8YO6ziVTEI6ooCV6c
yTxXdNpIiLQolKdwY9ufzo2PFEauwwbGR52CCGijCLd89m9ppAKiZp4ubGu/AZrca0U5zdqSO6uE
e22dcigcua2dAr4fZcK7y/lSutZXz/JmREXBDUKge7vaRhNkDENhzIAuzodHpa+/NLa/lzuRdkpY
LjFPk8XHHtS0R7ktoic3Q08lLvB+N+ChpPOMWVfGThfyBkOF5QOuxsHBZRMTHzliIABeUelwattY
F981KvZNfsCjBLY2Ua2KQMo/vb8KnAjK4oO4EoNzSCbBWp7p03edefn2a8MSe9TgRRBbpzQQzElY
vJwDeoKe+ULUv+zqN9vUE8f2Q1rcw8jhzbUbkk5kT3JMWw6BsXaXrys4ew2oi/NgUkKt+UDX0TXJ
VcbY0Ro9N0UovHPWt0BIlKWLM08ujwX+4oXdZBm/7q55qZbnUOTe/sfS3rf1v3rjZDNLwBaJ1alg
KY1X/WjSJ7eBmkvjTgAsXADooey5AFTikG1ERQCssAL2ojAv72MyGBJSrUq3BJJiuRavBK1IttmQ
5byEc4bex4Bj/LEn8P6KS7blcYajRW5m9CapwCqEuV6xnjLRij37w7EErJgCyvJ19Xvy4lsNEWwH
2Y2nJce4f68UjMnm1hb6krOKcrYxFhwevLH3rON8Dz6dtP+i1TUAkavDCZozNbz2mi5EPVHGd5wW
nZsCPDIRl23GoPJQsannfXbedbk624FqHt85a0L/9OptDWPJvbaGKN0sEZbWPFargLWWl27rKPq9
r9klUD1dNDkEb7UdeLRidjlWbswGAfSvCtSB9XmbE4kLMW2MJRjiMIJ11piIRCtdg/qcN3UOfwVt
G3PIIUY1V5wo5nmcbv7cXW8I240+2dw+rtOKlFaNMmCPW3PTrrtDBl8qkNveQv6Ka25y2pZ617mJ
NGgQXIlMrW/QWcaJHJkfyE4o2fotL87rSUywYl+uE9L4stvNnIG2TpLf3tkzmL+kDySI+entNMTs
1HTu3hUupALwLeT1SNxPZmO2gZOnH65cWu+YzE93PvxswQSGy0BTlNtV4j5k4aefhVryXvpunzp0
PHYi4/1SDkDTikY3A11s0vbh2VZ8QLUDV9DRLwJLCw5wWa18PLguY/MpI3xjthJFIYOhq4fRFycN
kWA7WFz2Tfw/p0hAFaWOTZx1SQZTgEe9kjKJOByYiUmmcX5VjsefEFMZh2TeVp7byNA0TTQrQb4a
8Hrkn1WYLMy/6LvEx1B7M1xYdLbJ52kakRjhWuQByQ9CFzePcJYASKgo/Vbgas+srLZx9Rit/URF
vq8Pc4UAqSSepXNDRLnEELP0opsQsDJTafNjTIVfvjsuMxAupU/SAHuuJF3AhZ+U4j0r8UsI6gpQ
CrsWECnTxeuYGU7h5fNFKbCxLDyhpzpmQfanTSlwcU1n4sU5GG+zmIDuMYKZAbAzUaUs7Bg+Ml+h
Dgs20+3Lgn8H5UfnZHsd9OZFdjJYDwisCapx2peDwYi59YzJksCH8A2IO2GBbGngjGkRtUG/hYd3
zQxhCID6AJcyC4OkHEFamCoRMveIV3aOwlBW10uNxbPqdFh/j7TrAIzbvSSPH4jjTIxhyz2gb3WF
V24GNG/Q7nEOPiaHkHQn4yNbaT6LFVSB6IcA+F5tzbYJBPLr7hrvNiHYLoGRu0wddgV+m8hO1jIX
IMD8FUf5OFrlkYf6Jld83Smps57NKRYX2JjdCb/WYFgAM+RZDaGfhPCQ3nCfqjvL8IGrHz24H89q
Mwk8CjPEt2621cz+dI+DCFbYQnV0B0NhQpSAaSUDcWPETNcRzEeW5RtuRIQ+hPxNj3YVSC/4B7CY
eOM5btTpjxslQnkpoBy+5SH81KkIH9Cb98pqO3tYvCtBAD1EYjS7KqRErEchut0QjsMjwW+jTWsh
lQ4RoM0kpPoL2eZV+ggnSMmrOuhnHy3d4Si6NqqudRjDD3DxuJRCDQTFPxnDbvL51XfjSPn1SFsV
ExXlok/X6DERWDuFdt6gccYuWLtX00Qt6KsWH9n+mQT2k4sT3TWFwa70kTaJBsYt1lgJrnVkwuuB
dII6PK74q6BHrv0e0yvGZUfenys1vbgq0Il+3FsvNJOWp01BLF7kHrCTfq4sTLkuriqgrnDcS5Px
WneoeCtXjiEt5MRMk7/V2wuqAck086MHTb88kNW/t7sLDjfu078pvAcbmABjoYbXmbFEweLbcw+W
nHth2t5kCIMNN5Cij64G7gwBYlNpwsTu3YRg0QAvVU9a15FE8qfgPJaXB0+gxN8ago8zAsYT4LDg
oLLWqAbyjIK9WYmor2RdQfGncT1XbDY0s0o9Lx13GfGtoRExAy/YIapNx20HMNyf+GgfK3DWH7cA
ugZb5vz22xr4sLDuvvqO0mgf4Vcza+8nUfJ9x/1rf7WigerW9h1ZTkNcvU90o+wlNydNU5Uu4H6T
jwVM7rQmkt4JyBoDeqPr9ymjVNJV5/npjV4Ip0JOEBKcS+g9/BIeB6h0Gm7CWtCpSiUWQ1qZcL4M
65S9WVIkVttFSoIJbR93SY+p+0r5Zxk+RwEdyuLrmi7wc7Q3bLWGBCT7y1vxEb3mBFReEATLVS4l
+CqOFivIJkAris8zRCwGVqt8b+Vap+Rlg6j7bhTZZH37XW6aYwNey8TYxc74lpDQ8ON28lAzA2xI
Kb9dBPJy7j/7DSAbi9tCKq2StSjgX2eK9cleGxEbfbND0fIry/+vgOSUX6gbl3/j6VEcHepjbbN0
IaBENvVZJO1jIQDtwBv2xUEhth/QeEK8GK6DrKQL5PHPpMpLUGfSO8sfkfBd92Myfv2JZ2Jigw5X
4MnQMhmNh1xrvexm7T68SGKPxmj6ow3sZThqtucQVtQVWs06gLKGRIQYwpnOuqc30XsPePP9ia+Z
wYVAs9t9zMiF8SeoMAKhBGz7h42AQhwj/BF6E2xyHxsmE8CYsrEscj7KmbdQF+6Nwv+KuyFIbSsN
syQPE6B3zmdknkx5fJvYwXE2u+bzMPZsCWAz3VdDLBYNRON6tmuMs5hiH37CbyClXBg9mgPzWOCv
nf4ZbgsZVTXu8gCC6cx4oDLAIj8ErbGI2L6s2luo7fHO0C70Akowj1Sb4jIBtPL6T7l6Pna92anD
8OCBT/YIhAnRHPiWbUJe0N7upjgcrIX9C+hLtJ6I8wJxGPVbLtV3a4pueefmq2+pbKc0TidRVnQW
uk4j/h/BbmiXId8QvCVl0ajLwamgXUF35S6r2WqjSXPjmbc/8oEO3oLEUdPcxBAH32tyXLjnWmKO
wyznMVgFp4rzn9dWcGjNerQsoaGfAR2d4Tvx4eMLMwp3utVhZZl3JWnNNseuFue5kRL8a6M7bPTv
rAJqa5IxSAkz55asg/Qcg7mh18ilR/25Xt3WDqmQzOSsIT28n5SMMTsarMInvnCRkvm08DWrJY5n
hEvBYrGRbRWtkXb+a/uJE10taq6EvraqFhVblm3s8plo8SH9aUY2TXry+uE37+qGIKo3fJRL/7lv
VpIUrjQ1jlCOlAqIgc8PMV0TjYonkjseKEJOW9sWThfUTcMg8miW4vtwsQUfq4e/7D9HjlH0a2L1
yywM8S0pPXe2Weq4jM3jmLIPMJER5aVO9NryAsqcVzEjNcKxclZD3WHVvVX+Vw+yX5c2BgBdbllH
mOIF8D0fK7M6Hu7w+qk35NiyGbqX+x+qZ+bvh3GDbJhBFX3QZRTqkJhR0zDAlnyR3jgYwjGEHHGH
Q9YPayMPsq59KMe6Ed0g+AkY3ZbNu2qFJLdMv4p/1r211gW1NU5ejs8E67Td/1W1dMWfWLvIxkAi
QWu38NAuwrWlrg9J4AyGeOtlyTNfbXresCD648gE5XCGPA4OifA+4TFT6dELn7CQNzVbMpIY6fyN
+tuHSUWlkjyzTczgsd0XWtg2b+ID5FPgTx/n1R4rpEvMrLfm0XpXvNpAQrCe4ADfKWMakfF8yYjv
K9YwbTBWSQpaYA59TNe2hT13M+wDz69k0zWydz1aQsacBsI3MSL2e7eXJT2fC8PL6CjnHyunrCbW
FS9qy1df2oYWLa4+IaePYu4cKvneXmLukpbphbkxy+lO1+iMs65+D42HHY3HssEC5CYa+aGj9Cwh
mmjMca6iNYP6ydgKCL96RQsF3MINcQ9Wld5G8JIT4YVkK0UJElsLZUR6+5xmNAIgnM0oqiBcGSU7
QWJ+e5DR3AtS2yE3i3oiy8u+20uARLWyyr8O97SIDw3lNNy/9VReDa1RonLEIKvGSG5fWVxpPYVN
B5tKnZvEAtxPITr1CCUZBe8EtcjfI4UUKzoaDkwe+ynV7UgHcGogKkQv9XDUnBm4JUBv60wse9d4
bBEQ6hxgZn0HBPQYWkm7ghxTwUIBCRXUwNgJ2UZ8C0ZwtdNbTN1S6nGDgBPMgzeRrBisHhMhn0yO
obNlbb28Hv9YPAArVxe3ZUzlCPnvjeTuz0pR/DPTh3xnmJvtNTeS0x8Q2CGyUa3IjlrnsvPkCuZe
t/mrU4a6jSl7ieiko5apLsaGXI7I2sf1AYlOTI18xWC/s0vDGW/gsEWiDsJdknPqyuD4aMhJQIsS
psb7wqiJ1m3PxIZeXB8OHNktn+izOntQeth6MAbArwYQO5TJUZ62qcKoSJDGDcKoqsQovjfTF9Rh
wQJRduiI714fnTNqYBk4u0rZaNmRzQHdK6HwX8hnmVExmYUiplREv34bq3xulQS/V4n0JVpVjpq4
Fe+WgW5t0rpNyklTdgnSxRBMMhGsz4kIXaEkIgecxmBvcqil1KhrYU9AOtUeR/lw9LeOZr/48FkT
pE/+cLzffuUzzZGzsb3N7qwSpT4+RF+KC7ds/zfAnV2nEsNsmhwLo2hk2CC67KfPu/FAOEnGvE1f
ET4/9pnBBmQcLPgO40c3zOt86JJD4U0AUBveVw2znv6OUfqUFy7/JVocZr0nP1d434CUrf+reabu
nQ9ubWMvtiTsAzNuHkJayv6l+FMhnMKr8IFxM7/g28IENiolzMbVXmmyzIkoD8KqiQNNvvNeY1/2
njmz/X1HlEqWFgtJOmaiJ16xGhTb8260W1k4SKCC9UpbIVjKTdnZZ7WMpGvGjDQn1Rc6H8Nef6RK
xq1oCprO44ShKuQRvjmjkqMALIZnExbnpVekfJuKpk71Eiyp8T7se74Tbaa4TUoz4HQbNdwqp86I
d9ExZTY2EvbHs1mYVpxB4GXxtniOaCu9tCzDkBLcj0SiMhSVRAM6zi6L2LyF3WZOoRWEB0khynbD
ajiNi7GaRf6Uyp+fhnHHEeOthYsHtKHJnL0qnNm2J396l9pP/cFF5ThicwKsZt8hIMiaAwUwvXd/
XTQoKXMFgztrMbLm9jrbFJgEbtsf00Wh1CC/tGdAXySMAnjxIAiapSlsihThhwZZ4Tc7Iz0qu6NW
csxjQwmzX5+ZadLf3JM/cSIP6UvBILG1zwNB0+2niFV364h4i+wEVShQtRLFphWti/8QygMC/0IA
JXcx+KJO3Nnj0E5h+kvAZWwHkEodwP82aOFt3dh+Dd5GyBpJsCWYSWexWrwFgeX+4nKjfDPVR+W/
4iDFxICvZZxVumFtvt/eWCGfNBWcovkuvQQGyLTDekhmSMz/IeU4Q70TBkEUiYKZenT9IILu0u/i
L6ElBEPW8UoGiMpTEvDDJcMPMP/prwyFDf2XMPdp9mCp9ur6MtA+62nlIKvwgvTjQDGum+QeJajb
Qw5AN87s3K7soQXaQr+cdq6MNwaBT2O3WyTq17jLGL4ojSgkNYgzrPLNQ+3LdnDjpSzUO+OptSvG
tMCehp3C0/NDXiL3NYgLN8VTsxdrbqTJx9MZ50yJAWuChk+nccHk5yoiz2MMJieFdE2IgEqsh3Ng
CeQ1FP6YWmg47rvYr2ZiO+qP8yjKL8CnhTuCRWKTfZ+touYLxcMv19JYkqRG9hM4My+RrQTVNYvc
08SJNYXoiQKtpnwovldforI224GQgaTHY1sCUeQH1RjrTZ+KrlGrm4YytgW37SY2feMv1k2+ejJr
/dDYLrQqMgg4C4UTHv/0/0iHvBuHhWNP3iSxGxdror/LtHIHtdgQj/cqXm0US3gl8RTH/e8+nGtV
AKezJlVww5Kfki9/EaKsP5fJdo/IwqZdivbj/NiPc7gPaM1fGQ83pDwj7cQuCx4HT6upnOViiKam
/yqXBqsXmnrE8mCJNh52UeERyUsAOUBqpgxPCqsozTEp+E7n09dZIBE8kTLWJp4B7iHp2N6KT01e
9Ifc0rz5x9kcY3Fu4oph9Fei68eumUmfLabboq+i+2EetRe4QsagDsT/ZNHYzy1KI4AC2LX8ndE8
Ti3EZQosNhzKxrTrk8+ZU3X21meMi1q8sHomjrYPLoMgyJScJSnmzVmFcppqVErI2dDwTWfHx90f
mIjygP+58Teq7CJeAts1N+KmIS2voLDU+QzPVF59VtlCY5Yb5s5u8Ucs5J46dWLLyaHGXmu2e2Fn
ipRGuEdbfS3M9HsdLrTtHCvhbuddiM2FwSS1wjKb95EgwUf6Tdc5BqLKc95j96YBDDONl+XeSY2H
Z8VI6A+57Be0E9NhZFkh8Rgp7mO9kQBjFIg8Ti36oK2o7eeKNRnaGWa5+0mdvtmFpc+Zs9VsygCC
IffYBww3BdBAm2iHOvldQX9aKJrDocuBWKoTrPF8t1J1JNHLtEtZXiltsUtNiS/CB/ZzGCuqhq6a
bNWfL40tPsXoAwrZ7BaeaZMvisq9sNlOlusFiRYeY7JcsgbejBkPraOgwQAqjhEXsR0HL7f/idVj
2GthEo9rNhw87zQT0JNf6HQBAV5jNjZ9slbfPapAOPys2wH9sAj3Zf2j0njNIJiAOZ0C4ALIUVQl
Rf6QBHqwoV7oFN/BdXXw63UHPSBb5ekJUMUTEJjNCeAMPLmHGv5cOQEOkCSoGbmMlwg9K294Zfr8
JCILZMh7YQmtS5NbnUWFJvvLG+Grr1OcOgoDoahLTYxWzfYlQoWeUFDAE1b8dJpXbhtqMfwHMFqV
XNOLkHRUyP5sdBqEh4bVVceqv++sAKsgo7X5aOoO1p9iO2CuAThswdckjypH5InIoNsEZ+Aostdo
LV8yLWaKHDWmRro9kUFtM/BHTe76hQk3Bzv9Oa9pjIbUjXGCk78tqP7av79U4+ryxsCeZOzS+Uew
1+LBxYve03i02McINbQEpz/Oq/5PGtph76TtmHVy6TYXUbiZTcxQoEpLF0bOMU4maiyRnygmtDb0
G3n4gQBj0+eBTB64BYsKBkDc07/3NNtnpnyQ/mVCunYVIT7iJA9h3FwS2CTiOKXG5qBSR+e7GaJR
nYv2nELV1fnXNPiT4vlHHZLofy07s5sucfksM6Z3wMl4x2d5PcgJz/p0mwLaqrtJgOwPef+fxsZD
THrKwm5CZB67YzsrZrFcsKPY6saWg2DKQXhaMtE48fcnQUXWQXmFqixtBTvl3FNRq6cdlNdrCEdR
klPt8VoYXG/FirhFIaUusRbTszOHk2McCkKhgoAtDjX/LURbX7mtqRMRy9BqkCazXZ3ipgsOKAcG
H1jZHGz5eESwGsmi5LVjqBIh1r3dzBGQvjrnGFZBgx/UoHXOtbq1pkHI+oZ/J8MPI+ZfvD0k6YjN
FEgnPf/sUjvRC3eh4FeZWifp0XbvEZbET2aGA5tcIrbOqPoaZ7ZtODKb1JbW8r+V3zb4G+8fywJx
7sa7md0aUwuIBUF4KtXq6evtDVyU5tD1t0kAcEg+q5JBfx6cMHf8RtiN7WL7KfENnvtq+TFLj76l
LYYg7ozgiFWFzYtIADTZFcjH7ZitKcpsnHem4rbIS0RGULey0wQIol3I92a0HXByN7l3iyf+HpA5
TuML6j6GxzOl7lu41iz5BpO9evDG2q+yxAxuh9TWBldmPu+ZL4asWpylVVlJz8fequnFZuzC3tiG
xWiVgcWH4pYZfATAAQpWxZhNHw+iIrdP+12XF4GT0Z/YgkBAEkn5qrJCW5EgHEb4z3wv4QXpuv0F
yr1nZeU0wFShwP8KiKO4zsMtG9rLzka7TAhop5mgDaaB8cLUy3G3e6NBKuDbZzuT1kR08/xC4q5m
5REfs7b2iowpvFMrwxhLuHADD4t6E7D0EwChGRf17B4LhnL0JPAjTEp99rTGU9bTNTzPIK8rBDtq
flUpIrftpw2Hbqs01kM1IVAIyeD/vflJcIfTHl77JUsA6qglQPzJeIFYrgyx6U+Gmd9i+vLY9SGA
wwHOcre9frtywLGIAMceAehcy0VwWxrhx2lOAenK52RO0IFSY9S+5brAVbHDeyWVezLbSinY8f1z
jMBbmCFhW1CgMreEnZ6iC8p1kxPLs5+zl6TCi8pXzNtOqeauqLax279HGlxxqiKT+z15pKdpJwYU
d+sBAlemj6GsRSvfQTz3OWbgc0fsiJ+FujPR0jJHz2DphHGGTNQfuy93rRXpXbRYTqqhm1Wq4A/L
QwFpLNmqYAtcyEi4qtIW4jA4UT2/blgKqbD79kjXRwyNFi6AOZ4n7O6+i8Vt1JIMi2FFhXCCmuWT
DZxNEqxS58k9OfFtKGb8s53cBTptmebP7vbr07BqLOS72DyQf7dvjwcwr+e063HgxigSCIJAyhDY
JtWT+x7CKcDGYVJyzODuvOPGLDHqH4YNgcaoUWHmi5Tq47N8oMZom9GHrD6ds77fIIMMB8WtuA3a
mx4BegzQMLOBf4wD2xYkPWl7VEq//6SaUwK9qrmhF+Y+4k/kSGR3OSl4GWg4VoIzJix8ZMpEJO+d
+74siJVHlQdLNyPCH+xRXyzPAXg7RPDKv/a/xZtRRd88DqaS4l1oH68WpFPYiZdlJFqO4lIlJ8Ls
Qd7RBCreC1/h+hS+sj61rlUbFdZGd45g0HO4bCOlkyFNOUOm5m6YHY42xPxRjdlWALTI1L4Xpb1u
rKaXFTzIMf5ZUzdDzRk2w9D4cShYAeubAeEnV+LIITo8K3ZqzqEuemTrVIhj/i+hf5zn48Ay2bQd
aZWxAiOBA8BhzHT1jG0sDgXSnM9Vuyx+LIPpAm7GrVYRNCYYTwGzsuGaDOo3EPTb9NtS5ODbtwCr
f2rX6I4/ixL8cbI2gC7FU4HpwyphBXh5zZS4K4Sh39SyNRM+jBI0j/vOZY8YDJD3yZQZVaNNpbTo
CWb8X+aFUZg4FMauL+aTBtnubiGPJNM++Ga8SGgniF9Do8zUVa0rU636bpxpHGlWs6XxIPSiaQF7
6ql9o3KFLB48338HE0NitDCPs35qE6SrLD4jD2yLQDD3Rw5VT5jqkMJbj6gBzwiQ01urXsUlpudf
diUTgt3BS/CSIJvY0E5Uaa1G/qAqAf8VCvx22qS5+T+zhfaKTWYXYz1+3OiJwn+QDFaZlvOQ1qKr
2O+kImiSM45ZXd1gV7NfyYrPdRruBje6dMHv97Y/CXWlxrrsLcBrAREpAx9MgvfApbJyHRxC0MHD
oQlD7Ztsbjiuj60WqRUNuzod3flUdqeXL9T0GrmTdJOtvdzjX7UhxocRjTR3GqZK7RA4kBL/run7
K9kdyG8WTvmJenRthw7Z4rhqQ9Eqb1Lh1E3jQ/rNxn4ElhiIkzPiOfVhnWiQMBcfb4CPhWhJqkfj
YkiR8HB/ODeXk53LHG+oq0L2N0OVlDQqCTBZKZDJvUlJM2st9HkErZwsTMdFyGrU5zKerhtic4gt
C6NHC3CHfUNxkQzxL2A6ysA/YOhLNpCAFPd8UT65Gj1u2Dy5/zZ/kf1tP6iP6Yazs5J6AqPiO2Qa
dNE0qvHZKcnjWSRwJBtLn3V02HKmQMdwY86I+X1qTHoc0dkIKkEcFNU623UUZrnIyR4sz374cO8f
LgR+ZQ+4uuvUnp01p3GEmjZqfssOh7R63N9SID/T22QUgDOIZs+WqcUu0KG4Hyj1H0sIaFVShfKx
C99bqKhvfh3IKBpog3ooP0GhejB5wU573F0bCWvbjtaUhDbAGYRVLYtKnatXZvbkQUPVJvMV0Q4J
+rNmUKwHmuC8CKqxI84kMr0aYBeolapUk7L76y6lZ/YiHQ+2Qrqk8HegqbNPeW04NKBrVMIRXkCu
Ua4NC76B8RpDwa/CmaHBeSHeZTaYT8ZMcoPQaLrfvd9NfIGOvNFGvc1Tn4/xEAHqXCfvvvj9DoG0
AixYJMAj67y+P91fVeNS/gqYA4Omwfqzd8vz4pbHIMqpN42/qjYnZKI7Fd9J/fpLKGTQ7BP5QF/t
NHNrG8La5f9VRetPPx1tcZx+FhSxy+WWhJiIpMU68ABfxAIZsQckVsQbyPc6/VT8PL162ULPUSlo
Wi5vu5uSo0QN2xtj2iDK57Ts2Ox+s+5UMwcFcFi4ECN0Iy33sDdLYtThghiL24DMrTQzWUWd4vDp
IZ1VlZ1v0/+w44Y96xrecqVq4TRZ1IcArtR0ayM2WlqyrZBLD+T6fCg3KGF8ghpKZXFElfeqONL+
R6zsEVg40wom54jOObe8bjuh5WM1rdq+oOdTcR/wZk++rE4K4ijP+qo0wX9Ot4+Fgcza/ngZNrvn
4tbY+7hulE/i8/41dRJKzL8S5EHL8QLVrzBnjO9XP/8sL3FbCN2YIwSUNz3zpS2U0YOa+d5L90SY
ty4yWQej2QnUhYdLTc7LvPI/vQwohhUjUujQpbUTDU7ZPv6AmpscfJLmJI79Qpl5vKvXf6b8NHag
EIByIhdKTC0PSqn49rsNSR+R0QzeIHn96gWxPZ9UKGIiJvCMFdwne51KNuf6ClCKfgVr2nZ4tlUV
TTd+MEFcHhzy4pZX9KPe6UFbaYLBVgqaPhy4/x4WyvXfkAux3iQ660AQb4qrFm3Yob4d0CibFGIy
5Zg6qwS/NF46cOFRAzhGEY5I9ReTAZKoJu81H5O1EuN8rcM0S/DFOYD5NF/ZEBm6gyh2xUfydHxy
uYNlC0UONdjWXPpmpVYLtqUC3EJVVwkt2fEfeKflpJXOfV/VAEVZa6gXl8gYAnElXoq+I8FJU85g
kV1mn92+7gAwOa5ZOzmUUCP9nFnmZ04ooB9XpqcGNyAdvifwwtHxZe+tSlxhPlXHUrufefokij9Z
4Sjeez9SrQjMv0GwSlOrLFT8QMxT/AlaTob6pyn6pwGmmV1OJ1TeXb0Ub56xCZ2TCkl2bzz9eNJ2
BI9bZapukFWDgqBKY0NcHuw6YcYpvcwZgki0SBcA+VPdfOFiO/Xm2U2jEZ3sCwRCfZRQjXCu9PRa
HBJpuq0/CLYHhsFDXtohAQrOMvmyIDIJQIngDyXxC6GRGXo6Xv0sKfYuIH7JDuKS0T/OKRf8ukBX
RcwefRjCfcZ5yZTJOphZUh5/ZGjpRIrce9PbOuVDi9TZHk/o49P/PmDW6BzNi1/Mo6RypKXgrufI
s/JCs4CTvNmyFuiQdj4fQxbQG2W0td1qbeJuDhcOHyqOGMyD3yaxTGwya5gTlv6kcp2kjKVCfxQu
FaN5zsgbUAmeaEAOxnDaMUX9kEyNbp10+FVFRXVWVtngaEpiBfr05bJOiW5FeYjuMFK0rcS/xWrE
3RwyE3tkSnq2vZOBTuB2jgvS2UJsbC8tR1aqzLZseIDX0VT9RVHEGTA7y3uiYcyiz6qV8I1a66p1
p8zwD/tBVD16+6ft8CxYfFzdfpztq9abd71YYiDKrGRSEbpYsvcfp2UwzmhegWaYKyoVjQO6O56r
g0wN70bJB+AoEWqzXtObAbBKKHMnPoosWLZoHssAki4bhgfwC0+gskfpx2cirfsTjCC18x7tv0zz
qVFpYfbqp+daFTrVmzfkYqTSpoAJ95fmqgT70VJtrt59L5WjgfdiaDkZ6I4D3nOhXwEKPhBSzru+
IELWe0j76jCzzRsFoWdDsICOXbGVnmtCjSsdzXP99T7zjTJSV42mRlauXXu9n3/iIX3iyl2LOUR0
YzKEH7oY8xpZ+kBW8cI37JL2n39QnTEhjNaQv5IXGLubPM7lrD/cLrh2ag/rz0RfzYYmjfmPCWR7
xUgs0rAX1WmOxFoGMvRbo/Jfe7uotPs6ptQjyPC4vxICTaMKOEkqZln9R4/SNTrzURQJequJqQSH
5q6/SiVXD1D/KJY77GLgMCmBoZtcCU4mEERt0I7istlgi454F5SybwDgBj0j73A0fCheCm5i8jm8
W8KwajcG4NC2VfjLlNXOF8/ikH2Cy4ujFVPGZyFoJWTNhnmMsGvXdrYR78BbZFGDn23sbDVtn8dH
f9pMyLhNkZgZf92vOnpfpNS2IV+7X+JpVNb1+OK4Wym69oO0Wtsc6VXtyut9ZqERcDbdJj5uweBX
8ft2Z8uqIFmPk1XhCEFAjDjQWt6nhXH1j6xBeycjTCOYG1Me3rZTYDovE2Tv+oODTAk45utUq/S3
guS+s/IztEYnaYq1QT4Qy8KDVk7V7UmbCR/N0PsPnvuaoKtugePz/4iEwmo5IzZCVgZuaco1fYg8
ReJ2gtTzeYFrjJjoOzHevpGR1VpBrFaFjUa37KO9ZhpgoWzJccvR5J2OZWl8duZ0DHX9drpAUrKX
lPCyp/WpiFnBsDyNwkkW27mv7DGNIOOlChKaN9qClNYzlsR3Tx3j9yU+nABJhyH+BcIDjhfNrxoU
5HSEjfwFA7XTvS42texn1TjoGlHdfLjUW4G5Yn3LhbqPhamx4DYqzs5UJhriB4kd2Pj29hkKmd3p
722FVD8sgQO056rssFnYAdEF/r0ve+pv/WRS7EGv3AqdPjZTiUVx8hWgf6Yxf0QjhfyFZYvQXZy5
mxKGx5dU9Tc8n5zrveNrwsUhz7NKJcAhE8oaKht/1Fu/6wE/v3QoxpdccOtMNd/G7Vv6oX4MgikA
x6DeRkWi7fI5ik+EqS+7H7R2Vyv/J49NG78/slegxp4ssifZQOVeIEIfffxB+/S2OLJOe5HKlDJq
NTDlTg7Rio87UD8YqkF/Gbs+RNFZCWIy3Hl9qlOVt3uK3/ncexXUwopaAEPdY3+9YDcHglFsIB+w
gcFIEQQqDkQrQZn0gqyA+R//2fn6EIDjFredYWYjJgFai5Cceqg2lWiiJ/0J4iIt0WO426Yvd+F6
8tRLFeRd0paj0Sis9oPqWuPO5+Bed3hY7jLX/6tciikvLO506p0mabWHqcHA1XZEgmlPsanqN5AC
oqdTwWtQm7Q96SBhnyjgdPtdwarDe3/+aqEb26CN3HdpUp1zIq3Vay7bYn0RzO9USjms/X9tTqBs
NTQamwt/dIdQpP/WXeYL8FwdS0MjP3mey/Yd2ICp01nWdbP5zIYw8SJZlgeNXt+DwVBynxfAV9BA
Q56IWlq5zDima5svbYjoYnS4WaAJEQ6py1euUBh7a706CVCZTa9Wjv54DbVVS8szgprBiYZ0Bu2c
0+/jIoIPPzLtliSs9ljDOWd07RWqtQ1ECmzieEP1IoQbml3QaGst66Xk9Ib/selGphLbd5449Pr6
D12/EfOT7HyDFIzUqKKuVmnRW4q1zgdc/5dxZkOViWMdeM0e/AyNJn47VlN4NycM6epHcNxco2Ay
It1fOxQ+reHVr2f7hMzoKFJxdFOO3u/n9g78U6Ktk/aBv3mEyQETPCs1eydqERQen7T3DHncAh7X
rDZKObjOFb/veqM2ftOrv6+Os9npPch3OBYDc/E0xR7tn+oSiR6GKYNvcU5euRScrcNyJbdShLeM
yi7akbcdqCyJXlciq1qexNoEMsByr8/YbOSENd5nkDUzj/ZeXMgUd134fO0J0QvKlDFmx1NLhlMh
pZrf68VSnrr15MyFxzhreL3ZsvEpqSf0ZyPQkcVhoux61YD3q6DVMLlGcumXoQLCdEHiSqoZyk+C
qr6m0D4SDADudIrPUSMNuZBRNXLeRjHlW+hk4rexuwYvVAfl91Q+4zCd9OUf6yHAWv0oseM4rQH8
25lcO9R6/kAL4dUopLdiDtkm+GNeOwM0Q6vCGjaj8+5LKLRg8+qjEDkRHsatICPepNul2bqv50cO
l6M6hW41oOWh0eJ7n7kr/Ah4h+tvPrkOalvE8xg3lKtZUy55c8CS9ZXgf/TPH3PpuRawrn2c9FRI
HcO1Ofz5zcSXWbdhyUF76AdScBj2bDdU9/6u702ej8/nCAi4BGzMk+x4w65EZZs7B7bYCKpaBUOX
ga4fB3brwseBEzyXGVPvjmzapMdxU3F6HzGEoNSSufUv4AIp+L4+eHybS6om8E8RkkTHk/U2oXg6
CqLoKZyXgfYiSW6hYss7ON6J9ydKuN/3h8a7D/5Xq2VoUyAqbs6xaiAVH9Nga6P6hX7k8L1eZJW8
Oc8eLvI90qVDZ2HJ/I6b1+4sslahlIe8Kp5GqLtKOJLCbzendj/ixTGUR5vj736PmPPHPCcE083L
sbX3Xrm6sG/p+esL9fePwJ+xNyd559mvqFrZ76RWVzdtk6HwHMF9gj+76hvolVRp+g/BHZLg9W0T
4BrZ/X3c1ZeTczIGdqmtqtTPB5EPROG1NwC2aB/mhl3KYLsr/skpmTdN0mmJdcwMdmWB7p6+kWEI
bMQtZRuntcGB5yOuaBzN7vckFRzQ9/L4GJG5bz4YOsa0KgAn7HqERTzA2pHMeLrJovA/i4pNWBaT
7Di4FhSGoHM/+/QqsB4dVjDFsu4309B6EHjgSq5LmjeOh33z+I1piAHWy1f0WpxEgqcMCFHrtrPs
wcgQxJbPzM6a+T56Q+R3ZOFCIx1T6qcT6XQMSXkzZGux0mxhTdfq6urf8oYKWDW3UoDyp3MBAnsk
kpqJGfkeX6hUAzOpuv5ACxKiKpQ8/w15zgwxYLfamJ8vXYHTLEaQps1zZreX3/BX2lVxYf/ZsDLF
mMp5xQoiuArSZjAsr1Ao8M7j7lTZl/PzVQuEcaERNSsNqio89LSbNCu26eKAni2GhNFPbRTS/sTX
B0wJvVndRx6NCrIaz+7+QiBznYEMohb9DYL06/wWsKVcjecV9tOMPVOR1F1H9bJiEmrdHYA0bOxB
IGKNbWjhetfVWH+FIKErA+fpQlE+JmKplixrzggM+9VCUEgCr/nJCf/N8mYzxrua4d0sa+LY3Id4
r03ytaseMzjm3l4bK79TkLmGtMyjpD5Xc3hQ27KY7nIaLhJHUdUYbeMcvhASYSsSHukSI+5g6RoO
LZ7Vce/m7mDhhl17Dpv6kbEA/yZFMZVecSd381GgQP7QysqBhxCrlKMjfQlELSWN3OgCGkvZKhqP
1aNNbuE1sRRt6MXjg0s7u5zV40H68wm7HD4132IKYgL6753nFLCPf2psP8KJrble1eN+FANYBWXV
w+adRMAplz0X5XoByBigJvEDjSoqRXn/EIsU1cHy+ZHLvkH6cNYfScTiYGb8xovz6WK8F0WXVeXn
yxBXW5IhJU5xl7UIflBijdBzwTRt5YCnft3nzZcgYlnzlXMYxEt7pXKvVj4rbDPOFLcgCF1CHlpX
DDhOC0P/G5Ma+kgZ8Vpi3s49hTwfXCCnrYRcPEY6g8ZPwAFzTsfUf/USjlVi1hSdsy5uDpOpeJ8e
pblClcxKnHKeen7LIjGJEcBQSaO0nErrEOIwj7v/mrPlDbjcDpWvTm8JtiBNvdIKXi4a1kknuY8c
L8MmUp07gD8FQP0tTr8+x9nK9o8DT4QL42Zhdjpej3SNahy6oVH+pb6CGf+4kTX24SqjlsI97m2A
xx2/8aln2fsTvdTXaQThasopToM4m0KBEnDpOk5fHy2wlx9zq7KTfup6iWEtJfVRNQWJJ3/gawZU
TR6a8CVTxuLrsh/4yt1lkhkx9aRZ4438wMJzy5bn1phQh3j+atNgj6ezF6TBn2s1v4PHOPaX1jwo
fQApFQfSF3X+8gqsvqf9D6K2jSah6eqPo4fUcxrhhfGk/tr9cPIfkMK6gZlR+pO1Bi6NGRl8vW4t
KS2VPsLSSSAWJN2Xx/XIwrxbWgOqESc7GSHH2o5hrYjCVT0A5qekEiPK7hMayULnFoqBD9yr50AI
2/EKd3popRj8hZB7vCWstR/pDnXbrSc8aaRr1HASs1k5G9sn7geBq7XqtpiF22pppR//mlchHUd2
gdlSnHJgnuCkwe76BUuzyTAZB+Ao0Q/VnP0GnCpRpvJD2NEEHG4O02j8w4hUo1N58iIOYGK3iU+Y
oJ+M4x3wnHaf0VvICZkzq3dLSKttf8cy6RPNUK/BZ3ewKa+POoTbaYkaRYvhW5z8cbokhjch8Bzy
DxU6RJu2ZWsCJEgPaY6VlRhjiA8WC4NnrOfQup45HJp1cq0OMzRcOKp6Z+qYk8DjtpLFbjqEKmNS
/fG+c+w5mngaBo0XeRE2U1HxQv1ycfuvoFNlQUVj1zuOJWoyadit4IifX9hD8q/0MUN6Ic/GAjVZ
rJGKQg3C3bEt4AJb80IAf2tCs0x3q2h1GKpYDGIdWaeK8mqg209WjJoB2pgT8f4NXVS28TbGEhTw
xMBl8cmvPblXSa2qDtCQQdPqrbboiqmnTXLyajWRxqsQ0vK56yndw60n7uoeDhmowptD4Md++cMg
ikxaJPEW2BuwwbzjwoQ6UKZjvaeLxZ21MkyqqYEa44xvAd/hHnlf8PBm6qJfRXapqIM0BVX5TPFH
FFzUX5Tgi1D9E5N8r4UKI72C5njsSY1mgNpxAM2XnaVwLKhBq+mnzPNRdtEojLu4nRb5fKWRiY7L
fqSv3WqOysJdI6o/NriE9ynk0IXWYjNY7E4qGvA6b3aQSLjqjrWkzraEWIwew6hSTbzrakS8zLCt
sisGAOsBHjbZw+QU7stjgLN/X7l/WrZ1m9jfCppd2ne+p3rJEMOFQvdzKkA1MNfbCYPppxrw+Woy
X1Rem+4HhDbIhYKPlpTtzsjGRmM+Z+r85I9ycgBYoM3Fwvfpq153z0ADIcJL5DMY6QXL0V39cBs7
2Tg7YRAkDVLwlCjVIyYBf8EnmZrDAjLdyLyFOFo3tR7D8p+XaCC2AuI51Ieb+5w6rXtAq97cpSkm
k2WZ9VJ0LQ1PZHEEe65CPDMCAfSgl46dzi93DB4y5PklHnNm+zGgRpHJDWz6GQHAPf/ahE2kO1mn
J7Fnzg5IBbSNZuE6YqtoFev4Mvc1lLIGNq0tX8mUcEZBxxaRYWFSAs3zXmptiNEaexoR0Geb5S69
n9aafrUuncBRelfVaZ3nrh+lRmtXhnhcr9JXAQJyn0iOAyK/yfH4XCDKn/YgCk2vnkXIdr5uBcJT
8Z3ca9v0/xY8HJ4OCr6K8vvNj1Ocihj4DQWyJ8intmXBrzMv2GBjeqwrLdlWyrL93j2hChagKdwz
RKSLOeOVfOU1bSlWhb9CNUh1LzddWr29fXP3KULGwXgTZtHSV2zQJPwA/cpCtvDuSAshegFG6FUN
NKgXTVT9S2faaoaLcbdBRnRr41qfyhA8wKP9kLBNCe1Ot+obsdrT/hNEhv7lsURVt+l8SHCn84RJ
a82NVjWFSP0i2fC50umdCTSJqDmoQYOPY/wz8uD0BAt3QNsAk9xI0g+g2L8mddbXZEwhGLTr8enV
KwmKQ8y8Ej7V4QvDWPASHDYKvaqQmPKGa7+Cg9W6I/7Ov86ORwBBXbv9vCt9Z44TU8tDQp5rPGdm
7YZujDIb9KHumrOHDlzGLe/0VfPxXXjvDvyYaNVjlisYeM1tgduz09/Wf187n5Hl6LDUfZKVQy4n
CJ8Bvu9kXLaAMaW9I6Koqj3TkI7gguQ70VscvR9NSrudS+HpWrx4EBdJjzJc5p+i3HiaXSU0ryWx
Fg1WBTS+Dg6dn2uSl9nHMgFpjfG7RTtTT+SujST1m97trtReiozIDCUihrKn42o+2Al7jig3EpmB
RCGY9mqlf4bGF47Liy9X24MvYStaXs7pV7PZcFxc4hDrGzCxBjtLnPxclb6437mKELSU6+EAD4Ee
Sbb2L720+sCzNYfNQCCLFmEJEm3PHgnWNXs6JmwdzJBWn9XlTnV5FbTIfzXYrM9MatjoUhD+sqAp
3MFLvNMzjr9B8Dxz2INGMDARsYIqOso9O30vG5vPPggZj6xkLCWSzi87OJCUc1XcXygOdnCLxu05
x9DMRpOp/9k1pb0gwBFEAP23syMl3rYbYjafqejPD3KzYvehjcPiWUqum83DzS5ZVHsCetFgKyyu
OgnZTLe33T5mmuSE/xUpeY0F6yY/8t5R/Osv/id1K0I2jPW1V5qkca/ZBM/8A4buWNu9mjjCQRN2
lKAHs9dccFPMF0wvgoyLYbYyjFFaJEO4kluaeJ+hZQGsAPaksSck505D4p02dSht/y6eHjuINxSJ
klCksrVKiG8PtQE0vPYsKLZxYoG/VnuKsFbeOS6/0pl+B2N94CZrVeHT9Wyl9pkwoWcPfEnnk4F/
gQEPVxeQ5TFxWnS/TT4BaGx0pu4J5WQkh5Xnu4Vfa7aDv5x0t4PKCwJLkDNa5J3YrEr4UQX4Wsb+
xlGvUVUeDMeNuIGN6dDa8ICOlMt8pWEWYqlFMxNa/U4/eQIBqKqCEcABwvdK7cX77KzYjya0D31R
HxqpFGD/S8/BfmHmDRlBUhbeb3t64SVb6fR2HoEIeL6w6PW6r7/TLSeS6ooCiChhTtvFb80K2XtA
qbue/Bf6S2XHI/r1ZTwQneYTiNKlS5kw/NKHi2t0cWx3aAQbAnjvohVT6Yv3BU3y9rG3sxVu1FI9
jzNnLJZP38gsd9kerJHxTaTLiXt/zsslLfYbDCi9xqLuLdaFuYO6dhp/xJwkkEbm3SyoaEEoytBx
8DGe5fQ/YFwG9MgiRe9VCh4yJFgCjUmm3mwLMfXM4akS+Om1TzAX92/NfoI0cpLvqGZ52l8amSLK
ue/BM4HRI/J9cYUXW0U8LkHuYz4EXy7biA4Tvaz/fOkW03kh3Cf9adv2vLVboWC1lYuyo3NBJA78
5O6BKI6ZzzKXQe8qIux7xwhTjPCM+IRiD4ZxtvU90d+9nS2bYbIbjzHOb3FRMDwjggkt8WmMG9YP
bWFYAcMlQk0ZJpCC51+i1ls0sirTi7GT2lkvPAJlUffp7Bj830807P3Mfs2JKo/RQrqZ/6ekQk8/
4fC1RoLHqEKfzYMeVq/yt1UFGp24NKrY01flBGZkzpU1/gfJoEZSM+LrKdfty944aHxkjcJhInTT
PAUChbICHey/yXX9VjTe+Qwt+MZYaNAT4GR5FN8SnvZA6iSacpCyWip5275mHsdEipVAQjTqbWDL
786u9jXOV3xh5QcssReGYkJrP0e7giFaidPM8tKiML3EsfixMRpDj0W8L2FpxphRvShgGUKia4nH
FzoKEpipThwdIBveIZQM6YQfHvHixbb59s6UgcWFAVMyV9JYGU8s9IDQn0GzXTNxJiLXYvLU2lx/
8Cz271oEsA6OOxk1hkCRz88uTLCZ0WBrfr8kzQtlfchNbPa2efKGzZ/YYTDGGw9LxIBGvbEdKOaM
HVvsVbFnS+ptzEQsEwIrf7cRKMnEq3HbgoAieGVUOuQBTPRZ9GOa6+5b9DLr3xefd5rCVjoBUJFG
Py9oMHXcQz6H/bCJnOnLcVzZ7c9y2ttgqkKAabIKJUVTHyKtMltqojjSpsaXnNLetSg+o6KupeRV
1lo7kRzs/e7vrKGBk2xCn9MmfcDQBVR05tN/RnQCjeI3EAU7pzyfxJJ2mWQXaMKwLv6mlzZNRE4T
vW42u/YJEui48p5kmk15Hv7hRL70gyGIilOmy9O1+oYlGAXIu5jjzxyM78YbUp7uUp7VB6V4iwPC
hTc9cvAFizt6+k95n5YWoMItH2CGaH8QNM5RtYCZU3yyBN8wTfEruSeLmNMrkL7kLKKAqx5hNmfh
4uW0unbPrnkl2HGl6KxyeSsEuchiicINRgYGjG7c26hozJlywS5Yehj+eGwQVEDx34Y2EdrF8rBu
8xJQUVBJVp3k7a6GZjM4hEvu318C7ifVXW1jY/Qft/M3VuGBCZ34NHk4/AhrXsgrDW7CIVmnOB2F
z6sD7YXVZXiVRmD2dl5VKD7DyFxRSUfdxT7iAER1ZdpKOGjVAmnulP7j8uam0rEOZGqu4GZk4jPZ
NcU0nAK1HYZPThqpgnaSGad1tbFA7Di6lk4frIm6LYzJro+Nkq6iK/zBjKd+gLw8mqRZWzhxJVBP
JkWdYbkke0dAUwG6J0yXTtzwq6DR05Donl3ZUwOS2XSEBGaNwKd9v3psp9dRuDrSh4LFjsQdRAxQ
5ylNE/1yOJzcTmav8vniFQV0glx+96bSn96eN6fb6D8amze49OESCf9e1Hr6Fg9OZ5aJwbB+Iv2J
kSLrl+IUpuc0WQJMw+NLaHXWvKqOgiQX3pzyPTz6EMyS/yPxQmcQBNG/rQz4GsTtzdCA9g4ORjNW
SVVdK4+h/7jbxC4ZPNdJa3laF7R4RooLPj2Im4FLEM5adQ6H43iOPL53XqIbu28fBzOVmtKEEYBg
bWjRKcXU74HQJSOXO5xcpldjjNi9OdTzYKZ7VQKrMKhwhB/P9vLJOKqyWAdhuKm7gbGDCJ5ufzsU
FhM07iacJBLoJsc+XqGc8pW/eEmwR4ie7o7DrT5THX+oI02rVYT+CRJXEjpul6dEklvpLFmUuOnF
AdiEiy0hCEFDJokz/pT3KkUcYkq1tOy9HstzAo7j3EELK0Us+AsJ6XlaSX2zeqHJj6FV8wrnIwIz
FADtv1oAOuU/X8OKZP08De3PUB4GVdPVhw1c5sfqodUHB3b6PneOfrze/JXUUF2Uk9XrWDsDTEnZ
edK4W29hHK2oNCylf9ZhV9IUyzp4lpjFW0j4zXntwfy/syAueOdZgmBiifeoLmxt8js+vBYG/Jc3
KA7gnXn/VxDDt1UKjYOfNJdHwy8RXFKLzJ1Fp487tkqeiN1So0zeojC+SWg5mK/0OXJu/xZ1AkGW
DetQ50BdU6p9CF+sxSRTHtC0vMUhBpm0LfsHbO+GOCd5l6Q8Q+L104zOoBXdKrztAgZr6fBCQ71F
ycaMWOD10O42rL0Pk0h8wlmr4lfowDLKQIHz6bjCcTBJvmjmId1c+So1WwUyNdFx328Oh7K3wzrZ
UYDMAGTHjCnpPTuwXmU6fuyNgcjMZhWTKqctLciSbQV3okCfX3YGpIF4xPweaYjCc8s5ULoLkSIW
2RpOtR4JSDIl9AJMJQw77HTR2OSe3VUnSFpbXFz7N6riYvlWA9WfsFazqnMUYa7pzIdF1N5t/m8r
jGOONtCPcU84BXLeqGzPjHHFh5fej5tmEFp8tf7zmmVJrChuodnMC7G5vnj6rmswYSP73ykwzRCN
thz/zHDMCTqiYF9/am0Em5q9kPrcYZ2fbPd6H+/fom3glS2XAd9JsN1+HcB0YD8xL3qnyycLlT6i
cV9r23XqMmSu0tIEbFfr5reZNKCr09OpYHGoWLtPXtv/1Ekr6NHf5W7nNB8xrllKXOI4Na7q7d4g
0uG0QxlZ4t2HZuMcs9IXzlIC/OtHb9DXlZ45yhNPEmdxLD1qazBS0bI3GtQOByjEM/na86merI4G
CWIMcIDKf6Mij9+WrI/tGIzo8WimAgGoGjHodp6PKRataao37xFxp3xrtlSwxGAIHxfYfrxxow/S
cXSL3963KIse/4NgOgOwruv6Wcky7/QrKHF6Bybr2GjZkOseobj1VGa9jxhLYTQcoMeFjGbb3yZu
Bms2DN1/TMUN0TLk/MRXYkX5Zq2zcwwcaLdSGVDuzMYhcTL4lL1LChfyk6nLjL3E6zryO1k009lC
oR6Po57A/q8sEJBGGlMOM0WjEaCZ0zC9prRl30I9IaX3Dj0QrFSeQxRlDOrtlJcvPKKVtGX2fIqa
w+FWNEtoaoFNAyAT2p7mZZ99PzNIuWUMNjkSqWsMwcOj1VdSiiKy+mqmnNi34aGCrViOrPhqM4hh
pbcdQJg6kQe9lqRrA7KhOiowKKdHbmlAznv5gvYqOii/qM1HyYv6r4/a4X7W0qN3KnPJpAF3iSyb
yoV4hP7Opbq2Ua0bhzrcmIrHryquCQkUK5p8xrjy4K3aC7WnGx0ZGv6GdHLku7U/i3uo85PzOCGR
C8oh1QPhcbMoQO6oVQokvv1Sza/UQ2xhMv189CgaRC98R1uOTWYd6XwXnq56CHznrZveXQgbTB5k
lN9s1NTrfJg1v0xNiTAzdcwgwB6pFqykPI1ZdU0JcNQ6f7cZcDHVBZJgezbFuFmRdJf0lHJ0m5Ma
yydp222vvFAAoKEGY5vKJqRandUxCVmQ+xH1MmVFaODiPGQs4S4h9F9x0r9t6NzCsIERsGMLBq5r
CVtarCHllIcx5xFvqvye7M0lpEuTLlo4fcYl/caBEOcMa9Oii/IhXcPQgshILr9hlyvI9il8Ju03
ur6HqKFSaq4Z7EiViC7U7AVxtelkOSXIY9izJqJz/tljeXZUJVtxTJTH4RQ/0qsm0w1FJuGzf3Vn
72ZaDvWA9RSyIgpu8U17tkFLaTKGZnqqUsxZUtXSXRdgETJCZ9pTHDyQQOv0apbMDQHkoQ1lcU9w
lDlG/wewMyitcEPp12vVduUmiOeFW0FfzfPTSlbsIN0stIVL/OtyOUFzSxR1tbNivbwNgFBTODLc
ynUJWR/kqrUEyVfyPK+PIuIyh4fnQ9dt6mts51f4VHfOMgtnqI3lYoeh7G6u3nODTwDDcKgz0CKc
RkqSl5rvxpQWpWdETy2YhJkCLJkQmScRW3hCfkNzKcczhGVKBqAYE/HvW8qLL+Alx1bhREoCh3yB
FLrK3fTXOuNzihZpRuTZuTcQEsiNkossYDYHfj6s43Q8Fd5EvOz+Eao8WdNHGACH2u7tK3YN2VCY
oE7fxHBMwMOApdoMVPyI23NHe0vz408kOJ7oMRslGpuTWo8uTRZeWHFIQ7AeYQoViVHYjqSlkMw/
1F/QpRll63kt4b0UJdEEPeDJ8rBm6ZY+yD6pc3ihSIBYm+Lrr0A/rl49m2WHBxhwfZUoQIsIppmT
qzjlmZHkVnaw/S2ZdBtNp3FEuAtaBW4mk3MPE57LG4snZRY7EHmgj9rUlb1SHA42JsR85WAV+30r
PAD9mXvRiB+sPGhncgV+vuMk3Am8pkokcvxLH9pi2oNduBuNKCsx97b+QqbUHW0i/BhesU8gqK5b
0/8rYYTBt9BqemAaZw0bIWjzGD/jlXtL+4NANCrnkt0Rn0q6UiE8ioELl+0CNNj2hQOvwsofHoB5
nXqsleoE4hhGDL5kMR7vJZr6XRa3Ck0ZpXXw+4l9dBk0/tkiXKbc2AgqJJ13+v2L5cXofny6bIyb
mTewdIG2b065FI3HFhaFIKAvCkCNED5w1ovwO/0fgt6uwze4HoBtLNxzxa41WCk0XUrpcPWfEpC5
jWMq9nJSrlDu1PzvGidlnR8LIJxk6V/EzZsG6LsgR+dC2du8pKM9Fk7x//VD0Hb1n2QReMO9ZS0B
vU5iiAJyyZUwf63qI86MXi/mDBqPy2N6GE3vMRnHo/PgdDCOZUZkSdZGbRi6/uGiK9loacbqL7KQ
LK/XEfqjTKKzCvQ7nBPLXzoN8eMaCphf5OAerqeMy2/mTBTi3xuY2Zjf5BUIx5RXHyz6fBiDvdSv
e2o1se/0u3P1CTO5ql7FoYUVHVw4jJwxKrAeTMsTFgHBJ0COyyY/Cz93+TSrHYv8/pw4NKUqC4xi
6sNQkewKHylPW+UhoHNTHeIqRyGtHMwQZZF+bPb6EZqLLEbxjz5A3Jb1/V4WjLf8RD5TeljAuNon
Pwsw07na0/uppUFnfjMxud+gDsqHcwOPRb1yCjgCN9Cy0JjAYuvh/voD/tHBC8OJxmFGDZr2uJPe
L2LVjcjF9DEgmNPkUnrzMKRaJJb2f5s6/rne69dIUTnZvgL1LgkyWY+4HACBNFGsIqc4QAn2J7+2
HMFATbXKBwq2/uLFKt6hCUp163et56foWx0GvHkvzC7RZiliaKkEXMm5C4WEIi47FwefH4mFuOS1
InAjDQ2jjsrECn9R+2DgR5SuFZCyIjq5aP6Bawwz716SWOEDEczw+TS5rDc5Dln2W8CoZrNblt+O
Z2LNn51eUK70BFtEGOnhBbnzxZL6m+K6/PKe9b6jN/8dNGh2x/5IL1fk96Ps3PikJktncGjPLigz
ANw/R/u4A2Lpd2ncElzD7QOQGBqY5BPcfarHpk6tZjgca40Q1QDGl+sPUsz2Xmeqw5dikP1ckZAq
M1x8GAHZOtF9zyzNhRvIi/eobVFN7PtCh8rOxPB67YxG8mRYtC2CA2rrPFTwb589E82KSJHHlIYM
IJ9EMJuYFKlp/PmCUrB9095o7dn0bN8PV6E5TneyKy+aMP6hXDQyA7USqlpCq1oHobqdUU4RF6ew
1mACz0LB3AMqfMJthAOgIUF+ZMFGGe7L9R2YLSltguFXnltbrA1VKX7U4WaGosXzQ68xJ0orA27K
pzPSTUVKDwlFzx/6TqXJ9OvIcFZt8WP13NxoBepTbkE3JKnf1q9XdQCAa1Tgz63bEtdDu6DPKcA6
BWIzzhL0roa9gBk5E+iMwCORMsZoI1swdgFxDgt0+Bb7j0sIWI50CUK/1o22UDOagp6I0DhxLLq+
LRbVX9egG6kb4hHKISTgkR2jL1KUPGEwBRT3hP6QTPeyeQ+VGZIgXFFb/xIKS2lRXZHX4LNOG/Uw
TlPkehkfvpLRxLrHy32FzH8TSJbVucOjKj7PWxxBP/qmubmp5dmKoPRjAh8wltCdfM4NnGaVUOTs
LI3U6GxrjMFI123GfIr3QtjQBoPdLDwkxhox7+wtZmVa3qLO4BhkdL76X9riM2LZFF8x6OQ9lj4/
XFa43G4nguRIJOB4U1hLy8yRlAu388EbdUHAyy1+UZeYYBP6+ritQ72S4vTtArYLkH8AN5OENnU+
Mua5D4Iy5Hjw2JDlLxC24fKJkgANbY2DF9rOuCXGpPPkavjJMyHx/2RuuMT1MYoc/GEY4edl/eqC
z2ov/r7ZeS/oovtGAzHTLQwWJhMDC7WMr/mU3DDHaHJntgNQuLPFmlgdI28TWLfT0a5Vd3dFU/3q
rzjVgq9QRwJEUr8sXrTGgMJ74Qn+F2KPhclioYqtn1zKb3PFGztLkIVtoQlR3NQqW5KKCy+OeBVo
MCxHglRSNi6HZAqhZQYTxZE37/fDCrLF5tts3b7WVG1dhFdES0ymHjeXtWQyZNIB9Vi21Ohi1EFe
5Pzn8L9mv8vQLAbgxx2E57X3YMYjOJwKsPaICjirTXhJ2H1ri1aeMHxIIdwV4YbA0ptxEs87z+TR
LjMd8WcUaBKgOBGHpwjASFeEDYYPJJ/uoqHSD9WB/tm06P7/XxODAQ53dAuCKH+qy4jmd8F8fkGz
CogV/3slmwYnbMq6j32+Fbp5mbMEoRLsai5NT1R8vei5MxXBbaBpZhn3VyzTI2v9CkZrIw9wMJ5P
YsBIBMXpFuucK8zQ1Jw6MtAKjgAtJ2sPxTjxD/oY6yyfIGAqSc39WOezKfZT5mCiwnNawh0LCDuf
QTUjAD52Z3IYmnb3kzZzvvm77H1ERRrnacossoviC/zqBqbn2JdGOSwmNT8t9sTeE8V0Gp7iGV0b
aRY2LRVpvvGLml240db1KsogaoNNJP+vi16y2EyoFn/bCIzMz6Qupp7/k/w3VFkHPsdfqmpf2zdO
V5B5OiSQgMU1WRrrGh2e119RsoJ6C3ERfuRvBzsVZPywOSfI/zn+sThRu+d1fFkW3BoNf0r1ueOF
U0vPEhN7CmT8xtG4oRYWIE/Q1DWWojBU37rc5YLyhTL9kbPtYJ+3SzAwII4LBI71KIggZ7Z6jAGC
d4FmmFkQasK8z87ZnndfA56VpdGnEKXrg9GQpeC7XLnQPKjHggkGEEmb5OCxViNzeEmDOASmvR7a
b0Nfh8qpQD8xM3ej04fLn+ytiDKOaO/Nk4E115oK57w1+YTEHEbiTNxxEeD+8VEU5QVv0GQ1GIvR
vjh+47BCu+b0MR2YEyuASetVcZTwbDsu32LM4qQczANLFYTTbrkx8G3vUE1WihUe2vFOokdOOR83
0Y7ENn0AzlEiLcb2t9RZnBu7kmE7cTE8WVlJIs0kAnRzi771qhO2mmNfnd24hJgW/GiAScuSg2/T
cHBmXIDUcuklV+KOqvQCyNAelzOQDpzWaBtyvSncbPHighsexXkV25H4ObokfEp+Kjsgd6dxhpub
W3vs0bSP5wB0kOU1qT6o6STtCS9P72g75pEGrI1mAzjLOr6o+Ac2jgiQKRVl787ng8+X0MfJ45FT
tNsa1yxOzHz7bR6/aOUOc1qnxS/oJWh0Oyfeki6U0dzd7OIBVzy/M1nmih5GfArL39/5/jG8bkvF
3w5ANHCjBJ1EBAXHZu/Jbnk4ltDkddYVB8P7/6P/49rx5I6rrQgc8DdGqlzEu5nTwewm0LMRdnqE
RLU4oyEs3NO9Km885SElKpIpseJ1vciGXR16wcEJAHKxKIuOKz7BjzkVvMXRIU3fTvuMOUDfWamS
alNdFRiQPA3E1W9DaikXGiSm6Ixb6Htw7NUJFnZy3WrES5EOLnDUvhwBxKQujkCMdPnO5aMTKvFI
jdgSTtVKu+tfw1xXHyEa6B/BKAyWHPdtQEespAnaV5I4A9wExa9P6gPpNiVRmxLLX18sM6fU2gGg
S+K0c4c5AQrAuliiHWvMsy+UrMXMww8ltt2sbQ5xKyrL6SCCOuu1FV3Cgn+EgFnmjfBhHQH2z7hC
fX09fr1ZPg3MqrrL1ng3LcfwDinOgGxdmTKeFAHguFrVme9M+mdZjzlIli/Y97vlZ8sCoMP7IvaX
xTwRE8PtApNJlWXBYCALhj1pHzQsrkvwOq/yCWQ0M0uVb8o/arkz9+HpYEhG6AiArwLEmY4LfeEs
hm7mNutxdyA7r6peoAV5tN/5DqUrwtN/RaE/muohOwBU1wG4ZCtPtkAeUBxnyBdlWu6/yyD860gL
6u5es5CYDWpF0+vlQR4siDNNTLqq9UqgutUJ7JXnIA4XUJ7sMwS/RWJm/QC0uHzWQypQgtYnqugj
H3xAKZu2ErFIXvAX2a9MLB6CY9NCCJ8AZfNFQWnRZq46ZfrUpHoVItjwsDMsGekI0jQEtqR4Bf8V
Eib8J+/7/iBtVuP4L1ryV3nVnlTbQldWeFMnPLywqKCesj67IFk1SjLXlEht5Q9WpZ2IJQl7bNQ/
j7JBdUVV3qZT4wkkduTSPts0vTgYtUa410Jt7MQuQmN36t5m8MRR0sJJUtOLu9iCtyjNHGhRAt61
vdRKdOUnodWGtKKTl2lKm70SpV6Nr4yit/XGg62cYrGLxAfKfK/V+J+EE5JULlabQjqsxQNatFIu
PU8GYkL3DirLEW8+Zu5aPY5zD90T0VBSeXDQYwj0Kds1Q2K/zdFgvn8q/tJOE6IxiHXSparX8lUK
RRMTDvuOiBcjghZPr0nXywPG+NorzneUZyFKuHCPpujrG/ahkWzGHc/phDJusMx7G5QUFYwYAZun
PYN4a/mepkhvY5Wnzh7+l1vSgor2BTqZdl/V8IqhqnDbkKLTAKeN+/qb4CM0q1zAkMKeK+gNBXgS
fCmrQgprzNm8ivAaTIxm/UQXZxK8QrRXb+kp8RWXONQ61QYmtbxjuxm2SGNnjfbzBOTeNqs2Bz+2
hv64blM58+MUAW1C/cvcgvYwaFnjbpxak8CidYwb8nbmADoiGduHKNMwwnfxLi5/zuBy4w0PTHp0
XRLk4lfK8yZqrxiJCqu3Pudgxm0lajQ9dKKXlG5PhR6qhYMi8gMHCjFebRgOTDBEbPyuXd9u6x6W
wCRsSldF0+ml1XckRnEc3DbfTm9JSNpgsxtWdeX1OREklmRqhdpEZbj4OAD4qvR3KSTVNMA2bB/H
1qZqDbBLfulQk3UcPMCgoWR0TeRgN3d3Mw8AOphmYscgGuBqDrv4R6GHTTsMvzGpZR0uTHwqJoFK
AX+RNLzLUL7fcgFBoUqFIqNHoxkxTjyHQ5cv/bUmMn3+Z7T1K666kxdyy64ncLNrqFIhbyHoZ4dM
DEzXxTIThKVDl4xX+uo62/OQamPKshboDySjIQcc0l19Y/GoLYuFlu7fPxmaSs8aACFvr23fiMRM
HPyt85Uk2K2LYBMl4v45m0ZIVjSE/DqHXVcwqIielsG+a37kpgpretyKjv33+iQOXwh6aXz3LbSv
A82bLOEC5JDppejQlo+CGoNiAeupN1hfctoWJqsH5yzn+xnZ+NJdNmzYlg2PWlO/uIZ4KT8sY0zl
UgfF6FFCjJGbqpX3ER2NzCNHV6ERHArpf3Z65NrcsmQgWkxfP5M0QhCIOoEJhzjx88Z74nqRUOMu
opQXoE6ooVapvSEgJNJg3riecQ5TE9ZkkrCGsfGVdCwMxEXeaiA71CaXPigCNCWqjSrJBD/KVahD
jsBEYOWloOzuO4l90ubDrrCFj6FAHmNzqUf9jPXeHH0lTZQ4a4PFsIo2duOSKM8Xirr9+sdsobTj
Q8V4TkoEjvY4kKdhE8L6aaY7dqfTvrWHxOuO0SB1WVJGkeVrkkJXohCjDxTaW1LlKfrboiEoioIX
fBtAVm5Zl6nC7qbvUfhcj9dPODkIe9NybYPLzfXMvfcLUd+s6BMjcFpLmzvz+osZah5T1BJjOBAp
x1jnbK+A3oJYHEzNETzOFSswYQ4YUklDY6nxoc6HTstQL85s6LpZpkOcMBPBUcfn4ZD71BuR0B7T
s7hFe/ZqxKOdfuuQNdL5twd9iQwfTFaapF/6ug4LDF5puHnb/FEJ9XPgwHLA66z5hgkdeV8bhY0b
F5Lhri6/QlgsAzKYiVbireUZa9B+xdvnBfAaTU9OJ360YAa3YFDMdEsR75F6DTT5mE2sCUphWdOj
ahIFQroRrnsk0SU0xGtiLTgdBSPBtdDguiGmGAse0bmFYBt4jLm2uANwPQ9GD53iOCBHHe3/A7SQ
4jfwduQxlEZqKO78vbio33+9+Pp1H5mfQ/drpS1THaoE3YvebV/EHl25sn89Vfc0FsxqPpXpoyMc
EOn9EuhmaeTP8z+ROxzipqQ83Q3T/Io7b9Q51nmZGWBRpPcLGm53n2L95C+NeSGSt/RF3CvOjRDe
t17h43XcX5PSlpx5sjjOLGtszN7UA3M/P3zIH3zY0rLLFqnuq//gzGPey9kT6cank5ze0Owf+/tv
efzf3KRAmz9QbAdsNtWzOuKt1ZvNeXxOFsPoaHGu/H35y3fj6G0LC75EAk5wEGqZAyKYyd7oa6i1
puc3Jhy0acBygnFZpfI/K6cH+BVek4H6cPCb1PWsIWOAeoXhufWKegHjZVygVpaCqZPayX3T3KyO
UKXUIADyu1IQ84fHOuUdvHXgWK+QL/QtJzmpSmrt0yJs22pwdE/U8zgkgAIOAvJu0WrkTi8wBsd2
UB3gtEY2yh4Hz2XZ/8BLcm6FTWJrq/QIo0LEpBr27HLm2+6oX6MCJ3ccO3adfRQxL1oBSy03KB3p
YvhTfm4R7o7VfC79UNo2SsEXid8KbB18DZMdpRXt3IogwKVApMUOEEr81jU8EXgzEUpXs0CD+hjG
ctH6Lf6kYA/Eb3hDJ5qdqreiu1xn8uxT2lDQmXof7VSZXlfWIe4yCIvH/9dSFfz81tKu6gUM3ak6
aYuh5apdUoQe4s4RYi3CoG4nDOZfdaVGMUVsQmM1xmvwbpjJSmAm+l5QUdGsJCIfpFCqVADJ/Err
iXnITtIwQeFsissX+v44MBu1iR4i/v/E7DVFMq3T6kZ25zbN9E9yre0edX4EifeGxhhqaF9SuBXm
AGUdzD5VNU8LbKmXQXW43zs/sKoIRECSrlgNZjHD/2v4LpKW87ij7/klkM/qtUr/LI3UbUb5Qx74
xZHk+J53yAdpz+K0IYJH7ZB53LuvJVpsaHKkH5H4h9UNMrR4grvj2uUxvQPbodqqY9O62KXsw8EM
hUmjb9DflVnWZDXhHwSXUwLf7WhOoi/iPSUMvvWYLsPsrran/JmXB276aEeYHSt8mbj3JEi2r5IM
3UhRep+/V3/TWS75DtmQk8GoAdsRsLe/K+KTIbKJx2atbs1H9tWAuryYFzfU0okSIb0mSQevyk+i
TH18lvYF2nWuCxIWcObCrj0jOycbzglYUiuzgbZ5Tw8/HIDQd3L/+V/DGuCjUDbuOv+CRdn7wJix
1SZ14u5KKvY2FaqfnGAq+xQeetlKFCgoagApWbmDgL13ukrw1ja8PKoB3ROXBBR2GvO2MvPEtS3K
Wdcr+qLX4MDXRDSzCCzUSJM6ylRHWnbeuFp9DPF7PJuEYi4+2T4X+DukYhdC5SFvJpf6p+zyeSb6
p+dCql/+yK5WZebrJJfoNJZP2nPTBOgl7XEpwIe++W5DgDGAgb1zatoD4OYMcHrSNo3df2kGooKt
bz/mnaNSXSpAdNwmysidMf+wu19Hknq9xFKdpO0fzBGN/YUAHrYkocVUprPX4uhCdELEpQ+E9fx3
lqxVpQSSe3jKwVHQHq57yYcFIYmiKmNGQxGQKA+GNGd9peeMHjdK6bTTWLGhg61GvulRMxl2UfCD
I7OZxAlb8gjGDvZarYTROWK6y6WDIpDHS2J3OO5yo7eTdcamhOpJdA3N0xRfkI/tYoXXmEcwQ2ce
urjcl+F+/l4PC3rBXl/xBgfn811CTissdgqrHr5vERVKhVuYCpAsPxLP9w4DxO7b514czQXDPxqv
q8MQ9bWrDVpAfDrxj8eSr1nUWVL7s+VxHbpu1qQCMJ9CBYjKpNlqpCR1o3YGsJleZr8iARuBV8QG
hnxMU5rCamHEganNe4rLKFvvP1aMUEwnVayzbDrpwdCAma5IpHYhG6IQpG8UqL0zz6xsIcNci8sR
SAFqX+LzHAUF9wMrS/yGM8n2SkbiW3aIFI/CUw2s9xBqZFSfxXTVR0UHMHK2KRdmAPcUwze88Mdo
aVK6qZBX9WfH6/c//tEzrIOVTPnRPJwO4rt15E6u9uM468zi2LOIaQjepnhdLUfglpod2Y7T1rN3
kYCKd+zAoriq15w1RRygXQNzx4/mvPDo+eWz5BUUfbNqvz16adY474UjxR12c1ac1Z9/3A2tC8aa
MUE2+B3fFDTXjr9gkJrIU0F33WSmGdZxXQvbMCtHbl+MHUp61oA38PJ79HnLegXImescYe6XIswF
gHGcW3uSN2tmkn6eWGeY4Yxth69eLs3oJoe06bj8tUGs11CLkpgmQhc1VAVVnJVFXLRzLsai3c/F
D15y74s2ppOQud19Yw2wxTzn7f+n1iaO2Zqu54AArpfK7UWax1oatgHFMQxPXZ4ftt0JXytjVxtI
KaabihXJZMBkaCFeSLnjZMxAAULcpPizBnvVOUZQxuxKe4rqO4zFFAcNEtn/VEpai+4CNF3+JcJQ
0yyNCSPLaaN8pnSqqHiWO1BNGz/qhsr3OAuT7y5FH6Dgd2XVTLQBPa2fJiFEksiF6amiLXyZR/U7
AV//z9oX/4OGWTSNeXjNtCm6PTO/JLUhU9ytmvVIE0uOklbvqyEpmNqL1+Nq77t2ZyWdxrfl0W9h
38eHSRUjBEnOrjr9KzGCYixZj/Wx9McvUxyFICdcX4k8TjXIiD1MpejIXZfdRAjDsvk3SA5RdSEq
nocS6DPr7CQToaAHyuBBSFV1OF4zIuokZer7oXvA4mAzWh3sibDZYY3r351u/9Hu69GJUpE1IMlG
S6MmM3KD4ntjwZoNxgRhNfvYHeBDSnDXat8iqBTeN2zDCTJ7Xsf7TyV6ukyx2Kz9a35AZoFkI9Wx
8sBRY0XlHzXZ8AuVzT7I2tKUeCQcVAmcD8LW0KEaHcYuCgcih9B2PjT5YVDtTgF+8cfQqLrxgHsS
obyrCenuR3jNxGbK4IxaKH4vjHHm5nYU9bVHmyLkweu188oZeiZhw9cRFdDqSb7VVsyoOk8Fm5Jp
ZGMxIa/JWAYZXXCz1lESWaafoBHwtKskmp91TWjxhtdWApRfQ2d/kyle/MCZ4N98iIDy7Ut/SfGk
jI86TqR4nEKw4A/d1snedXzVVwE6ELhFei8OuNJAN34jvQkP6oHMR8yjMrRwYlDpvYOlDR3M7Q3v
7sq4dXlZb3AELm2TNe7n9xIHl/3XOs9KpkvKBErKae0MH24vSGhovdfYPwv3YgfSJR9BemTT3eZd
vflTxD+J4ICDi1/aWVhGWW0AQZLGoWHFIqmavzOQMT7OnHOgdDK8gfkxIwzt159RTlNvBosUtL0b
CedNoBgRAlyQg0OU8r/jbIcB5Jdddf2qRo8xYbksSxVadNofr4M+Hy52R3I52xzXc2/UhcDqcU9c
tU919xrCvaf4WPaGzkspbkaYqy/NcLkba2Rnnnp2zYcUu+tavk3SphM4NN+6UBpjCl+qYH55gpAt
39hbwl7ELgoKAPBksEfUNnG/R063bsDE62qhZ0AU9YX87MCEENarGrPiqtsO5tb3vgnuc0zAOrrw
L1XsdMfQQlXzdaD555Xo0LOzB9P5z7wkhDPVLp81F7ADCBd5xtoN66dojDHtcvT0nsDHXbvaJ3Yd
WVvitfcCPCHRZH6A46uOJC6UFWyo3cIgugb6W/2ABmaC4DHfDRHMtDNf1PIN554kw5Sa8rXfaU3Y
bEZJnRH7sB5ohAlFcp3LY9r/1YnE8EdNpVoWAI+ga7avWjQzbR1jzOJXBUVdBfHqgX/Ti5MAyQ0H
086MbS+wQpYggwEMf8UjQJQapHAvfU844PVK32HX/mnoOG9cR5+bL1VeAwJR+6PHbv0ZlxsjiURj
y7R4tubI3jOLuRX80NM1uDuIYTIGmNIvMm2l5DZ9MKUAJljPYQUuVI35G3uGsC3jGhVb02LUrP7J
YxZM1cly4bceiOha3LmIyRGSQFeOoiG+6zVytvBx+bL09471dW7qohk6HZufRN4JelG4QK0xk35J
u/5Jf4JIkHYd2FDnGR3HgEEXfzdQpqmCsGYC1tRGC2MQMheN8kUCkiqektunrnaz6qwwcXpJNAaR
j2UZukU47+zKusK/CAx+oe48hi1IEP8rkyZHshVAdIIrPZ72SF+kpqAbk+/E3OTzAQZLEkiSB0Hf
/Oo+cXkVi7PJ22Vy7vkcDxCoLi98Y76sAUHHTrFWfpeBCD8ve+AY7v9o/NISmNt/Ol0d6yGvW+6v
KQVA+TMpJi8hvcwZtHFf2W2gvbfroSPC4mpmblvtn6Qtdg1vFUCji9SQyKMo2B+AC/0OmTba2oOt
0B0FvOuOceXcG2jGldjrXGoTiq/pu9K7tz39JnKkE83o9Uy8SCxM/P3J/u2Vv5Htq1kKiN2mFEV3
Y4+sRaghsfaZ24/H+ppR6fnNxOTEdJeKT2svd2DyImk0LwCJ4NbMi/9P4DWgeu+FNW/L/MxKQ+u3
AiGABRBA4O9IyazJaYckmSJAP6GOUz8HJNQ7Tlz1h2boZ/HgOFBCwXnra1Ee2VpyUM7atG6P0GrY
gZQNd1Qo4masshBVC+LohiaQBc6qDggqNCXl1SrbnO/+qR1A2oWelHZpaCCFsIwMhh/atIUYUPIv
oucG9ejvnt5/j5Dhmu14oTUzxYoKzsn85QXpUbB5typ/AqsFNXXe4MjDb7tqy/2CaWPCqjp7CQja
xtmVUPJKMwhlpLUWgie1APGfPaaW99xu17jk2CIOM8TOcn1ttQb6Q0AmxRZzZq3yjbolUY/Shpik
lSvCLfkZszDnC9pjFwTuTbTG5jKYygX6X+id3X71+k/tdKrHbxnwz2GABHRYNCBrGPbHhCb3SDY1
A0G57z72KeQfRUx/9KonWzBRSAyHorUe8EH49TvINzE5fvEoVyiZI5JDvvhofXMGPyfJK4CN9QdB
4yTfnMobZpvoMI+0Xf9mBJuHV3Pxprs5umPSSnt/dQDnsRBYMi9c9hffqtEJLFZGmCX/aNxeinlV
OXGZVZg7o8BwPVKyb9ywKzJRyD+UNjwjDtG3gVVQUe+VhN1yzyuGn6ATdDm5ZGKP+CjZBYMsArPB
yeou7UanCLneqHYQsShDM9qEw270XfJS1aIwuVEpd1t0A30U0DGY5fSxy/uuY6ZjRZSqJmPhLlPl
RdnNIJVBVfGwevMsulhCDpVd7eBNK7cVBo06DRCteJ8YKo60giBcGDVoR9sHsWcxXkn9fpJYzKXi
foHXz4OKgt5abo20+kzcDEvmKGQ2artWr9OmT/xRveG9WQIyu5PZnMmtBwqRxpNJvsQRlTDpiUlS
5yhgBALvP5rEESpxwEvNu0SNZSGAQ8zoUoR/qSbVu7bl1iTTTFqVe6HZU7XHyj+oN2X6qD1Jkj4d
DDHNEdUqi7fbfR+VTiNuRkxA5HePsWVcg5+oCqnMMj89OZFPwosztCh478s4x6oEnE2oomIS17Yw
BFJFdd95KoORzoRhu6WNooVhWiNIbtEPSM0veeCJ9TtGUStsd8FLb7x7DesDUpoKwMLh8JrzYcZZ
8Kv8oWoA9S44y0Nxn/hClvAG5Jmtvkiw9R9/pyPpwkyPyX4bwWub316Z6Dbm8gv9o829OxbHJswo
KvRn3/h9D3gBFUU8LPP4Zo5z0fiCxiZu2yfnMhAnEainyR0W7D98fSWWdnPD54dAyjS0VXWuaZhP
i6Te8Fr0MDSeEdqbVzFnIngXn2ox+c8MTOYpX76X6G9KObRbEJWw2wyjLLkbq4MsAjAJuMEA8MXD
jGqoEbH3sXYC0SH9A95pjxHsi7VmIRfKbdJid52GWjP3LFnMB2UN2eMx+wIQhy8mib5cYtv5JnZE
5ps5W3VeFV5wtNSjF/9Lu1Ky9tfPcWNmzLL60WWbfV2Kpbs41IAx+aBOrUM/yPCCaKgVimQKhnmm
je6Do01KVl4zebCiuTauwnZFygo4dQ/AOOQ1wl/aK67lihZAMHFUY1vvczYaGdrub1eEdx3vmjun
nZbkYVIIMsHi1n4HQ0azpoS2WVNfqIR9SQsMAo5y46opGr0l2UvCUaG5LoelJVrbw4NsKUlnBPHa
1ti3qHk7XiCzIRxu3zag339nMmTXHAM3oPLv9pThnEdxOQFEKK1Yyq8Vpz/NKSjQ7C6FiVBnkrsX
g/M4RIAoSAsuLsBG5LrWEVBA+0z6o1IVhFTFuS9lcaky+5lsfikTeFRci8qTm//Nor4qMh2Eh1vS
oDqRc3tQXuMsZO8BYgiM2O2GB58wZN5EHtwgz+isOVJ+P1xJqGO/8Gt+1/L2NB6v00r43Hf5yO1v
6nxbMyOHsMVGt54hgIBA+KfMvjGOrmn5Wum3HP0HsrxflBoThsm171kyRPUOqpmjsSkZXQhzAaHy
XMh2PxzVui9hOWrS+0AB515mq08DLUN/XryheyIiQTySKnRK/Q4I2BBfdZ/w34nrytHIj4mxH9c6
twHrKi3rb4ib8zVy2sOTVOFkEk7c6Zxjn9J9UrBstiQ1BAw/JMIvQ4jqBIHSsTi1M27XdfRTE9XK
YeA+9a6zcyjRH+V50R53ICv04+xesSn513yQdn4nCNHAEYs1HcSMvZNWTYjgJI4oV4kRkPRuBqI/
wjvbAkHL4EaFl2PADE5JVR85YrXoh3XQgwrqr55wToIp+0Z3PQUqeU6GRrn5jozfYv1/JGmk80w3
8k8i/I4B+/h3BZGReaT8UHdedh5bV8CX94MFTVPOsk5uNk701b7t/I1MNTG22sGJCnlsIB2XoYet
TQ4LxsGcfu91MynxyGqmeFYRWeWADCZPwX0G7ucAFZhpIoVoid0vRfIDnjkCYNGnnLySr4pX64Wx
VUbwtrv8LsO8CkuYZcJ11kKDRxkz0OjXU9w35hzZ06Z2VZkXlQ1Vg1/DwnFZpBZjXsN0Dj34N1r0
f/DsHQwpMh9ssVAXXwPY8qhomDNY+3nt8FsbZctAPckvejttsfifO0NHbEC5Va3yrVuFe2k/Xauu
FBjkmIgppxml5qqtczLwcn540i8o6Uaki1PgNwiJz3VyPULAWg4Xngk0q/WrBfP5YgMwa0JnX+Os
rR6mov6OtohRM7wmYeKtRHSvRP2XLxdpKJeUYNKCIX+8IMxPJzNOM8VWe37GARmggnMoJlbsGGxa
VYbIEuTJ2qb3klFkJyJY1AAVs7KROVA8oID/KiQBQDKmWTjhISSLo9CXE9+zeMfLj1zgPcxtCMPo
jfOtlLZq8FDx+V/5RqNGDP48jQo6HC8FSquFaXsS7Sz8c0VpYDzGHLAysRBKniB/FdXCsZyvA8TA
BmrUhrDfOs1XsKWXKfub3kLNTwzbDqVKPSATrANMFhhHMj4ZF+jf4ovlndpckkD3jhP0kIdOTJ4s
d32el/1T/eq3BbOVUg+GRFnBfI8YBwfk7WmxeH2HKkJzoWIIKpz7H80VenD7548px9dL2rjlnFvP
J60oafQKW7bX9iFxvzmk+AwZRFiti6acuy5kiv8eEKmu2Q5bLAhCnnguHyHOY7hn1HoZJvgRN98i
Vkx90FI3g2UXYDuhqwC4lo+9apoIFiSX2mZ+brdrfdNZKpZWCe84H3WAD1kGnqVsrrrbAC/BsA+U
+lhSheORZFZy75XqO7xCc3QbaoOeLHbgQTtlf0LSjf5EEb58pMqhPDUfXgKr49nei2Yu4XbQe38z
LQStfykRiwvWHR0YoGzNtLlGi1CXV62rl0RQnhZGcJNn/oCjm9A4rSiDdsCbGxnvP9q+RMSijtzg
T9KobNpFyCBRECJhWGnD6nCefXjH466qNzAisNstNmi+7OkiVEHLdXMgVJUFctyEtZLceHTPkCSz
QDtd7CFeYUOv67MiBfOdL7giSfTyP5HpwvqsL5B4s4zMm87ijyN5owd8E2qZTJIEL/6Q3Fe3SwiR
HH+VUuev5jy++BbXwzmDNx2QnsBTYnur20zbIRBg5o6Ja3msoCONRsul7NDqSQjjK2inD2FvOkQu
HIuJSTtRag1seVJgR0e3F9NojAlYrrmxDzqWgITSos2/Tnqc70jP96ijl5n4TaemtYU0DSDJh1cY
P5aIqECILGIx5pDF35lCmzCLvixGSYdos7IkdPuFLUBa5cPijCxnVQEUhm81kfeqtsJyE2X7utas
8+MQDCRFIlMadlBn0VaOBrAen+S03dYefQXE8iDbUHKnEZi2+6LUJF5PN8YMJRCI9HMNAM3IfuRA
kHReHd22dNYB4VZAMugDv3/PmNreDtIuow/snDWZPzWZ796Y91NqukJgmHH3M6FQ0RiKx27466Uo
frD/qNC0uKhyiGGtvVfaYxLoKF4AhlkiwuQu++zbTpah9WHvXTLfNC1oS7FuHAnw0xiXHK5Hjtmk
RkEHWcb8J209dhhPzVGNahhjliixVyO2FNLTqJXwEz2jSysK0DnYyVhFR80q85vLuZyKXpH1VurE
ZRX6DMkX1DHFnkKFiT4mna4EzdiH1RQwDgIYa4cLkozncxDbaVbPw1JEAmTMkcAjdJ4NzkU7vurV
q70EHptEdhsUmzj9h8wPDFZeAG+qF9jfR1iWEAfjKez6NhCaDTdk62NNovNUGReWH5Oo6TifLnVg
LBfkK673taR6RHisdNvRD9aZxwl9MbM3+C4VvTDOLsd8g+IqEm+04BMI2NjYEo9COSu6qFgddvlp
EQ6jfDcPc2mbHdfCFbXS8UqILlcvG4C8zIWW/RpoqYfgg401MBybMhasyqOS3LjN982F3rsORMtf
VkgJdNUDXiuZ3/0EgmAsT/9Mn2UPJ15R0bmgHRC0EIAVV0EYiR7kqss0ryz96P7ImKVEc2YWS2Lm
6EYrI3eomx2J8E5HcXTC1pEt+G4WzjWJDWG9jQp940z/j5fCOBmLMm4YG7lISZDSG9Osm1MxxITL
LtY1/bITIYlwyGSFSsJt5bCM9iG33XxSjP4ACbS4x4x5H3h97qHC44o9cKTf/2fylUJ40/dbn3Dt
UHCbm5HVeyXcGuZTLVHEO4O7y6OH5HOtLvIu8z7mAAPGh6UNz+18arqyhxK8+pfOMgXwByrSFnSB
EcidiiiN+PhqfNRsob+/qlGTu/ZAGbnpWTOBx3EoQW5rF+yZV/hYA0Ybfwepg98riTCBv0E4gQ0n
NzR0xxtfEHPgKzXQdu4l5Dod1N5bJ9/uvjdymas62NwH5360NWMcOel/Tah9gc0RofHpsd8m2H/s
2BLZSza0jPlCZdzOK7/UyG3fn+pf3drxpUIrt5tmQD4GJKnBAXMcH9XV2br8QBXp6D1duhawLqzj
JpNV/+uNOJQP74bApJDb1RU1br1FXtxNz5m/C0L1zKeVm2KI8BJVgGLGF2dcqW4l/jYppQZQi2ZA
KvYldpTDIhsoHwHt5UkVm8lnBzLLMXnxfzL6qoWgHEmTfGcilyUVzsgRWkQni/CzGf27wnAfbgF9
H9mV8aL5dhbmrx+artXZqMzWGXQbyxjBxjDlEU+FPnIblhSVZ2q08/rnrTbted6gyOJtFN4j1xGt
iW5GsK5T+x+Qa6M6V8NsnYHoRC3fJM9KsYuoLDrgen7G3KSb7NGal/WOrA5N4rDLsdnu/K0xqV+1
+ib9b/PM90OeVfcCwM3NsZDjs9nx43fRtw2U5Cs0i0fIOAJ7NowgofdDzYlAENLj+xhQH8qucY1z
FXLz3b9Y2fSn8My8llmMAteCgnNIrHsNLLCF7H0rPNcDLNw6yQWm5pIreBPgVYXrmiinUBrS/BEP
wQnJzQvsOLMlaHWkbAzJ4LNZgVoqBb/AtyaBuPcB/JHCvBA5ETWO8rO626eakpgw8W7XCCpkSwHk
UZVTaJpYvP9qYqnwir8mO30dEUvcfQw0w0sfl21g+KUyxjzc5pLOujoDKJIFej23moRPfqRLmGeg
qVIJRKQOufUPyft/58yuC6GJWPfDt8s1M4KPGUlDismQKBuruGCdcivvAGJUrpRMzn0HbYK7aHFQ
bkc1Z3IgvbIMnd7oJ5LFJBLpSVkQmW0+8fV5hCO77IUt5hs7anauneESmFMIq78FM5FYGaOwtt3S
DjDsMx2/KOklgnSdd24bqZKfRyMWN4DhY5T9GAjZMr78rPmOFhX9ON4eM5dGsiavxZNxKXn/PkpX
X22jDnr/WNWuTOF40IRy/TjrPAuBObVqP6YipOYWCEWmnhUqH9l0sKGVHH2mUeumwJbL8ZJ/HFy0
tr0Oxi3zlXXMiaDdggkw3uGQK2aARoj88DLOvp6h6iTBCgW3gtQb5PRWC692TBoC/ZVspU+vnB02
K/NjTPD+tRVo6qzNOsp+JIBHmS9/bvH2y8Az9BpL2PI37zUWhDo9ZRuwZwflma2ZnRNkRbFqzD6q
++GjBwQPP028z5UVGPwfQqQ333n3bmypvwqTMylXQDZfhVsPcM64GfM1Ff1Ci/FNdOakRulbVOLJ
EFE+coyIybEsv7r7QYDQRoy1bXP9SSnkIFz/RUr+HHxsjlRfGIPRVls/LvAcMH/MZjIYyi4yCnMw
oluAGkMqQJ4LIcsDVkoMKsHvJTXsjPIG2VNeafo33O/aMczflOvT6J0OoGSfhIKXA7e0e+aWMgTg
6ttXW6t7jIZtvR8QAgC4LL8BkhmM0nUXwgKIlOQQdrmXgJhekIOrmJdYHSw9EAG/cIUanGbiikhn
oO/IN4GoxxTeKKB41rbqQHW8PyY9HwXtmvv0jonJvpQUPRdt785ZlLwPyn11bTHI/BeQ81Qv/fmP
9DsOQEBolGwl1F4v0ETSrlBs8RdpmeLj3RLD8qVqdpXKXrKEW9PvlDTon5R9C7nbEHwsQFRQ6nV3
03/bQVJH3XNQDLppp3oCshJ3VLNoOxvbXQnp5dRJeKDQGQdE4wmxFqgBydQ6AzoqN3az0TpM+cSf
tOne44BX6YH9tNtgT7lyTLTgYovoPlji3qUnmRDEz4Mx3nGqdo3rT3sJduFD7WmUwwTn8lkBtSD7
QZ1SOaEEFa+YHHV4tX+vbVxFS00HEKPxhk9eVdrewNBe+V/K13zxg07geJ/7biN5tJjHsSKPM2YW
rsbx95rRFb0STJ+M/8bE6IhYOTc6QFvPFG9YnCraJvImjgA1SjRZpq9CAyIG9mWOqc7BK8f65FSK
vmwUXixStMhP5L8jOQMLGyVLwi8uLt00JzLu/2uNK19Lo4v2wBsyFu7SiE0RZzcOxa84Rii/j7dJ
99GLYAC4p42sjhUs8d/F6P2NRQqD549PdQ/33eJ6PUhYgUmYakUy1URpp1IjQLvYvKIA3ZPSIvZl
6ZHBYKHoEE9aPrcZDhptzgOKqxwi3ZlEn99NvW7YQBxUE8WX4GyDtV8qoQjG5NJBJbic7vr6O7b6
qjEqlLZK0xpXbqeXk8yHX+Zr3fWSssosw2VLNt07sxGLgG1QpsnlOmiP47BTlt2ArotLJxkj3yAw
6DiSNALoIFcpkuwIJcOtVp9Im4pJ39lxCD7/MQpHtmlFidWoYA6xC57Do4TlCl0KWYviylDJqsO/
GziniJ0n1Geg0ZJl0xnZJbfxHUAEYinvndFrrSlWFTg0F2ZvrXoDIFi0ML9H/egDB6y5tEkkHWeM
fKXq1CmnCeddpVCt8Bfl4bM4+qfeevhu09Xs+45BOe5rkE87GRcc2MeD/9WdF+eoI5clD8Gcogae
4T6/dO7unB/KU4tcGB6jk0kX+UrYVtgGBiUUBURKO2A/0Tbpxe0imuM1EdA7ICrUuDvc13khagIC
96kX9L7LfbX6Iq03X5OgmqomzQkTvE8DGEJEe83A2ghLB9i/vqFgBAZiDWvGoXHkExlPbTlrtA+a
/YxBd/RMDGUzphXJnnGDQd4931HJ1G1gldi7AoGlYQoY1w91HfuvvgEMym+mqRekeCGlgCTigzRv
PAP0iFPYsowF7MI1RJuR/e5dsZPoI0we1jyhuCv9h7eGzQOJz98qbtK9ODQO27JFwPvH20+Iw84w
MuK3krfrY3b5KH0/VgZlA5BDw192DLG4z+zD08l6TejQHq2Oh2YL0acKLr07bjqlijUsV/RMu7SF
cG/VERtbX3POSCBVXxvXOXGIy6TcHQu9QPcFaCFAj2Ag1GIST2KAwWTLBIl3gxdaHaWc7H64eJeq
+ZRnxqZbnfIfVbe0YgeKDtvm+zezk9GDnyn+aj5VUZ2YBaNvRz73JlqwBmC6/0d2p19+VB0RoUO0
p7ilq4BP+xkKMhLgpP+2bXBTdSc7vLiBdP5zWP/j7c0kNtFBrXOHCqd22WEs/gO5aoQ5XDcyo5zU
7muHXvnsE5yjG8JNZlMrdBYzjkCDrxhXiOPqtoQ7WGYxON3K3jGe56o/jkhApH/yfoJ0P1VmRwxX
wkf1ksxwRd88qDdAbWN5TgevpWK8TC6uH4qxEJAIhqq05p8qBJUj00exFJh2CBTdB5rtQtlHWD44
tgogJNpAW4Xwl5c0Ac1AgM7Bre0DR+z1xkpwACcASg+ty/s0UQvcs4NOgNSnNFj3Y0i4EhWVNcvj
XMVYgb1T9+bg4PIO2hsxo4qkV+iAY77fhsQzFR0025vUEvM4/R+1tLYcO1Q9AUqsR4sQXe2xMTnc
z2miBQIRdlyJnbYi/1ux438e44uPKWyctWXN3BgEKgp1Q1nM6At7Eiu8zcJ6uOdyxcCljzhUKo/p
/qAm7hNDv5XfX0qszzEPJ3FbYcBE+IjtIu+U9B8lNlfPHGZUCIIui4xXC+GExVz/KSLvb1xKRxDn
37tdpGxf4o+o+mYHR92FEOf5xmBGX4qX+b1MTJcW8iEduigpjs4F8gdvt5t4GVUi5l6qr0Ph7vRk
fGjDxhzvECM3KC5db0B6GBy+k0WxikTryEjEvT5mCL3X9y5kx+sBZJDGitTmmnGvjow5/NP/s2GQ
yI37ZABI75W7sZjbOfWJ1MkN/mqwJ7eBEPeAposUXFrRQ0YAeJ1zZVPK+8zhDm3x8ObGfoFzIfwf
fGo11U1MJotzk0F6laYyR7hao/PhO1H6EcXoFRfot7o8JHb/WQbWl+421nc59ImqwCtnk3eOD+Nw
zZ4HSyLqCROhsvQ3M+7O1rjq3+uFPNR9QAwvyWqaOunsRPpH0t+LuNz0/RvXxfE8oJujcAGS/lWq
vO4y7jvH/6jHTxl9PuW+X4gTDyVVjnYskPRx8koYWVMxxrT8IIOVxNn5qA3pid7fgUA+dWF88fM0
7FDk3uYIU20cbYwW03ATS3FTyniHZinDFuqjBGi1rzCLJK/udAHNT2GOGGoKL6U1xKjbbbO8CGx7
3m6yJcD5LVtM+wXW1paLR/twPMrwFfzw3QgIyBKr6mYcPtoirpwEdV+erGX0746EuTmKdK/qK002
fgvBMntNmHCsp5VKOwPCUDgl9Zwe2JQaZ4iK9aLHUrmpp00neDqqC1zg2C3738dlXMjQjPcy6FUp
Eb9UbuOoaiiRk5C0WHp+MvAtWbLVKrGXQq0gE5dOdcMSkoTna59Q/ws0ZulAUAJdDObfKaelEotT
QYVF0G+EMm0pyaK5XY3/mbQYDroNF5DZhpeUX6/VtxAJvL+Or1+9isUYfkGHonQdzYlb7DdU+Bk+
7KWJaigxCsZC85nStKEu8cKKpLlNjXEn9U6mhMis+LHBrDxdLAsCunsl57zVT8P2rSwMhL56XDUI
9YIKAqnZpJuJYbIsn05fq3pXhhNYqAhWOddNE3yUFYAxDzmGxY9k94KQfG4IA3Lz66j6odfB6PpX
vpnLB2svUjvJ3vNivGWUv6rMqqFGLIQlB9RDOhaKUMkyLKIv14Yb8OeFDuhYXP/jwFKjLQVKRKSf
NBpIdD0EZthlEDQ0yPBLJ0dFTzou4otDk68ohUaaNtlh3fJhWWc90bZR+LXes4Aybj7k4DkM0ASz
NkFiRpuMKb+ANAhT1jMFPSzoFxxludSNFAdsZufJq9gsBWToqwICdmfbWWp7NHC8Ky5YZOUgLYDX
u3tKE5tYDpMUqkTUK+eDrUR5mA1sqgkXiRSDBZDgMqm2zTcTny91KW6+V4lNur411uUm+tlrH2yA
S3RUcNwwW/Y2d98ThUFzP+MqUJ3QRkbAUUmaDqICjSKMUVaprW8dV2awZoe+vjLMqTXwhTLhenm5
3IpOk4DR8tvv6sGD7ZxDLOUTTm90ogcF0OIzNELwElhbHeIhVzabJQIJyIvSv5UUONP8gxQi2Ad5
9AuDSAYx9yzXYuWrWn+QsvFzz+8Qvm6JSsBEB1fA7WtPOkkYIUWsbA3RTHRoa1pYRFhejSYnN2Rn
UyxA69SVitOLZIu5X53yEWncGoP8Mw+Bc4mwgvhuwYVIEd7uXaA6G9FcegOHF5eyPEZ7kZ0mnt1r
LcBUqMp5D/a3s/wlQkp/cwmtzEobtIVhBN/agdpd/Vzey577sXRH4s7+ADahcGA2Zaa8d7v2Zsbx
ugJagm98r9cj7bdAxXeiVzTj2PoRLkiomUqWLuv7gHXt+47uRgvSBYL8Gl/miHkbM6TuDJGPh4jO
mEaIfewZUDf1z708LjLzJXGqwtcatqo/fGsnHLvYUY4XcUNIuNrNrv46jLJZ3ZONZhszkQhHqirR
M4OwQBABl/9R2xyy3BfZTCTfpDRKvslcX18qXKpd7gTtJzb3sliJNBvKAVOUjTjm5m777UtBm84r
WPHgiWjfT+P/oNv0r35V82fbHPMJFSrFmXCIDAWcO6yRZZ1r2g8+XwbRsGllvl5ts/UV8/2oK+yB
F/vcA4GrEYG4xo7m0xu16c4P0z+T52rnRj5BgJdNEOJHBbJk34kIcjnQCyKxp4uH4KNRfS1Yv/kw
0Q2hyvfo+CT4/MRsu5TfIKTDj4AS+ma+iQbro5PG/lRhBkyM5YAbzPPbV16iTW9T7BzTEyTXeRI3
vvY6SvY9IQbgjCG9/uODu1loYsvewHYv+nUNHgycBuSq3vd7Jsqw57U+u+f/nZ+oUEDYQ/bD1RMH
4wOdl8+vBhhJl81ZTMSXEympkVPpg6JN5F/MomyPCwUul/h15+m6zQabLUqBKQBj8stP4eKK8HSG
o7MKs/B2WxOGXMX9hwKIwou+cIb5wVFrNn1iHKVh2o2jh7HLgXZIu3TpqyWFJfPhzr5yjb6txKa7
jmM9z0rbmH69isobByhbNcLwHXS6DVMFVgktEIs1OO/gmXoCIQqnJUV1PzPw1mnsKItH9zJExrZs
qmWSMMV1qOCGciPlqiMx9zMRZQ5FUka5QsBO+Iwunbycjeh6YRi7E/4wYEaSqfbWzNHIYNA0hTU7
mplmFlfTF9RIki6dy9yjem1FQMrCzwTkUwMM8si5tpcWaYo/4hFwoasUBlz/WcSwGz26kBo8/Fes
uExjXxDkcOjG3dqq0zsyyXpgVEDuxSMJUZ/YqWzw7r2NW9vXipvEw2pOUoJnfjNl233XS1Oz7cN6
s3qfXvLjt6p17EC0Q2pPinVrPhSYp3WoT23sfNtP8BnWb1ifU02RFA7MI2+L5zVhc23jivk32Pte
efJHtUT4zFwZ/AMtFOROnTa2YR9O2jMAe74rofuEQTVAgcujS4Q0d7PM9z9EAMDobS0MhArBR/0S
99zoyjqgxjYU3qB6ZjcujoPiUbAPYf/mRDcRpeKED3KxmJadfQMivaGzy1MFTzxkMwjU42klq3su
TIKIDNa0fRFfBib+FfdrMBMekI1BGe1g/j/BbhOiziEXCLs4lt3RqA393b0afY8xT+6n+JeY9PDy
BKBj2Gygpq06Uztk1Rm+cmC7C8AF2U7c8sT6LA13U6N5rHGNLPYOGPqHJyuWzFFI7GueWn3OVAXZ
uqfF4oudc6ohmdmfllIUmOnPxI+enhqKZOY5K5DZKpOWvpbdqY2jjkcB3NnZOFN9FcyPWRcON2hl
dBUfh+TTiFnDUHG5QiKzbztzkepSfg4/uYZ1uTQ13JgWtB6iFVjLb9G9gFoQPfZLEblfEgqaoBwn
paQVSwB95Idk0OsINszx0xHZJzpjzFwUhtvD1AKeXj7LY1I9TmuJehjD61euO0WkA60NM9qq80yQ
+eE236v9+ZUwAHAV/o3wV2u66nH1Eze7+I+oFsvlgz3PTd6w9KhX3HMmlqJ6Ey7eWdNyJxR2fw+j
7LvxlvS80tIiGCPFWyePSMKHrNTmS2dhz/OuiMJBC2w7GCRad7Y9U4RCYfM9q6yEBhJ6UoHzHqoV
TY5oqVkKQkZWBms0qb4E+rpX1ARlq95SCHymDOU8YncuO8fUz73N9Gp0XBZ5bIkNMJpiLeCoxk++
38OQWVyX8Nr8qEJLDEmmeATi9k2NCIMAYHG53UhNbU/5IleV/OTseBkz5brGI6n2q2EUD4D0y30P
3Bh9D/NNU8TaYGuDtqSu/lXSRI2u3zVZkPOqsHhHAkT3wVJ//FzU7uohHd0/ECox+T9kAbSLBe+8
cXxtvmfEMHrVbt6X7ley20Pypje44MBvS/snSPcnm6zqSa8YZmBNwwhq09QWHSa5g3C5SlFhvgQf
VcrNaAXgtdz4X8a9XvC+vHC2sMgma0pxTNe36QsEocU9WK8qU+8bpo5PGUsipmFRh4GLaDjWWzml
fB10/MZQ17TOMDc3Xbsv+GxuhFkqXT4cHB6NyESiOvHiRvsW+kPcO3n8FA7HG4Qr6ThvSFyiShcN
F33hxAxciU+C+KjO8rzwVc3mCF/DinlgJN3nUafA4ja4BkmTyMZW5oij9lAaHMyvnl7F9DPjgUqj
9E64dcBeQ73BZWggAo8Vr2ucMlVX13MD/AqXTyC7qENg2NvpOb4WcqoD5h11BFvPk78Cck7I5v5g
Sx4htmK53xGic6qOFOBhNrcw+APd1m6R6KG5c6KUJL2NGDdbMab5gc7Nq2Ytmsn5CQbSja8d2Dyq
ib9YZLt2jQYU9PlyDLr4otZGxhlzYZeqf5PzVX51+o71XTsiaFSit6kPwaJZTNknYBikYGG2ezqe
B2I6DxJ/g2oDbjFMZitbESjCu9OT99qzTeJguQgubvulMpsF4TlI+tF7Yre8VoVRbKDkPipBjNJk
Uw6gVR3U5SH36c5ah9dJShVOy98Sy2u0bjSw6ByXkIriJfOaVnPnzXKQbzxgjjw3BWLChsnfhK4i
uXsudoPQaDPAMIHllJRf4I79rGWOtSFSKFz5E8IOrYyNV3XJudghLByq5j600BCsxas24Bsuyf+J
3/CUpC2Lo3wAco/FQOISJj1WNyZkeYw44Tts5mBVqEuwDlkEvdNURJvuDJYY9NhUScigzn27m/xY
jV8zGjF1dOg4Ur/iFaJJLoSzigIQYRnDv/b65x2TSCrV1Kccy7nNuD91CyMgVkIgcmYJVLMf9v4B
s7vlrN7h5cvzH1tXcR9UsrNkhKnxUZWAgxZscP9rP4t/PsUiRBSZp19Psv7HDh6nvENlY8+biNVN
Oqt2eUnGwW5usVEZiuEhyqDVLYhKcahqcwRMjyrFeTZq9Q4wBT3UBbed91CAVDhmRK/d0MX8UMC0
DdSPV6uXe6+UnwVNSdi3O4tlKTbF7fTBk+46eMqJzCNkC3rQGsTLxzf72Ad6zf6GbdCcl6uX8Z00
j14T1ZGNOBnUOKWnzc+GZApkRuEiGN7c/eS9L6e3KDPLzXqFoAngnl3cBaClPoiKcWFRGy72Q9UL
57Hb9togB05+5JlV4ODTKxYCef+jrTvaph59XhpHs2yH/by4xejIvTMqsn1+xmw/RmUZpWlVYrSG
5zxM3QUbV5Ax0ZuBmBXSVcKsBKRb6PKkTr7PqUNmHH3BE6fCvgur/2EqFZiCtI5ZpaFEyrAAiIba
DK7hmjgRkJtuphOJALYhUt3DGRPVVXRe0C7MHGuvPRr2Rt4TYtehVxDiUYUGVFZzrBoQOlrpRoUE
K2dHcO6tBK9QAJz6mOOnBl1JetSZ+GWw8Vs2Lm8DOHa8axmHAHMd+wmWiuitX7BBSgWAEqv8axXO
V7/iDi27I/vd2sPlxLdllGBVC5pq6qXnZ3JU+sMn3oYZORaOlz2+KKtYTcv+zyNNhqtVuKhviSDF
z21OizAjc4HMERVOPOFTHkrfGUV/LDC5kjU4lEv6kl23W58IOKK9XVJOuZLRLA036iaCp+MYrWjQ
Ei0ZMuUVuPRS7hHcDstrBSEHBwN31rpbswoNYBqPNrH+/Wkah6IA1s+hquWC7zNLQEmEAO0bPMcB
2qm7Fm0WQaZai6CI3jeUnrNgxYZDB7fy3JIlEuILh0Uj9hOOTuKQuIsheYCUp7v+XG3d5JExgWI9
SI05WZanre6nCok2b+ii7N1fX+7e/amJqQm4rojdthupDy2pqKaakek8NsLer+XhEg4VjKFQkvyV
k1S/Vu+iOLxJzY9r2dXwxgGNZSRwY4YvbHdqOZqz+knKMRsYk+aGZiXA8VWn0CXGkK4h4sUKymdb
85EX9llvN7EhCfpYC1qmvCQxAKk6PsNLZgfAZYI6X6fd1dqZvhAb/c1cSeKAd45rZV0EGhZtCTW3
zVSiNr26r0OshJXaSOfb2YN+b2vt8dFH2tWj/dUfo3yMwi1R7VQRDQEZ3oM6sI0Hihr5x5Ug3dT+
09jz8X/26zTxbw/1J/oaEv14ZJvx09SqhgqM61wmXLqkRAF2MV3P2vY0TRRj+vfsmgctE6LGWuyM
+IKpShffdEEw4V/DZEtA0xoMtAJS5cwD4Xk3Pbeizd81VUzRuoSATGdrHbVjBINxyvphcBgB+B6L
6SZuo0VOcJab6Y7iS+X9mw63LiNpr9MBpfSbtajSDtNBX9OgsWUAoz6Ql4BvlbqX+IXwv81lSUP6
fdUMQFpFYrmbQIXqszT+m8kSIxw1qU7Q80D3PL1Zf5mzjmGwkPP9w1DUdYK33whGnYZJgOK/wPL2
4AjFcc8nUPe/JuuIzeo/K5e7/tVn+FPSw+wcv3Zn9S/1VSGvsi211JqayrXmrsnc318RbWUKX8uT
KUXI6+sT8br4tTu8PArdWzvj4FdlcDVRTqASszlGwk97bZFtXIiEiCRyA338W4EXcIoNNnlgbMtr
OnHaD7dLVRBPfarOR/CCJHIo/Jdoh8zj2lyY5xYlDJqSQJvDLyhdTzn8TV9Kzg7xUNgA+WboRN01
V5F7hmuHf5KZBocT8QExSGraahLgZg5tXYQS0IUF0qmvKouFEB/+1mfXtPZkMAdxuN4Sxmdob5uL
pBxtxZl0cqG2WxIrhSDrNLXfsw0ya6fQXXpZ4tWduuafxrJzUunCXnRuqxRQNS1gj4DermEx9Kdx
R+yM0XrwE0Z3JA3G4MxZGWrUqbTixM3XlXKG7bws+Co+BUOIOQ2IqxEez4iVdUsieuXK0Rl1mmzj
zPg+v4GJovDVzF5M/OCC+IQKsMM44PyXhhg89xb8+Kyclr5md6qzEHZNHEmW1h1EkiFWrx+AdWPW
tUoYNMbu/oYqBKsQzk4Zh7dCTwMwYRxs0oMKe1bP4PY58QoY6nsYzslOxTj9JGNuaKAw8K9EBZMf
XwVUEs0iTL59bMwGhNUooDOwVWrcNokV3bnua8rGbJbMMNZjJC5x2R9l3Az7TNeu6ZLWdEQuRhBe
E0/PT8WooDUdqaSck09sUKjFqatIHHPHVtth4tl6ziJAfUSqtHscm5U7sMeuHAs89byhHNEbtcls
SOiVfR0Ip0/nskwtOP721tsH57uh1VcqLMdsSp77y+Qt/xmX2Y3+IMOxeQr48yN2e9wXoMCpSVm9
aWeZL4Z51QeIlfLaehPM7dJmAjMg6GS1SToWuKnofrc8BXUnpXpQJ/vvZ59QZpN8yv2az1RBIGBj
vcgOKcmD3ep2nd5KssJ68641xzR/Rug5k6jxVkmfJliOFSzS1rBZJrqvHVa0//Om8+LcjmfVlbbQ
fPaQV7rOZsziwtGLddg3TE9GYdwXz2jqGUynmTxi0i7JiYrUgCYdnl1yaPupphP5yMpUveFLY+Xz
/b9SXEUOP1qkF/EzyRz6OD4n0IvPRocLdzQA80HKZxDg78dV72xWEjajxefRQyS8n5Z5KIiW7rSw
QerF+7rV5E4hlT/4yZhupSnHtUSXUiLU1R81FkmH5EcRtBHBJPhfxrHZUBp7+c3BVxVN2isVFXJM
ju1cGeWyEe6IKQuSbuvMS4Ph9/ixqECrOKuNWKE3G23z68yAMhk2visoa7dCKq4qB6ttvpOwOnlW
7wz5bw9BeynAo+Xf1i63HmY/su/+/D1b1gHbh35sAG/Lr5f7Mn9yta0rO3STbTW4jb/5J59wSC3N
go0ZH4MtSklTGCk574QlcrAJ2XxGAYW/OgTXCCg2lvJ25wCb1rtdUVbJNqsW/XYB0IfopR+3Q+WC
LmltoxMbjxYb2fIc2nMOcPO1eLn4J/1uv+98Ip/lFXOK7pI9BkeE18VFlXPzRHG+F/Dbe4mVg094
PmsUI7WEt/6TJLASRsuZApJDCkpna3o5f3fuScn+X6J23Z/K0ezqvBQxfHslssNatVG6ZNVqpkVI
/jBc2MKjGiBoZjiKR+Eyq4ZA6IbagsAM0VQM2d7Mf6uXyFYKqazz3CBLuVRLA9zA8R6EooklFGry
572fKnVpU2hB6pxFod899MubXDWbg9dSteIDb8l7CxRRn192KIlyWaMekyeB9/RTmKJtSA6ZH256
IKqNW5p3EKfKI3j1iq2rHB9FZueH9U2f69jtJN6BoucrOWOwlNMorLmNZsNUOqwklYzjxW8/GUvY
S6XLbYhnm6wbUT6TrcZd0c1wyfPHfXL/L+uL0JBfr5BTv+D+rVdfCSslQZ8MW9K7rLRGuexNxLmc
wHRFIPgEHajiK8dQxOtGtjFFj73AbVdXvuR84uGLZCEPfDd/0Nprq7LVx6yWzFa9u5eiU0VQJIIB
5h6FFUf5EGEv4qHoNTDuL5XOfdwsHYd/krFuRmErGBstbcut46do1Soc7sHXllm0oBfkmFUdK4l8
xzIWazXa3Yl+re3sWZeLf3NukDo/ecEUGX0j7AhvQrHSDtBAF9HnHqAwFef6hbhjyoAoNxnkVzSc
p2X0Sz3j3ICDy5aAFD/ZdIfUCzeAgDC2I9DffJJMp0UsUk3KpEiBrn/jFXeLvJIlnSHwYxIF8SQI
7tn5obliakEr5bOP/Ln40TjE4hY/m4bZUutmFIUkvV762WGYnzpcpW+Nxu9Rah8dDT1eQNkSA3Gw
xECImUOynmRxowLjLYEuoz8KfkWkVbIu3R+01CqSz9HDq5UbYC0tCAdk5ArEQYm1pfyo3ODRhbqj
vQqgrzizlSaJYOkUEE0mJKl0CoazrdOBfx8yXdZdbgOzmubIQhbUq4ExRMiwr3jyo1iypFONMLp4
aQtGFoD6gK0woivZwY65VnXYKw8cCmwCuc2vXdJcSQwFIqeUxrBpkGlX7YefYFYM7DSvZTrfvTTR
pfMFbM4d94kf+GYICwCGUybQNpNy+j9f87B0gRBoSm5gj9pNlA4bEwhpIOzWaO7NCcRa55nsSk/e
lvmy0lkhYRZ1s/bIbWDp7tK+6d77t/8O34mYgoG3SWzCv13wmUIER48/IefMjb2iX2bgjAXFikSc
u/d9Ct3Ujymud3mvfQi1ev31jodzn0zd1dZCqJqqnYtAOZzJE0fgkLhyYrRWuYqPraz0RG8myFgT
SsGzMKqrGid1CKNmZIVvn2lD9z+n16GEeLhF9daXJ59i2ONXZ8kdb3xhNRe9wNNuju2787ocCxc9
AVWzVztAWdxnVYKRI91UsOFWB1vUazzFGizhIFp5xrr1n29Rldfs6OArPOLIqEG+13ZeGXJSV6+V
8If3sK5Mww2U51WfbrmvFAmy49bZDDDfiR4BHH5vNA4DkKEUl1LFJ569mEaBtH+5/gs3VzpOCH/i
bMV2Qlw3ArK89P0nPWhKVgGAMW1q07ucuNqbsocRUd+dOYgaB7RCek8m50LNk+AhB6IzTmyFvlR4
pRGanAVruFqH9dVwD0QL3MWOq/75KLuodynMDUt8GJuVoSs15+wTt9/d0QCiYxn8Ys40kW5jeGS2
b1Mcdl7M54UfY5aBb5R3FnlxwHmLHF66yjyVCOC1+Bp0bnHnneUcwy9vmERgOexHMkVPzce6pAHp
m93t5zS2SgOzF8n2OlR8XXzrO3qyOALKV4zDmePOulN3exm3Zr05nQ8LJT7fxIBdotMTPbZ8VnbQ
dLZJczjUkjZjUJ0+7fo8cD2IGjC5Uz4Wdgafl2Dp7plsGHkAQ4wYDROyzUUHZk1xzGR0tgi6IY/F
q5Ten3tpODOcmHW/2SEoqk8pmMhgmItHPLlp4qWWXxYcEZCgsWFucdDJavp1HOw1qNVlGKGhrD92
4O4nfQ0P864itEsASCMZF7agoJQmoBNZgDM6F8EUK0MAdMAXPJ5uMOVAVJ8pauujiBFegpYvN833
zxac8QJJak5Vr/GeLwv+NaI/hY91vTQeyJ8JFqcZ5s3yyuIk+O3ct901oKCyEPLC49bXi7jsrIm5
h5tNBqOGRyvu13RHezr2HwxIKCLHzTF7BzkEZ+0JuKUakEQLx+SjnxKCfps6/kr00MaOK8jwdpub
KH6KOyQjTheZhZtlc1GbijMH2MJg8ysCkOImFTd2EWdC7FI0JCpgYj1taR4Cr+2dlzaup6vAT9fP
wC/AH1Kq2O1oQd6VPsTwXahm5xqLR3TCNNpEKXjVdJQIYCWPzAW6YAZqSXwIYk3KNO1OlQ8w8k1Y
QiimaH1m6oVTDK0Zxky4mm4gzHlXLjWYze8J9R7MIhP5+tqmNz661NYQJI5ITpkE1BDKgwx3rbrM
9pYabzKzt6DsNn7AwrNcML5yJ9+HS8lI/77YqpdRTDfEvYsWGjMuoISj5yp0+IbhnVmUTGxPfvJW
Kfyjg371YXSOavris9V3CgcIcxsd3l29RoSZi+H43fdtiXl6grviF40D3rd1hBwF/+jElWGItjFA
ksfGh5L3OxNYA8bSBeHB7NcPeaqE0JKb0w5zC9Uo2PnpUhHS/cOB4QqEZ9tQndG0YTCcONS56A2S
l1TbuS+FaKUP0wMd0cl4ThD+IebloLcFfuujKWWge8EN9mQgSnfyfK1o5nYSoW1KEabwL0cAyHMN
7OWxbGpv8GA4stbibMNNVnWNBEG5JUyj++iNoUOKxgtkQFiJykURIcGnJI+vPColnmXjQedKsOOh
NNgg5pORWPSU5Vknm7aQI3XemApbWBZu38wTbUBez7us6jWGFtM3c850Qlm9r8VEuKj4GnxmFTgd
wq+GjPmlOx6TqHUFLa5O6kKJ2tqBfFC4mezygqjpgS/kDQk9n1c7fhuAy1k2fVAl7WmqIhV+4nyE
mwlYJ+DkuTO/mm/S+Yn3dfUvfNBTXAeK+tvt8xRp4SCEEfiY1ePc1Zh6eUTgjf5y5rrh5LyJXfkS
VxaqG9ITQcjts7slpdXA7K8qjz1wO1f06qI9WGuC97EdYeTJX5w6qREi9TtZ8NvaRiGwC5JD87Bv
3rmlfmR45OrSQnsTQy2Qb7o/VWoA+49rX4YiLCQtftomBG/6docp8uLmKrqdJI1OtKWcmY7il99/
AtUUdVtfZquusQ==
`protect end_protected

