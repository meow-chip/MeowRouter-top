

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
oYYUZ0MeKqJUJoI7DJiuvSB+q5Ix+Iwj9N3EwG3d9aznfrZuw1+Fc2PVy4cVNiksbh9EhD023m7N
/1rZI7UBsA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BmgMGlUziZwp4Aeom40PM0gFb+Lk4HIg7NJ8Ke6/iR/nzJgqwxvBOYZHlsOO/Hp8XOgAeNb9Zd4o
mPFcvStSgKrLqxBJrTC4jOtTOOUVOGECik9X7RElVDiKeZuCTuuYfKks1rnTANMNKsXOPeJj6Svr
YyXA9D2NRP6YkUNuPRY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
1jtnTjcMZBAylJ3gewlkrSdkM4rrC/SF7w+2Gpl8C9SK/D8Tzq+D0qrZVMnmX2MWMKbqqYu6bkIj
sy7Xox+kttnLUyhBRsrBNs6gr3T0xsxsJ7Gnyco/P3Bde80gstdJ+PNfjg9uJOXa0R4ym9WtfNGf
swawtPDRNO3XB4oPqX/YBORxc12Z2+Xzlc5kJQDf1WM1UoKUm0j7+JBzjmig2WrmokL853BM29jT
4Ht91JL1B2bOy9A+fEpZnVLxL5NzuQ9svrSJluHfL94vaMxePXlPq6InH4B+XQp0TAFlIitjElNz
4mBAF7U6zb9GPz8ite7f9+Ofg2sCbTc7qhRaHA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gQeqr96ZiBT2MmGHCpbhB9Ma/ONapmaS0FJH16GFlg7E/VRDUjqbqiiC9oovpVsOBnNDQZNmXNgv
dI/YoLxA/mPd3NXizDTj33SvvwJdHC+sPFJrC6pT5rNUHqY3WkLW4EktYj3xtwACazlM0R3H+N1W
ZL2jtTv4hCIZZw83DISHIwGMevxP0unAXWFpAlJTyOmzC5wsjnlwvjA6I18++KC1ECVIFCC+grSL
XEAA1xdZCU131f12m2UaGi1yGaQH3scoEe37TXsoGUkWCMAn3jD7PddNt1X5zhoSRxPsOfUDmtSO
kCNVtrnPznMY8kVS/SdMToJlnwH2sKbHJZ6YoQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aYbz66wynlNa4RYsWnE11uoqAUkMOGD1rK3oC0qHnHAmOdMhPdz4cV/CAQENwbN3ryQY7/k4qEBR
2l3bOqYxA0+CBRl+jt8CXXxWU8WE2qwf32lPVes4/pVAbKANmE02/Ysj4IR7MGLvUvtr934XOsBK
cCc/KqvEbWgnnzkEdl16nzyz9Je6iY7Ni836+/z9BA/OYPszoNI5lKgO/06ni9esrcL9aCuvKXjM
Vplsu70i86fjOGURYjM2YFmCk8Xng1M6ROF+0KD+TufNMvK1W5if6MPJr/BsB83OF/hzcDKyULpB
p2+Eliq8StuhC0n7jUXEo6ZGATEY2a8DWEYVhQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
B8e2xR5DNyjb6SEEOPCOnfB9/yUC8O8izWpzVz5s4/hfcHkvr1SHS13gqMQDj1DN3uSpaoGxcSIv
a3uLHDL4nIDztAAEPOvl5rp/eCLKhGUauWJKGzgIaInIPCBXw0hsptiyzlIicQEO3rsxoS+LR4e9
ltN4asLfvR5i5+Aru5E=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o08P3wLx4KXr1Q02DiaLH2vPxf0H1jXIwF3rbwsiMxYgYGWIJGF4/mxUFC7J/WeIjcsQFoTUns3o
ZlNZWWRR36HJ1r2GmZoMunV8HAWjNjCUrk6RBWvB/4dYllizQVzRhb+3YUjmiSEMr4rkGsWsR9/t
W+i6luLQskwMDbMnn7puINFUehSDaOzDytgvFigNs9cj7haJi7XjPeMPUBa/JbbTJGFnxz8xzl03
55+BSHF5m9JHUn2eN7uDkExSgYolpcYI1EQnoCH8U6Zfcweg7A+n5SfklkTKUeWInYHoz9tHbIHA
y9aJwNoT7f6uxEt4GVf7oKjEfFlxUe/yajXHuw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 132672)
`protect data_block
/Bqfza+AKUAUEZjfatwXaX5t1IU7wnAEtG8gOmFQCufXzDlsqm+nYnFqa/EWW5E2lHoeoKa2VeMB
OVvenCbCMf8J8ES8IjFiuoGurovIGECg4OluRhSbPnClLPnnLZwni6Ykl+uFlFjQxVaqiP9X6u2u
zAVlUtuJArxVpVIfvm84VkuSxBkVzRg89N/JF2OBwflxaLOf1ZU/5A4b0JENlolqIOIjTjzvWdBJ
4ltMqfoaSPjGyNpWaUJcV0s2JzJl1cWPU9/U//dhYP3V1f1SovPj31lcFS8kRlphMcYtZWRseRvv
mWq0qmSAZJGRnu0AqVeodgXBZSnGoyB+GeA4UiPN2dGSksELF0BriNLpAnJ34N6bNgNxuJ65XzHQ
fqNc4dZv5qPROASA4Xr8smBjW/q+8yZ3W/31CGw2SQXCsvc65ReKo8gejhFolXeJb2B4LL3nnc99
rSzRm692Yj/mcQKwVM765D3fuzW/DDHYIiH1l/972lVZ62g2Ttb2TwQzsPJBjLh5g5nmqfbY95sn
Fok2/TkyPnnjwuFR3iP16jMLiORIAMx7DzPurhu5uEVQIxjU3MM0XoqINtkc6PBkBcoI8WX/TvBt
Ci3h1h8B7V7k3SL3Fg3Wlr66FjDTdPRY/UNBjTI2VqZ6nPBcD6ki0Dd2fBd3lLemYZ6h4ANg0JAq
I72R8r2EKJqpNO5uLjGxXByH1fostHYMrKjjcm3GvrVP2Dowd2TBIYCGH/IO+BWrsDmWIueJcHCL
Co6CZ09PI3+pb5B/584xHR1FsI6lcKXZUigAZiLDp4Qri/aKt/luTrtsAdS5XXTJxIVYxIH47pOo
sCSlfLQpF2QnG3dGiSBDHnv+aEFIxpwCc4rYmHwEyWiMpChlYRW0gRYtdk9sIAR2jNkc8ZJ/sp6U
X//90bieBO5gfQyCtoDQJpOlIqatzGHNIVj8OB8Lg1Y9T1+/aTpIl0rRsEyFBJ9dK5/Qtg91XIOJ
4K5QrdkfmPfUzlNiC4exOSFLIZ0RjobuJRSUFHX9oEOzbcUluPc/GBF7t9p4AMrGLAFc6F/WAchg
gP+9IgE47louJ0M2xX/JnTFWuXzdX+FXXg1xnfCbCpMJXflnYwVovNge/Kcq/7lK4y9ugrNcnFJ6
1FoETQa75oqb2ScUffE1BZlPPRTw6W2FdApJ9Rv6ajHvRVTyojEqtKGoDT6XvJCxPzbhJQvP+HvT
2P01YmPNmZNzvl446r7SUmNVD5KShM1cVikQv47kYRZHL0YkvQ/84UUeXEVN/lNs+P+Ps+pYJtVT
d6AGiC2J+dghip7u93xmS5Zu3fNHBa7+wEvjv3RDcmV0tGFMHSJ73nIh/jvZ2IayBUtWMO2bVz+F
7rvVCs6DSAalY8KaRvOwreJhRNmvqxxlMUFt219QC2JVF8q02zfkKvNTApCky0Lkt8qX/Wl+CyFh
oZlpUiLWKkhi/N0iDSzJRp9EuEtbMCkgqCCkXbB5Zv+tpBkrumeQChTPjr3WOa0fJlq2idQC3fvr
TxeC+IsKXa3fCp0BvXImCLX4+yQV6Lx4lxZb4X0A7YuIZ5OyPpHAzr1mvWkCbaWsA2CrIvVnqgJS
51eXNcW+JdLR2kuaeZltr6eHSrUQM6dMMvkl93+qVGs2tGZLlZdg5pF4bShRsyq8zStWqD6e+TcO
OcctTFxpebBW1QjiBerapR0tqMwiowgkcTA0RfZzHGdWQq2DL6F5U8Wy6GedMArxIEy9tXMlZxH6
wDfXkRHPTTvqMPQX7Qy/oJyVe75vr06d3kKx4+evDtJYDrHbCdAl7oLKyu+ARukPep7nNH/YMvsd
as7Xr3e7nJ77uQrOmdpC+YHquvEI8/6s9n6pSmc0ZgbbIxkGfxVfO4T+wEuF76zL7LfkwbGdee+R
u6jhENmMMlry0+b6ynkWebiQdifOdTdSUnf5/He/X9T4cQLGD6aro4NdchtNXlsxv7S6FEQuaLd7
tEuRcOni5owAxm42AN/JsL/Cu06FBI7nvXmIJIVaOdWDjJSf/HRpAF2U3RDRahzZgrPKWSI6wQxu
T05hnu6SGZWDxSE/JX+oXmIl2sYnjVKWaWQsrXpe8yJLWbhUsJGg2bKXYiXDj0CKe9sJKaf8IGM3
x6Z5+xaOUkx870FQEABOLcaBIJDQZ7+jUbdkEBCYTHG7cZkxe5+IczkgCxhnYe75f0tY0hgX0le5
H2YqmBJ6wPtudsprWDuGe9LhP3gD4bO0/6PO7pFrwdS4CDjR3jzuxvkDaRB9tspdGuWpuy9wQnOB
RoGBJH9lPNCI0jMe9pA7LjevoQWNM9AIN42AzbEPuBtZ48IJANa68DKBaxYnnrY8mmvxKhy5wA1C
7Cmxfq8EQ2DiR7/y22eKJWogEaFRjPsjdaA+u5hjdHqy9kklvZK63af/tc/ke4hl7h3D53yfjtn4
NcjbA74uvXYHvKGbBydhvKeiMVmQsspCM7ptYlhoXxm2GppGEIIUHBPr2KxWGlXqvpnziQ1U6zIG
fU0xXKazwmXAACWxHq4H83jlNcnw8OjJcCBSXT6lMI4gMa+lpFRIevluCn/umIbSfpLv7QBe1sjW
NHJrC9Uue5RVMyYjFH7JiQ+MD2Q6GlOms6tBj+Cl0c0TAQ0kl8RAU03Whhdxyfi7GQ47hEQ7wt0z
/asb447tw6gkBaYbxiN6NM8+GZA4lqqJ07dpvY/dbNfwQLcAxsWNsAyj+ZDOPYUrFxNdQ1otcPvw
LeQyOHxuET/814BgGPH0fVnLqb3pxNz34aMeW1zNvGRZRrR+5WJ40jxKp9hG3Kem+Z7yXc3QnPx7
DIwKBOTtnoIjpPw1SR3QmKh4s6PqcKv5k1E/9M0f5e1JdwhzoIkwTCDBOJ+B4BG7qHhVFIinc2AK
RCBc8D2a0qYWT/nkJtJMA1VvXpjLcX78RlAryst1fosOCosj+cj2dzZVSuXoo0YJFpVSO9yq6osr
gfUMxbSifvqjdyx/1kNAmRehHD2u8K1Zo15guX7MfJeIwczFiX4NNaAFdVz3T98ZXwnX5PbyiwMu
yu1q2uqxsRb9eTNwhGLWabxcevEuD/wLzW4ppPNBGP+12UwXVH7RA5LkdY3nYTwITFN8xwBB3z4Z
shiJJImyzFlekdFEgOpqL+t1oBZ9DjKf7GXX7UuAZHCgck6stWE4OGtT58O0UaqilUQVwUN1kBWY
Ld09Tq8DN3zkwdJqruEx6VtRF8v3kfLcnoVT7JiaXnouLgzOWSnIooPO81CD9N0/BPxJGy9mJ++N
+AVE9A3ReZOsfSYt0H9uIJ+MoCD24huJsa/runMxaLN/cCMOa2Pn4iKtW8dpFIU1sO9Z9pmeaB2H
B1F86gJdt1c8mKSWQ8Ac0lZqdclbL8SbcB971vKD4KlP8V4XosuM37mitfw4MhHS5Oz5CRUnm+uG
yuDQRIM8TQ4lmVY7GTrN+sA27BuzqpzC9u1y6OG4tUWHY9fqcnhOYeC+nLpj3wAoQGtvd4LtmPrf
+xCoX9I4TOX9FNShPEKnkKOaJ0OClv0wLqj/iAH7vnYtYvdxztkQpDvnqYgTuTWm2G0O6uX9odCN
t0hexN8/U0VC2zMT23NhZXhCbwkCEqDXaQV2jhMKg9+PWSd3+6l2ZGybhjgYqkrQXp5clN+cnfoQ
icQTVXUrYQ2+H1vgri4WEMPQze9JMsb00RLRWaO53sHLilydtSJF/DXZQgkxBE0dwLEBSOq5QRQ2
HbKUkeZ3J6222P4DepcW2Ct3rNchv7pRpbLDiovNIoLQibyVuDlQ1bpUAHs7Rl6mG77qm7dkh78Y
Da7KHeMjhUO4vLagrqvKI6GDKuqrknclKCH+i69uGYv4JNjtDPxbEdw6Qrmjq4uA9gYWu8oTqsQe
vkiFHWF/Q88JHwoV+ldCqJSnBvJfrt6o6haE3+LAfSaLwe1ge/Fx+nF6BvQRbMnR1ozCHNBprXUo
f2AOQiJ/eUYwoJBoTj3t/KOfjtbpDV655uDLCkGJtNy7CHyzW/f2ilFPpra5n8QP7YfrWbUH8YBx
LEx5q7LzHYO6P+/xEOMiQQM6Ax9EZQNBi98hr4ifvTDUJrUVscUWLfOBWHbDN9pYqTIYW13uoUXT
P4dvd8kROlLH1cE5bosmD5qbGJip6y3y2FJdu2k7QOJSDFumYxUzkoU0vZPEad9LzCmqrv2Mw6Jy
M0Avfz3aGYbNITkeTdxYttAAvuoHN2+9C00nMupurDymI5mNl6VQcUi4TLVEiFw1EKZZq1Ybn8GJ
koJbfXpC1MbpI5xSGsOApdc+v64FotwVaHq43mVEofu3ccL7n+/jhO1y5sjtz/Q7b+adzhRIo4yw
WiJtF8nTnGa+OEXnuamaNBBuPZOmbStXUVMvhMdX5miIasF4IskgSAwdP2cbQZjdFQ36D5dB5mf/
w/lvBIYgkjuuwpVU6ylZU8o+TECmocE0Nm2N0MPzjYcu8mtgKqlzHblc0Qwmikib4KMsBwgZJRtW
QiDdjyOVXPkcMDwMdFb0JqryPlBAQlf2TA1KUj3GgoE2nwLY2XGdyUlP5ujBdWgpB64cLp7Tcwcy
NmrT54Ug40lQfcGt+aUWdF9kaXJxXqus27awUEVLfXC6G7Jei0Rrxv3RPBXX1IjPQZxgdZqEcdQv
aGoNdbZXiA6VMoiiQGhj9dis/VY0842pERhOjKEIMadXPQ1Qfd7n/j2Avmg670SJVYquN89K7LCY
H+VCO0C6jmTcIliRc3HzkSi45JV0CSNYtBFw/JjCSchLsZxEUqYYzKPrRsiAGFKy011njdYp9n+I
NY+LETjhk9S/pt0aNzxTj9AUDHvQeb7t2o2UW+QCBSm5QlsqSK2oa9vvguMI5PuFhac/qNAjN23J
86zsZETCGD6zKgmlAz652Z4uddON4u4FThJ4HOdK1Vdb+RURQaR9x4WJ96sAiD6uEp/n39XBez8I
y8s5aMkxJMK4R+CQywWFRp3d2adHmQlVKL2Qid9HniA8lbmbUyg3xOm7J8IhqEzK9odYJcLaHx9u
BjxLsfyl37tggLl+MA3gOzRpFDjZ+4tqXMpWgj/h3Asd5oE5K1uzU9zF5T3Dm9CS3g1HEencMbYs
pd8tXoQMd7EC1ubpkTuKTqRFpwlaP1RogqHUI47cjxjwFdMoya4C//hT7vJcBm41UHbwEWpbzYFc
CyLYt8DdHtwiQTCDl/08DyaaAcSMv9zoi2WV5l4OCj4WeId03a1hZbl3rIPAaAj5kSgJF5MpIyJE
naLr0uHCqgOOuAT38IwGHiGVRvcsS/Tsp6YkY54YUA25ippDMW20xtrCzSH7QTuIDrwGy4swabhg
Adic3tB9fbXUYZ+Zb+xCdNADywLTpAuPQ4fEap/8EA2+jcWn3jKGcGvGaCV6iOepXZ8CLwBYJsfk
3/sXhlWoT3VuJU3G/VuPiKkLwPBGjO/hzkHbhfsvv3nE6J9cnsTGh7FTqYAU7XKqkRoM4pnp/xwo
hJqSWrT2Mg/NcbM0CrzF/L8L8t605peUjY6zN4UHP5lDGynKQUDlCoRdjVM0EUTMKQCyu0HabKnl
z9Nel5TC17n4/GCtQfoAnFHtSAigwQW+KFihKh57zFWYe4L12vPdE1ksCQ6wX1kkQgbfaJ3kjolN
BPqyMWd2YdnHcvtCEIUW4CKTSIYS4C13ZV/jUZWABjTZYxAW+wbHwfcvq4y205VS+MTkgjN0Nk6b
WFRtAlrBDjyoJeVN3Pb8EoobzsfhcN7MeSdg0ftBkWa0CcL8kUi4o4voDQOwC1jzPpboBZrRGx5w
Fxchz3Vc+erkF0rB4kZ+NHFYfVJ6/C00qYVZPtdHPziveZXRxJx8TZcIK96I42hbclBYp4Y4Sm65
0qsoLQSgWF0uvE2mwbCVsACYh7Bb6z0GkVdVNOfaN8dTNv+sBP+HUkBOqqPwcJ9PAZ1irdVrUhhG
NG9i+9VyFppytnEuEARvdZQhvhkMNVFCk/NHpY/f4adn+1SQbuKoDJQf7NatjoqH1jpaVN/FXmav
jrmn1+Haa/c5m+N2lPpFaDJe1iVot8vx1hI+wJ2Z8lF8Kl1JkYBrc4HBuax5Q1mOCDhhIVgxIUKQ
Co1AX5zn6dpVVNAkFLyf9XDVhBmJc84s+iQzRDOWE0nA1dPXpsHtzHcNUflu2FtFFLGFB9xK0mvg
2FVXVHj7wuchpfecaqMo6BgBycgn2cUvBKkTfcjqaJ3Mh4kCTLk/ns8qivZRHsCSPCnAAckx6aNq
MhDumt3g/iTgKSQ0gsSY4ulfnU5wC45Gttp+GwB3M7JBbT/MfLo9l9iexWcJHWL6Aovp7fP0j6tP
cyJFetSRCjQNpeNvMXGxWSn22mZ6q/Ih6E/wvWkFnweEoELIdUH/sUTWl2ZkX+FzuE8lM5Kik8JN
L+MHe31S/UFbfwegowWEpxvGKzK2h0Ajl80+hf5pEFPzrTNfmfdFCRcbntJf1odnGTmHSQc1Rpkh
0Jxnh12xBmcZ6wmCr36MRwRrw97Dr3H5JopizmeyalaN6sx3cIuhgHm0R9v1JHKNkFWShNMLC5XC
Y1nN8dLvNfpINEPyz6DNHnpr6WXq/ugd8fdskmR/2AP3R7jq0PpnCTxXZKuK/hexAhL3Iyd3bPue
h3oN2ny+IUlhc6K5SBzJtyE4S5CFl2LiecTBiN3RaWfLHkSTEYoB6ct7Z3kUTQ1t+hk1mwK3+wTT
o7lOgKhVakCDE2BOuVsenEAhJH0u7E5doH8qQyLHKr4EkrMfekNfn8GLN/su7f2Br4Srn3bzLlDc
M9ygpXUPqNe/hCf4p8Ui9PbKta8IwAO+9LW8QE8KnLaIDnv4i9/1LEMnhltkAUZiVB5xgJ3QviOL
fwOVFqskHvdPT2BfAmsrfUX6VuwihLOm/Sg1G1AW6HNP0Xo8aE3fszQ8Ci45heyuTdzWQYx1aYvf
/uJrvijJ/D4on9nnFrMbERVeoD8MpBJaB4w4xbM5KVfha1LaOkBGzss4AERkKpeWaplh2gZuGJgG
ZC0aPno8/swDqZMrXdUGbF2xCK81gx7eQcdf2a5pD8myBsQRTM21JEWEuFrT1HD5Nk5WKpIwE1zl
eRy5XTZ0L+UTj2H3aNFciKfzQZi1cPByIrup8asARdhUz6oesEnQN3T6/hPuZa3r3IJktaHZ+h7v
lq05Vp+ROZR0iGKA220ekrnIQ4de7Z853GRGtIlGD7pTCfbGop6tgqOh6zaY5fBMGCMOs1wtrgJt
0/yNm2DQHfRWOB+8VaREadT06mQphXEpYwQm64m5o1XjudK3qNhShQXS4Sy1IErjRyePne/TGhrK
9pDmtAELva0ezhZ14SmLAa5Nzb92U+wgTjpplFuSFt3k2xfIPB/B5c8txIYjqUE4JWAJlMIb0ZoE
8xg9rEOfmLLzQzN0pLOS8EFWJ9LZjikKj5cs1LWH2JMlHeoOzkHYaU7u6yMGNe/fK++DLVJcVp1l
eYFpHtoWCCf8wIbLrJEw65QSt/BZ61HRD59HwAwPWA1d2tF5MmsgTIHDzzlzS9pKzIJe/zd3N9NM
JDBKJvrZmF0BLmr9HlkYV8D0DAQ7PGMNovjMCsODtUSsvP4rHVl2Z6tfntr7iE7zQEiqgXC85pCr
alD08HllKdL4/H6bg5YxeiXvAIrGU1qQ8hAZQ6+EEnYKi6dOGk6yu69TbEWNy0gKdw4joOAxayNv
P6pY0Nl64XkHxcj/9HWUfMcZgvoLgAbL2NHEfd+wiEeWuZOK9GQ50PnqwxUsFSff7QYY6hLk8mFy
sVhrwxjLaulIbLE1vp7kRHohaJQ9Rr6Z1Ef69AG/jku4A6dx8qIJoT2a6yuQEFOnEy+SfcLGAzwt
3dVU578ZYSOF6ElLjrap8XaxTmvh574yTW4pN7nk/h+2YxBMaPFoakEINHY+D607hEhSeAM2xAdI
VE3wU77tadkEqOgpJ7RwUBElYq0vF03B3SeUxBdiYQmQKNbeTQVKvEp8Qce6cYEQlZckTuPL0MLi
+iv2KekGTseMpXlN2PvdCwyGed6dVi/9t2Fjil4UKNywxyIdkLwmvdzhfoyvBcyNTA/B5/deuOFP
xgTZ3WlgJAn0jmxhdmUaCDdjsamIZHafmrNROxGFaTzhR525O1cjG6DjNy3tovB47NiSd4fO6uxV
5e07aFxjkSobZWy65qwXc5lessCdxnwiSZMAr0EjVriD3uZR/4U7ZXUD7cvpPRzF/ORP/eZDU5BD
rw4NL/j4nrUVjZauu++6YocjqvdXaih+jr3z6sxh2/AfkPOXoRKwAYibq0d0DebW7kmy6UvXCk8y
fQUAHXTQMkOOZi6G20Q7ylzsWRm2n+GFkTQ8MhuwVJLlyFJPXPvypNCwvIXI5NietIhF5CkaGGzO
so4Qrh8VamC+tKU3YMLedILTX2CbTusZW3A5QmvkKZijpV4vOz2H7JkGy0EqvJJkwIFrx5fnI4Gf
GZGZomv2pTIfxIx4UftXyU7jGDUSz1QzGrnawvgf5DIcKaBlxT2OOwtuo+UaL0OiOVIb//sOLI72
SPZ+6x3B0b7gJX9FrmsXESayUusCM+lckWRGemFouFjexN20sGAGtfI5eE+HKnq5M6zY8MasgqC+
Zj5tuYnan9y4Hz+5y9GB3lPzksKIcInPJ6UkWdMzfILTAwcktk+tDCMITTATewTlgLrQdZio0xCb
fTJzsn2FW0kov0IiUu7x6zS61ioFQqfEInEmE7Z1qRepq1JXyEVakeXZyOjADgRsIqaRj2qw82qz
zsuczPI7tyQNnO0SrV+30hGAjwKByqE+k5K9GW8dRyWEFspKC9f8FxdI9CaOYWJ6fAAszepvLpFm
ozR9VcyEXN6lJOT24YmrnzeW2NKuJV57l/yk0sdvYiBE6LgL+WFXg2Jd+5wrFnkSgCp0mnrPQJ/y
wizHpjCyb5OKcuJKCZyARUWIhM053i+M2+uxY80Kosp0EXZPu+5swL1TMaPfCViWzWKPkCWNdIsA
e4vyUYBGKnjwefDYv2EgdzRi6UxOShqjziskz+5Zmx/1rSXk91ksClWWpUV64gFng6ECoLX3blKQ
+PaWjHt/b5Avs2KQtYSejLDJl6AsgLZNjjo/7V+dvIrb8t8NXc+DU+SwGU/k9+apOkaHIeiysH6n
1V//mv9EfoW6dcXAjxdX9oQIUd3laOxN/9p0bwWlClJQ5r6wOto2OUCnRQAbs+JO3WUuxHokbHr2
AfBxCWtRS6CA4qlKMDnbeXB/h0F02WLJ9Baf8RjsEqIv383wpD6ZzAMTWRwo0BMkW3NlnhTM4eVk
vOG/nvXtGOcVabl97NfJIuCWX9GSMjyG+TpC8l9jKXGITaUDJ/sCr6pN5Ra7+k7OnG0TDC6pRN6y
+3teJl9eWyZD57LYN+CS2WptjV0KZUFiOqoFlz7+y1VvP+kA0oWZo2ZCAJzPuPuCjzLo9W8uIFso
/x0lKPCCNB+yhfRcPMyzOt6jqh6+BOl6uGmAuQ5C30UcKt8+ZIqmrk69FyWSrhtkcIz0O9zTAyCZ
tdpNsUjubUf1TIU7GDQ/l18JVT3a+i5N55b3g0rg/lWmBc+Pva6HR7xsDVgVmPISr1u+Y+z5uiZe
mCzn2gyV+eYw0gwXFmdqE7E5VSG4XcFkLTGcCGaQt6iwv5U13Tohm4f+FywC+QXhHvO46EYpGR2J
uPt5Wu3xOOpZfnPv23nZoJUpLrDc6576B11o0MzUqAUX4mKj4bLa2WK92vGx30yvIimALUEBCcce
SH7FxheTmz9fjTvx1Z4WrzVWfA48gMqoDXvx8rwBxnqElmGpUzzgW3Ngm9UhaNZRaXL4nC91IzvH
RFgyFijQicYGoxCTDFkun0q4FSFjZjqul/HLf20kCJSZAhjBoFX70oF1jM7Me2XH/1EcoPbJYLbI
ukLuILA+ubOKm0PE9Y20Y66OdNqDxpuqlvV5Jz0difRnFOi+qbY6hAx6M3RgwC3ODjltKAHz6sxw
SNGVvY0NWXc1S6x57nfn99KdQ2THNVycjUDHiZ7ubdlEC9TM/y/sP4VTEFdXaAfM+BELz0jEduvl
ygHjGC1erUeK1DFvD8YtBUxkPSAiUBwy9by01XvmZg8g4a0C+Qv4sO+NjPC2lmXN7pOxCgrTOlXR
VnoOtFR/lIPn2vepjFSycpE2mmdJQoKT1dc74Pig4nUmHKAPlLDYKPl0AsupQrBr0k6ONy5yMqLf
RBfbfZpDQNV3NSDrg0ZmT0RHKazwsUOzyxAqtSRlmZZWynT8hh+24xshGgDA4JIgf8hSq/RO4Kgc
9grI2x4iCalzO78YNvL4+E3ojCAsUa67rYCeHWfHPbORWOAFmIDd1cyg4jUtqU1wk4IpPGxHirfI
xXFIX0egCN/6bozSQawCY7LRVCmEP+l0OVbIrr0hS1FwUzj57ElwrdTt46t77L/EbM7mtghIRy9+
5YEaAufeZ5g1SdEdn5oqXaFflXrTZoil01sSbEdQQL+LW9OW5FpzxcuWsCsa9LWk0o9EFfDTiLbX
Xv5hBuK+kZQATy1XTc/FqopC2a/CidkgwLHJbQntrXNHoYh6IF+7Ziw6UzHXK0Fzbsxpo0sUlBz+
+GnJD0I+lyLyOjuWnfcasMXlZvHnkeih09Z2iAfmunqCdoAy8Z27b2529CWMJ66s6cfZEYoVdI13
JBZG3dvZMQpL8NyFqvZEmA6Afu6TUw2Ak1WZEjmeIyTVeh/1g11ak7R7bUmHHX6cLaY5FF5X1dq7
KYr9YJEedya8EXW3Lt/dXAOiL65mCunnz04SLOyCV3R0niMO4dKrmKAOvR940qOTp5oHJ40h0iKZ
6VtlBCaoFMRQ8wgXl4FhSYpsldOAsRXyl4h/BcKqC8aYBInln4aDG0pSpj2Mi9j42N0jWw9oto4P
yf9p3E91awBVyT9d49HaI4MkWIp8RY+dZHqLExKYF4ZJvSSlFy7hqefDE6voVSBsAsr1LAk4ywBl
9kHuxQgzT+yIEPUFPW4zHF7fVGe0IjF1oS7D3W857UvR59RLob1pyv+1j/ypKUEBcCocUR2L6BpZ
9JJbmUkZiJwtVOrKd4aCZ2j7Xm8Mi3BqpdP/Z2XkC+nFpFzdMaY2OouoeAVpgbvKXgBiYuBqvDfE
pVMizwDUyoD/imYunzI6KGxIb3X+yo1gpvLmmqgW8gcdxG+cFjjASPbk8bUqvGTCaLnGKwPJeZjX
pLDrNH+rP9urVm9dctiYUnZvbnnq9zcdXYmRLkMOXhbmMmlQX4fTSrP1u3Sp64OhjiU5LCgj6jGR
JtVJzyxnyoswzGlsAMcDtNmI5J45TxKX65GM9Ii61qIIQUDKjoHxlY+RF++qXplL68TEuuHLIGvE
iElqQGxS/SzcjWDBY8fgnJPKuutUKmsEHXKCkphEHFaaQbYM1aJprqqIznSDElWwXUP9Giw+NgdA
OPNObSNIZV+QEiUld5GsDoYf/PeJ4xsNQUPQSTeth9dk1YBNNe+6Y4n9jrOd94RWr3yJVL2iPIL5
j9/KV2qawLM7VHRxTUG3IHDcK9BNVW5iW/PVcbTmrLyHNIOGeyU+H4N+pXDt5gMyl3RyG++GqFqW
B6nnjj9S8XIaWZau63Zt3Y34CUg68iX/xytPisPgOFja8SE+hw/aLxqPE/PfSiZefiGgKe0nEMvY
655NEo2PAcx4HK1fAhEa/kpd/fOPQNWDBowr7Kb51niDW0VO3McM9MdCjtyJATEa0d6wY8h7lb+k
AGYXX2u9jrnmkXasd90oh3LlKXkDxhUliKJxeBuQh9qAPxjuHOq7f5kkJeoxeHoe1xAqbYv3enta
GOToZ6wmDXh0lGtfX94DR7H009D5kMSWn5QiwobSh6FOVg0vNnmljm66LGyJFDyAFMRoGpdM9l9g
fm/Aa7ktYFZAfBnO8lhu1hjIGEflSFMI+aGEc4sAOj1WvKLAsVi+IZkUhep9lhXwZdOOIuBXuW1C
/sjMUMEVARKyl1xxuPl+QrF4dHWa1qamNAs5wxuCvPykgCo2wMesX519UIJhpJm/vKzO+DXU72g7
zG/YC4cI76Wg2scNWWYeEcH7pe1tdBCMgH8BBRSOvnT5DSHjxDWQ247WFGxG/v7qmWoj1kEaij6Q
iu6/dgySUWwEaruGWxQ8jaFDLa+pNTMN2zsVnQt3BFeEmCV94cC8Ud/cYT5gvBNchMk0icE59LN+
fi2srkPRgi2lxDc42ucF4SEd1NLvJFOfo5FVQszAcfxhAVHOXcXIyMTJ1TJghq+x9T9ebTjaprVe
6QZMO6AwWdsV1ebJxSW8giQ3WILbPvqPYl932W3pjDE1auuhj+VgXXILkTTSFduCMuSS9fNzRlCd
F3dBba18bQDsgqrT3YOSxl/YBTesxPlvle5NBRH98gzG8yzsbOk3MBrBnP2oGV5X82jn5KPYcA00
JOWr+UnMrk4b8xJY1Xn03twoUn83I9fxHq1fuZlTDSrAotfbjGAn/oYcA5MHFPyM6mKcH7tmG24G
hxbmagw4SjY9DNS+Xu25DeBHyc1lix9GEBahnvQEud5+PTpStEP86vWgSOvODvQ7cZgwlikF478a
IsfAevnYvncKVNJGp0rEyhiipEpJz4rEJa3oZE/Y29GOakq1zrflZxmQ02KGbR8Xd+VPyo3sObKs
n0pma45sjceDnPQDxl2K6kLTv+X5Bq073n12d45nzT0PCTyHevAUHlZEzduTP7wKCRkj0YcU7GNU
IDeQ9ED4C4ej5Bbt1NzkwH6ns8bhkwbq43zu4e4lCaKqECJePu+wsbUyodt2FEJxG8n8uhA4SKcZ
gGy6niSa7OCnvZzYCgtabNDHGicuDD30QQmKHODozUtGcg/vzqqOcSsYZ2gqZdBXErFVUoAp6vmh
IaiY28ucRxLlD1Wo9d8FNrKvsTrUSLIyq6yORJME7lj9dmDbvO5wuWR/hGW5yim/Cn/rwE/R3iiD
Wg3wiDNJrhD4vaJFm0zY6Gcn0ZeEB4SFj/zkYMyvXSTPQ0bx+7pHoIMbiW8ZW9F3grOdiu/Gayrk
7SY4MIA1hE5K6D/cClp/fMyrIh6HgpNq86bBhp03gqvsX26nMufI1GK+K66y60c4qwSTkdBjIHOC
tx5mLfwLONo0oOLEqY+h1XE/TUeZDRT1ZlmabjWhKI6oZc7VtYRiJEiNVxq5rbmFsIP6pGgtK035
0RqL2DPCC2SMY6EOw6I+8mrygjfYRw6OxiwSwvVbBX4sl7UxRq+OpLzfDGbS/h/VXND9AgHHMoIw
lO77JLydCNAq0KLtjrYgaYnEbTWwEa9WehKQ8AiC/sA5tdKJ29eRHLEdafUQSDYObpYBwwRfz+PH
HrELcfUh5lKxvFCIk7ewPGe0CcTwIkh2S5gd+gmj+zxEYRyLQNwjaEazxKqoo0xJ2DDJcH1bFMk+
rJDyuwYJHS4Pk6/6zNoSiG1lI0au5ILBj3YUv15pSYf6sw6InNTOQirr1uTVB7vdTC2eJ47wJIeH
S93xTRi3qf9bYu6FQHVQ6kQaKrbe4850el3NcITiFRtFZpQzCvnflkBTuMOC/nor+ukdZCK/5LWV
wg50ztRKcGAoLA0iSqhqTx4F15Z7NBdgUTLMokl1zKSk6mQavYux/EWpel2zJMXhnb8lN8pRWfgd
9jp8D7WivOZb9avZBbDMdBFu/pY+mjuc8YWh71gdUMKA+UK9qhJF7PLsgX5EXZAd3NHdNtu68mRm
UWTpLpjEO7N0JI9ttNhAnZOPufRUIRJgHWFxAA8ZZdq/96DurFMICL14Z0l0ersAK+XIa0xl1sJi
t6vJfnhm3yeBCaA+sRCNoJ7fOsMEab1KXBr7Suc+KKs65Q7mDooiXyyASLbl1yCUcUn0fiD7EHC5
W37Ta/HJv7Zz8uJlWIwR/kbpmXla08viXmk02oqm4jV+/JQYkzKcwSi7lLmdaGSVMfykTVoZ2BY6
tCP+fcsP0v2ZNtVr5RCw9mO89JSagG+4qLh0WI8VWpB6Lm7WmeTbI864NBuxpbWYHIgSf/SirFaI
mNBktG7W0RpvYs0lJ/MrRxDxKOe6rkn+7fwhweZ6CnUaqzgHFz/d8QVgIEYfpPLGGSYwpc5k6gTa
hCqt2o81yGEnZv5Bh/ot1BEv0o0B4wwIXsdD4AEGRjrVk650DXzGwCbSk1cqR2IwET7VoWk8D+ix
oqwt64+69foug/PtVaMTFY98wPgcgwwBEul6gh5vUJRyRArnDyBP9PgSfuGwj5Wxc6RmfnC7fjdz
KE8wh4+/gi3CITj6DDhK70l/4lqlgVHu6HLFujhmdSluZalNuZnSdiebuoz7SZMNNpzqJ0IMok52
nDIXr7CN/h4MiQlirMyCz1LPQOGQRwHwOc2QZFaYABHwVIbWsm/tT8tl8G4yCOzhu4b1HcaSLyWf
lLqmSfFtgT8GKu9Kqicydr3jSTrBOtJnLnsicHqSFmA9X5ZArlHtZNksfSR+1/P3JNoWQoPahk7j
t4soZdmnNEuhk9SrWApj2NMhvj1DQpnfwKjLs0IcKP5h07zWNYX69gDwJACSWtXV3xY10BPiJCX8
UXdEAUP5A4MwzBOvnjU427CWJOVtR2mQsFBeCoek1xARvKlmeFpl8PLchZBa2/WRTHRCcq1EKk5m
9VTi4a/ua/RBV3Q5bxWSjol3vFbqBe7AVcmfkzA2oMeuqjA1JVAK/1mFSBKbxkkhsSuX4hjK6CqW
SIQM4L7ypk7ySXVQI8f0qe5zG1C/e5iuKcGPzn5JG95/fmo3EcTbgPaoplfqHvKUMMF0eqW+U0fB
E5osM+D79kBiRz55H1Il+q6UsBlhNb9p/OWl8FTq8Xt6yRBLlyUC+iISiNTmX/13k9Rv+H81ptRT
JhJeZe3JjpF8FqWjhA9MrEG+q1r1gMk90rdkoSxqawNZ510XkhNsulU5yq13Q+39KG+SoG7dCJAx
Pb8kFRP8UJ5dRUxcJc+FiE0CWON+mZNPz7TQr3Xo/3vd/f8DYlJep7Y/x6tbOdZSyWhRXRe1Y+bu
0brmtmQNbr5ikRbpetF/kTjOyqKE2sgU+peEx3aaEPYmrVDoyDksedbCg22MS3WR9TnF+duPExwz
wltQXksNa6liFW4O4h6/Jo4qNjQB6CfkqNwXaw+oaXJxabtleOItIaMlYGkQIC4oJqqKGEC65qgT
MEuMbRqinb77gkrrrJ85BLzTETFcayfXahnNWQ68Q+ck2J1wpdPP5fUAS0CIMXANNewdXBpZzAfU
J/4GUhQk1NV0vHE+icnwkZuZdO2Omvj25YgmNHUsFBdETZEaNRMcptpJOiF9l8YlFokq5DB27Qb2
15+l2S9X9BLLwVAeJsKNyf5kg0smMuVHxyp/o3zkRWloTcJvkwUL2hLTBDQwqB15+tJILCbyIL9B
N5BBR6r2RmqTmGsMqgPd+ojlUjwWF9p39+shSyqxbn9y1eAyUDNwkJvOdzIYlCFi49EGvtWAt10Y
cjNXTV18Qf0Q/DO4+FlOJwNdH5JCpR0FA9mqR7U/hSKirXSuOcUBqob8xuPCw/Qy4jfyS5Tr3e12
cXfcJW/iD3DEf57pN/G2wHc84N5IzebB5cv6OgAC8g0ifIcAnBhnRFSncXZPtS88MSwyfeKOkv96
BrqqBPNznH38pvrwqnvJaz3cMrnAg4T6HdjX5xsCGGUjFUw32j6v3bK8RkYDcJpny/GtbXps809n
W34nu/DBcD0IyXr1mefUJ2g72JwxalZpOdKXbwl3VjISVg+XxLR8X2JExQw6Htg2zRz13+OXhERy
bpDr6XqPACu6qLzWQYCFSuXzl1hQ0DITo5kZiZRYiPoYJ4lfNHiWUP6qnJNpTeI1B2DnlU0rkznk
YbiKlLblM/6LadwkgxjUMkemYTlF5+TtVZHJoejyUpe6Y2NZ1lxSQ7AT1WTuAwcjdmpJht/QnyMh
nhEZEdOxto3fC4pKhDuQdw5uyneezyFpegdwLYl7tTPAOXLk5v4BgA83NRVHnV4PUGHtGbyd/xO2
TyToeHZxchFast5QkyuoHMZa24RMi0TPylksK2Dhh99JfePU/zbmx5Ff0SsH/EhJ6/uXxDW/lVWJ
raW0eS2aEkdTFGfhPz9H/ADVUdhurgNhLssLrRAi9MJ/e1vb1BQMw3mdtpP+hc/A+5EQhGaHWqpN
Bn5TaR+BhEahKx0w/A4UAOzbp3n59ZqWSOhXLOmhu5jxZTbQdOn3VZFDzhjuNSZj4kXbtVXniXH2
d00onfPTs44c1uQ5cKHahwb3iRBfoZWb0q9UfAIpY+2HUcHO+zyZjRFhKU7GedaNulKk2sp0Ni3v
LUmq7gy5V2RYksdhut+EMQnKK7lvU2nZe70y2MaDwJ0RvLdJHzfwHmfwcRSekc2zTZEwotfI9HM7
UnTnrAQEfOKrDHHJQD8/3VN6/yRKtkvIUkjwepTFj2kFvwOO2O0C3LTQrs0BnUilfugpgUVmjCAI
kBQu1pIcjvNtthuuKwA5/NV5Nvf3YubPmuIcCAC6k8EqYun0ApdVhrKkQgkf0eyStS5NZrQ5QtxS
Ri8uWCnaGdQtbo1NKnjJ7RxcPrpDkD7oGnLFjSgIyzyZfXz2OuVeoAC7/nL2CpZFq4fC/VcdJ/TW
pEQIfpFRr/IkYVRR14FTQJRma1DMPM3r2rYbiopi1koFSeYK1UvZzP87DTbAeN5QGVjblFrNB/Yf
Oz2roYShQKOGiaF5NX/ZhGsjI+W17jTxg2MlxxEoiEm0pnYoLWT7ezz6nx8xzrJmdm2zs1ckR9tV
gkC8dkvlzQvHEf4R7dKjnn1ylG2Iuo4XSMfX1A7j0Dw3iQV/LOTsjFwzX6TojE6BrjFZGLmxtfrs
RTbOJNToasUgxRAusVB3lLWUZeE33ua4pqwGbhKjnc40gA4S6L93sQFzl78zSku4Cyjw5Br+bqWZ
nkYiEoUmJPeMIJy+datfGlY4GGVyVjJhyLKv7c+vGQmenSeu7J7eXTbYWs4OqYZ2XWQ2FAKrp4SF
5THjYkW36xNSKEx1wEB48+tqqm1Sq0PH1c/S5JR56hM0Aq5gyHcVWctUxqtL65qKNpxzXtU2Znnb
mmPrgdquY3WzjdBBcK1Y7f6TB0D7fQXttnRS1Ky09dujFQv09VFYBVEfTFp53GZmuvY+f82moy6Y
xkVIvXu03vBcKjKQp9f/YK0aToAjkO+E05F3f9tm7FJdC4KpVOIrVanYJ4NEh7BSr9j9LgHiouaV
PhNLt9X+ozB3KFU4EZInMIalpGJDgJ/CemwlnChUV1LdtxPoN18SwzNKOHuL2/bFA655lrE4NKhW
U/wi0Ayfs3ODM6BAv5z+YMy35gNjF5vct/MT/1k2n5iGRsH2uovwCjk8idh/g1DY3Nqp5JpQI5Fk
z4pNK47f01r0bvwjxyj+SnXxQJSYJGkW/+nAn6rvA/Qj4xwey1+Wbpj9ulWWSYz06dbUbZflalVV
W4kFiJu/dnFbIkYx65FGJXfPdWmSBHLnOYpWaoF3ZWjHexsySzkQMfEqbwuqE6HFb38Efjq8ZdGl
orZyPO/H87ETv1axlp0/PFLcn9QfctAZz7Ijm3iMQMznAR0HkaM96k0gQwGgA38Hkq7Urs225SOt
jvosRr7LRsU0FYknTjRS518JrBA66ncKTuyPQjl/4PsFJLidwS/GcsuePFQ4JQYdlAfEmBuQxnF7
N/TrtKydKGjfZ7RiWIc/XRudRQynnsbCluuJrwbVrsbzItmqfxLjiRRcfstFn/hu0Kb1vBJpU41R
Bi5DglrT5R5d7XK1G76J2XSfJmA7RobpCWwPx46G64kwMinKacRcg62A0daOL4ODlbxYeF1Udywz
R9Ek5YbFWE3YGb+niym3sdLkr7Tw2BzXTEYYg9TWPNMUoERzKEAdgklmxfFAR8vjborTSMfJdUnL
4+4Jt4nUW3khu65JB3hjH+7t7bl6NJCyLtbIfxzaQloLAoahaofyLwhv8lQXjubJa9eOM3sqkxdj
U32FC1CIFr8J/esKKdSu3y5NO/y5N4UeRB4Xu7enPMehVZ8Z1lpYglauDm2txnove5RwqFihzcG1
h3pURsDIg2As/6XwgdNnZhNGQ39JiQs7ws1CHXLMPy5Yy9Q8Bl+lGDtXo9/wCqsxLXBLtTklrIOi
onCIXmlJPSvLfUft8AR1UCxUzPPrHBjML2hUsx/osNKV+AcyqvijiDX0U0WMLfgnco+2ZAMIJosf
Hke8SQIUv0tswwihI+7IJEkBTfnn/Gzg7z7KuhibGsPGWunLjja0s3srI0TG4tb+Iq/jZ6c7oYxM
XSKAf1X92pbZvckSh3p4ZcyA246Bj5MQu/8wmVvpn+0VznHvkZMieYbt9WlU5dfGWtc/T0c8JCTU
h0dmsVEb2KPvQeAr6HKV5jUCFZ9C1dkR5J34Ydu+1ciC23jEQjQ5zFT9xon+PyzbQtI3m/bwAPXA
6NQq7uCmmn+zoFuKhZQk2LtHKtEJK9B6sbWje0xOhxCsNE4ntgaoDCGiouE8CJxJNnzrsywpHpov
AK+luXpCZjVHwfVy0HgXngr3UM0KNK8T5sYHRiWxItcWfutDjNwL1K6cEJJQxEPYRls5oToi3XSQ
L4LktkywdIgOlBPc3tjY9KZi6Rd72AxoaLWF7j2rAqBDG9mS2klRF6KzLnh+yZCPRDgYi3GbUsrj
BXqlSTzfLmGIdko7pkcoOhb3WcjvAvrFQ40TH1bi4YPsNkdEoorlJ5Uir8myT/4raYAOciTcURzQ
p/SggKR7bakpzuO4x4qIOgIEB/KLEcd/UiB8Mq447NJ1cyk2rt/bXsfnhflzbLIOoL+kTLzppBWO
xI6z1uufVriJ391Au7xkRbRig4MnRd9mHOab6yZUc2RV/wQN5yfnuHOepwqUqf4kObCgp/zxVSNl
6UtkqTw/nvgJsjZWFkNW5qcf0M2Xa+SvGHQgqFyzzBtkmC6q3u+TjMu90iDfQdnWx8yrMDvRmuOM
9FifPS3zaO17kPvLjvkIpARBuzycRHzjqJWQy9wQ3YF1cEfhjz3xCzTRYA+5LUD1A+qBlgR9GTR/
X7NwlVoLtUC7kbR2ptpSVYlW7Kz775oKfDmtG2PmSPEnQiM2ZaFL76fbr4VdBWqZFltXubPuAnGW
rhWEnETcSAuLfzjZJSlLoNijuSxdt8vyM9Rd0EPlI4MprAdSuHZEWumUrWJ2nrKhezX7+865/w91
yE/WZpM6Xnh9nejr9MuMIzJURq0V349ZfBNV1Gw6PAy5NgLW0baN5XLoI/IcqXTRnocsehqqAa3b
ZvCkeg+OhMrMHywgSAzeHd551ibkr1mAd1HIxqUloeyszw+ZdBY+cjxFyRtt3Zis45ERpxRFIxx3
R+LWc/pZLloJufmPWkwxsfcVRdWnidcJP3kxfqk1ipSDf0EQfVHS5uTsz9CcDZM4fAV46BDH3eBz
V6V6JFBv0XVS2Sxoe8wBBvvqjUuad9nAF4lNKzKXq9949RGWZL5qmhjZn2BItx4aQsZUX5pPnGaf
qPOXxTZ9WvD7hx4cPzTcQ/4wv6QkK0k7sSy412Vfgf4jDJPtcJJ7Ng8G3+sSo3Q1N6yrLLUnHzl9
MFLQpw6REUjPb6wQtcE9giSDDDanruHIiD2yQKLarBhj5EcsmmFP7lBjcAVpyZJ+rfIlkNEDje+w
7lw6OAXxVvicJxgR8VtDrIrMOQtSL5OqOyO4/d+H56rl5x4qDwMW8GgTBb37OD6jDXDuGSPu5WUr
YwUedgUMlBPZkqCu9xI6mdT8vmWDd1iU3VhJtvggKGzQHcdxwXV0Bpx4W8eS+KC7MnbmmbLvBnTh
iPj1fHs75LBD5gmnaWME7yekc/8egXW9P3Yhf9VgGebwGtlVs5i88sImg+lBSgRoC/xyVfqyNbF4
cmVNZR4o9tEjwaxLOWV82MzYO7VOvBQ0voEHLncPMmCoc7WL5lt+Lcpp2yHi/yRaEbalH9EDPw7W
wu9W4rPUHexRQZ2/3lYCxljYybW8K2ecHESbSlfDpellQ20VFPFbR/LdmkXvZ5MnIgiZmn2pf8FG
DrO1YwVs+zhFewWq5tO7pQglBbX6EDnQfoufTdbSBhCaYJPdb5Fs0gw3AxS5skugd+adrpmNfuT+
dT1EDgKVzocfn8P2U5yHjOPPJcctmZexNFYBlnirWsB/7MS5QY3ymUVHI/wlOoQzBbg4jq2GpjGi
5yq6951Nd1/baMsveLeGpShZXmNEimZzKRZ5rlKpODHIDwByCDR+1XUhVdP/TN2mrlGbl2yDepKl
Ifu/bz3m8o9fCvCOJ/mZEjsjBDzesIUJvJupapQXpZblI1BU9p4r0oee9k5ZDSnhwBkg18r9skMv
Vxv6VdxWbvAcb18BEgGTv48aOrRjoOEjpe2xmJME/lSoSlaVJpIiTPcCi4VsCvf8govbvOygvDoF
xZi2kGe+3BjwmCR+t2f3QntiFzPnVLsNN8zhLdNubJUz/1W3SgttkX63MbqArMlyxv4k/htiPYfB
y9/ZHUGzNoKo+qLNu0XU7ptFITY1TvoIjZ7xfzbyWq14GyDSfNFbVF8muIMHlJsn3J5mRhFA48BW
ie65uDXs+P/glYONQ3IL9w80DERzBHvh1yvfOjinU8/Y/e7K+ZMXyXhL1dQUKLfChJ22jFg6anVC
e9ZmV2cyomTyq+05wH704RJsR4gFzlYi0O3ddYbdOfwcPpD5shq7LmApJBMDwhUM+1J91+WC6Ghj
K4XhNDxVUeVQCPsykEyN35unLY5XkGUaYm4wV672dJPU9iaN/l1lsv5/UILUQfKSzotyhQOACvGi
itOgI8zJmUfF+YARgV+zOUXeUcaGiQUNEZnzMbDwnYA3sOZ4TZ9v3x60TfTKDDAepIWEcA+tpPmh
N1vqtnr07qwgo0AO6Obr4Lq3233hdrEyO35Q7R5bzCZOw3J4mlgWFAUhDmgmt+gCb2ZdXlOcVABB
aIQuK+ZUvSqHBCJOGsQJi1efPOn7m+1h4rKs67EdeLfTdOX+QoUbKJPb3Sk2wj+VWRFOPjMztX6P
AaiRFgF/LqxzT3eN1ZLR7jNcGHHsVz4Ljx7Wqqsn1boIlXzj1/tBwLkUo966pVjzuWt6Vs3HgZXA
ClQJI/Ynf7xGphI+G3yxj2bV/TLbUL21YZcYxB/HyG2VZ76/GWYi1QDMPBzdXktRMyqCMia5OVYq
Tz8dAWAeM+cVK/lWhNV1qC9aA8RJRdgrtIAU06FaoECzFLya8uLBzwxvNhWkMQkyJx78ynm/Af3L
QESxX+FdUL8g0W/8es2aqS+xppZsyWDQ1gNw6k2roOaYGw0zccXwrmgQQTrfog1M2YlzyDEgh1EN
4SaACSSJp9iMmtGVIlCMXTOgpc8huhYkWolcUGirjXqL0KuBKfSkNdbQxlH+502f6RF3vqGVYSIa
EmU/wFkOwhRrv/GZ6xCBcsbYc+eK/onWJAgADP2sQg3tgwd8g0w+yj1eoV6xYGGxO0TVDyRF00/O
BDHonf/KbWN24M+1R8LzN06mzyOprDGn7yaeLfzfAqkOUGEWSe2xx/o1moY8C/u+60PZxOfBaxB7
YuvimnAwxME60HJ5j/HdjaDiQw+6T7XZ7YIgz8oxJzxd5407hcQpb9QkqWGyCIIZtpScxujbgx92
tE7789c/HuVAtKSX0kVJfYPtsFqVpD5VVOjnILWJILakQs8i6IJxx3CBShliltNgpo9Bmcr2ub4f
QvoFFirKjsWpm24CVCX4m3IsazWHHYR2BEZDQP3xkHG1/z8DRb1NPsYlMupoXOjRjJG9lSISvlMI
7LU3/m5tbEGlkjhRVGxeUTFSLB73F4nRUWUQjhuzeGLvFX16D85mBTQZyXB8CldmXHwYOiAvM9LR
5maD61K44Mo0b29FCmfbHYOvz+YtwlRcVT9h5iaSk/8K5RIV4VdbHZWOvChiBQlix/WBBHSqSKDu
wIs/11PKXFKd5yCa+1jpBf92nOkKLtGnDtCypyHVFYHPF0p9M5ad2ALv+PqZquj/Ezz3Y84HkdlG
YFY7V0xqI+cwQ1jpVn72HqOImzSEGjnSaKrWY+45xexb2AXiA0mFSyRXvAFjfaoutu51RkfGFXUv
PJiXF/VO7lBxbTIavPKm8LaaB+5yG7/2ji1ANJwQEh3N2w0S99epeQxVHhDUM6XYepkdokatdgGd
w2KiLCVad5b1KfdZCBf7qt3m2DtoByRziLtPX8K2ZD3D8NV53Z71Zimhi/iSv8/Pti1ZHSRv0KhF
z63RI2i454I0ExVbbTZ2o4CQ7BlQc+W03YP9uKCatr6Rk/dW9LIX+HcuS14977BpPy8dBkNMMXpZ
MxLtI6O3NACPAAm3Q7MC117CVr1Ul2ZDT/cLsY96V1JobVhKFZ9rnNgI47QsGGGcb6RcmMarSmxI
GfPl5HPEm3ApGbi/xQirtfeBFfTmy2sBDivP0gQ046FBjd242DdcRdmbYjSH9fW5Y/grldA3Hr31
DxptkW7uxEnEf+slYDVx9BKXzP/+LpRW823+xtfRNZ4ACEkjA6lC+6UzW1Rfc7QEjVwBBCzKScO5
c1iNBj6mrd9zrgsodfxlhFBvJkAgm5CSs/hb2Km/X9veUehE/qZEWnqyykLqSojnE5YI0FOIhGNl
sr7hQNf4HZf9fa9ygKdt/POIUC1fX2nnL6FY7TB4BGz9bxP14qZRhyj7pgEzrGvi7z/r224q+/Vl
sDmp56+7Y0jr5/Lc4qrTuV4/OaT7LtrebWGTXz1AjoNOCH6VZV4ZLwsMzsKPeI4i29hG/8BjRN13
r6wTWIuUWZDhC30wGZGkZA2ExJQdxiwES/xkCpy1ZqVWaOf8rkHAaShhMAHcvX2ccRJjTLAY3CEo
Hxaz+ynVRwyYq+5mMcVoFt/0J5P4oXu7dZPqU2pdxEPIx98o+0cwdeQ/DU7FcBxjYevAEy9gGhBN
iTlZZqLK/d+pXbb179EABrZLf24PIQRlGMEJAOjG5O50MfdguulFTitBKCFocS2X6B2xwfh2n2JH
htl9TtfD5QzhPZxsw6kmrQUd+UyXGx72xZSKx0mXuHNNlFbt0URp8NYNZsV/3sKNcL9QjazDTwDl
i6waGz4Oz0hurMKa7FQg3Si1pGdvvSW/SFS9tElJpgi+FMzp9ByczYepul8IBzfj+5sNDyl5rtbO
1dVyaTxwQ8l0ZqpU2kvPOQk0N00I4CrAOvaUN1y17sVRgwm9KSlgLLnJllniVEflzbZcQIfa2nIg
7/yEZ9WN1t19UkknlYAD+nXymbGzPKtfFXOMlCRkefoLtcY/SIHU0jTtbKzrgVRvTMQ8stHxe0ob
Q4qlsCq4kAoq2siQ7c5kC5NbMtVuqF+DYgsTdDG4wAbsWtcgkMA4+J0LRvwvbZbGtKjOvFXJLXC2
sfyXMbuTeGc47lXhA3+7EEfsbAmgJ/L00iPRRQ5nS9G9+6yDmZuQwZzG2kE4ao6fCY6JUsHBO7Ut
LfTeX4EJG/rIWIa4qqyQHCNffV2YXiT8UT6DuB8iocwENeZb3f1VEZrdHSkJUzOdF2+Sc8hh5o4x
5xnZ+ZYZqXub50DZNZJ2pYHeXmRn2k5G6DEtKoo34fS1ClTmG99LKFdNP0ufzD8T4zlsjTR+aCa1
Yq5kG6K0p49glpfl37QWp/PuGs8kzMiAJdMHnAUWcJ2i3OrIxwXfmmsH3rl/n4mrxUD9rrEjsdeH
ImDmFPGWZRffNwqgPIm85VCWxeAx2wR5DWdihX9c+wRcuzD+CbmdfcM9xjM3IT5Yz1jLD+U2K13p
jT4DxWsWoEJD4WQGKqR8crTJ9RMbPrlCVg3oRnEAgOHM8HuSArJH5otwnQsh8U3VyVzJX+kgMcWH
ynm2zvfsPSA/Y5jWUoKDy9Zon3RKzk/mG5OTvCs7h6fTr269aiWp5xB1cI7e+UXPegKK1pPnxk43
xhXiCjS2V6JwktuO9taks0aGEPgElSAUPamND/sHzRtA+GaSDF1zlmN4CUyHzrGftl9oL+ICDIR2
XxCEblj85KypllNAjXjfNbdHXGQVc5DW3RdSIJmqY+yMayO1ufPowuxL8yNhqzuBVp0p4oTk6OHt
p4R48sfdS58Y/L6XZJvujK617+CvCNZVJkLl+B206RMKx+VwW6aulQ/uBEu1wqASW1swtQJZ8kfu
jayDjSSPc1YtqO6gpuGXHe1rDs4rW1p9LcHF9rfSQ/UrR6h3Dnp6t2N6SW+FTKUFgXTF0Sr7ef4F
A8KSmA7/ARq7L8rOtD0I2mGeOePyYbKlkjZwFXwbaUiFnImZFUGiGoJtupJ8/bppr1uYJm9herCa
HhjQnEhpD3ag8GyVxh3KQBjzyEcDFM+w8Goi5kLsV2OQBMRhLTi730Pe4vSuc3qiCKqHH1ms91S8
LK3SICzM8wuGEFuL8TbR3Vbiw7Rw9TlMegAw82ZzjfGMtP2oWOH2l8uCqX780g7ERPi/HSLV+kee
SoGNnw1IAmLe1qAW49jktP/NBzeWgxbs/5L3D4cSPu4tx/X3lvIap1knuNVymySEp9YXTwjygBZc
qbKluwIZT/uispiAA8hCGX9vah1P6iuLeusFRCw1ZBf+9k+vJqw2UBU+sEJDdfZ8NI2IGuBXAmz1
k9rOMnbLb/MPXbCQWCktRjbThdZUeJFsKX8OnEIkUEz4yIF1sE3Vne6p10+SauL4Wanhrc/QyCns
1vfdDUM/CAsk1YzUoVvrVxcfpw1NokywpV/HFFAKEC4/lY0AVjp0s+DwZFVDmOuBKhlS3tOXIlr1
A61tcqf10IHtmIvaw0vm0SkXHuTnPkgTPuZopz0f0KczBpiosbTOWU8gFi7M0VRj5fctqgZDev54
EBITzy3uEtlEXsVEA6SXTwGGMJt0ApWCbPUdFu15b+yo/UeT+FnUpdWm0PLcy0ZVaa9bjXPXa6Qh
2jXagOxAr7ZgTsLewYcUmgq/2uvfcqfUkcKUm6F48RvjAqanSQA60tt4m2TZoFyD/2ya1/9pSJwJ
Mq2N3GVtoukk7xESfzVlDvVBTOWUi1klPYEIgRsjt4XYRf4IP1TZtXzNMotmjwktqKeKKneBb0ss
IyYDwg0nnBRyLorTlOgyamn8D92iWPfjwefdV2gn+bd2m4tFEJoy+TDsraeYDgrwGLZRqxfIf66R
gN4ii1hbBdozlvSFwXTIdJUQ5umb90LRDHt/w3NlEmZu3IBRgYp6Mu8YRoHzbvVK1SLcWfr4KSFL
cnQyt6qGFfs1+EBEWl5XUxSWMlCOOBj2Y+NGN4IwUJ7NA+VtV231obozRQztZpv/CCzJ9XERUYDt
03JgSgVWBF20wW0AwvABov3yjOYHY0b45tWhevM2A8/Y6EctJhk8qls25buS87GPODzJIWUBngJn
pPoIdBlFZPhl7Eci8jzbOCC9dEFsfPQpmBys5BeRhZ/73KQWG+v/mOXTz4bFlPXwc0kuYwjnkGog
+gs1jMfaMikenJ62KyVpvDSUP0GBt8E+KVmdKoSjRNvCKYUUSeuKOYPy8zx4f6RcMwn0J9sOXaJ3
Z/G+UcMb0mMx7Wai1gfEF4/8b2gJXBmaMXKnOr8brElhom5jV/u2DKqS1UUhxi0YirpjezYtX5oM
9rqOLU6q9Bc+Gi/IRK0VSuk77kgkVky/syDfg2c4usKIEnl1BPwQr7+Ia3yjLZbn5+pYtcnhxNwu
SnBa+mDFAt3DwSNJ50sCFuSDsoNoZ/uywRwZHXpsKRfQwzFG/lKdxJ8neAOo16tvpUbA89mhCWZa
uBxtkbYHrVhZWdFbpTYFvYh6h6xt3I66R0fjdCG/khDGK9TZTt6bkvDUBO7gqJgCiIshMkaEG1Kn
ddCeE9KzKYY+KEb+66JvPXAVw4lDAlqEEM8Nv1e02CLGNcGVZG7ayCP71qW+s0mUpdRYtu4WZBpR
wvV7w3tQdzlG9os8wSCRtKsftPDqRdMWg1yOyWM4Idh3DszD/LjZ9rDesAx6tuJKRiFZAX27ypRy
5TZIYH0jhvlU1JkKuKS6Ua0xtEvobUJh6UlczPaPyppG5/O8sp/C92J5LyEiSr5/QoHrbIB78sbH
wvcvM7THowUDCE+si0kaG3fi3Aw4FHGGCZrVi7p2f6M4uVuf/Px0uzmJTEaCObAKv3DZGzV+3wh8
czjzx9qEkj87hN/uPwyuAxovezm7/FrwGPp/SPlkDYKlh6Upn1JyiwqKiCtxPoRLCnF6JCd7GEKh
qahSYiBwSdD05SBJssFhXo6jmMaUJMKQBPw0JVwzRmr/xsiajC9fSAuEtmweZufzpZpEXc+Mj2/+
0R2PLYiigBTNEn8p4w4Pl7gDZiOAouAZKbZr1flEz2bIqwlHT5aQ99KAKAOqiNOFuTGfxC9XLgjc
blnu/rpAG8EasvWzk1zFtELlGU0s5LmVQ8d1bzWXPzir1TBlZJXFuthg+ZaO4YW4kf9qUwo1KUyP
okl9m+fY+bVkPpZv6Er2ju7du4hIhDLelcOTKwRnBdESxajbqE5nEwjLLkgJIuioSNohnGYqF5MS
IrK3XhR1qlIJKIXavWydF1yzymhEofNVbN/xCdH5lxSijfh5j6C7Dn45B5L9L2npUmtctoSKXMX4
7Na3wHcoisrk4ds/1dWmFgJKYGEW2eioqGbiS+30iaKvPbB19yE8TIPzSbQfr1U6U7RVNdK21IeN
Eda0Y9IqbJOA5S+TfcOrMEoTvds2yAS41kH19xGiJx6NTHFedLn7i2MG2XpEHNS1Okac4XTMMGJu
T4Gq9eBo3euH9aMxnjahOk9JMJ9UR4stZH/XfObcjkBCaKGP9AVe/8Ejjv6ov3Yu69TBk5rswmw7
985GipV9tn70bQjSP6UpGxOSRSbg5M9te2/SrHEGoWu/d6/SCryiUwC2FqsFApRGVshl0HOk18e+
afdktSpW+ImKck2RUeD0AdMdY8zxZb+16CBLM9+lATHxSMOwbmxdHzrzjk3Ui4MrmSasnso8GfKQ
vzaSYcMMrbZjpK1+82VRkUYu5BJGX0A4DRX/J2UrXS2m09DeBtp7fZ6M0pnpTezy5SsxAZQly76n
hxcz7s8yoVketvmtxwsBSVtMdlGrLIShZg2sOXVwIgXHUx8/sisyb7YUBioL9SMhch0tSoFHMIkQ
j30poEjLr1jOoOnGcZVIHmWTULWePZ3anQu6GAEKn6CYvb/PI2BJcuc8OPsVbdKqqr9dEmV8V7o5
yCwYzq2IVwmzc+hay1hrqCAULvXBtWsTRC86aJZt2huUIeePaJjKMbX+zeC0heZOAYnni7eGh+lu
uAWwlnONrKyhQo28DzqB3Q6nhC6pBTg4CnbD93m7PxVCWTX44fVkweoDFG8nW/2FIwlBu+UWxuGB
jgUnXx2lzrQYwz0SimLLuImE+u89wD7VYI12LMqwfmWqcRDqnST6HcoVzJlv/ckAhj07rB4QzYMP
mCOFjPY0A4VBp6RZ4y3S78hmAFHq/dAcF4crxx0RZTgw2klbwVWvZKAQeEj8Tkgpl9Xed9GdbavF
qs14xI9fPfNO41hmwKTO72h2J685KyfEoysLwd2J2Qc/W8UooXQ0187Vvyid72KkRm1vWZQz0S3m
v5vaLH/Amlt+rj6Okiu4/EalLzoGDhw47QfyMlSAg9ytbHH5mKh2kQDk6NPfeT0zCdyVwu+wqBbZ
jbmo09vgaz4DiM3oRbnZgsb/rhiNFdVydoZVTiFdpLchHPf3YTydIDlmXEZqEok3pxOlZ9A8ncrO
2CNjp1pCSsx76YI5mqa6MoG5KqF39WqJTXGCWbSNNz+Ish/QsdNSIvWckLL82UgSf8f6+lf4dSiV
lLvTUFBWwC+uKH95ZlCRZDAE92S1NGUBVCyApFRrwXCvTCOYA1epEGTwbiJmRkhCXppjPtGH1e4o
TnCpr21IjABO3zV67sviOafmB5bsA9+rBUJ8Rjp2CEf1uENQS3nsDSnMsNLr6UsRaEF/IJsCtVi5
MFYmLNtIVo71gInp3JamARNZLCat8K9Q2LvE5JPKs8lIl9GT3PksodwCPMQXlkUyPRhHoCRjIK6+
qc87z++G3NKB2JL/Oc+5LTcz6rHQHZAfoEKecDPEytB5886VA5umbPuf2upWy6tCnXNkhZqpxJYw
sdlFvd7M2nTD2PqzwDEEkOkhfuE99WxwMvG5w9JRkRGT5IR4JqgyaADLCGYqEIT1vR62nA/qSVVN
Se6LFpDkBLRMEyO9MIWD24D1Tza4y8LJr6YMxhY/HhkbaUpHjuZe+mVu63WKKJGXM6gRVKSosAa6
D1TVE0aQCOMXhdE7wt2lJ4ubcQlLSWZJSVPLAPvEuWjv0gRZgPkrHOZt6CXhwrBPuenCOhtS75dk
utePQNTYQN1oNZdCcQ6t5esgENNrBK2kX2eC1spWjYNnnluDcunWNdPGXTJ9tWg5B7aOHG5ngZeU
9QRe6+MHsRxZ0JMBpUXr/KOgEg69lGkXHcddZDBgvYLRvrgx6ajFmHh310xkJ7hny6K9VjnW7bqU
aUOrzaADBL2i4wcpdPYA1pzRPlmCZmIsxsEhAI1CorPLr4NAs4BjBG9BsD8Xz+BhDklrbRTITUjs
yP4Em6uuAkr/O2mZK0rLbwt+CPcrPRbqsc8LYtBXx1K0iTHKfYIcK+9LAqEfEOwy1ImLdsXoDL1k
5j2FHg3MxamdPUAXWLaHH1YtAHw29U4FxZasSbN7ohnEqK0TO2UAuLvfRqIw4pub//1DZZOEi8F4
+11fCTq/xiS0BB/vVAA454eXnvWZioK1pHF8vXX9r/myc2yJG1TxzHNBueT0EhnkKQuyFeEowCcP
cDNJ1ZaJxywG8OoidSSa+bAHnAAPpwLtj+xApHrGWwP1YYz7iOhHWL9zDfSeOahOcrI5QoaepIHA
NKIJcdh4KISrYEJhpnwF9lrzutcH2qGtCnbJnutVjkVdxGqdQuhSLRNUdS18GOh07DSFNqc19Jk0
eAHkrnQVdbNjTo3BlCD45grgdDr8+A3ldzZ7OwPNtdgvoOSQfIuDHHQDDFDzvcKFUR+B1f0y0IZs
zQ1sgEl++OaDF39wT+m7KR3pOwmCHwantLHXI7jNjZkN8ZJYs01agxRSpLEN0QUqLjhN1SEIvvGn
RpmMImrmaeEEKuO6xrZS44xbyplG0BhfQiJ6SZWe9ZSp2tRT1Y5bPO46gGLtbz48QDPcI0p9G2L7
fUoSq+7/eL4U4Z+7180kF+JGv/i2LTrcFcNzTze8GnJtVdTfkJcjHnyAWF03Q5ApO07p6fHiJ0JV
KQmU+gtfqwkdI5MjFblIailFS8y5kFy1VtsOIhhxhR7bpfnS/xVo8miYDfa4BWeQLAv663R5UHCc
VMcEqqF8F9xvbI6todUOuybG2zNfKivz1/hQd2vp2sAfjWT+/ZuLDKLJESPgxCDlpmCl/smappjv
u8CqX/GKd4SI2Z95Gk4P4KTkOSdZAuikTTITbkNfUgwIaOopVZNGqLc42Is0/yUZ8gU86FfaF3Vb
Nzje0yCQtAWSc04hfnTWwjOVXTsxIe/nEef92EmDgwka8/r5qBkFy7bOxCg53LeGFGb/VOsVSmjL
M1KeuZh5MQCky/ZhgtN2MFhPLm8CKPpCKZM4Yn8h8orl7vsmg8qoj9Px/2tSg9v86eQXsXfOqlTM
XJHXVKwHgX4+Q84e2xQ9cG/17Kio3RKawRaDPcZNd7XuYu0pogeIBIMEdXN/1FiHpQFfRg2zgJed
WVd1ZkYa9YAfT19aLr3G5O5rudhNcSSJp77CsWMIAlKB5ht9jIl60JaxeBuhl9b/bGmI0wwTb3SH
ZQ4MY8bFGzvUiBLIvhOflVlbD5nohopvucZxQvZD4F/BQM0DLi9Xso4aI5BmW8ZMHF84VqP0TnmY
cdAsPgFcpL6XqGzsmVMBiXd9ZQUBwHAE8QPphZLjPrAYZNAPekaHoO6aP/PlVwGuk3UKzJzsIOtu
wamiA3aXwrW6HeAyMO7kvmxSVoOipZOxiM5+pz41LQ21WIuKSh3uegrnTm4viAGtC28uOQ3kLRW2
84yTXBM6Pz6jCnK+IxtwIZO1nVmbNTXJITp0BfwGchXXwTc1mfjoYNlQjvOMldWYH5u1EC0VrVGY
YPz42Q4Gpt5MsT0xagXqV8oY19mKcf/qqekq7BM/ZTLIQBfnKeSjSiP6MSsOzYmalFos96GxIk2L
gdTHJDXNRsaWQFaldD25uvT/kWuHNfJOAyDClRIwjZnurxWNBcdjIJSabiR4+PG6JC2oE3gFq7j0
SKYEYvopoCKvlnn5CpEkr3pPZCohdnTs3MTOFiJoSGH3f3tMjnd96Ys9E+lKrPkNkCqeIFiE8fj4
7ALO90qYI0Hh4APc+O0mK+atH6mbnyb47ox7gCpBUBWN6mDK411a9B9pvgV/lm2HmrFGfr0akukB
P/QEExMJJp0TyHe6p7RH7Rh1HhIvnGUq5ZqaPCqI1VH+BmxRdme+Wx3WmhA+fATjvitYMvcduNta
kIWmLaCC4WOW/84wXDH5zbEEioJCjRZ0GerQ3MAxXS03IVEIuyOJu5xo/4eanF3URtPC6kE32hJ6
z5nmHtNg1iwmI71V2tetATMgCH/xGszrbsO+Z9MNYadUGZDFbWDVem9Px8/3tb+NLBHUZXMUNr21
//CksZnXuaBsEhHlmLeDMEgSldYX7ZCJhZjPIj9BOIjEuUpXrdheoU5aOS+5/40yFJjPPtKeKeOF
454KV2GFZ5EOxFqqcN0J5N9LkVVAWf7DV3e34Q0zs/T5mm4PHl9Gp5aBMfAz4mczWIDBFmV2WOkc
1PTOC3M+GBRCUZICmHb2W3huMoucWK/J7N4bmBZqdrkqCwGy73A1EIZMRSDkAff9zZpUrOf5VFbR
vIg/mrEkenc7bma8+/4+OXYsB7FF+/wA4ece4hQlEXVub8tKJo9tqkpxj0FnhoiE3eKWM5lmRVN5
DBiiDesIS2Qee2Tv6B0ZDDxW0kiSAJXrVLfzYaUCPmNE4RWucvIUNub9iRI7XB0grixzFTxhhVJJ
5qjaia3fVCNYlNQJX8EAClt3qUTk+fWIzDLC2EczVkuL5aAGK8yen1ueAcdiuY+TFy7ZeMht0CUv
6lRe7+CIxUx4oyqfwMAZZyKtthH6DXYB4DEQnPGeWacxeMOwChKq9uJ0XgB+w44yRO/lfqlpMr/8
NA6qODJMSPG49+FvzqFUo4vNYT1T5vIwIJqLqirFZ5gh+YUmyaPqOQol5fK1R+XE8NCZqqYuwPi2
222yvQKPi1Gpwt/PZGvwYjJHUlovlBDCkh5XHoKD2nolWsMpFZrjL0c/aA0eSS+ZcBhLvoaOncBu
aGa/moRllKkVUuJWJ3d53130AnxD3AIekTlxWq+/RU9Ys4dQUHcp+3zINJ4Yzd7YfgeoFb++rsN2
0WQa2n54ggUbrGF/70yWUf7tIS4lSrYKyzUx8o16726fXll6PbeZ6BaRMZCb6BJsIKxq3fZ5PBde
QTm4lCSMqveTv6Fn84o26KHgP4qTgAYvDQl/DCGFJowJpfiOBMyzbqKxOpIruS+zs4PKKKCzhZWx
KhC9uNUQt5JONy7clY7cpmwdz6M+n7ZztLL1niaoDbuFd03LNiotzCcb2pE6r9MM9Ng/vctq02LU
zeSBLooH3S7nSdIwam5UVZpkkUUgflkhDHj33FBuWwc0+wGoBJgbY4/axH66ZG0qJuJxtkQNyXpC
DbbR1NZffFSPBoGEQwZUD3kC2oilaFboYKLwLY6nglfPsA7JPtN8QMuI6T1bExWrmVDDp0f7gi6R
GVdGM0jY6sF6SeNQsA/3st6nV+6zqZV9qlhRxqB8oI4SJQEpBxEBcwh9c3awZyEY8ZwF486KvJXc
lnZJdKbGCYryEQW/alYLmcTa3tcM9Vf5jZIeJQQGPMuE6Qu93S1ysPFc8d5Kn1At+zqUYbE+pp8v
NrJaxrvvsge/8lGKpGd5mAjfMb1CA4mSd+QVVPayitT5nt/tf9TpXl4G3JBYmulAdg4HkxbCeedn
YLVgxyS4gbci2kTiAaYz/4cjhHy7iU/2DbE9eokp/Xt7k031Hjf6RZrErDrJarWNHa3dqV8biLT+
zyWuQdeusnmus74EZsVYjz8nf2P+lgXBCehRHnth4xpgizRBbmm1v865HbDSdOSfT6jvKVM22KxT
A7oqJSaljnNqCRjPEbbyhd7IsfSesgWX+W8kiAbP6wFgc0OI8k2Yn+THn5eqLrBszoF1WRcZEfA/
GRmmQuAXjRmKVjudnvVd4vrRq3+JPghy3QhJKseRZ7Q4tTDmlLG54ibQ8KNJ2usNWnw6UAP7s1ll
9N92Lnfnx5EfncsAaDGWyNL+iyikN97szripkTxIn8c9BctX+Lozp77aluYp+ow6fcbvu4DfRol8
wjYE/uzpTkSDPps9vxCDQ1Ig2TgQrwtP8qENoh8PXQh68LtlFgoTtjFdqgI/LuU1LH/pAWytDlpy
yECgVh8jIFlt2MS6IP+Yk3gm1cTm0Ws4WywkYuTof1lirUl/+PlT70yXvQFl3T3XYNLGlfN4kxVR
Pt2qythUyheOnP7gqL3ddErPJVTZJxwG+wUiFD6ZOvw1i9AWoPbAre/7i5V8FTlpG5gjteUuCDuq
7H83+9A/7KE2DO5+A0oJ5qwE78pJDvyreNspHYW3fEuQx5AJN1WmiC6YfQAd76wjlDkWg1i6OjQS
+kaMyWUIEPNnEPak713bzkMcxx1yR4PuomeoPi7VQ2oDYGNytr7RlOpnjxyC2kGCE7+z2wgW6xC4
pYZ3gDrdA9uQGBXNSuvEkjNm0vb3cdIkp0WFWvb+EjwJ46SPWThwsJ2wSt1JJYRzvptlX4bvBf7o
OOSfpXt3HWRyhHoOto4g0nUlWmcQbfd29UjGeFSBmzZF76HKf2+RhcuvC1fxhBiB7I1usSvBRj44
SXh+Ov2s7bwGlPhZJZXTlQ8/6KkE84hoEjEgBLRI3Fq5ELEAWBisxsE9zmRUyh9Z1ie/S5LVtKLl
yZNPcCkX4RIfnQwqPDyC3vItKqCb7koFYoFGPlYCCGl0ohMkz3d5yUm4S0oIuS4LjurBAOv4nb7K
nS5bqEzZy/EteTuUvF8rjQ15hmkesG9m3IVhQW1Hi8ADe+flxXXdMLoObwW1/bh8YaYN8p+MEL0v
xzbJ415iJKGMaiGa2mI/PceNE5f5eTSYWKVzjNPgGaird8cR71h/fSvRHYDkFcWzCl8lg1QlQBfr
YC3qVmdTopMnZ2SHcTvsT8JkFyrjN2UTWSfTr8cugyMgkgT82+uDQYKRGpke9MTbDtcqVQQvKryv
LBzqljHDNm4nR5yfjJXbmC4rRy4/h2kVyGezmUiBpYpXZZCHp7HQE1HGOjyvLWbk3Qik7IxY55O3
eKkh852q53IvbLp64k5EmHuGWP180KiKtAI5VZ5QmsNBVVnBasOXYby6xbB7YQdoTFq5LRYwwp/Y
rO7A2GUAjZwsHsvBKeXM01tWusvyg7In4zp5SAF/yYTO14Fj4S19SLmp6ZUVQx/a1nm/lQxJyELo
+DRlT7m7UNeDZAL9N5LI4rYGFVYYiN+YzRJ3Ht/b4I6EQK9Q4ow3aFe6RoSrxIm3Sfoncjlvynti
W1HHU5MFGJcMlkFzJj7sYBcFt5kYMtAsVrj8bOd6gjtgxPwq+lBLcnvnHL89k+9SHyGzWRLM/lln
YFnDImMjpPDtDa5S6MWNZJr+cXYJ/GH3phZnqICpLYpH0a5EtRkC6ISwsAImXhOSqVTULElaOaw2
W7gJz3UvN9KCSvXDpZU22d+MShJi/JjwnSLoCAd4FQ4/iKt1zaGQwx2MoNr5ZsOUOL03SXOm0mMF
fxlH/OuA3DcognGmrlCBRkXOg+YrtxqVtMn5mnH/VtNSPbRe0BdOrkhN0gHUb6BhaIRBR8DygqZg
27YALO7120iJFgChORSZZbPKLlq+2SGAOIQClut16Bsp5zzFnFgG94mEhCW8gBoj35cylHvQqUYK
ZydO8uQj3cX7vVRID2wWh3yLjviqyK9zq812dcM3kJjHUE/5zqsZyIf1OToj/EdJ2QRl3siMcZzJ
dZvWT4ZbaiotbSfySMQPJUZIWHv2b7LZ13bswXzwo/57SdRUjgYPuUrrYhcKlcEmUew/oZbXJ08w
/5axRZUItNOuremkz7ca/VB1CSA7J2sm0420gZ9K/BXd55LfAEWfC10l0YmMU3GO5eyGDI0+LWdR
vv9K2gNyRwUTCwUtXrabSHP5rOJ9Ec9dybNu/hoo8D+xTHYgtbTV8g3QCLo0DpHxpWmLTZAyYjIC
IuF6p/TUWSTMtN8iF1hZ4j281hgjXF8YBrua0CaEE7Ds/PFCzJecmZCo2OwrPyL/pGDE+syc9Cat
eCQCMcJaDPLSpaiV4IaBhgIOP6VJSRXsDRwcreRVLaEZxnhs3+E3TtgR04X6ISRL6O6XOof4LjEe
ecwYYiuwgaMVk1Wql2YI9F4QhS7AKGenrHFjosK6qxdMcH5C4vwJcUkpXdVreEL6pwyjpJ0gNDSW
bZpZaEhsY+TF3zSEKZU8QMkc07zwbzFk+WRzLtopr7nXDcfaf8x/QEXZjUIFdy2SbFwE6mn1KXjF
Ty+YS1+sJEp2fk9yFTBMpCEMZxpDEWjXBrJaekWkS3Ab3gyBwnqFT13z4guGtvFnhqoMj9fpb2DU
L+2YMZux4+5kGrYOHBnlf8z1aaRZpjJanLtRqQcAiTaSuq8fPGVoHoB4g26WzmHuy7nk4+dWIu5G
KxaiDzoPIngZNDRFr8v+V4VryGeCx9I5FaXlRiH9X4oOvkGaqbcjxmMcxbhYSGV/Qfn/+8RLKNPl
yyXLKJQebv2SruL9fvcptDMjs+yVwzfw8EkE3uFDzcJwgNT39A++hZ7j0lQaS3U0DDTTq+FNHG/p
RO9jMPWJ4IwpEpTjKr16aNVp4Z0jTPKZv6pjMHw3FZAKbjkqXewT/ZpDWix5G8rZ/Q1Y6qTR3svA
q3tTeDpQFieRCjVP1qlyIn6YhCrX4o2bRyT496RtdYGjSIAGIoSC0FLpBUSoscbpqlY4DMFGJ3sI
gUoPVTZfpjjWFbZCGhWYfJzTLE7qbA9d2v72RfwoJr9T8kiQYSkd0qzQ0CQJGwN19p9HFZJIdi22
URZI2BOFJDOSQGDdNgi0ad1AFCdkK9oWocdB5ORNWqQLschSRQxa+zb4BcxrHTEynxPfbjUIKTQ5
7tPI9LioxkPGUkIopsy01vnXXXVxWzdFy19BhGu5tVqjVGAmvMiF5/M0MYJvZN+tlIpedbS1iDmd
KsnJMjrFpO9LwzBgOdmeDs6kdjqd2YYwREZPLlJNrKQDz9JYGj9YUga5ujyP7CHWD6AIPamf1DDG
ntNv9yRDEzGS9yFt28tBNj2uI8E2SxstgryKLAp72klebtQAjkoWD9tWUuEopSd8TUWXBsQH62hw
Jz4GvuoaiV3vBa0d+IdPC8nwvqf5emlqD3j2S6g/qIwBuV3r/0ihbMNhQ9LpUJfkwySrBZon9I4e
oTL0KKreFsgZrEOPsNq8EPt8xmrkYZlw8HlxxmdmXAMs4pbSz1yFXZDbdpFXe/FW2ZB2ux+Wis1z
dKuJJm/d18yAQqpv2J9POmMXONCxz/lG6WIHQtBd5ro14b/C59+6Ad9oR8hB6p72xlu7cSgvj37M
ufa0yKC1lUAV3YxpUWNw3RpGgEylFTK1KEWPvJkq9PTxvm8p5KcnhMxjSTo2MxuGs2A2F5uPJ5Da
CE7P9TWTyVKiKrcVCROr4NqwK8WwPSjGv9QblakJf48EAp9bd3oUD+L7U329Z1eaMUXOuRW1bn/k
r+nRmwKT/JBDpnxq00QDctzNv7sikQINe/vbqIYb4H2ucLgYlhCes9JxHaZKD15YOcFtT+BVruil
HvP/hZNuSSINNaPwj8WqjrGKzBoSBE/kicUMEtXQVa3poKuH2GSSnyBCO2A0lmUXCPqg6GH6DWIO
kgM9ZU7J00/kUJHQ2QhhHmRL8ttLORZwVHpgoSM4b4u7m3YgVM1H/NkAUwM3WOlO2109qLyVG2Nj
sx+D2kppGjtaiepRDH2Zth5wCS2bCylODufpw85UhzDFxO00qiwTKeBhe5TLsukwGLew87lc5NdG
XSTUlm0U0lx+1kZz/8+u5YDi/JU3OW5Zzv+hKGEeHH/7xMnNoi5DIwlopc+GHNE02Eetf4TJl47r
YAccyZstR/KSOLKiVUn3r9284meW3Nx4K8+Hwpims2AqZT8rlH7CYSZDfU7LYQSWQPwGjHs84xoZ
tK2JAkSFBATmC3k25avEhLKmsr61peNOpQx19xgbMfdREmW1MPUpvkpCXGwpj6PJu68qXL+6kJ0z
4fHJlGrcsL6M/XlKxFYEcKEr5DEq0hIKT3CJ/VTLsFki6NnCszJfwFMdrP6AMwDW7dPGLkJZ75lT
yjFymwPPSyAYcBIC2y2OFJwIBrCqNs4HE1eoYG4XjG/vj8rRUDZUQ2MdgFhKF/iOBWPFxU+Wf+dv
hsF4KuPSiMPyi3Ekl7nDddwn/ezQtLRVnKBJBRlwQIRtcBIPFIh0xA9IuYvumQStXEgGYHLhJjVc
cZpglMwuGxrGkrs62VEjfXfKTmpLMhCe7gpq2zuaZz1oyLNVrQXOd3vqJwgp2EPq5aoy3dQuRgJi
gDEpmRo0QGcU1I88crZSdebB+QsKrd5PdyiSVfT1gZN1YUQGAFlYZAvgTN1JrW7BMnc4WDaKl6LN
RrWRm0zJpotSiemSZMSm9m5SQ/Tu9SgSTxTEkZYrm/6US5QHJYjgwJaEy0mWaZT5pd2LWH4M3SSJ
SXV/C3tmmdE2NYtPUB0vwM6fcviEQRLMQZN/0sHPJ1/hqqJn4WD2WIKpn9lQgtwZmIlVtj7ehX0L
OLG0N1OBAG2bQk1AlqPq72P+MaoebfWX2xdG3HmfCpB4ORJU3zxgZdegfoi+a/6g3bFoeTF39Sad
0quaNHng8vWZlYYRow4oHrcK1ZZH7o1jv23nY6689nBXq9ATJFbshZ23GZqCRmwXhuIcmoRc0iIx
/XE9n8SF4/mRSKp6V9piyyj3J6+D8JYr6weGwsZpPklUQeXprXRUdfNU2xbfW+yjy/iltR3VBbZP
dp9OdSvWM578uu6Lj8bCdC2oAQMtJd1gsZlUI46Qku6F3u/t/+1ZdTCftw22E9LNueGSiw9IcDLr
Hc4IRR3tjFf0tm35RGzxs9ZKpq5BUxCaTwvPCmEi+qEnJUSmIGs2vEmEHT+y3S9aaezjnuIO9o+j
N22fbG6mRNi+aaa+xZLlVaZixv0s9NQigJbiMl/lEAK21Q9zKA+hb9mkpMcvzR1Lh7vo3Vh6phDy
bRuMy1mhKgadVGJsI8FCciOZiE7IE+cDQUPjGOhDH3qpxrpUSsPF5d6p1RIEH+X16hhxsYSfcdtr
1+8R7zw8Vo4irMBIuZVRmlzHK1qOuUbxUqMbUVhXCmg6isuQ0+TeseNYH8X/ODHF+NmZzgdyhlR1
x8733WjIskLrkr6IPUKspJFCRB1PrlctAfo/+DbHb2EvkkYv8s07ozu0dlL7+yPOFt76L1yPIyBT
KByeLJrILug0odWSsZ+KGNsWCVyZticdwXLJxFeSmONnmnrVXMMTdsVUSlV7DLSkXVxJfzdodtpz
Z1x5y5FKhEX+neG2wc86K8lG5gnT0reTylZcSdEu0SSjR01c37go9mUC/Rz9Nl5fBEs1PvbDz38b
zxJFgV7IPoabv3DyNRNumGTsJMaI5Oph5+4NK0m3tRHPG0uBJ2UBAMVDDF1YkxS7ti7bnTsj0M4X
PstvrIPj6OKaekQO0zeiDTdfuZK8nUMQOP/KFEA8p4xk3wT3fb4XeNGRtYjviv/BSt9ubIOyXEdu
h8HqYQaEw+w0kcu0BTSi8tsUOo/xsRN4BLb4pEpfDDyriNc9QEUfRb8qzj7eZZB4xacFFlbyQIu7
uN1SEDiFVe9ezXxJbu8Xz0um2uoDZsPyMHHn1aYCCtMiF/ZDqzPoAmDjhAMfkrMuukUxYtYvtP2/
jgYPlVP732LQRGJ8jYOYwGV7xRNXbpi9e0/NZ16nP6x/FAURKhU6/+BCIcAmsoKIPbQZKst0Fm2v
uGQVAK62B1dwiPGDABQu6HGwjwcd84+uWzCjKYl1NtvOiNGfoNPdLGs0cx+s4Po62QzwOgdAqClt
WuTmIeSPJPUBvsvKZH7xF+16gqjfqoozESXhIMgS43F2UbFDaRRekqJYt7MLbRhC35ZV67NGy5rF
K0bFkvnp2Uqi2sAJmUK13Dr42YdMvN9N64dm+ZkqW00aeEURTwc70t9HbtdJY/+Go9GMrIWs39gy
YebZbBZNTYAchhcvNje0nTY+8KEg+pM8q4O7m3ThbjXL1ua74uZXCigkxN/gcfNlzxRJKwjyuV5d
L+BJHTS8702qAMXEgOYuV9TvWVvUimKqAftQcA9hhCBuQrouNOD2Coj4v2QP1ar3HlFSrDuFGTp4
R9yPji3IIEUkgbnoKXjuhM0FdmjPMLMAZYkZSrKYeq1oppEj7buENlCmxZGjWlD35fcoV89h7emq
UVpWQu/Xe/MWr9EOT5vr4VPVljFIBs3G4hP1NyD4qRqVuEgdQXDRQJqyDmgqqbG4M3XYtFfyQrCk
lYNWs//SZhhsaE6MBaVfErRzrgL2QYNcr5Ba0oe2AKYc5F9NHdsCIGF29dQsv1z/e1ihVfxRD4qn
LndwHZWvka/rn5xsQFhtKq5CihzE2gU+uFxv70q1E0nnVmDpn+5mBoKlV9FY4WdpXIUSGoBlOXml
grQymWhtKB7SmJFQmaYptzwZU9KZcw/jK1E7vpfsZa3cD1+Hc2uS92653m8VkfUxezl4q97Q0zrq
CkwwwSCsnej3LBOQdCu734ONwbW6jWdfedINhlgvVPvnqkoLalkj5tEE0yz0eTOas3iRulRu3RPd
stdqw3Z0Qejdy3CBfT5xT8nKzJbS3ebSOXafmqE52n2cCR4wqBzukHOnlD2Mvz5EaxA1btVWpCsz
3wvvOr3xkygGMWUkloG9/jHmxlCfFQXHwScfcm99XCLkLRUCNheS73KXqXXeBAAi29eAmcb3SR9/
I1eChkopEsHrMiVag+WLWGgLTxAh/Os2lidEP5ojcY+1Ng4qDzp76C3BbAAIqbNVDQI08T2MkTHF
t5gRIO88kciczlqHLbQXBQNEDdHwGwhEiWvtkf1Z5CrPme2sDN5oSiKKT8OWHzIQllDMbKLK4fRO
GM+exvdqAlHFRD/aT3eDHvPPDywwnvft7Q4YprIIM6G9FTn0uqxtiKb+0hyM8+pmZEOuEUggB6Kg
z6WEAIsXK9dOHF70HJlMURpM0iK/f0MfmTVOAv2nhYCsvxe6LMaC98bzTNCVC0O0zs3WsYHwYrK4
vxvF9UPYonE9ktY8XH3gSGN5ieVEICxV3SzI7S0JZjPzJ07qph7He80vJ8cEtU9abKebNUP/tO+j
hlZdngPMB4e8UX1c/fM/hioG1SfndkNeIPwH3VAcjjz6ogVpdr71gdjROFLSEWtIpyIxBYguELcN
UYntE3cUu4xyXT4lUYz/dVd1L/xa5I+k8bvo2o5Yry0Pawg4ABe0bmNPUfTXY7IlCtjCQQye6XHh
uXuNh01Vfi/iRkxClNw6rfO3qG688nNLxb+rb69PUGx1DpDZjYfIXfkkDPZ0IRit+WdQM5ouEHhU
SU7zDBvxo488RrDZMLa4g7iPBtWgaH2JVo2jgjCLhWTZ/e7or27m/SbvqO+f/IlPkeL+vSBFQEbJ
agkgfC6DZCSYV/CZYsUzreahNMUPqZ9EvOP2wr3nQLxeTPjRWyn8nLT7qPZtqlzWRhCm4iiIrfJv
4tFzRY/kdj4xkKLfGBHXFHaPBgPN1L/7ma29Y58xeC+QG1Nd+hUzA0xLysDNkrM4Nmv37pIiqdbF
vjntzsLzoeY4vOZgxshsIcdMosDQ6wsIT35QrFAmxEo2T3bE0iYzirSRzNDnPmIiEOJS9dqj2Skw
jtZlTCCdv2bFI50KMlSNsePwrajDEedaQ+nvdo5jDSVHXaqS0+nqqRhVrkx5PsdbUHzXvklC6CHz
Lszi/sMi34oUhnL4y9uFWIXZvmzSK8FyIsmqLTHFejD4+ytyW5B2r2qfOD5NDF/1TxZ3SussoizL
a6l0D3T5EILoKKT0e7w3fVVvuRR/U7mLhDBIm7CdwwPbzSjw92eeAKz5tKOTYsJTKONmd/LdyI8m
OqFi5HoakA4dNoD6fTPM+pGYVDRIrLN0UqEzZmS/NPd64pLe54iGOpihWxXs2TK1MwNQ9udiIara
9EkXK4C0ryAfJDC0N2+gMbiuyDqODsGGZmai8XBMcsmXFzEetopTYVQVGOVrl51EzN61XnjSsH0W
PNsF+CorENL0kpsh0a5IOn1+R/5ZxAOtJwcdPMyVtfCHHavocoxlL6GNZNg0pGPNHBqU/1pzXGrk
0PiezvySyh2dweS2JeLRD04IXM165W97WHcll9FiTnJJRhvjZXvi9sZSNpuxjrAUAZmcSZBPbHKz
D9gDA5od/i08JXMP4v+2wBSRGcaCaisJS/zUV5hxIwN6/djEpLX8cLNw8+Dn9y6dAgB4FsS+Xv0e
St/o8A+Jz2HGyGcQPKH0HVcULNNetU8sXI+WyAWItrJetXAQ7LTqbl6X75Dmg3BWWyah3p5p1hxy
0OFQUGUhWTn6L3TAsL9k/2ADpo1u3abEOLnTExOmpKUNFvr4mpNnyhhhB89SRc4LWUYejE+HgNXc
i6fwWcY023tyY1PUpTNnthiSFh6jKf7BxcjOS6/Cxwzl/CCGzcsokVN/PDtJSzCsjXf8AeufBsuJ
emRKo1y132snkGCuH30+Mypf1nQg2z6ET6BA/glU5c5p4uM1i1tvMjt2RAfeFsCSAiSa2UFwZScc
N9geAYidQI7CCzD5Hh99Oe7idsbrh5HqNlQEAQpGgXTnHMnDeb4R3gcf80nkmgixBi9xU3yAc0FZ
0DecLokG4LpPWP6ZVSJTAgmDPu0dW7kN6eWc9sOkoGc6p7c22DU9LMN5xtY6G+wTKoIqCVVqpQRd
YRk379y0LhI2jyvyGfbxUwWY8R132qaYXm4TcBj9k6QQcNiY+d2joSrljiuui3rP+kQ3F8whMEEZ
5EgMhAoVAVDIyln3QkudgWmu/BZo9oEHxMVv/LrTJz5Gm1dtpbPXlX4VzbRj5/wd5Hc6IMxe20LH
WWFvoKhfoFSIIj2LSvOY4GNeLQCZ/mriiuZUbsHudoupHb/hjxPW4EkOeSONavgSncFnFD/gQhNX
0ZPM0s4pwOTEBVtGS1A5YFrj147LIM3WN2G4lxINXlkiD3Ahyv9g5t305GckmP68QLsNujoatiWj
IMh36v2lHu9bOwS5J7jrQmPTXwQQP01jxvC1AtlG9h0kLz0EVMQnTWsYpFLWTf6phnl/b9M9RNFj
qL8mjwbv+ASwuV3KzzwaqpZxhs2WeylhHldnw+mzoyPGPt1qS19uTax3eE0zqOORmkcjbKinkMrm
GfWB8/2j2aA1VP6QayZUNMy/3LFQa8HhqYYLVtRPozlfrC5/qRCZJvzwqnmdCNzKHGheRpfUqvKb
RXTgqcpnpn8VL4Ttfrtc1DdoL0s4B71eT1/Cjylr92wUwZrN+90CNDq2jpQuqs8wZW0X2N3fPkGI
nWGqT2/Ez3rk0FGqS3daMT9f2HE1X7vYF/ZkJqk8SnU84KGNo0HTddezxEHF75CwCEOf0Lwwwd/f
A2BMuSStms+t0JMdfJTngFdyhTAvMjohGi5yVj9LowrXOf83/vp0g5fDbEScIAQS7v4/Qs3D70Ee
p6Ff10wHMnBMg5Rr0W4kqjPykbfl57gsBkgFmFdrAP71xGL1t63ja/etwQI9hAIL3v/kPLKD+oMm
4blTRXEDCkzNdzRdfdoeqUsdi7uL61WT6kKgNIS5jrjyPbCNeN40bVDSncrDioZv5MpbYmML11AE
HQF/giBUIQScfHTniDfRrPQgoU68+RsAD+jlhNazQ9h31fiSdn9IH22TjnZNExysurgwt4Ri/0lv
+iJVqXm8ZkN1BRoxzOMMQSaMveti7GXDIWriQ5b6sm3ODW99A0lDLKGMAxvoiH/Iv/NgDeASiIUJ
pgF4/8qC4VyFaeAQa1DaRQmv0YLkWqMv13ZK2wH9xpAwGMu+XjIUHNtB8Dmhj4WSPqQFuomVEbx5
6GWZRuKIPWXuZav1+EoKausMyuZ62zVD2D0Th6WYWUpk+HkbRbn1+NCT8HxY9asw+dryZZrIFNEk
T6ca+sP5EqWcRsX7cLQOml24ALFN817/Oy16wOoUQljLpu+aoBBAZ0/OiRPOFfIJad8EEXIKWv3A
kRA/A++FPFMmaSmbAjIOCSAP9tMKlzBGWsP8kJQI9R/E6gw0u1j5c8PMpkSz3AFIe1z6Tfh7/a35
v40mO5BBxGv2pHlA96+TV2pGyddAaIv8TUSOHLkR9QNt7OL5uNQYPJjiq2JWyAGKgk49T/wGtpr6
tjMY3tbtD1j+FZ8BaEtchreVx9XP/eoqI7IjTW/sGK2qfZjocMP7V3Qs3h69E/kGwortobPAdk80
Aq38dDZ9DkvA7N6sveN0kozwyv/BUG1m7q6kgRCTd6LiElwxXZNjqF7dlAAGxbKHuFFT/lgZ35CE
mgDmm+6UNccPlRhagTKyBYa3if+piLCG5KCtCYg0OpFACBl68iXtj20w3oZvsQEReBojws6GeENd
HOpckgYmteKQBalnwuFhf1whxZbemAYvBFGYHpm0gHXyi0xtYJ24m0vrHtPoYeZmVnfWJqdfNMLA
sW4zaYVlEDaWERTzyl4qr8hGB/qKdP0A8nwW4xcnj2aWjMwphDGC6gkkpuT3p1UKvKoZK1rWaPEW
BDsWX9sJUhzHJDw1Rn/KeLfr4jEzEqvNb6Con9NK0pE61AW8b2UHABXWZRsZGsU9wv6837Jl50T/
VKr5jIehb5olLUeAxcrbwFVwg/nNcN51UiwhsOnJBKne4HVS9NYBsAPB7UpV2+3hYkOhzbXlvnE5
C9x8cRus7abQdmvYersuCeBIFB5Hr7xxU4KRnT80wu4A7EP9x+nqKnq3nZGDalUX0lGB2QN3mQnf
Y5EnRJHMvURQqqomP1FhrOK3umDUrv1G/pHWcWTca0EsBPO5Oqik7g2Gjsb4BWsfPoiaPJJqn7hP
hSZDnpsoHl8fuJchquC6MoBFvbf7h8ACntVVxM5IUMEHTfgYlrpW0uW1IKif60lGUddMq5fTa8Sv
onSdQLw4niNlQfC0EuG0ViNs07IWaaghGT5usPvDZ4NZNq3NzqRpSSiT2wPbRIHeN8hVJu8Bnlej
Eq15/LY2vXXzLUQSZ0ykvvlMutjErDVVfA5G4N/xGtoTpMb0lNqkR/9T/4R4AHhb05bYp2UM+pj0
KiPpUTNIJ8svnjMnjA+vHKHXhksR0T/Hloe98emlictewGxLJXxI9sFOb2tOkq6NNUtTwURLgjuM
b3tM+/tp6y5l8msUnQci1WISsTHRWiufA4m/fvnHZiAJnkjfPQ8lqv2Ivst1yuAP3yMfA0S9FKH4
wufbQ1R164g6vC6TPQvlRx03l5Vli0k2QlZe0Y8Wartn8SXlQpcDtj85h4QfRWinapxzL9bC0Z1x
+jJs031ZuWz9L9VJvM3H9s5fks4WouPrDkH44M9yubfKZH2cV46mTijiWPG9afSFDAUtVaF+hQRy
FKgo+W8Bz2K9JmuVojkj6yHnF1yMwK0jBNbjcTBsw2izvAJwFDw3VMfOVYVJmdb4vbwuIX40Fjwf
wBv5a7zfgWknVfJ5rMQbGz2P0zfD6lkOJW/0HaQ/9ViBflizIQOmZxejIt/uQ9oDUknMTJWWLrIY
9AqzSxOApTaoARq0QnxrV/2WR7gdMs3wZieh1YuuDdnqU2dnpdHaDIDRDe9TJngNDFm3MT8zBj0Y
bO0ghVrrWCQ2s1Rq6wWsEyPslcNUrTEpIEYNif5ylDfSn2pYod0O7940PnqBXnGAnjigRFdp1GsM
dR2E5lg5KGRqr6Fgqe3XyrCnvcHI8FRuO7oB9eaps3tMqziHOXzKSyOOqsidHTaDx2nXBXe9MEpf
YEZdo/BEa7JOO8ncDEHKqmlKsESHZhHI7np8LMp3xav57ioIfOs+rhnKegJP8C3cZCrFPw4U5pFW
/ytD4pgLW1BaZvEbDLH7sUyIUSbXbWa+2iKUhfG0cGh/SWIMJ36cQXyW609TVSKgOXATocwIJIGk
KhyWVhdRa1HdPUGdLaFr72k+0NF/tqwUqz7z7qp6YB8f4VzdhHNu25b6ToXZbYPi1EM7zit1/oiN
yUpvjIj1o4JNy9FsqTYbKkLimxpSjjrnm7lU9pE3qwJ+Vk5KRvt6crJzAQIhJd9ZTFzoTwIlKAD2
ytyCElJZXaq2LyhH1c9yXKMNVFvlDXdb8iah7w9UyDedaD+u49KSNl+dBsbUK8t7m82MCLF+0RMs
mL6Z4GdPEesKBEVO//n6ELPGCbGmjasEkf7WNbWTpKB4pxLMG4j4BsrygaXVlm/h+sXrlZV/YZ0j
9mft+lv2ISy7EjKlekQl6aRwiWk9gSWuECWMMyc/flvVsB3VH8+m/8O3YHE6JJ2YqfjzmkKP2pl4
P9a8zU4QCBVAehglsuocFdLroWD9SigDlYNHyY/uttPzOZXxA8mR3EGN+xuaOaWUaRH62+dNQT/m
LaYNIajwYXIqpy7QcdtQt6JRAF8tIVzrknMY/S4Hfu/2UnfwnIbYvHAzsUATK1sxjLa0Dx/uCssL
06c6MufgaQ/Tq02XrCNbmw21d+9vx4pdjjLaiUACA+8yR+1YvbJWtVaJt3uvVgD+1SP+uunYHSiW
VjK8zs9lLM8OzrgdkDsDleMIWazatAZmjL8iQIsmhba56bPOpQkVMDUw+6A8IbmbfuIfViZuwGKP
utCED/I6InTyCW4sjZR+udGWLTRMDIYqfPUcaBhlJqqAhOSL/rx1xZxJSFirUxMCGf332w3nf+Ir
Ko6mblLd+jWPF6vnZ80/et66oCYhZ1pXlKn99D2F1ofWCvvirc3TNhzvTNHYuzOzFOKtJzLdf/Ju
4iR+kXXkq7zNcgz+2jTJcr2fH2PAVu3A3QFOHS79uYfPvHDKoiFWDQYuDlltCaZd3tW6OqMfAoin
iHuHR7Rw4M5PEl1C2frEIM9GGqaqA9WHQFA8iP4vHdsk3TI0b3O8UzoRLaJfL1CeO2UY+yLJ0a3R
ib8WQak972LyAB+c/bFWfY+Wr/FeDc511p9oxbWjiCsH5t+JzRChyMOZ61hPuBPd5sfsYenFX/QB
h9rhAmgydj9+rr/X0PAoAWljfUNW9xkoHD2cgzF8Ko3ScgBSJp5emrX3rUbyUKB56jKhY4NpKTh7
aHPPdyLIhJdAkbuORjNCzC0cXHm4R6Hc7bWFd6Lw4GWc9zm7GCdN7xwWnbQbKhh3u9xgROG6CcY5
8pytDoCfOZm/Vgm1iq2t58HrqtXimLe3tGXecg5OdhjhJxVMI/+Zpg25hL6YiGZVIqo7Q7RQEsXf
mTW+QKaMgFtPXjIpPUauohItqm/bD+faBm3RdQZ8qnrE+igbhgWmpTTlPuuC0MY+Fiaq9tGWAEjh
yE80xE8FRYSYGFc1VQrv5BuLgtdHQLxdigsLM/s5Vq/+ZgNYGIX6GYgbgGNOuiPI4/88KzzopvDh
/p7bfaC/AHSsELgrrDkHrczsjqRCgd7+LMC2tFWifK8OOEXAIu4qBuhcPimeYoQfnCwmjLpStVd6
gw9/ZwJOckZUSkFlGQKLLK/WvcJWLcHnXL0KY3GCgrF7Ac+HbE4+1m03K5ZpN1mYuxIaYPeS9NTK
fHg8bSbsfJdBLNa3J6PQQvjPWi6WWgvnoqw/LKUCrIkVmXK2V9Y+0De8c3AFLzygaClwfcX0b1yw
inaGUZuiuA5CvVUYk3Yh2vyTd0UCJw0MPbYB13tykSuza769PRC3LQ+ibaOIY1xSc2CjlmpWXpD0
BhEbVS7V83AWESdjiXszDXRUTo+u9yp495lr1/IGMttF2eDN3gdjZeOfYlSotOXsFlfLyTOYKa2b
KNXazOuJDyoBUK00zqgvDvOd+ZnftMcDkJgeYTWsfd4Wn/2MQ9tedTGTxGDGdBUOLN80wnw7I56s
sW8gcpTBAvsm2zYQc4maQWzNUxYXh/2ARXpPXECzjo/sYq8A65+vwJVeeBnR8R5UBLyiQwe1LGbo
9GwMWNd7qQUWHsI4Dra6jwn1xrQPq5ulrf8BbJSu0POZ6/x+7jIeGSFrgUw+WhqLyi1FQz9dJhZF
pf/ZjQiLD5krzivfCpBTgbzT2JUlPwTipcDD3SF7pQOgcHPXXLmMLxFGhdpDbq9KwHcD1HZjDT7P
19QEf6cAQOpBVIDUgVf4p/xLx0B+smUWKv78q38AqcEzu37WrrI3p42Kh/d+aNv4cNOktjCD7Oeg
Sn9YO12gYpgBIWGEVbQR4GyrFC53Q2rrH21h4rEPpyzJEln5J0KYJEtADZNjQ50pwTOBwuc5X4jZ
tEW/PxFaVPu6FLZB+6oz/tiMrx5+Vr63x6sisPhMhY1Czt2OwYGrYUKwmT5w+cmUkmcdRfoDp+WN
ez0jkqymTc5/i72zg3zBAQG41rzz/QtRF1kykS/JN+dW8XscrHYMZGmoOLtFUjMvhjek3N2Pfg2P
rGLEw5lit7Iujd9E317pbIx4RpD7oqIdx33c1x6ZEstE/9OHYKyr0d/m6IKBehCZruPxptFSxX6f
n0MtJs7MVPrXPaB9SJkZoTPLjiVK4Kxv4YFtZuuVSLazdAS9m1eHV8O+y01zeMda2hNB/SoFdNm7
/HV6HTbL1+9vHn11HFcezsw8SADV6yYMJ34OV6iPJgyxKgdS/AxCLYSHAG1EAkgDBnICWfLo/6AY
x3g9Qgt3WQLWteun3a5RdBqW+pEqNr0yTxcqiXqawfHvb1Md05U1dgkeHAGGSu8bxLLbHsSL6oBg
DuBchIXxBbXrfGOQhxs712BaewyFY8R8zukst95/8otiRxNaveQOVIxfVK6CqJHbs2nQXcBMQiOO
3d56YDslZt7nS8GGuP3oI78dI/7IwMEkoZWYr6UyYs/u/2A/2GcbCBJPp/lY535D4MhyRcD7n3ly
YikUp+WHcxTH4ZnA90Rjw2dd28XWulMP5DQKYwtymzuM87pTn1dy+ne7LwcfyB8V2MQI2swT5O2r
b72AiOJDM32nVIvxXdqnr1XKqpzmuXk8SDPO0YLrezVQwXNKFy0E/ObKYBdwicBFnFrT10GEHaO+
vMtiqu2g1RR1+OQ9z6p8tqyw3LSWeIcmCaNwMOVS6o37DMT7LGt5JX6mUm3dh+1jzJwBsTtJeHwf
EDfneghe6NbSRD74s/hA1ABE3G1539Htvd4EiSARJNVVN3DSW42ujP0hcaYNiT6NQrhB3VqdE0QC
7AZ05nUPEKy6DEdFH2pDVmoZg12Bj8zs+rSvkcCDAU6THK2FguZ0PqvuxvS//PYKWS8raWf9bcmu
2fWlRqJbCe8/yAJtIIL6n/yI34IzR9yD2mrr8sd6ig6u6qJNyDop0wmegCl73ynvMeU0lEdVBa4f
j4mZYlesGKAGGrXxHwaTkGpn+HSdj95OcNm9GVQIzLBx9SUhVt4pfIdQuwGH6oeJQgiqXpcPrVXp
iMVkrVvGphbVRJd4qobOwYmhidfAcmyxGPVBgGTNUAfWAdgz/jNLRbDKOj2D+mzxlJudBCbHEuFR
9DqTpGY7C9ynhCp6XZAb/OP/mFm8gK+bBdSbYjJJECD45M96+7c8Kz3t3BnJe7MD2xLW5q/UjtbB
hxhjz/u8FEb4SACAwmUJv8VUvdZMaCHGGX1Gc5i/rZlEKKDoupbXTNs05PjRg6h5nRdZZBcihNiS
n8cwO8c4NybgquO9aNxYWeDLShJxER03RsKGdMU5HDqbGAY4LnLkvetj0TJWoVViymjmx/h4aAxq
DvvtWAbsQOH2ioDzXuC+OTQlUx9vfKipIOLJ53TuZjCynlkrvBf6yJ3Qp6WDZ36qyqkIpFVPl+oP
JVAJhGTY0pz2z+yQYOwAHOd++ggQvmzSEvdsvyhe5Sd0L7RcM/cYCeFxbK76zqf4njezY5N5HvJX
n48vFOly9q8IEGE+YC4JwyIXng1f+0JconSQbQ0Rr9hUnFaILR3LNvd8S2VgHNZTG1rFNeASB1de
afG6QT8P42TAb7s6GZILoZc9C5wm7A7K579sHGrJtEtnFlbGXJWyI2pcLMnVb2JK1YsWDDLag9De
TpfMRJZU8yXYlAyQ9w76Bx0b3dAWYSfu889g6oFpgzJWr7SKnJ1IKrmUetQzDqe1/Z2SSs8gT3xy
7TdRS1p+DVoGH9EF2IHuH8b2EHdbxRam/jzFsCrlRqWoDyekon4JXztPZnFMM92gciMDb4nJQUAI
Ez+6kOX6xIKfzD8rYsQnzAZ07QkX/cPjC0LxptAEw+FxiqpNgycd3gZ5v+4xyDAYQYbUjFLhfof3
r/tgUmXXraOXpbacIrEKIpbA1OS9kaORtqR0Qdfq7ORl9W3o6CfcBzxf7aOccPPtUzq0zABffPzF
xA05ADPL5sqN2YxRFg0wE1t6loPqIT/87Q8mlYgwAvwFC7hwzdrwzEWDOMWkNcjHdcb9p4i1PCDq
IZLgsFCf4IZrrxHundMS9Xe+WBKBySH97rT5oP/kJPsI7D+NUqNNbdI2t0EK6/vMypZ5q8d0B+Cq
rA1e4YoUaRvgLauJfnX8Us1V48ozU2xYSDqUcqMKQOz5ZNFQmpHuFdjvY2e6nNWb8sSZV4PFlH1k
l5IotvlDGe0HFQXOGyTfi4wPRLeRVVJEs0M6MWohuDxY0xvbVLC2Zl0Hh8CtTaiJuLFglQQAJF34
sCd1Gfd8NM2iAhS/2jvccwj0qfxjy+2tqawmGbR6X+2oAF0BTMLCS+5GPJ85Ce9cqjjG5OMdT58d
Tczmbto04MSVEm23qmdXlyCf8umNExf4HdmWpoTZaWRNPJ3PSRfRXSAmK3AQjdp/q1qUj+IvgUWh
BMFHSPWdR2ubmW8mUr/Zvq9ulWMR3XtF7/d2nGWjm9sBmq/oUyNWLJ2rOXaZAPrUD2+mS2PtLko+
6gmqlKnfvBJ379QwG0zKihypuCjw+2I2QxEeZxmg29I+CSaFlsruCoQZrdulUv7GUwNgv67CLSNZ
8w9nIcMG6iN77qYYLIpBRT3gw9r8FHZ++RhulHpZo1eoEDhaSpzhZm4NzFHbzbtshaTvWX2IGWY4
ivIQlTfhsnKsivrR/l9aKr43ppjjIdrS+GKeyp4/nWIadwpo0nPcXfKP9p3+bSHZVGeT1twMldg9
KxwiB0YwIW28psm2iv+1thQZR/jzoAxQ9+KYhg12jZhjBgmB/fWDvjzJo6GQvY9cSHXgkr3uFBvm
JCDG7ZPb35D/XW29zlHXptu3wah4YpxdTpVKLiBcHOEKCaRxhWnXagG+xzKoYW18d2dEr85GfKNs
I00n+JHIvFrSRi6gmGPwhoUztbNWLJom3oBGp9c2dyG5eaUFjPMY4lvMjN11ISR4rp9GQDgf9zKb
8BWizTRkuMoRlHag2EtA8GLuDny8cHGjD3T2BlcwQH7xWhmgz960+npqte66riY2g8QXeLUKpx8v
Rv9EqXBtUfPjwIDhVA4ts9bkx9D+TlcFeb+z+1cmH2XiYFSa00l2vlDYGuhY4rueqMMLA5pa1JAa
HkgLamkzSVgEqGKkb8ycbWvFG1TrHad3jN7KWobR+3j2erbFjyNF8iGgR8/+Eu5ewez/YbujxJFz
RRjBf4vr/Z0Y1bbDiVm5QAi/jb4VLjjTKaaS+5WPmaZXYkNcjWlANMiUGMJgPP/4b4wBHj2KlArE
wbYwRXyB/FRztHx9C1SdOG9dkoMsw4rONPLTPn3tFd4WS9FFpCGVtm36AEr+XoXFnh/ZSUHmxEXY
l2U0xTn623OUgntrA0Az8JY5LGaFiqAxJaTkco6ZwOy+nw5+Flpe7XW03KmX49gRxiABoWDQZlN6
BPhgUDd8EfjG19pwH65fJJ5DE4BVvtY83FCXTk+3hmCORD/Mr52C6vn6d+hf8KwpL4F9/9SMz1Cl
biyL6KBGflEVceteYSylOC5KumbKDiUV1RUFAkFJRht1mPsxP6EZGhmQt1ydBNPIEH6hlHXQy543
ZDvuJWSxbuqRqBfiKu0BZJhYokx4p+Od7yON0G05s9+TPkB4YYfQA5oIbocpkvQWtzLujwBekKmi
aOYxeDs/F30ClOobzmAtQoZsk+aySxTB2DZC2pO/SiyaZU5B508RPUa6/Ibf3hG3cudqCS3ldoUN
Y79r57tdJvBbs36hi7L8EwE1sDENFgYQtIfRT+qCXDA3JvmZMPEMefEYnw92OK4+lcHY0DJ21EAk
1pr3DJaYtORXb/tAOi3yGEQHK1A+KNxhDg/0ldCTKsike+TAoOkMSvfE2BPzI25Z7zKLAf9jDw2D
HnZIyJNg2Mq8gJgzXaZSa2efkT1col+/XwvsphfrbHpybSDBj3+f6oyonkuTJ90xxu51CBApLYdF
yPVLFdrM7/e3pNX/7fW0gK/wRI2ZRJrwp9PHVIbK1wd74z+Nqx6fNEDb5CKpXOLziKLS/tn6c8L1
oRLUJtlv55Ms7L6SiAMojAOKXZILmdEtFl9t5GAVsOGBFQUmQbvXhJeYC403RWTl+z78vffNyRmr
fj6FZavPfj23Yj5gZLbehZDPxzQkP3ldsjXrZ9jKI2KVRvaJUW7YgdxiQgEAj5lYtWvyVtkr5et2
yEB5aEpngIi3+kuH2Tbde54zSq6pgq9KOMBTVKwwkUoCp+jcR7e5aghcE4H/qMtQS3qQ2UMvp02r
sGbQ4Zgz4KW99s+dyLWcvJHW1SIkC+wLsy08nwE7D4M4wNoVodmQZ61sbyrX1cphQrVSWWQo1iHL
P5zqUlf7/26JNXikwZKIB5bIPxotXHOEQ7kZtEMq4uqH1W8raFWIZd17nN4JLf3emJhoIX6DhRY5
D+DYkLlKbVwGoYgF3GGn58PKoBYNvuyyQnKDnPkdlPNHg8misdhTUo1+9Pt/wF/YzGAhw6IoLgFk
aOOE+Epw8S36je4L7hUbhh7DhJWMu1X3MfV3lOgspyaMwJ4XWbceB/zXNDcJg9EIdzkCCeX0+cp4
HPEYs6tbX1VR86H2sxLzIdrgQsgKAuR58VVtk4eH3SthDQjrGZkySiBOXLAHCApHUS7KoWRDCqFU
WZFNXYbka/5xiu5fUisrMw3rhtFlgmtg3gdwkoPDQMu/KKlRgqVOhewa94I4xdEJCDrYBlYo9nNR
Kq6jLqgU5l86SIVszMhxJ055hPlk4yvRLuKUOJvhULHYj80HDxKlkRoB79aE/A84fIMIfnlpJkhT
uxyw91tXrC1MmOyoVGH89j/3Da1XXO1o/P0SmOU3ScCubZ7cGjI1HDgzQ9e7TqKo3CY8/X8HPpXu
P/OQbgf5nDS4LDwQ0rpwVKQBx+MJQw5EHLzA5q/VIQoS7658YV9/k5NOSzOionG6PO0VEHdgN4lq
+zRJ6+vSFp71BUs2rNV8Myk1AyRPSRu3iNwuFeBXZQYN66q3Mh3Q2l5SiWa/pkw+rK7+gux+FjhN
9JhDEPIk6lrw+7AWZ8Ws+CS5drREm+3WZOOeBGNhJjPmGcIuzxyPkUWDE9008shPuIS2Z7O9W1PQ
hrYtkryrL6iSsbemaFiWio3IP9rgUrIgP3jMTHqVjyIrW3wd6S+76sHp039KxlG/17ftYLvBf8ya
mZyYAMq1uWYRDsOEJhWNMzj4k9aHOPyzJRtfqik3+y5l0PSueLl+LBHdIAEVJL2BoRiYj1AMwt54
YyvGKXJc+hrHHO+fUxLjGZPcmlzOUIi3tWO4FgEceCK+FE3zz74LlA2LHhrRM2TLmL9tcxGXAHTy
8c0ydS9j5vmpkycHKvKVR8XYDVj6UGo+CEtAg++ta93rc/B11HN8RUwSdxk3phA+qQl9cfjFeO3m
NegGA0iP47alT8c/xo/mHhRNKjHyKU2YEOCK3xwc7Nc3dXr8TYs2bM6KQNQWhiI6fVR5POPQeU0g
77ce3l5YBnrxsxtSh6VNKzGBO3mpbUv25tJk0SLgOU3Zop3cThlgVm48fjvbPrJlvjwL+nDDigSB
JFrwqzSwSxbedYvYDXfr1RXW97nXbIMu7F3Sqi/ipsVfc4J8c1ljQCkLyt+5pMvskGBIwNVjDmt9
NVanhL2rnisfy7e9dV48sRuG3bnXnzwCB0me0+835vbdO0pMhvVEmQOs0bbOMvH9KcBcxrHMWB/6
XDTjlV5ZlPtXMarsdhn9x8q4RHtQ1GQeR1clJohwkJBndvlNADop8bNDHdmOw9D2yWcR3/9+dt4+
RlroFx8mLQJoOCJt0iqKpjhqLgMTUPLdX1VQTYq+fwpq7J1javyhYQgAj6wthb1bOL/SVF3Z0P6h
Jq8G3GepDOH3SRAxnHBUahbPMCf7iX2gOydDvYiJfLyPQusW9q0MP9gyYsUft+LD7bjwX2z/VOkL
qeP7NjxaUGdIDZRsuYeccRupjEavZKM05DEGh6veGDl1k507bQ5jfax6UcUiW7zE0d13TbK0utsR
+yt3033SuxJinvAc6SEdqndEBTbNGGGZFx2p0gcfqBbki92TbOQTm5ZlNZaRePqhLoSQ5UBYU8Gv
6b53ZVXYeBq1vbqiynbGnwM3uQLkOMlFxoHn57g+t0JNcvoN3vhfSsyeVAA5UGD7M6wgxgkyF6cD
dWHDKNv6pfkWHSOdSRav6dtrlbmCZqf0A7Yk3DyShysSvPe2wk8U8Kk0gzw85qcT429nKRZsJh6/
JhWtHDLF+kKB50bwOFOzkqnxCWpz5ofRDEqIh1eu1Cp/o3zYeaPxxU/RndrpQa6CA3LkBJBKWMoz
AgzMi8OogsXTdRe18Hy3qOKpEaorUgSvdlHGTt85zWhaCgG2amfJSKqPT7BEu1Di+LsELTKeU4b8
q7/EBvRCmQ26JI0KYlOX0MBiysnhxFhRspw+nlDT/R82FVr1HF6ZpY01piQiWFl/7K5hR7RAS1Tu
iMSb5NMiYoULWXaYz4WySRuM86Ld/PQTuDC09trZKu6m2Cfa6a44404i5CZxMumMQUeM5B4yMmyH
p1OiPZjylp6c+eIaDKdAuijAwiBQ1viUBuFXeGbZtDAVj46DRJYMBAw0Ycd8V3+p6HLr4QwmI/KE
rpbA1hdsM0AT+9SP/FEsRxkTUfT0e9z0uONY258Vh3Eq2Ea77r7wcw/DpJVWDfWiuKtRgB+n2Z0U
wQX2oDe2EC/94QVPcRUtxzcaE3BhFHePRgiInWhgo+llWm2DIDrQ5fgBfEKtZuSGw2TJDjG7AhvO
qU+yRqGZhvPkrmOmEzVNRt+TZWsnimEMfiCgvdHJ0Wr2Xxjy76k0a/iLZfm9QV2mxlzjSv3V3Fxw
XxqB17z7KL5TcOwD+vgjKXaR7IjQTzfGCAtOoNMs5E2FlpLyOrhooD9U4ZS1f1BL0DbtRZ+8ZdU7
DnfBXTRB5bfvj4lBz+dI9Yv0CY4kzsw+QX95UW8ZOvya+SCcANftHueEvA4WlErMfR+qHrPy+pVh
81lRunRz0mH4oBjwaH6ywZzSkjkr5796A05C7ipqL1Vt0lavCxWbVRFJ+Vjqms+IW6bNoXQ3NM2j
CUFtKOVQxJS1AGKtV9T3+Hh7a8+Xgr9PPIwz04PuyMZHvDtchkx75wByuS0n6nvhUX9/8+4/z2YA
BT/2NQg1RXQX1vOLfAblFBNSWaSvJ3yo/GRVoSHtxQroWVWNmw84Y3cwlRzG1debO09a01o1T32Y
Yszxmsw+BCTEveoVm80wPA59qWIqutMDzQHaNaxcaCXZnU8MEOoBG2OQumizB4dyz4XoqMWde8gY
s3KOZh4oBOlVtez+fD2H/VWPGRnJ8EQ4rNnzOy+6RwXdjG7wEdcHAStWuED2D02r+WD6IZCNtSsb
OOq9sN8Ew57nTxG4B9Nk3fjKYxLsGcSW+Bql5o8MELeZ2y4lc+wNzRwvwQe4+L+rkObP674suxgo
PJrZ8d2nXqQzoNxhawWkA/d925jD6NX9rl8X6rE2OlC5n/cdhbDIik/0Q1LQEGtIIHdsIM3RRs76
x7VqkwEmHRz1CDFeAVvlX4J3kWDRSeYwES/fJBZe7oZVMbmCRfcci96iwyDGLkGNNzhzMVfA8aW6
YdJPxPsNRBh1XZLmmF1zlfn/zqP67MMPtBbH7eyZbi07VaogbCkmHEc9xxDbRFKJPrXcWs5l8xD0
X+Ebu99sCd3DRPOseax3L/h10GrR3U7ZP9Hy6UEbvfdkBlTVLFV4GhsWEdXBKYKNLNJaPClF09c2
59g6un9iwHBa4f9/YSbx1E+Tfx3QcpVOKdf0BeQ3z+ZJBICnJ98kdXTWbD3a61J3Xn+a3zSPnTjn
QeVITQVJodxWo/sa9QDhGBnTXxNkfcYBavds4XiXuFtQ5RadwI1zyglGpW+Xy7pPyj8LErsFqKQ0
HRUyrBLpxuVFdeLby83BqtGpNaLbu1dbXgKN7Pe28lTWZrzS49Zhtz7UmZX6LsKddxdpCKseooM5
oQLeDgo03jPDk9U7hN/4vvfRUTYsk0sLmTJQXop4MXQ/f6E+0fm/QkXx4ZLJeW/UsR3sNDC4MdCC
q+vJfO3kRsAlOdHGdw/bDQ17FLGQTWKtilXxzONRLlBQ8FWtDxmrMumLEKrB7PNxlHkxTaKd4TeX
xo9jfo6Xt0urJIbCHrMQOAgleZrPJSe3CPjRnZBzIyaNOmA7U6Ti+aLBPIJj0abWFLy6yCrJ6DDI
fmXMh25CIrrghcz/snf2xobc01P5bm70w0iNEkyIp/sJCrriHpgNyb3p4B55tusQ8E13j65GizUN
2l8mueEYGlJdhXRAvkhIiFCe6eb4ixP5VrZSRLeIFEUJKefi86rodY6s3l78wDnR10sAIOWqgyjw
TiVqvQbV8XbTSiC+YqWcHCnXPxLAhcNHhlf2HGwpYb0sJCFaxx+QE20EtXIfcSBGjrqSjneJmEon
5iM1P3qUL2vbaZH8Og6tNI6gUFe95stdGQXk5AJPDdqwoxKHmEfsv1AxT1n5LXyDgElSN1l/2mtq
zhXLuMhcTq3Pt5WqtSP4nK1CC4Q/LsXdjMUHdpagulZuvgeFpnVYHCUrwvwmHKJS28+UhVh9Xg6a
czWYElKBRQmBW9jEIeWwWSVmI8cZC5YHoTEZylMJLPXGx3wvYlB/Hu68KR7bKaF7yu4TrRsCqV6k
s8FQ7kC1b25c0jB7MY1evO2pC4DwqOnAnUCMiwew5s7jLrjx0L5OjHj+3G5Lrzry16uAuQCB96Nx
9qWEghzqyRq9RR+EgDxHK1Ba312OVKJqKeJzCx9iVvdEzMDprBwxijR8QEmzKI6BzaQ4FFHDQGp6
8iDCLsHzQWyVaGcTzOWpHt7KqW7b6dGtPRAtkAul8ZHJfuKCsYSUQpaC01fpl8C4hWSqN3A+4krb
Z9ocY8va6LVEmQYH+QbrvQOQjFsm3YQiwvfsCGXSimVlSQdUTGuuYGASaSD01OnINr2lWAz1XLgV
yyFD5VjoIKorR6FS5PJv3ea5QEQl2OlAwAOx4ZU0oSll1mnUh7fHuMdrZ9ow06PUCpLu3CAk+BBL
PA133IyNvO03W3F8KAmhjZ/SEeNC8n7lT6dHHhoQM0R2YuxYb5y7vJDg/4P0++92Fs8YzBv0kwzn
OQRqFA6VaJfUEE7gBs+QDIJhND5SyfKXlQiT33O38gJR43cU2bszGkor0KwggsGhi5SRFUOu+BLF
GE0vXZqDvtp1AWE6HO0iuHzbW85KylqUjpF1SaHP/HRmIKTbC/DlWntl/z91sZedzvYBgTmSYR7S
38e6AW4VCXJWCDjg8asxpSs+uJ6MKGm4KyVzBvvxQxIdh+ssLLjOBwUUY7qChG7iwHmALNprvMYh
1QIcV0xQnLEC/bwJskL5W7avV0WO8ILMTyMuEUp715tyG6kALOa/GZop0T3nhK8AwGdxINr3i2uo
mpWAXT6ZdBVEAzuov2xg32XM7MJBCEvEuELwpKcbvTDrenCsDTuuAnEUxLB+s/WyAHQB/OavXhrL
sobo2eTrXSGQLLnTesKQGo+K5RkZiUoo34Uwh6kI/1vW2IIiHdf37g92otuGUjx2Ajv3sMIcnTJ3
1vvm7N5zhj/+Gme8Tm76l5g/GDxY6O+glsL3nFCZo5iB2PK4JdV8kZi447+19per8mtI2COwtsvS
7gWeolJ0Monu4uD6/+FcteQKtGV7ai8yo5y6yXqkX7kXO12oMAMLwhND+IYa6m7auH0iCbHiDTFK
2W0/uTwNeYx1u2yd0Tu5K5249b0QKOgevFFtPTdSJEmvka1fulDOGWWARn2L2H8o74lvi0jTrd3b
MixDs5fztUCb05n8Jmgl/u/A30DeTRNB1ohLyonIJqvyIGYa1TFfFLk4mjQduGpuucYM8+N2sg6H
K3ydE/FgCom2kvyTSA6cgWtJV/C4Q2RjKKF+vO/WTbp2S6dwbLGT8EwQX4ujlxW2rNcihNrXGGwt
He132oq9TNM1+Q11tuSARd8SJBH449VVnGLgeWzQuEi7mO+93ElGI+tvr9JYsTQ9/7nUhIYl/61P
9z0AiD5fPI4ixcCovXC1FaMkGyGONxxHIIDPbGpeAUKLXoe3W78Czu5L2l1efo2pbiR7dYjmZpJ0
10PT7dX0YNkAlbZ9Ryko/yemm9qjObXNDx9M7Zu4nNyIpy6CurPZh3Ma2dwhVOefXKgDZHbwfyBy
Iu+il60C5PdlocsYG+NVi1ChSeZqfxedRVjNOohSO0uPn8BzodWFLMOzSh0rKJVyyjn3KgFL5B+T
Fof7EqP/YEMo61yNLlA/aiXSKL2a9/JBeuQ+MLBFz0gEGvcb9kMQ+c35QCX+0r29bqx0qyPjc9h7
9QSX5QHzXP2g/w7UOxOlZME4KVvW+J6+yT8dsCPD6Kv+K153MVifmx/XqkFJ2htS0pnawz8GlrG8
4b4YbrtuZ6WOfHSrQi7zozv9ntuVTkJmvZmoCeCBgE0RP8MpbfLO+vAB/X81DtkHk29zxPZF6f1e
LFqr0MQWxWi79Uv4R/POVKD8+PDq74fIA10M+FIFtQy2atc2ZA+BD8P6Aki5p/Ld3xzKGpPWy4rn
eUUHjbXYfo1/YxlqYxZR5uZkf/DELDMf5MGlNvoxe+hyavlW8US975xdLOIoh2x5gylbSDGHZJh9
2XxqRnlKCy0x/53s70+HzqAvhkGZcacA6weg+38gFzCVesWd2wZLM8c3UeJxDj6KILEU7lp1YEXz
C3Kqx8WaQ270N5PjHE07OjCaIm3UGc2aa/JNB1X2459itqzQcvuWyClK5jo31MjGPeZijVl4Xda6
7ScHjNlNn0PW9dHa7v/8p5SeTfue1FBn1bSwj9NrMlpviJvnZ93Q+W+5QzsaDYIWX69ixYx/K0Az
Ws2gc6aAdJTIIuNysw+LNwGipeXkiA6NjczpPAHtmENCHUH0Ycb8Ee7z+VuyDLghYTEPw6mwS4UC
MvsaswXcuB0q32MzUDWxSc3YnJVDP9VuxWNUVvV6uuFfvcpxYyeCXWF4aLfj5+JnGQ7XlAnEsHa+
I3kVsy3a1KzSQD/DmmrCsq+lxHQ3hoG5aUX5/CSpP5M/1Th9LRCMRnPA6jQJpUIBDk6r6Ba/qzdD
eBzQHZ6uvi4VC7jkUY6Dn7+wLsp5kLfCez9WW3Vh33SLJnBB/Y9jcySCwvBe10N/SI9SMbQDWIF5
XFhxvc574KRnuVkCOVCXlGBjqy+qQCPVCzKTuwmysn8K8cUZjvQbZ3zAclYEkrp9rTwogbkHFyUe
e2Z+ti9qfLZxMjZ6HV8HzcyShDPy1NFaoACkLnnIP4O3LvthBa4dtnEJ8MmMzInzjPp8EyggeMLF
5FWBhGhfm3ATG8boXExUJ8Ck19/e4DrztNn9HQuF1WDqLjDWNBRPWqE+PhH4exBpmZIGlHishsG8
cv5mzLUr3nHIt0HOvRa2Oa4N+up0OzqtQWfDN7zbWp+aGER0iDkd4Uh1G5SYLf5PUPqRrMQtdHZu
vwrt+E+9urcXQActb+EMU8YYM4c6yfQmbs6sgoFcb1uyJwRX39QwfJP4HJdfkjX4kSsYYuJzYod7
OEZyexNK3+izKU9XxBpOhCUz8Ux8yhJBTSEJAV89W/4sIYtQ534pzwqrG6FN/bWQN0yMcdHI5ta0
VpYfaKBgimY1zMpD+yKrJzPqo4S++LDWIR0xFT4eTralTcC1KBNa7KDG9WVBbLTNoxFhTUhdjP7v
7aCaxd3YBboVgCzSynNPvhV1Z4jA6yOvceJ5I6b3KrUltO2XadC72Cf1RqcaRtrfy2Hx9v2DTM5D
kxHY+TQfG8Hq1z5VXMdcUsxjZfIURLVBJCyCqQMPwt4P47pvmPRPoS9sqm6WXNS46oNuvcHmXVTE
VDXe1hVq/UTx6cH7cp6axZpmyINaEweXwE4As5Fbw0EakHD4DZKLteM1aVo1kv0gTM+iXf9pnfuX
GnnBBqvgmyyHSBoaZCComEiS6iJiGKDZHbl4lkN8W6gEMK5wXm5mDiO37freAyqBvkvVHy8UuJVl
qTBU1NbEkkf3ZvwKJyiZxkx8EdKH9c1zDfBojNiAvqigIiSENq7xODeKXp8gAmqmfkEczTTXR0tl
NJqo/aMihYaSY05+BzIUHbgMWk15/pnpi0YniAG80pVzje4uohF6VWNrsAyoNSWUTOCP8SX/s6l3
/1yAucogXeZd+smWo1MHfzNfQnPLa5uiMnLVrK5gcS+Yh87bn09pii1fzM7gjnbFVbbHoxapoMiQ
a5H2vO3Yj/jN5S4G1lbPOHGElP4kQKZUyCBJiDrklE5SUZOTUDE6TnElEY0JQDLH9EyePt2j3/7R
7kh2VTZFtD+m0yOl6GeFr3hkU79WYNWGSXxevBKONUxF3bjIBH+aDanhNzlwM+IMtGRTIPhJpk7R
2UiNkwAxpzc8qvmPO+vTALKlnk/zmpnAONIRK73rglTb56kCifkkU9/vVlWHKkz4zGIFec7QxHUt
HLOz8CaAq9k96BrMJZaxuv1hy1sx+syqLQkaW8d8nx46J86jGzAnvp5qxI+Ih+7cGU+9WodXWv5W
UtJ9LN/afUE5SSYyMpF5mgKBIgnRNGvnDtx7LuaJlaDpdoJWzn4x/V/XKYkyeG8yr7FWU46iHV25
BioVM+l9rYweiO8/2frXqxlOPMJe3CeZ9bDJjZ/6ZjMPI0q7CtrX1hqadmkUAcem77e8n/oMzr49
WFrhnuJXMMVtGn8jXABf0uXZPFwWt9bOlCv0zmq/JzBxK9b77iOSA1Z8GLyBd27WVmTMQdnKi1YU
5tQVxIy8K7fhepDmlHE1Il3zZ0Z9tep0IJ9jVroWrHTyX4WQVgJ3uBgpEimo1qCC1liudJ3UvzHo
Vdr4FPuEyikNBPFd95NR5ESdxAqc91TMGSkaWuLBF6iNZkA1JQkAh5G8XMAQZWVya1ypYPMwCL7O
UZ2zeAfXIy+687R4AsOoZsG5Bo9mgIv1JbFenoGnh0GdLpk3blJIbLx0LmRjQwWZDruzgY5ZIEIc
I3ve/ev0RFsf8zPYKvhc8wxgosme+kkB/m+XfmUUlgCjDvzrffa8cHH45ugWPstLQNKCIBQ9OjiC
BKW1BSPCEr21GJUT3s9wiNRDRWJtxveX8bc/QupRLPbhheCEM+Q9gpgYeGRSApasBOsmmKsKM9lK
AQABJmgHcSkuqJib2HcZK+1koVsFnV0m8HD5QCm62cucYr1LiCM5PtFJEwHFGoqUqIAVfUwTul6X
+988bgbMXdGAaupwBUYqtvz9mEMbUR+HhC2N00zcRXMGuZpHaMNgz5A/Y7QFeX/7bTivv5PnOXfc
vxkBlvjh7dBnjUUMI6q+zbAxXTb+RFt4975L3k3dRcjkx3V4Zd5gjsLZT8VTqb0X+tKBSHO30d2r
WkvQwJLQFmXDGFRy0ns/pt5ebqAYNB7bzXNU/SUWSmXkFPbZXcIBYf+fR6OTrqr3hPxLV98gRn1Z
aLad++MnNaGJgUZv56fwoVus1Cfgk7nnQ9etYhrrH7jXhWHYdpYotrls9Cw76wnBppTAKv24C37V
eG/3sEy3Yn6c6CTG4EPXAjZ36Fl+Ec/rVY1q9qdxkaCsjpo1AGO2zz+7PGhfbXVA0WYH0MWWVUnB
shUsGERUkvhTEnhVquKwBqdTHSpQSUgl+sVvFI35IZJ/RS3uFfQc52JE1+wx6EQLehOXMDB/LD3G
N/FwS/d0FmG4/g3b3ExXOshJ9L3DWH7CnatIOz7/EheWXs7V9TPKT1O17NT1ldQSM94bSp2OSQM5
0pyTOymdrxB6+eIHoOjqZPKcYrv50xLY+U5knm2AOgkzfU4l+RCVp1iJbbzw8c6EtOk+PY+KdHy0
0To486g2E7mwF/hgiGnfyk2oeT01hLFQFiH5W/5h3X3hj6k0Oxv3wYRCZOmSPJlT4UDNJA3hcaS9
zJpEd2EFPPLofzRt+WeDm1havdad7OW61qtVTA6m/mUg+OeoRNSPoju/auTCx0rmBkWxhCdw46gB
+nooU4MsHARijEPkM8q/euiM8xqHoqpEVU/dHn6jlFl7vJx45HjmHasqSG1ywRx8o8A2Hg1ZfDn5
HRQ0xUC0q9kQhRBwn9Ed+SXzML6EXJO1fdD3vygQ1WlCqlD/DTAQflVAmLMC8qgBPmFxu9sAKGZJ
Lm4LqB41EWeM1Z6eCaH0V2FdbXnRYui5yUyqjMiatNfDBMBy/Cp9q73GBTSyJQORAp4S8AYPxNDd
05feHneb2bHs7T2Bfgr/pZ6NGKbEPuOr2ERFLk2RR8e6deo0llIG7gKNK1wz4cVPY1i3DpTKGyE/
kNuUAnU1AEwNWw/EBHmEZwI7iSdsy2IrCvDFjzy3IXDlYbVAI2hjjUnTa+oC7A9xogiwU2S0C01j
zJ+BObFBNEbBgmq/rLlXEHYz9iBHLco2c4k6cQ4hBygbVmJdnLKcsauywexrNNoCVgnpzvdyrc8w
MtS4lziv7+o3aq6egwa0ulEbL86sZZmGj/tz3Gf8b0ZqPZROsj9snPptl/6rS86ldCqD6jv1gGY7
V8Uo8oCYOkl4AEUcWCXV1po88CuwJdZ1WvOSKVPt2iRBTnqWK+C77j8rrIQTCeEtCZpN8SZZD9t0
MkWUIjWQ+sNhGFdzFT5eRLj3iy4sYh6aF9gEOq0DuuJ2bHcxuLbhb1jcY3kSzjAdEMsyqGkYufac
oi0vNQB1OkwCGJ4z18IDAvAuPtcuV+Dt/fKrNjkMioVFAskP1rrQaAr/SU6jt3Y/6FM/mVi4j/9R
4MhZuSxhO0U3+iHMo1L5ZGt10dsBVOLeIc7K3AXeJNzH2zzNKpHrhfTmlG2Oyh0IoZu2VRMmN6KG
0D/YpWfUoYqwq2QFWUDqA+9RNdikLAOcA5OEsu3kUConZjCNTnEkeTHSe9JaUPd11jKFVWXN0wto
jjG27eZe57gicfyB2R8Z8rKC1eQ2rKbFE6YIXAYKrztCBV8frCxRvF8kIYSF7a1whoyIRAUNVGzf
N/FLezOTiNHqtoGVs9N77m50AgQGSRePBzr+HtpqkN8iyoJt9lPWK96Rv3EIPlZxSueMm4DtYrLt
/KCHFyPGITyrv9Ofz/9HZG5dGMCJRr0EqpMWLCMHQ//GKjMVVfX0cdmcdLCHCTaAUQas04OwUOfG
Gf3pL45cJdfnex0aKD46kZ1Tcch6IQLZeKkToeTb+gJfR0LkP/o2nMh+KEe9xI68gpDRar1w3JGS
5aoeG60CdE/st30ndHpp7a7YMpJo+D5rV6zsatgo/G6tiRzrDS+537/pOynU9uhVj8d0NRQh6wRg
r88h6ztJ9XasbPVDLWqHHl5noGvHacqbg0ZKbkzK2U5HJDqIqVM2Y3MUN5rcht2bbOdfDVm/kYfI
TkrfyAJIRYW9mgZwPLL43AsIB733HF1BwJntzsT3Trf9JSjjoPOg78t7YBZhwfqNzRD3OO/b4lJo
+axC7Nw0tBTMFBSllPZ3ZRggIRojm/XvpcmQQ7KRJRrSBsJTDQp5qRooSeOy5eHkohK1ZnFtIVcs
7g008SRvB45a0TF8YTB9a7IrS6HoQexqtlxIJPrlxbfTIkbuwcRDh2mcO6VLBmxmwChJiKIslbRh
s8xKZnE9nMIzX8Y1O1j2XuUqRlzRTljvs1QmenE2yOzVX6KAuk2gtlajcoHy7V6H1venhHUNWPl5
ISdQNX+AYEPi8LkUQkqRRIQPGKp4GURSkkBUwrXVprkM6rj8lOs0qgxjx+CN8GhFupjE3HV2MdpJ
e2pEUkvD3AfmF9atbMpOB4KTpVEDdGzL7m3b2su1DmKhcTu3iCfhLn2qc4J9XCl2g+WPE1bOgWd0
ittHv0ebin61d5yMIMs4Y9lUWb1X7TOl6VuywGV8ZxQOfQn4whusCD7WAzJUCPhx6uzQ3L5bcPce
p6NUywcBjMMWKVytJaK7kMKYYVo5Ki3i/pTismuVCDDxIAUuxNf6q5c4t95AlwTgLlMmOFQiEXWG
XWlcFIzePkAEytZQUNGANLmDqMOe8GtcSIFT343RbYmD5Q3EWm5JiSDiHh24gDed4heCMoB9hH6O
DoQpBoTy7/ESKGYQY3g5pG1jT4SXT38NSK6/Q5x2N0ayYJo+IdvSmTVeMRd1+9crj8F/rhVummHA
Brfoakv6UFisdiCsksWb3qRCpNZdF0jIVvqlabvGSC59ffIV/RNk12lEy/8ETj4v/1uQHuAiQkwM
bhUskdfWfOHFDiyM/4nxVvCcm10V3uG4OgbHUXPJ1hgKgtLTs1X5jcx5WwJTOg3IbE2yokiuL/F/
0KWzhHF85nEHQiVhNuHnbfqQ6MvqQd6goDhh6OKJY920k66W7rj3aYCT+AFPTGKxv7nhR+VLVr1T
BdKq4q0tz2pFJoKA3dd0q+zaBMUnoSkrpQhFWlBG9JwFMmF4zPY44EXuFDb1Ss0Mqj1M0XN9xJEY
Mm/nHt1YIuluYRAOMzuj2g1tEymbr/xtTkthg5C9UkpTF9h4mtOnrswHq1UtX985B1OCGMU7XLnd
D3lonITMGoFUtttEaeh9245iWod4kSVWJNIZIzrXlNPKzPCUrfRKkirznLe6athspE9KvA5kUyF5
0SBuTOvuB+QKQRjwX38+nReiFH0jW9+JmpA7/xwo5Sp76R1d4SA0C4d/+tSAs4vMGaRQ9aPhfdLv
gcTjALhbNIyDVUaZ/ADhR84gztj/LEuVSo6O9x0ygA9pWT0hr5dh2DZY+fFL/b+mMbUKebd5h4jZ
Kj7aiwNfCbWgleyHI/Vs16UvC9PmKw+fULna6pkYiwcgr9KGgkeQKZJ2UMmg0/cn3xDGsfiB2YbD
XjiHB0GmczTWmWNqiz8AIhgItNG0lrVxbW5JWxgGV5SiNKSX5inRyMqo85hLbk6NUtp5Dv5GMjDw
44uqOSH/oTattZSsgtdLs3TxSDohEyJ7v3mNk1BpiqMcng56YlsG381DUjuMrMdMGf5zl5qbbfRY
n+oZjpIcyDw8AFYro08Yj5HiDkWiGTYrQHrT+0gq4MDnFqoU3Sqro4MJl7m+wYykchWOWlT91TZ8
YMFpKakxAUoY4qlrB84DxlCtDt+DqE2chkemAv7gkBqiWYpX0tp8t4JyucIkR9JSHCuiab9MvzMY
YaLarCyQUiaAbNRK+GsFz+TOvNrmFjhaoPgF3Q4T5oORB3ayGXyXREBnPaNfJURPY8ChH7/YtVbl
kXbw8z2jqJxTdCxpjofiecD9lRZUdlCWQQZPEh8zARvOPB0g78aGOX5nF8cAJEuEsoBamNPgzU87
OmlGy9pCT15WqJ9uCTR2ssASlbFb1wxvZtcQGUJbsbyB0IDmk/y8RGvPP3b1eT4L3AE4L8KJ5Fkf
iU1EjNRuLLD+2WaEbkDIyLQtEqYtBVOgSRgwvUJVY6ghvkQ/lHhMAIVEfwNt4fX6iaoR7k2kAEQK
PPvXmxFbRpmgIWTWRQO3nLuFfeBmBr8ysbPFIaiemlSNXvCOLQekm8RXnEHIMSXln0Lb16mb4sql
58qO83tXJUVRIm3yzUCV2neJ+XvXnS3HILIE7uHgyFLIxRMh254gsKEb6C34rmqqvXNIZXOymtmk
Gjbrv0T5UU+idX31Athfmn+AuQBVaWyEvR12syynSbZcXkxemDroPgPHk+DpN9kP5uVO0j+4nOl2
q9YjUkP0MZ7RCsSMucwhKG4LSP8NEcU9WRFMm+V/pZ4xElG0iuuSiUyo2ftEh2XYw3Ypg2Js1FrL
Ky8IEpU1rnpIX1hqRbiXDTjjw0H+EMg27vW3k+PVhdNgUDQMpXmfCNsWSpNBWDIEF+xM33dhehYD
ee9lTtJLBiU+K1cBwZMpWQI2/BSQz9Eod+QsIX0/RfTtxGfefmJKqJIyiJmT/AWyt0x/gr2ayNpc
jlO2h7VZnilNuv5K1d2GANnSRoA/kquwHKInIFUPMQ/xlt4QwbcXCZ+b1BxLHMhYBVagHkzW0lhE
z0SeoJmR3+Hs/r2x7Xg5GUo7j2j6V3lTAGMbix5IWziLmqvSUsHiG68IR3ghuSYVtoMF4avD6fqB
QQMS3aONlna+o3VGVfMkRxOnzDrvtb56NZHdT/Qgil49FPZZxzuEhgNWU0fpOz4VfqjEAbN5qIrh
NDK4bPteTCM6j9FZYJAJvC5wr6ywneCv3aLaPMJzfgS6k9cH5iF95XutP45SVMiMCUqlma9rFxlI
r63W7KoG1PNW/eTu013hC/q81qgfvIyvX+3njk8LpDd8K104mPsTOyJQOvcvlqLqraQmDmYgy3Sz
FPAe6K/uCYPNc4u65jZqqxWu4pPVHXacv9YZnbKvy2EulSGyY0c17OO/p4aOMtLxqoO11WAVjjSs
7I3bNaIavfoIgngkiywQWhszbPuCEHgErfrsZ5AiKV5KOqQPWzlUMFSEu4FZfl3oBqfS8fQ1XZfy
GflizO96rcJ3BSwhseq+j6Bopuv+xdXH/XZEvPzcq9BZwUwmKU+tzbkDhi0M+E8hgi/Hq92Rnfrw
IkXAu7592fwN/MnQm2xEbBkEtTvT4ma9toHFesUjxMZKw3neRZdYPTnno+Fb4b2B9gpDC/dV5osp
Qk+neavEEWJpbXpNxSW1+Q37fzaHdF21ilthFs5oyp/QNLtcIgRuFnZSkQ6Qtf9q+Rb0LlQfzS0T
W4YVEuzijJ0ELDBZjrly7YubjdBkz5G3pzOSNImj+HcFH9sxt1vNNf1WsN907VjmmqR59r1tKqHI
jj9H3pc+d3r7RKNvkCAAmNvdh8SVzOOptJTavXlqoXwB9hSud6wIQkoxhX98r0w7S1NnTJmE3SRY
Ctik6Z8WTfhmWHiWaZf/6x9kcH4E+fZtk6B/Icn49FhgXS0T881D1AHDKlMd0dL6o5AuP5W2FHPV
5GlKwJID/ilnYid7ygn7IqDmkP5Db5rXw3EZHzJYkadb/18L4h/sCdh2bp+cnDNk/3X2gJiWZC9T
2YOl0VLcxHrGhKB2/hGaH9qCtdJhPk763Bv4tE4Z6E5aIkpNtR29JColIWcH8du2YK+MtQ9KxKVq
ezKEu6zCcfG2T+9J0aFNV6oJ0DQ/nAA4BkN2NmRlQZDk6lzXC9WWsLxDQJOo7oLmAhX6AVMoy55Y
2QwBTUcLpRpL2EY50SD7kEPIXVPmVxxD01e9bMrQmN1DIDS92nOox+DkYfWXc9yLRGM31YYOEVIK
syaIOgi7KO+7r6wpTY8AruoREYVDnFw3bXrMHe23HrB3VLeU39AkAEjv/q066JElaAot4onRJDms
wXbrxWLmqc6OseNN9yNByauI2TJlyqULA2HPajRUriFIx7X1XBvf5pauhtBcm0S/xlbo9ZqV9Rhr
+22ebnzr7JjMjcESsHtfqqkTeqF/HlUD5W1OIec0/lD/kMZBJgcdNDBVqcRFrnvOpeHM2zcyF5Zo
dBXhXWcd2DEI8SNba2XZHEJrpnQrSgw0D5qQ296bSGLzKm9ENuMEOB4l9PmGQvNszXY2S08RCLLr
zecabWWfUQIgvFg0Ti0Yc2GWwUgqJSOu79F3c4JcFGYMr8Ml8ZWJdGsefQMB7Os47g6vjzifKIdN
DwIOMwGQr4+zyN9yNoMoiXUYsDe3q/eyPTgEhEOewt6iqOia08b3G2GzYljvEY0C3EYF24SGAsKC
K3KmxNBQDHWFsI7XH3sOv0P4wrRZ8kCbvPHYKxGqq46+12JYx3SEmiNV0HIeTKkGACWHfeJo2pXz
8cQr1NB3izZkStJ/gH7Scv85oVuyR+9l0qzn+vW+ykvC4Tlkp6yhozGqu7MsMqgF9rX+ImYAxJwf
aYeUmc1jLETdg5sqos5N0AGWtEiDh9wygfNWjYtmZIiMem2H6gV29ROcJ/BxEN9f7i0/jUaLn2ZR
t3KYPhwOG0DoSuC9qHyD3Y8i++o00jHbG4M+YXqAHo8SAMdrNQIybfIMTv14pKoWX9g1OyKhy762
0DAgbmpPz3YloiDbTFNkSnDrb++h3KougT/tcZhanpk/x8Gs2x81SYgx3222Jm0IOS+sKJ8Tj9C1
65deDrxkRyHRdb3epJqbKzs7Bc1c/oV3Y0XRyDah7kSgW+IKx+DOc80OwfbWMjbXkD/0rlpSJkQo
JhVZMuGtgKP6YUPEEgNsK2tMyoxEvETTpqoNWWmwOBoiBwxQ+Ld3wSHAG2CTC09XBgGWzxE1zNp/
bUSht8lJiG3JOs5DtHt9KN/yMMx+bY/81kaQx6P1CyvvATtd9Z86JJkoLj1OogossLxKS86Ue/4/
JDoiuQtnQR26p1tniU3i5m+MFInFVDOnUOIViIKfIe0WrPoypTy5wOb5Fetro54RE5nG2Zj4Tfwi
jN92erKIiWpV1nzwV9bmj12sYKs92/2x/YTsPVH7Y7FpR7sXU/+RxfJlSTInaGA5qAZXnxI6EgMb
G5pEFPiRRWu/MRLeQTU59HqLhFtGmRl+FvXLEOdx8qE0dOXh1mVOyE0D/ALelYZzwMsrdTEdVHK+
pnIqxpo1C58E8tZfUXlr7sy4uJUcGFSZ+B76ujI8gLfJm4EMJU8LCX0UUdyyuL+ytAxS6CWiqFJf
fuRsUGPUTOuAtno/+su3QQbLrKseG5/Plcb4EVh1TyN7/brCSpiJuXwsam7JDEyV82L+pPDM42L/
3MlVyDwc5zpiwaNVF6+M2lM0yvO0ucDHAB0QVQ174OrTyTYUSRYNaeH5TUBRgJDOud0pFAvd0iMc
psvKu0ILQICY6eugNGL8xRmLTAAYHwNFN6gx7+wiTE6Tg2DxQa+eomwUIaKzyo8CT5k+aKMZ7yww
p2t42hOUijwwEObv9tiEBQOaHeovlt1RgdyFHScI7REAVZ9jJ/vO/YHvK62c2OMwRB2swVH9jfWC
4m5yGSiCiMb8S2Gcn73n0hMiau6cVRkgIxkIZ5mWxf2um2em8L1pjEjeOhpXYKKXjWVs0BHVQS1q
yPwg6kBqJ6JeU2C38tyDAkXOR4qJmuRxFqcD2K8dQypQ/uXGA0XkBRvcUh0ed41pS6SNyMpqEDDS
ts2TIcMEPieFBlpliKICQsZULszNSwljVeFDBT1dAMNj0zJYuApAvR4vyACg5JFRp9G/eWNVdBk8
DbT69cZlZJQR3mu0+KJe4Uo3QuFobZBSce5+CH4070aKd8aWjb74wOXp/Iae7Xy3UAAyEp2u2DpP
DRPU0qHuwQSlspXHwSxQqaNO0wZgxBBPl0OwDuEtEpZNocBmd7plLpId5cMfqUeeQgGw1vzF79lZ
n81bsNSC0HaRw17TGsG3G6LsQiX0jGo2apl2c+eHMPuX4+GK9FtHWD8k8kClCKsZknVFeI3qdyK5
5s7BV0NL1c7XRBPmkhghVnElw6grzYlA9GmkGUhinhozb4GegHiqx44zA+MoxWUwvGdVSk0rY39k
ZImuKwnTnSsqHtyr78O78U4ARhkIJW/8R8EUP2rWkDaIQU1JjIfJdoiEDX8qknIqsywNDHhJ6w3A
Am/X/YqXbwVpPjj1s1yDH4140MVOVaIKTYPrc5G40uuMJoeftPRZbsfY/73Wr7KOuxGMD8LumfF/
QxjD7vmBhT5uIhVLkZcbQMiK5OIohJfKmnG7v8bNXKWeUfORc77vWXpbvXLwM/eZJeAWmA92CVxI
o0VYn2r6YGIOx0ZZuLNngU+tyw8F6b/64zHgKIT50s0YoiyQEf8Od5ikhSwYWlV4v7acLAjyS+f4
DP25Yj+9HOdcSzI40ge2L21Zwx6Jb1g6nX4A614fytdlb+zTxuv6JP2pMAnUhTjxVbHqMdTs6n25
Nqz0eIxbZYV3UpA+y97P3R7nF8xcusm3ZpXqbkaWs297EGDiTqUTOsNC/Xueqnc3zci1JWuZj7oS
PGeacaa2uooyNszZ7LodWxT1Xu6f2map1Xy26B8iFe1dFiAqk2zIGYaYIoWQueuYXSgFgTQm1X6V
Us3CCGUqrKZQXYfbzDQRueb66LGOXTnGx6Sqob4WL967Bxj/WYvAzWTyQpBlZ3/xchz+GH4EQKx2
DgpFZK7clFlcRGTaxAPHOD3zw9eyiohB4MBGtQKVVwUnIq+d0OkuQugV8IpJRNhNkqY2/qbFhenw
is4mNexQRyCShwdfeZSSdfzDrifyQzQKF8loHGgrLRhmdwRPFQpgoWOCEW5PhuQNFtrek5rEPEdC
vsKSdGt5cOQ+lXmPVzPxWcWcikE4yxNWsxsAWNRaMoji3GdDpbOpQZHD3dTVhe1hP/wKB+N6504K
qqe06eNHY7qd0okKVVJ1WHs7eGZbQJlSnlG/9iKA3jfLtylJP4IsoHTnbn6BldV6DzVqhYDs0lqS
q5uyheDN47TszgOAH7T5vKtbsflty9cf6iRB2S2FJE71Yg4x3O6WRikS6lUB7q/W5wTPyTTcn9em
25lf/HERTmNmWSgvakCYYEceymF/GPuQ+tSnkKAgEsLVPhuttjR0pGbsDY7HDT8O7kd+ojIooqKe
427ftBdt3K6udpSmpSgEhVt1yLEAiMgY2ZA5cHIA07kU0FGzaOxyZ9dkVQ4Gfc5CVRW5vKkGR3gP
46QebbCTZnJqxFiJPE20CKS/FcqAg9bCPIWMVOhs2/SE5txEnrPbjM9K4Dx5G/uoscKnPATA8iNR
5321FjFqTWVZ6GXJGy14VGdpZ0U7dny3XhhZFmr7YLKOaRNA/GVNB5XqjCbMAVgs76cADugtzEqj
iXR25ELRxFZOfS8sqQk7Woirh1ijPVugS5hq2kNDAiV/dpbA32o6rP5y5eSXXh+1OTaCGpNO7mGl
W3ZbSU8u4TaTywjrLQT8oqg4qVVGMfX31VYB+a5scVkp6PRmc7trqu5OJ7QpAZX+1QVm3jk+BUDV
uXdmcc2iWoq4cwJ4WH4JI5iAVGwct8euUAZ1i5HlGbK9w9iFIoOC/IxEAV1XPTauUMk01w2IZ8VH
J5fQauPsTWswvvTyJG7a7JRy8YqGbqAQk2qJzRpUHFEq0pC6Av3ffLZrhiO9cXdAO56c6d2nfKss
Ku3Mud2wV5AnsuGsyd7O30oSBUkWgKtF+RoNr1D80ApYPFj1wOake1mwb8EA/bI0FP13LhHgiUj9
Vhxz1MotVNpGyiGT1CxMp9FJ8lWHpNOeThmIHS85/FEVGOamG6oRZu8peZqXIT7W144TU2QIYuQ1
YULjeJI+tO63K+9TVcUNjR/w9wnPjt0Oa+V9KpGZRguvW9Gcsdqz+xMUPk+6ftYXcJvDfuIUQ1BP
A/OL8H4LTedThipTy+EuM/1sdAGZfmW8Ks6QWqTtx4JBaEqzu9Uxz03XgiFGdZWGH0X9DCbGYANN
mt61Hf+new7Y7pXMtQwV+0uy7UFeXesa7aHoxLSboPiOZALIXBEkzlPwaBIYX4iTfE35V/DJc9in
9PMHIAJ4XdqYcUBtnd4VvmT9yNYvPPSMqy1KQya5G70omRQqNy+oXQ633z2hQ3jYzPqz4jUrYJSR
/D8yDOK81H4z1vKLSL/actFWEy3YGx07swqIoImzCnFMJgWvy025u0yi5OYfDMEJ0svcWsOWg0hM
oTCBlaJKlzN8qE4Wx5lxWJ/ChoCHIfRZB56Ga3LdWdJ4E0ZqqywaDO3uA/kiVe0DBEMB/CS5/fXO
HFhQpJ0NotVOXJqcvZHDMVfxVlYiiOx+wG8GI9P5L4kGWwuxDNymeGy+fKzHqytAOI/sE1GLnJWZ
PV3mRxE94uHou8KIKnuev9LgfEHHbM7zvQA0Z4axUOu99BZ6R0cVBgeOi1ZpqzKkG5LBElbegAnj
IWYqlMaYrlAgA8X4SQuuLCg9s3BrKkhDxXiQ3DLgQ7hoh5KVLX91yAZbmla4Ub6hwJ0narz+dx5i
5I+09GeoDc7DmbtwIKNpPFJl2IKtpNUMpe10MXUaBTOJ05JxvDvTTiXrbn0Ql+FzQ9HhO74nv4XY
hDMR3hyFJ/eyYnIHD8S7yeEkoTFOXLu3wLRMeB7WRL8aC8+kU/MDNV+/VEJ4WOnU0EbGaQxzlWWd
8eE/e1StqWZlYM2i1f7jbEanb7pfG8YVmlhDxbxbLFKmSCQNDp2Mn357CgI/7afm+5/X9mk7G0Og
AtJKzJevZiiYsNW5Hi5MZsQ7TEDDDjcNvDTDykyohuHB/h+//bd8J3moKVQ59qBHkkjzi4PALEsg
JBlX3T3rpEA5eexs/U8I84Ll5EnwkKJUVKBsIVG66o86esEageY+gb59DDJgoq7K3XNeyC+2NwZx
d4scE0FaEym5r3bCDULmzoJrfegSegrWYLQkZWqWGKUKZF46f7TO1I7VyUrZTVQkraJ3YRgkf3RD
Hb5C+LKlTDgl/wbUu0ovoP9up0bi/OGPxfZBY6lFM6Sg056WTK+zna1I7fNawH9YKsxy3cJB7S29
Bbd1xHcm6VuVkAo7av11w+fJvhtuqcoNPyFynbaCopKbn5B7FNylaIZy97TJIpVDm9T3JIbK8QSn
adyu9v86gMy3x8H3kbnxZqe+uINJtJOKUJqdfRRC8MhFXBOU6lwYTX1mPnWUJPAQRi4ipwAiMbS4
JJxVwkUS7HLraZEwuIbi+ZNQLLLj72830XeNz4jeDZ0PZ7Fzq7csymG+VBoab4qXiUuqvL2BJ/V8
DYmlR+wTju7gnHMorjdhUB4m87IKc1fDuvkxHuduuWU84N4YvzUNHCd6pSX4zCJx5mSHSkgSL9dr
uenNlbhxfBW+GjqX2uygBrWN6z+c7g/V6qOO3KuhQuhgaJP1cnvxWT77NxiKpIfbs0iV3zoG/lpR
chGLvn5V2TlAviZtLzYajTPeE2LE2hdKyhBfOrczzRqqm22SZlSbHxWlD5ky00DRk8hm3ILrRG3g
A6W0pYO8iw5qZ77pRzYf98cvSPqaxcJFMx8hKtCTZF9KJe5nDU67r1ZksZ0YwfTy+ACR1+bw0u6U
xVWAJ8ba9k0rRIxIJ2YBSboedz5PFnx/rPU3Mb6qlmzeu5y3YC5xO9YBkJ/muU3sTJMLyl6KVros
at3dlme0g4Mzfgxrzu4y1oLrwpsf6jH/fu/FEhwVpc9IvJVFOEWSuBWVmXmTS9zwUtRXGdQ+1/nc
0R2BPp+fQksZIt962ZkZp9U1gloRxYcMQjoden43Q5T8EhfdBHiKf6RJJrykR1KTkexrwcQtm+sL
eilXdbWaKC75NVr5Ufo5ZKhxPYPZ+F5murgS6fit0XdqrwR3hyafeI6tdNI3uVBiTl0o8IheCzFr
l2W5iqIylHtm+S3Sj/NUe+6EAMN6zQhNivJ8NsjqgaAx+NuoZplX0BGNKXsinGMC3d+cf2NTCP7V
wUiADd5TWky6O8PKGb9tvHQH3eH2pVhxDguImxS1SHd8lzl0f6hKTRBe9wT0q93tOouWHaqOHxP1
40rN72CYOm5woiJt1lAu6HVMzjW0O9HKNJb3tux8BAi28OquUJn82A1MjQD38kGxZhaSIWxvIEeu
gLvM+6WwFDDNISkCXl2izj4S8/TPYWbcXq671KlAj7ERI6I/hzWON8HmCfQv5vei3TXvCfQDluZO
xmKo3shMpV/i/2szc4n8bvrp36hxjWLtjbxduObuh8E6lHv1NU9h7dsQAVkkIaqrh5q+QIik9lZp
uY6HpKeSXTQWmpojuxJw5YWJVIV0iWUFYObAyH8Bj28yx4xit5ZwWQlJ/cGLg86M0fy8NKfHy8ML
yA1dyVp0mPEQ95JfRjxjuRIWr/A4THAAi8nehjdWA1nzHXgiXVlZyrclp4wSs/6FCtR5Op9eyP17
wv5XFa6TLVca/FQzheqHiSjQr0nyE8aTa3X1czrfOoA/UJHevhvJ38TuU7eVLjqHc6THBH2y8yaF
m+iKXU8frFpj981GT/VNp0l28yBlPMOFTGIfa6Kwb1e8uvKLsHmIkrvxIWMG8qhkk6kauDqofkF4
RZJZXvbA2N2bDNe58vxrBL+8cGOtFaGqs7oV/zgaxI8rCfBYk0EuEFRLhhxlQ2h8SbAfhS7elhO2
HKRBiDUfmSSmUcmehRiBy7p15Hhfigqg8DidLCa2amSbpnCHFk6oLxPDCrb+jYyDCNy1rf0V+kSN
38/ScEkeZoD4dkdV/IatGmsNWhIzGf2d4gi6soY+PkSbwL0OU7O50OqQCHddDpq7woLYVCpQD7uI
EG2WD7MoPUWb+wJWAz7yPRsyrLgFLPXLJOsnffE6z+smx3fZA/J/n86UYEBRjRMJSTJUZykeQzZ5
Ap+Tq1ZaEODWPMZuFdfLJ9hUb8+d/VxmZjGzJbJ0c2G/9ZPJDtjMyLd0/FT6VGlaynM5C34LVprc
7avB+KO02PbXtQj6TxudNzmJ7j4DSNzVWWd8gg3qFMg4AKVL54EDw3U6GKzTURcoBizNSb8Eyrxw
/B10ml2A/Kg9f7t49Yz4w3bmgekC0B0hA4xavhY2YHGwsRsQ0SdkeseOhOeyAaufUSX9OpvBU2ws
iMS1v7cp4csO9jq8g2hvuazmJPkcyZeEUOiZkol5hSr/QHy3gYB+7z5P7Vyjv+5779WYuB3tLKnF
LeyNtqmDCJ/Pni0ol3nDHUdp/TH2TPApYpke3XJDAaBF9bENJApYAaRUk5dp7+INMY8q5GVMXqDp
bTHJqFcD+srVafEqzvYzR3TVWg3fJAaQo9TfYKEsRd68iyi5/ZtnLde/P1GSfWXWafeNfNWwlZHi
+QhSKp3axzi0xgkkE7Nz7bBx0Jr4iO6y7MUAQWmmb35tIfebNNt1QjxDnLz8BhNZTe2Uh9fWWLkl
bkKZKHBdGZMt6G4/LBreF0eljMufrAm0e7FIJL8NMj6uZandETyKsQ6DN2HbvskFt1QfVYAgWe6+
H3jdhw4y3kNTXzYxuWG2d7aE9830CoEVcnkCFNGcPWLt1/vhynWkDspV9HbphVOyUU3hqxSfoORf
NKrftvFGzI2DChRezgVWimVgoEAxVgGcR2Y8xuUdIJsFN+jTVb+rqj0esKCRcsuZG6uwkBlbhkRX
uUGT4F3pZ/uIV3+ruvrXD4ZKeOWc/uBqRpBXXdTzhAdH9P2JsYYzf5HIRo6Fu9uLSzPXwzvgr3Ij
EITgP6AKG857FzvTlyg+tgKLTOgYbH8t85kcWdrK5xCTgrEjeVGc94sAUwPy/RQ7HK4ZSTRYFPBP
ICzIMmP/Sh1P2HkVAF7Rbbz6tWCaKTfECA6KP1JlB7Gr1Np+EshVN3EEcr03MctKjnkHqhDwLRO/
4X76XTwveyt9KUpszSJWfJ/JcsaShYh7lpxWRQwZvM4xHv3Csp+4ogF4C1gXAcCJN9mhvTNzSrM2
lh3vNLg+1Bc3t52zGX50BXsHi0b1xBZtsI6CXkvKZzX7/ef7xcPjMfGOxZVXBa9PJWBSzCOyDMYJ
BDFVJtkmMw2vE6Zn49+FQ0T+pC0LouRKgb9aX3Zt9qLYrhWKjQq4Hm4pwyBub1KW7V3G7W390ujx
HANcne2DLBreR8/HvlMiSewvDdjIxXU7bi81ghWuOeWI8HvXzoWXNdmXUqoJT+uYg5TXNH+cF3If
czcopKwN3dVVeOCP5X/9Spw9M+E0u/ZsUx3qcxmZALNIeUXIdMPtxVbXo1Za/iGK4/8n5USdsY6j
8hb1uHLBz6hmNSh9a9Y2qcZ+vtrNf4bLODOahfb6NXHBomhaZnMFxHuDgetxwYUYPxqmUBQAItqu
pLVXVFOCTuPlAQsS8pNHzXN62FXgQhx5YixzeKlWfnJSr7YCHdqKyuOwc70tj0B3AP4Sj1HOyBvx
HNKfmPuJ3z/+YC71imki4MW0xUjHTwPIYnGJ9DFNFNySTL6FLlvm8NXpvnCl57eh+9NHvZxA6EQi
xpdWNzh5333J2CgJEk+OX4KMt8ZO9ccabU0lYvdZI4lKnPJ2+kUpxPGtbHCclG3bGC/e2cYffuBd
WJXLJ9lc6Pmsha3wVGDp71fUdDxyTmG12tsaUVlvWBEoHUdraGh2aOZ2viCDG4OqB3B2BCNOuPT1
hsS6ohUUxOIm1acmuf0ljAGyshyCw+zsCbIcYhl48GSiTzaCsM/G6jqUYwvxKMpFQR/7cFhPSUSa
2MENMVqCJJLyPCzQKs2kxpD9OG2OyG7kkO9AGlYFpe2hHc3G2we/qEPkj1VwKk0BjGn8Dsy/pPLH
RWNsSJnOSlOW6blNUjtGvf99c8E3Pp/FOQbGfECwJMIJluTVg40VVMvV3zehbcyq424+knkWAtfy
dECFCC9auiL4DXoT3BqihmC9nrzLzbKZpJH+9Pgg/A/8r8jSv3+m/6cg4mhjp6xrO9dkpAGeyDZW
AQ2E+DNhclNio2stAoyzW6W/I+Dpy2hpMm+FVM1k2XUnvK1Q1QiiAT8BAv6IJ/Czpb6sT1fxwPqR
iCyw/rfpTudgaL8/Iz7WWzxKAuEA3GGLzDgcWUgpLdr84ogP8Y0J2TUMLmJRLvcvquKsrEAJ4MHp
kZ11YLJeXnYUmW3J8oVLhaVUNPWId0UFtQNHiIa/SUXyPLZu0Jo/6pGko/hYqLAY7wf8Ve+AUsaC
Xjfp8D7goOnluYM6Vjh+Qo6IzjX8AjhLWu0VwS29QFcwvIg43A9Y7rd3BS7Ah9oPFz+XLWQM7TFQ
54ZwNHwFWpN6iscTFURdim+B88/A0hCvC9JNSrHFimLLyQMTNfPVq6gSQ5MqRc1rdPnqE5pXqJzy
0sb9AY8VS/MurhqWef0lMDUgtg1FxQnxDJ36qvC1Gc3KnPYDPz7Udkc59lH2xKTQPnWi3rWF4ne9
0WLezZ+nVg0c0X28l5sGj/D/V7lfwBeN0QBnz8GOgCtOnl0TZezJN59Itp7kq2pJl3DisKtAdS0v
/CNniLxjzkWR3fFnywAdne17WLD0KLTL6jD6QsvyhXC4k7ezXJ4jU2dGZkdUbkFfDZYlLtNYMhSh
flZ06ULPaUsRSF381So5M4rX0/Jiv2ll56/uz7ZjZtSrB643se2hmynsIhPxOhGE+3rBfez/EnXA
63kTzj4HPxoX8w6OeeXfZ4zSbO6DxLYGBwWoVFkZQOYLHKjir1lq9YOMztrpd7bCSroqqAs0ZP2L
YH4BBt6MzVelZhet3t/WtEZhpWJ5fVVOxC/799Znp3yyEv6TrxTKujnNP2N5yIWQQ39sDy5xrGFW
GVXwiITDImVnI2iW2Err3ZuBudpODdNhTrqyce8Q3xNMLtl0xvR3KPZnfm7lPNqAXMLekLYPQ1w0
O8uRxTHR4Wf/gmEQroaOEOiEVNmNFpNQlbkFRVLatd7R2WOw+r7nSSAjX2Y89TrHtbWpgy4nHPwE
OXLnxDf6DxC8JM4ctrHyOillVLYF1Wz5WYeH0o7P/F6GO5cZLo0p8P+xCK19dloeell9I3EEPcA6
v4YDC12mbFrsIsvL0bXiC5UgrtVTqPSkH+lTKNrTKPCZ9DsK2vJRM3fgYEBBHr5K2vJPORaHhC3r
k6+VabR1JmRztahWCGvJt1l4FIwBJqHh18CYDrd9fl1JrBuL2ELHppvwD4MnSeXizSk6ZpZ4hrG9
w4d/N+N/kHF6JpPQgpjY+dxqdJq4NtZd44ZdcJuWhgJBiW6ObtAwTFK6CMTHHi7gbcFVr01QF97f
2kX6LhxVmYYLViaPX79+Bysl5fxCOIBnf4Ja8BB80cymIUCCp+LpW2A0SPl9tA1c75xCZdvAjldA
0DMj9uPEvUBIKsQl5Sz2Q0J4zABlD4AMdrPraXw+W7p7i7/bJD6D70obKEtWpe+vQWVSQXZ3V6Ai
FER81VOjGEWBJB5LPKEQsTumozqs8bZBALp+PNe0PqhUi7pV4poezUNWJ9Dq34S2V6seCihXHMFH
amhbmpySICR4uXQjGeei5Stri5E3Um48n7zypc6UBJQLMApIXzBxWYtHzyESAmapYFQErm22KcLF
9UQKuYwXUHxHZL9P2Xb+9zFTcBZJSJxapi5TnEHVrw1wInXmYm+WYyAX8MTL41CCknS7tYA6g3CH
ZEehauD9bPbPiwlIqkcSvVO89JmuYfiAM40xqvIYjQcA1uL20ulGuwT9R0YO/k06X2xQgbzQHNkK
m8e/RSpPyhMvybWARuAYnD92/Sim0YiC0dE8LnSDVjnuyjfqycYM67yks2d5T+5KWHhEu6WyB7WA
OPC25iGGNeWN8PxytxR3WrS6fjTFjIdiV/L04Zg77cz0lfR4hXQXSpi/iFEejNRvbfnBssmmWDzD
fI316Ha82eAgAQ6eNIpCCqBMUXSPpFleRR3Xt+EvIAQ1oy2SPBxf+saPQeenQ14nOwcwL+lxyRig
5sU+bTaow2T2tqf+eRZdlFkyPmj3MSbRY+1+u6geZqCBHAwn7L+supT+CNztQvHaU+ARtD81yIEs
3uBpII8M/Vn4ZzdPn8YPgiLRd1fHFNGWXTtIjgrGXFYmAGxbMsHdCsmTPinc2RNp22G4sgwMPXWn
jTEz3vgTJayIW4GYXjC3EWxSGGJaewDZMfxnm1PEnpacgTCNlLx9F+zpwAtMqH8ChRQjTozN1I+C
EuAqPTiFsLj9+6q4hl55kvsd7pZWLJT5xcIaWFvdQrA2wLWBBvTgRTrK0w89kQoOuuwPdfTQiMpr
r+OvgvR5xMELxJxHZ1sWwfRIsDF37nOswubQ8dUOLbwGNf+QPUtgKVrE2B4cE9m7VRD7WJ6osY0I
ju26ZJRuFzS5hVJ0x6NI/1rF70pK0iQNkGIMXPx59+nVKnWGisrfYhmYtHRzu9y6l9m8dvhEYyIg
Mfjmv6uFN3zProaZXTsgXq0gJ8Y1dmigEyX3OgnWNv17FTZubjMz7INyPbmub5PmYsCvjz4p7uh/
fJbybISP8C7Fcp0Odj5MoQgirIx+4MpOczisGaVDdRyqEAShMgjptFmpF3qZmQK22HFMSN+awvQt
cVAf6aqPZ1Mro151yyEEHcQ8gpBPcZGOmqUKL915w5jMujY8p4VQ2SAVeWr7LxnHuu1RP7aFnJh/
4d5gsDTFRVYquk2MMdZMfId4XZR/Ak2gCaOaveN7GrxR0Z3Pti005DhNWC0ZHBU5mxA51AQGEX3U
MrlMsT23mVZguk6Fq8BoyMaZO3qpaYqJD1cB2v0cja+cSwNhs8+nRTnUWIasa9xxgbkHriX4GGnO
3k9F//FyDzejVyBXtdg99WIXXxO9ruOEopn6Vaxc8oT57vW9JnThI8NzD0uJBionFS3/HDJAHDpe
6qmOO1XqLVomKRm8rNL+K7rSfHPrUpdBuyIf+iMHxsKMsj+ftwoKlVCJgD5WKCt+eScU85mG2ixM
nZFoMrnoISluLXyd9u/Zpc3eYJ6Q0kN2/x845/ftq4C6sQQyXm3UOV0oxttUQgECfmKh8ghaaetR
uo3fDVevt/upU4Yft1R8YI71JJlhN+75MPsRp5JpDaugxR6uyXpaJrbUv+Q+jvy6Vv65lygR9y/b
o7cr65h1km/h2K2lwyROe6Kt9dHTJHdzRvYqA5qoRO5w6Ris8xXKTXq+x8VgOsY34vLvgbe9X8dl
uV3Jxu9GTMCNGZ8h3yEyXmtHIhxFJ+ED1ra0PCQ73NFFtcLxf43iyKoy2m0OGJt2b8W269KGOZLS
NbXGlllv7D31QZvBHuROaV+seUHNUvk/41wPecU8BHF1cORrUoeem4vNlPik4NX/VVdE+kUPGrRA
VfBzzdRUOxtFi0yDaRBBcP8p/raMHZVRRWpkRBL2V8XLCNjnxLymmBgp1xQgjHRwW13v8sXGI5lC
xxRSlpqzBy8H42cY8vbF6w/LcImkOcv7F6wPxHVvgrF/POuuwoYdWH1U7SadDjutOM+592Z3AieR
HgpE289U0nzGi3+d2CQlVKzR5Og8YCkos9O6gbG7hqOG4eS7yJilOlLWJ7tBS5PszqSNC2ihiuRN
0Q+M8BEumEz/J2/kkmAAFCfvZAJJ8c0KKLrBONy6tbSLis2/UzX6UHvqcxGlHEs8+iZ6CsCOMdxj
IERnWaLVypULFffDv8oYJe4E74dhwdKdIU49jFjshjErwqtnsyrv7CzyeqVdJM81e8utK0JFWqDh
lMs0GSOSYnKZQVW2I3YkAx5bQbMrwaOacmw7XHA4KXnXs1qTZPi52hakZrfFuwFsoo0O5/RGifQZ
Lp69XafsdwYtT4FhhqSBz22obUvhgBRyvJ/x80whkatt12V5gUuUUxYONGDoRptWjGgtmDgGUttV
fEY1qxu7mmHNSptY2qiFNTEOs5q7JAM/QPhaCHtwota7ivBacdlU7UzOQoa4gk8AsqNBogwVhy9U
tn4WMTP72ZY2/m73XPn+xhhw4FdeTa9/KPGBmWvKY7/NIXJfDxoJxCre5Yax2NN3TyMHJlj6XkIl
k0kXUXwAKitEyHxcudhnEBIUOfLIO1f1HZ9Qft/Hzc8LhF31871z+RIIUo2p4mkC/cwIpwhiJ4Ya
FSBzyyjE/EnuMe3tDt5a+f8ecPdLI6PLK4UqiLEVO1ha7lC8Yr89JR0KGmuGlXv7LwuVNwY2dBuu
srlBPoIPedGmRr7OY4xkQTPZQ6Zv9YNSxi9/rLSonf2AL/4CiUexK+C9y3oZIZViVJYRIRr7RCUo
5IHXUHHW/4Xl0cC7JPYTsL3Gh7sUktSw08l609i6PqpBcgxgG5FEWtaz6sTOU0xxFIMQtfHkZX83
oDVTQhOIFURzVTKYf9i87PQX7qNCA0gr0eFukvYfGIuIgMard6lqTDrMcAcId0/9u1uvJNVe0e7w
lT6geN3g0XGJIrdxqoziq7MNTxDOKhqIfxvD2LcFIxGjR4YRkR99WxkdhmNSYrNAnC7m3ef6ETQV
lS3Tw0J7zzwP3n+IhDAI89LzQEoeupz26zBeTIU82t8AbcLGX+SmjiUQfOuVk08aCmMpzdpAwWZK
9Aixk8wmeYuuvUVH9w55sDb9Zt/2qPalLhgm0tiPli++fRL+MFJwYCgefJZRfg7afOE6JARYQgiG
5wVGx3sm6WLCKZ7A8p40lxL5O6qGp67S9s0A4DZ7sGslPsQNK1ywuUDwxu4nKFQWdpLV1us1EL76
OifAg8VdjpdtVglGM/+Z6A8/nNBl2YDtnF1S8EYkmOKYNqi/VcFn4d7XJvOBdITlTI9JbD8P6unL
FJqqrVnl5zY+r7ljE5l5IQixbfrxbJzjpT6BRhPzWfVZCxQnwl6n/R+R9xr9IB+5N4lvrWpP13Hy
eQLnIGFulQGorJBGepG5kXEFZHsf3GIw/i7ialliqwk5yo/1/eCW8cKqClgDH1h/TZSbXEt+qij5
ZjuRvzPJCiERpx+n9t3cUFT1zNZzZfCyyUPVBC3F0IWOwh7lAsS8StxXJikVuuVLBiY4AXm4zmxl
u6CxHo8YRZs7eHErn0W04FMQaVAbgL2wjPWXunS15q+exa/3h7vP9xUVFH9Tr+i/PFri8NJNli8I
yoRhPfkG6anWva/QqlIYGMSlCJwmCrGw+BP21q5bNrWnaQ9fSq6JvFhyS4N5WmoSzPtI50Xcf2pV
+kzyUC+QETePx3P97clntadRc9dHPRGrzQ/aJWQZ/EtmXcapdG1CyFR5hgbXTlDRYWen4w8XuNcV
HtQeXd4qQfl5LOL6ZVV80HpbbUdhXtc5rLzLaKRiML40/nktBUd68PiFJC40F0m3wcmOPKM91JYL
vCidRKzZf2xF04DkFrZmMZTcBbmsWk8UbkfKKvoL/38P91HoxaLHDymQ2tl7fi5XlF46G3JrjraR
xXK4/Wqd5Xz1XXT6jsIqj0UlrsngiKgDtJTu9k+XzqL62UsGnGFFeF8Vdj/ol+yzUU//dRm5m9N3
v2Jtqp/YUQlaq15FBGmU6d3WVkOijLEisfNREdRxLyATHolpHjr5WxdO5KhKGL9E8fV8tK3Ns+vF
i0WWn7H37+B5Pf8QqFm8CAmmfwIHXEB+b1j9SEEmij8eduJnOhP1pMqjFCXgplTO25vdCRpd90Ok
LPp55Fz1JM8n0u3QK1KltcYIZtcnDP82E2Y46dg3IXDahkhNx2LOfIUK4+x9w6yAfXRoc2Xjq/VZ
b3Au1TjjnMkeFDhT3jbOui0IiJagyUyaYS3746ar0nrOAlULurP4XoNzjMKwHwQTCJy9lDXbx96c
tYtRH0ahLUwPGCMcV3lF+NttA1GDJDq/cnW5B8qgPmWrp7Ocd6AUIJl32H/0OZgwqJNYocDGhoMh
fWVFlsLSbx2zC38jVhEwzAH3Vvn94zT6jSRitihmPSxy++/wSiOrz3lN5GBtYlSEcFxDzrD09RUY
BK0uGsmUkM67hf5CVltCcQUlUrB2dmyUbVjWbafegHsr0VWr7J3yMAM9EW1ebVsSSOmyIBXsWmEs
ZPv+rnObNlty5EmoJ8wkjwYWscWYaIiLqQYUIJqIjrQiWmX23L2TefnxeNgm0IcluesKNZRIxDS+
rfz4L1I7/JbCPBvJB0/L22sZKxLXPzJ7w8cV8NzvSiyQoQ7f/+1XPWE+QA5SUAnnVQMIDSEeW50k
zWEkpYcHa/lPyrsxgKjavYFGHwmJY38keU29onqOHPGXMJMeuOOKorYN67iBFDG0Im2ySXRK83p+
qww27UtkKuz17i/mFa94X50sakCLbmcnvZepKuAEkYQiqWh9Tn6Hw0bVnynkctlwceJHfuqC3xPt
JMtMv9czQcbE8LGo9MJGYblYnRYM3oQZj9N5oG7CkIgjqSxBvT4YCzFIjQe34IwYAMk8OJt0zmmk
g6Edk6NPmS453urMAXlVKHuqd1adBZwf/jl7MMvvKNi1o4jObzDYTc/SEeIWgPEm6+f5/ytgXJb0
hZsF6euKs0E7Y+YtFFKbHZjCR1bwX5/6OeLP4tjFPddXGvbVfNkz6n+srZ8Q8JJtKoUmqpgUHuzh
rL2d8Rsm0kSwJce4mbvvkPIpK22gGO7xmZNwSnnaWNosx1IOgd3bgTCYh1ZDeqgDOiCtf4EdpxaK
l7BJ0r91uTaX58AvmNJO7kXuihA7ezxla/z1IYjlA6KRYdJKk2Ml0gkGXJEQJuWtkNyRmCMS5KF8
UaGT00EQzwpKqzxcfj3seQ4QL27Vnjb+7IoC3Ttb5EH1PADblRTtjpdHxbdAEnXJADPeJMaY+wVh
Y/ALg6AIb2Yc2+lucGSdIBtOQvgNDj1mm0aKTCUgqNsx+tRaghWIvLoVJKb4iGpSp6uQGLyza4l1
U9HktTvB1Xxz2oVN4tQZPXxHgAVxydEnbiRPbOXkYM9nzg9HqqP3kUdqTuuY2uHASmoFZ+3N/wBP
qsupQc82DbTrxhbEatNGf03vOSAFz02q/RAZXIvkBlJ0M816KwB/+2jfpN4ddhYRTpu0FSogGj7n
gdjOO4Bi8Ugrc8IcT0lGk/BmP1XajzWfZ0s0etEkatfuZdZiKoY53irG8GJJEAQxEKLOUEMvj5e2
TdPbDh+bz+EZHObQxy3v8kI8JWEoeGSj7EA6z87VS0Yr6cyMHKeoGt9DGG7BLC2AeZ0Zud5t7Of/
D81nW4/b6uC/4NAEXfthEzEJBB+SYuttXzzfvH9GfkWgw5Y6tdxy4f1Toe6yAO7PwXKH1ovNrNRb
Iz5cfmbg4CVldKPVL2znKz0esNm2a30QsX6TVj1vipEovmEwim/iU2/UKycFhTjG5K/zsOhJZiaq
FiAGZ0Mvihrl4Zc41kS3AcaaV/BMtAbPVC2f4fRImoN6vQLJ2DSLj9FY4vL4mxyZiHUMeQrGeuah
shF6yNcM15/v//Kz3nJtvQWGnmSTWlehzrhXytIFBT8EzSZ8B1SbpaAiCBBAVTqTaa1VR7kN64j7
UMuWCWn2BHeGlNF+TBsUdGv+SlOyYzjEXwpfelFnNu74F/U7Xt4KqOGgEMumLa2AuzlMeQaxnJSt
CrezO9CJQixm6k8A7M6usUHOPrOTZtCc8pJ+3NF2/u/DPPTd7He1MU8NPx8JbqJoh3qI6FD/Ww7z
EAm8qxW+DNDxXd9P60I/XSkFh+JfhNqtj6qnZXs/2chHVRkEFuq808jP2Wu81UQeyzbsiqVsnfJp
a5PUWkXmsXKO/3Jcx5IiinajFzawgkHRLeQNM04gaf//hLEi0e1CEMR1oh1u2y4jB0YlP/K9Wx41
E2RVxfHex27vp0qrMnuOAt2DpvHrSsGIjFT0z+9UcHKrkCB1b7eVusde/ltqjqtlxoXs9RA2TGvo
yC3Zfu7vLj0zs4bC4Ka0tPWufylfYMmrUanGPPPe9drDuaEgmsTB+hYTCvl0vAwg62KNHzPZlsMf
J+sVRhRGNqjQSLAzzRan0MtE8sFKmve9xE1mS7IIvEW0zhXH3N/dY0wFq9y+saz/JVcF3MmBr0Dl
qGVftTpZ03MHTA8u3GAyDn344iQkAQE0QSbwfOxoyIVakjOOODgX266jFYDtYQHG1EtgeOyJ8hDK
qPUtJVWtXfFQIRhLuPVpjBqBsWsTtDphZG3/L0dRr1ozBp/okioMs80COI3Zx72gesbJIkhdLZQw
nC0FW5PnU4TvcMZHn+ZHMS4fjJwbfiri2f2YGc6dsIrqvTdsX8kz0d11lSydqgJjJZBOlAhtGQO4
ZsZeWZLR5QOZXDNR8pZiEbbXIPdMmg2XYkU2weSODtqfBHRQ/YDSsW6vJkdBrPDICDkansyDM9b+
lTzCQ3HJMUHv0c7Rl96PVfW6IxyW9T/tN1QJJGJ6WTv0Ttt0vRv0kOIGtOi4Vs0FIvLgFyV6AnUC
kluDgi7EpiTrxvwLGRnkXjauGbtkieM0N4VB/KSPXk++94cEAIauWAioWGhyXDmLI30+8/dukCjq
yQUAS8HpxBABGBiZaNzNQIM7wM0u+zBz+JXRyulz5J4dUOGU55qzRc5D2ZGPfGDofRrfpi27p/2z
0RAOuK781a/RnxmSLcqQHlWxtum5Gw1kj/OiajZHQyoC/k3wtdhR2ZmwXYel+sSVftbgV7M6Tt4s
DtcDSabdnxfL59PjBw4tHNrWAqqlk47XPSMQRkryVAClI26IrYS8KSzs/yNop72+n+FhomL4KLIu
D6rsFVcro6KlekySsAR4IdlTsfMJLTAmljbJokoJkpf6YfGGwICyXwGVFvpNZOVLKBJBHsIoLYIV
wv0+qjN0WpI2w9+k1VuwPQnWG/1uUgvSqN8IFhG5M+dFNO2NcIjgdvzSFYKxJRLnciDmyimOMsiN
J5NJs3q3CbP1IKm3XIKO3U1ylD3xA6iyUPGvuVJVspz3regJEgOvF60Gz1TgckX52vrlWhPRcbso
XJdZ6COTT6nW3pwHvgNGbH6DnR/AbbxanjuiQzAktOvm4aB0plb61LCtWdYOxGieDW8QLKljfudS
2e3S0jhyO+2eKEDbanKb0Cyq1A6pcqK99CqH08Ubr1oA/otdgyEXMeGLd2hfrVgiwvBHyTrNVLW9
aicNz8fnV+L6KF/iuEQbogom64cC/AXLUixTyiL07EcKfqp/DOxLAjh+98FZ5SxavBJDvAKu6kl6
g55XgRFu0IzURX+4kEKhb2sFXY9Kb+HHLNyi9rrSik4s2iH2QCvS5DGUUQs4gyJqame9gJCGVEwG
2OH7LmLx3Veuhnk/GiB9YWeNrlpt6yOLTcRGpkCv3dhrzkoDF8PeF/hOyzrMRwvzo3B/qcoA35fw
f7XQ7M/goq1Ud+01ozJya9cKILzqlSLta5bYaeoUL7cPt22zw/vXA+NKKRpCO2AGEE9G5yWrs1Cn
jdK8rkSoPyG4l4/El+zqtgCHMhbXK0wZuD1EF1y7Mj6jSPDl50mgoqFfJ2JIfU0vQLP7YYbo4Fm1
92jPvpw1hvX4oBLB53s1ZVzfuVHGH2JcIwJN8Tg0urQaV5NilAO6ABlJXEQ0tUwMHa9X7j1803pp
M2uWRz9yOD9yl/L0vCdacwrhutPFkoCoEFIW0W51cQRthukQa807cMh8w6wznB684j5eju3FzWJ7
SR2F7IDmzftmQQ/Fi8RFvGP0VG8nc2WGfwR0JR6SjtIuV0Qt2P6pXo/c0pjVS0Q0U9GH/faMeoAZ
HMR1Q9x2JjdBwgJOfKwmCb30lUQFzj6TodjOYi8MO/YfbcbuoZNMKU1YoJ6tlOWo+MFssp9JaXzS
gaTzkOZUmuFrZEzcHnNIHJFf79lInNfJlvqaPnRy/wHvbf8+zP2sUlXkD8cM9ePaSiaC8rqqH1TK
gekwxn9ecOGQesQbgnTKI8230UUypagDy92Fq5QiuWH4tS8ApJPiOVPZGnuOykVqpw7zkB1oeI0u
jhidhC43kuGmoZN1tvz+KAZW2LUX82sLqzf9Xr5ADFpCb17otVbt6bVcVFcEHPxUdKJakYG3jrcD
CEUrQatzCR3E8m8KDLC4bZgW8JZw4z7mq+QEmp/TFErHFbSX8ILqssKUh+5h+mW/lNN2l98A77cp
vAA5syPSOM03Hudsn3YEHUr1cByL5My0QF865AP9Csfvlow15ZUvctnVpSyBdtmdyaYaAS8jrXsY
z9mOgdqaTZP+8pimWXJRPqJpRJ3fBNlXdAcymxqRg+UzxvT69bhCGBSNdsT5mdxMwkDXRxXx/AUn
oEapshViOzL2CVyeiZ3woVh6q+MUyGQM2hzerk3nJa1MXN9ocjKyIDK7JzBD1XcUtxC/dfSznDwU
ukz8xprLk02v0O7gt4wYC/5s6fFwbk5l7gptQWNhz9qegKDEio5EMKFHQGC2AD5iIRMYKr2Ka/cK
ce4f6jPvhIQVe1frS5EI5fQW14LHGXCKUQ2h/9uVEcZaXqI7czwJa9EuQlHwrmemqUsgz4zb7qA2
T4RCD0wUOph8g4vgyN6cE4nrXwDFm0dhP+qqYgVgQ8A52Sflr9WM1GTr5D06l4D6xOMuzftZvAl0
Kkgrn6v85bRga5v0A32i+1kJ1okAvwWswlBr3MpT8M3kGiALIW4qLPekyslE1pa2hoQomgUIulWt
r1GpbU6b7hO/H27g5Ok9POMbDK5cX8TQ9ObN3yG1uFG0wURFjiCQcssNv+NMy8GowdmGlBrplI62
UGDtaMbNbBIBL5ZQOWFhZqesyEh8KCeK1NIIiEO70MdB3mXCbBoUVXaVVfSaMR/nHpNFO6A+0ARK
KH4Y7QNrJB32rrPAo1UIg5QQhfD4syVQqkovXVD4gupHW0GUwKFW2hGbeiu8DYe0eKDIpcxuLTJy
rhoNBGHEC6cpwNbgA+yEpI2R0Mzgtg32Cva9V/oFXNgo/WZKs44s06dVgH8HSQ6igc/f/vaFtsn6
PaElfNukHEOemwYYHu2GrsyOWuDXfkylykOso7M24RWI1EA3NgWEuxiAANoB9ElyVXWvXpH3CV88
ulSYfamaf+FzdAG+sfhnCfU1by0kffBJX/C1Myfj821NP+ZEvc2ORBdq6Sh37yRKEOglsmcox3aO
LHFMlWgJpM7XJEQrQfFyuf9vGGQchWtZNDAZTc00fz6+C44o4WSVLSY9ABtB80yU4l9ge+4hooag
CI3yVBgY7dHhgAWrhELPrnRRffbDzKjRWhailnk90oC1GpubQkaU0TCNUdOtmXyEJ3J8d2ojehbL
7ikZzdBM/j6QZXAFY7y60mthgmtUlevcTv0URZva4IkBA1472lr3KxXnVCd2Y1DFm30vTk7unll/
S/dKDQS6AKEESwim1sDgL8+mgBkyUP4XcI+r52ku+FWwpgq+Kf7t9YzY7ga2giAfhqaAEl2xNJ5+
QHqg64Id6kN7CJoTEVG2DTU7Y2t322iWKebaoQUFTAw9LKJpnpZO5Iom3lWdWWslsSKJ6IsAsNJ6
L8M9afodM5fz+CZ15miJLLbZYXc3YeSTdTapT2q6ZBqSts1rEVhxyPyAe0EezDyRmR0uOZtCKBpX
zSn+F9bfrPs9N8ftCQkKw4SKXSxMTxGE2iD9IKyOkoNu5PhSKQRuOjrVRX15irIn4EpRq/+FE+p2
i+trOBFQAunhC3oFw5qGI8cnPcMXKHqj0gq6TWWEH8Er6tPwM4S/uPMwLcBkhyc6qR58p8D/FAQE
x/ymh1UanCfVMKE5HV1Q33qRKpMXqhOW0uly93h68jh+pCnz7+D50jWNCKkAHjCJX8c9Nxku4I0r
AWmc67gDQnM0pavZWv02wkdfh98nX2Uf8+fX7EsFM+vOsmKiZaHt+IwT0hhYm3pKVnyLxgAfb4Nz
AEC374ofisDtn0sX3aHvgbxAxhwymywL803jK8IXwQaAq5mY8fcIRooxbTUVj4gDRHjJD0bOjnyX
t6B4QbC6Bu4ZtEIWCEJ18N1wWZuD+9rbrtT3earNRIBaMFKp29hlrRoheraGdBaGDFXXmWi11bJY
shuhcIRQpZv6u96c4tjxPzMQ9o1rxP6MueSmj+IIDzgfdZBbHUhHdnmWJuFFE8a/mo4czZwxBsxu
iNdk9G14qdThnrEAFcHXhStrJ7pkMe/6TjSzEpW3zJ3SjWboGAmt7rO3uEi4acs6pSXmFXb996jM
r28ddg2HlMTCFZRzh1u0Kt6A9mL6D+c5Y+GtjQRzJlMyuB2EEXH+vWEvVxyh724jjpP0IWmgpj3v
NyFqvQGtA3PunR8FtcokimVcp4oDWvRmfZO8o6z2oLJk8cptCs3fawxTfeWugygy72fRIGYqz/EJ
wpkf4Pck/Lu3PT4n6vxZQzcaJpryfp//snfDdEK9y2TRKykiBQkNTb/BCkoe5ntmRz/VlQP2C3vN
9fF9DStl1hdxY+lxzeHrJtyY3BVsDaBo2cFQEoCbPTUDnMzfy3ld8P2blJNPnQ+IzC6uEYmzoykO
uPizEFdThGQsDYrZ7ckOjP5OP/9AnwXiRlWgfpqpc3n7oMkQyG++5HZtaXbh5zaboG2cHW1WNh3+
+z7fBq+vGwnu3yOm7xmPtPj8G7gXqe/xpYKD+Eaj34fjLH0j9S4T1leP98GofQpGlOuhEwnvXjtl
jW1K94muBV5WUEIKLvDvtTP6IDbbyynqgrR9V3qPXDUH+fug5NsdWLRrH8AdezZDVvSlK8vajbdz
emBOSrQqzWnmeK7wkxPnF/RzL0l70jZNiU87bysTwhHxAeGHcQAMoIKvRLCb/zCfmUaTwre/Nv5Q
NI2hxje/zlT46ZJf5vgcp6mSB46wVTvTDv2B6IoN2sVi2PxQKRnTI72WAO+m9sPYzTKRROx9qyxh
TrFbkEPPBJmTanUOxrMGQn1js6JNZO0ZiDJzTkol/4R6cBt1WHawb422pSobmI3qpDPPLXmd/t16
anNUnjjGTxwFd5KJxCRWY2ehLRXUeEPu6hWOZpgbxhqR8HplFncjnSU0vsQla8pyFEtcsyN1y1GG
/88ZMvIMBW9Z/PfV6G2Vnzru6DwJqFd/1lThC0Bge+7p+8Rq6xe+hsvN83nsz2n4JXnZuJWn9KW/
rgWlxhiDsa9S0uCXKxulHiGzn+r7Gm6j8D5K3t/q7Qi+Fmr5LS9xXbULonQPWQJfBvtogpvKYdZj
yVQtt8tLHVOs5TCGI0kxzQC8mb1QGqtmr2O+UNEuBNXQUuTYCQyq7sLfgWmtmwxSOEkty9clK/Wn
w/7nLHYug42UdgqF9/u61n+9qpUwP5x8ealZwgFLB87tkDDfHXAmByveOtmxIhLhGm/gNtDf/Axw
KLpEvutYSLsr+NMjB3uMMVSi2Xy9QL62RRwyOXSCsyO+3xNUNCzU+XrrH/1kUjmOk+L9GPDv0X3P
Q7IkpTFfXDqWEI4bukkd6k/5rPKf5aHKSw6E4IAqJ3t6rCbRRZ7z/+Ulgk8pk8yhKUWGayJpzDw4
v7hKC0HWVdY8AUpkltoaTP9OCxuyvefc6Ogw+ppbavRVvJ0yB6pw+iRVvubVq52WjpOaK0lNfN27
ihFtcrFD1fh9rpBdy5eanIRp+1RrvDiR/QyaZLEDjMShnJNCZOwbqlP6ImYCkeQ7xztewIYwZqPF
FPXAv2XrvRQJzfEJF2O+3boghEHY3mKKUwHtG90Xd4dTbaZJK5NqzgPJZ3kVEX4M9KXkMJqUNM9/
uGH8rMG39VfBg47z/iK0SxnHi5oCZQtrmAjyXcjOubcwFAwsdw7XsQAB5usrjxID1NCx0U2gnnTB
ZNOfmedAn+0kcc04UoSXKd7tE8DqQ09VmGtM6sLkuTq3XJNHqBNEfFxiNAZ/sAlBkOpX8BuFe+An
cctyWnu1mb+c7uv+XMer3DFaNunlw+bMPvuh6WvzmhJjmaEXZAAVO5GhrbhKHb797cp78ZeaUSIR
yiMf+KHDtUVj7yEGxrxkF3xPoXr5JALK5CBP2X9cEPz2JpOwO8k2Bw5//FnNwzbWZaE7x463BYt0
JO6PtPZcyxCarJq6h2J62Bek1GrUwp9ZQUaqt0jiuMNkuWUGsrLU/BwkcKQmucyhjnonenfL/5S+
oKimdUdnpC5QcPBiAiI+KpBjzbs5PTF6CAmkIG/XippkITcu+J4eA1ttzRmjXK48Gy1OmasfVL4E
Dr0MnBunEJ083zNK/xJ8aOH4apTaTh1SSu5ffld+vEFI98cjPt3fl3Wc5UoUKSyj6r1a+VOmb82d
m75izbD4bhBA257napdruJArapl5iaPsm6DLjhzY7GSioBFYt24VJs3NoiD/lOrunKlxSFjIb91N
lEVGElHSGxq44zL66Lwf0Ck5gWMbXEkoBSqvzU1jeBmiTfzYZS1oXXRIRKdbllvCt7/Eo9vWWZmq
vUsFGu9b34N2bboJHyQHf1nma2sMcrubpipkGwXaMZjRfegDOIZzoPxh++k++aJxDOFIweB7TVqp
cTP58vpjciyaXJROUa7zlX6XSXvUc2DLKK25BUuz++Kphxpvg0Qm5iEM8T1+5Y2JDsSenJeB+NvN
PBry5SEjlUCyxcudFViKaZ28kY+LB4hqwpmUz9IfZYCDQeHVySX+DCYLGmrW819SghSR+OdPjt0h
5QrzRwo884cpoMgflw8o/iQDttLNsWrsgz9+IcvfZSCuCiIzyP8wiWa3UWaYNhtL8h5l7lC0Q5pR
YQMSe70yPyQsSFpgd/VE8p4npehiZpEVJGOoK2JcAc0MN9lk6ypYvMht6l850afjGHchwBBAErxW
1SJMp0hzmmI8tP8RPmTAxDzX4MdoZPW1bhKoPnHFaToPFnRCzo3U3qiaW6TnyckDtAWvLhn+/N6e
TfsuMXQMsGqldtLz2MESSH52ONgbOLN6aiAI4flOOg7pQzwgiHOQ1P0eXfGC+9NcjlCfwboXcSO5
knLCU/9/VtE8n+Gk+VEM7H2FxeIVHOTyn25ZbL4ngo8SpQGy4l290G4exuf+3sGeA4uPBWka62Wa
iLZ2dJRwz/InFKWZsbhhHCNmatSCQbQxrZoajO0X1UkFgNz9xjeOaCCDLgHjA+U3v7GGM1rSiT0I
QovLAOTaTjTY7T5KiqmVnBxPKSA+umFifO7/7JZf8JvyI2207b/Go7UPh62Gr6tTA/vd0aWic1C4
9+nMvM0cOy708x2bTkt0FDePVHmw8mJBOl//S+n1A6o/Q6Ul3yF0O6lOZ43LnZ4FZZyuqtlfWQZy
NpAuaQOC4bAkXDvOge53LwnPPHQqMkWVHB31yCEqksrTZEQbHtMEq3PAhFystsvtTr19hzAX3uUL
eFnZHcUuRz56Hy7epFVwZPe00vmSsr1GZXeLh4WIrCwCpExQmB4/Bmmi8TzD9Aynkj9IXnj+Fz2F
2XquHtIYF9hb6FVNFLdHQkR0DAwKCtGYIUQ73yBBoMo2RNe0FMwN99d8vLXjnVm27uigSiIUnxux
jo+VfkVzTHhRakeK/DpCZYKnpUpkmBzH3TK4EB8WSBPNLFinvqUg3LBKjOv6sYwQ4C15RWwtUo3y
X0b4by9kLZ7i3buHVZaNSSlkaoRAs8JIPHMFhv1DDvOc4I33dFqYEOALyid2vtj3onlHocP06hy9
TEPJRk55viGC5XP4bbcboCcJmIG2yTcVdhBA0xyOVTbRDE1+NceQgYmn0NukQYFsO95CPDH1P2wh
znR0RFEJ66SphDeYqd6s4SM/s8i856kIAu1W61c76SzQ8HukDez62LrC3dHXcmLWSk+j/nFP4N4g
pkN836yIuDmgLvhvgWj45CtptOvcFXCZsJzrf0+EIJ5tRebewARIMF1or4wuSgiSd1UrGxTsVPAl
1+hkxP9elMaHPDTFuW6vknZWinHcLCKjX690OInThb83YQUvILnL8ATemnEEjUuViq4Z3aFxZ2X8
wQMV6ZycetByzNy/WU8rkEhU+2dS3K1Jr9KK9JLJXgQxhwI/cXVaQ3mFIeyxIi1e1uMDOnDR2QsZ
a8qqOVPtIqBFIje4zf5o74PHmZH8vISWD++XTlTdm5LtKg01HJbtsWUTq73zjKmXa1XbT75QJeP7
fbSKepzM/hUm57cdkSyixb75NcmSmgQ3asAXHHZi74pluL7l8iUg+RERhuiFqBNdl3vhcAzyh5ra
0qWoklhqE4qj+YM678rKFHgDB+UwDFYNRyGHaKnOJnj66Yu6u3zuzGKVG6ri1tw5FuTWpd5bzvem
m/6LTt/qFgJWTUTl666XlUYhXS41MM3K8UsYtVrCThdNHNj1kgIXYGBCjF+y4Nc4+I4i2V2hNZ3E
REfz11uMkUMPIY13/jMuiiopioViSZ/sCbTva0RccHkyEfnihigOSRXHPny1lMujOcZi+IeFYs5t
W7RVsM3kYZ7UFGX7z7aXjoph05uuHrqO7A4Rl7u0uUHod5CxgyUpTvJPwoCB6p0AKY17rNbAEnfJ
P6ZDVGs1aYj+1mJJ1rZ9CnqoQ7WMuABdTCxNtYiBGKJ1Bz7HgJWQylGsU8vG/rOnopvSr/c5YbPE
UgbI4vB6GUd7bao0wZRtsu+KUvn4NIP0WvbO0NHjW600xZutqcJJptI7v/lBdt4riIs79stxXXYZ
aHUq2n6NuY2NRSbxZtmff+zSddU3E3hvBCJFpYaEYPjKY6miYgLFzgVkuy3+5af7anGeZPA0Fdi5
0/wMt8SrzEHIw/Pv9c7UAmRavptbQSF9ChsUFn0Vcn4WvfGqfQsCa4hPRd5Y6EEfHEJQHy+aSeod
WQj+MMxmIy35vzGBzBOx/UQXyvIAqm4EPtKbQZtRws/TpnqVI2wC+ZaMumh22SwQl/ql0NF6Fkfk
cKTDSK3H1+TmjlBRoccBt8+yqqVKFKu7h0Og0/kbJG7Gu8NEz5DHO0GpabvmD7xbi9nYmSYyKVKq
utO0RSDASDkWIngGSry3olM9DvpNhbSqGPXke5GmR13IU7OXRAMLrhuPu/1QKEYyZil41/IqMLNE
nZKDhTy1YqcA+xgKAy2hBdQtJeGQZs/PhoLI69FAlT/vozZfQAfs9mP8TdsBmleXwJ9LIAu1jy7P
fuAWO+uNV6vltPB5manPi60Rdyc9J4f6MD4oxSbiO7aBDYJVX9ttJ3zSho6kXXM+YmOuKX3egEv0
6aOM63tYsw9O7RdMb0V9Ixb2y0vPcy2/d0F+sluFSJ5LHzIdAvDY5wZo2tEdMVyWzLW0fJRKXv01
Kkj5n6/1IBD2uuxh+AxsIIXHOeScnalD8Yi1HnC/KTGbMB2iwmi6jSni6uQL8J4+g0bxXsWqG87d
vbs9rD6b5ZOrOZkfZPZrCu9sXH2NVtMEgrXpH/m8PjJH6OoSuz0XJkzAOIqcg9rKC1iFyg345CyX
1pV/SmQnsdYt7Db0gpkgpfxeZnqvWT4rM38s2dMaG+Zmwl4elTW3QkWKsdXyySblIyiDIKuvHLME
+b2W7MVkAIjtEEd3TyWBRzG1VnWFBLnpmThePAv8mEvEV84M+AhSK1zovdIQuiMlh6oNrWDG857m
+evvK/ZUJPI8hk698zkMeoQBPRWRQyMO3Dj76zXyYnP0iIxaSZ1Ay5Iy6+nXdnw+kZo1jvUOMhK3
im18yCwiHF2AFtDbFcjvXx1VIfhq9KQlppUHxg6z7rDFOrAlFb782V0TLlzTPfVPnJwEkVMOE22i
fV/7VlARLJP/It0yMDQiAa/ElKARzwMJ9TqUi4Ph0R/WRnwFcu2uuAZ7wAm//J06M3PkXmAirZYN
1udEXkxVZRZIn3AUpEFUTVq9j5k/i0hryACUsmgpn0Ol8CBf9+9gk5Ik7AcVZYnfiCX04ymG8BDp
ChVvTpf05tqn1U+AdidIhuJ5pR6UoloaQ/r4Nl6pcQwDzh7z6vjJxe4Yj/XzvJoawTOj6F5kkVkK
uMpZtldbR+mBcDuAerh9cAxBrSoabDz+B3RIENAS/DjrGcyAx7infLhm0cVBjr0kpybqkmdP0UbL
EYwanlCEcsEHhQg17026P49wncuMeLoA1CtVMRyQvf7X/aYROHZeCRYjlsK0LvZbyxCFsbA1aBzo
YQvCvuyk+u7nnqFbUXiDk9UGIOyjYHWRYcuXGCK50XyroDXDRncoRSgvNR5ZO35PelTVWQu8x58J
y3JQcUyCyOBLD3z0nXuTta3YZWjn0cwlGKoP1RUDSnToMr3DoGYX4fYDRHiw2YqiMn88EI5Nv4e/
Ut0ups/EhyCmteHFIcAx4UjicyqY4ODCGPtSLXVsfJUxqUhJgZd1hwmJ5OpVw5OzY9LOS6QM6c15
YdW8OvudmTIPT9mZLMb7wPVXUnW+jRZ6BqvJHsNFZrdVJheWDa8Tap9LQ/D3ycgjcfaAmYYVjhDz
VKOJ//qzVFfjGtJjsGQmLPdlyTYRzlPFeRgoSg3uk22mh7wmhVzyVQi9PbZGhD8XnU5P9hD/e9Jn
W4jrXYt1FF9sjocmM4+K/cf2TcVF1/iWuIoFTVaqteWFmrtroQI4s4VQCKHymx7aVe8oaoznSLdF
wrhrgpuFg5XbEYMsRRqvECBkcdfls9p3hLAecnFXQeS8+CQDdXD90hXWe3IrU6DTNnOCnst+VNha
1rZ7lNkyZ86itBwQXTwhzyStgNlGWOKFjG0hKqGbswAYf7ccWKcTXHsfZgs9tRkSeqAJt60D8gWd
6weZZL4uLWq5sq/QPxM72Dj+R1Kvd7rTVRwTBVmcG+idxPvkxFFvVTG2YgREp/18Fu+fenBxy0nR
7KmDIu0kE4WOr3gQ3jkcfaYZvwpwwGdY0VgszENdHoaVMf2rpjo/Z5qDlJxx9dR7TIOZhsyFt19D
e6XTcrxFtP0rk3oJ9c1nvR/qctasQpVhgifYnJXqX9yGds3fQwpKgObyq/9sf873Gy9PYwJWbHmX
koVOB9InNYDt3KLm46uvR4cDSFxcSJ/uKyy7iYolCb62SU6UR4QOG1WLlACglEM8D/Q2Nf8+QSBH
jEQlA4yLgEQto3OgPCYowhzZLrhJ6OCQRxlI4WmU3ydtD7ymb6tccnkV8RxcWFkRDav7/ih4iAHf
fKIWpeXwaLzTn9997zSnkKokc5xm12bnrpvd8GbbokYsOUguzY2OC42rkVlNuNJxxpaTsY9sSeR0
AYYV+7ts2Zwfn0AVwXrYJ1YFnKFs+WhWRbg+yMGIgHfRYqMwPB9S2hB7w9asEix5Es99tPGpLuQb
U56Iu5wozxbMC/elDCzz+m2g1OAEx+DiLxNikCq4oNdsaUKt4nR8jaeQlMAKiRQPBWf8ubYJrQQX
czgQSkPIuOiW7lkHnDK9w5oPt2cR+DOT8o5XtpI2yYV/lziAK4QDWN2p3NTtF7tvFuLlepRCxp2n
pBwhf22lvvMGDQiDbsoJ/HVhSe8DlQFPhGTTfsx0XPydIC8IlrdybbBMI7bqQcNhk6NdDTJeXIZ0
WldYcnTTgVrGAmhZaeUxpp8yYESpe7c8SnpV6EM7+EKaqjTkOBQtg/FkPCwqch+Ya3V2rqDFYsui
qRWiYcS8LzGMQcyeyUb7PZnxZed1M0DH/bbn+Dkfr6t0JDqAVRm+S4fF198We4GoSg0peWkAZ66I
eD+keuNA2iVCIFX2m5QK1BNZR9QxlCnJqWN8FqBWuB6/2nQgsMiLIJde4BneoPp0O8v4M55sPqNY
GnEn0AQliPRfcEMulzYz5NMUbgR7ax1iPI35vThU06935nh0fw1xaKYNV3zcG9ihyKDKiNPiZs+O
T1JbKKr7/Z122fbctfRKedBq7fyLSkTRF/mLj6X+Eydi36/CylMMTJv+Yy119uNJ9tAcNG8fGM0U
bOLXAatuo0sMOe1d/2OR8095gC+xUfTzvBqX35EX2CwQ9Swlz0BiD0VvgQi2WpOQj8Eabs90hhPf
qJzZKcaLDA807aqwDM4MzAaXLJveDTvfQFusJe7cQRhI1i9/t8tN8yxn+Ta/8pdkS8M5YaPmOjkx
D7wgA2wTNOVA0Tlo1sdzASz6EXJbjEHwR7c0eDofnLK7fT164kMdKGUH4+KD3r6sh19HHezD+DJT
/CmRek219VSiv4yooF5yU4QOS2G4/y8aoyZoGkuuLrcAR/6rechusTP+5HAmw2RlY0Q0FcP+yrNE
cv1CjjDct/fRxRXzqEMVrcEyBgWBC3okmv7OnGXzH4nNcgotF2+wY7fLaJFNzLbr5IRdVvGG5GvO
grf6F2agTvmn96r75uQWFNZV4Iu0cw8jtcCoBKYAuhicv+tHN+nE+YtbzZl2d8ibICxhLKP6iyb4
D21xwuBP2sv3rRH8SvDDez88/ovYS6+/11nzg/27nnBzWngSWuxxKXe90Futq5/D1nivZZIKsQhV
v4QyNjgVKUsLs3Xe4S+YmwSYMto+AT0+82GHb7iyuINXv+Yac4pm4dkpcBdh86vQJo+1qZO9nsSk
lCZjhNwVRWYH3yV1eLG/RlBufB3Ke1B8Pa7I5h9SXkpdRew8DbnWhh26H6yteavINljtbgfiia+c
w/1FZFU0D8P9qRsJGcyalOK0a1iNlXUnWMDvHM9f/GjlxyizBIULP0jx7T54+7aEVBdecCSdaxxk
gq0DzxhxjC6SvRWQ849rFm7NWec/kNWjqEfHp5AJihzxg1jm2QGnafBW+a1TjHDJeyEb4scnm1Vt
rZvNWMx7Ritiq3uU3wtfMvIdR5GX/LBZ0agx8emFsn8Mf58EiJj6pZxLuDYV6ugx04HoUWFr0tT4
D7hKT8nRUOE1/qnJtXRaKekp+XylletlJj57AZNDV4IfpeDjq/p7GOSiTo5DlsuyeLVhuZfcLKm6
bn4PRcZmpfDcJZRRjTIRD8uVACe1xbmIJK6OyBiMb3CWukQlnVcsvyBlo3KXVQbNTdQt9peWTMuS
cAF1vZJ8chHhI+q/KHJYHCWU8oaCMhwBgskx8ZRyw5s5PS1QsRiq14M7VQe5s1cMLLsbg16jf9Za
i7wD2Ar9LlCKGnyNVtOOLvm4118Ho4O9awfElbjiE5XFinmDMekjsVaNRMfaOOduC02KsJlctOfl
u49pN9yX+Xpl7JRpBVZ5JnRfj1llPp4KKFlC5/WLMbaPO04JI31MXL/5w2D3KiDeZc6sv9dvBdyv
FlIaUAQ9HeGQYaa9vTGmKwT1mZXgOoU0eypNPpY5p8FeaqJkXz+/wr2wMQoYZyBPwnomx33sJmfS
Wr6qUZf63hnT2yhhhS+NAult+RM+qZhZOxQVA1pMlAjCMLd55TMJU7EFMaH61TxeuFeppBNfyWER
ycn09+Rvau0hkZiXaVRD5J+SklsekU19mlKPg/wLGlqzQV9ovHQngW3GEHq4D0ym1SvSQz0Hm789
azBBV1ypYpXtwKwsGfO+puK9P2WmOgxsYDjLvZYvK+vG+Yf0xFSCljxAxGW0AvQD2Zd0yr5/uxxL
ziqnq+411vCJm4k7KBGKyuCTtZqKUH3ADufLiMxz6Ix7SJd7bb6zP66U+R6zlOtv9eJ/MCnfsb/2
pKhO6USskRhMTBuIUADEp9ioXSHxbC0dp1sIEHqQDiHyPD9/zsoaKV6ZT0yCLu5aJunrZlCRarc2
+GIFBlY1uAmzdJVytLNzTlKAOuzKVjeDjGUHvUIqZjjgHqmn7U1Bi4ZKBIT46npo1XUvvj0kRjsl
Sehh393Yn5rNZRN9hSCvYmdkIotRIVY/CgTpbaWgNQtK8/0YhE2VEtWSdxIdMGHb2yPNNAPXIxOk
BlJHsTVOz2sEjnCnXOobeaViQv/rKUA4le6ALY64KtWZYZC1SYp9vMuIjyo/IhXSqLLU9FV9fLZ+
W+xWLtZZErfCPnhV0Kf55E/44c2USVuWimp0nyPyCJGpNBL8ySV+VYAuU5i0+Vo3+bpb8PicsPG3
RqwcDh25ZsiafPhkTaXAqOk+Q0XvGt/SfUmF9HpXq0fScgCb+LpVunoucnSIIcwC26e02RdtW44x
LDa2JSBE4q8bzHx7H/G+Ue8GOILfYCS7EIDI1MSXUWSYxj3HSJl/Z+JaypWY4tk5lxAsjyjMoHiV
sk2hMCPYCdwcvTotYvsnGPniDIA9L7VJ2FTjRLCNn/s5HPoZtihBcWIZtv7DHMCkrOV5QsE6bQiD
BaVytSiWG0pz3GxBNePJLRZz8pvgoevQgNjV7c4a6vUVedPH2DWzMb/opq7T8X2JEODfEbJV5Eiu
zqHj5K0cYo7UvYCVnESVlIqjw31ZW6SaopLbFVP9ai4Lq1XW60dC5bYnIb07SyzKlHB/dIGzaEwr
w/Wc+z9YFQpaVR2oaYTIqajLvjcS+AalGUOlmkWh+a7NdhwdUKhmteeDftAlXbF5LYJkExwHelvE
rURJOdTHrVXAtluEInBTSZuH87LBAanCHCEGtOSA0ZPeSv8Dm15SQ4RDyrEsirExtzXK2nGgO9T6
X4Iw038fg9EW67LZqTT2GcvJC8U8xg3785kbBcXfAde2H7qyjHODkjO8YT26BYU+x9xWO9fut5t2
18RqaTtm+UzlmLpmKCXS6OyttmoOoi257bq+Bwd5iffzVp/gjbbyNtNGiwdAOtmbdTX12z34qQVZ
EW3QH9FNaFMWXxFEvpgbQrFm7MYBLrUd52VgBcvSElK6EHEZ2Ub3+IG0nqcLJg1LWKINTrZhTDhw
muddq9WvdHDmBBTMHViueKU6iXp5IBISCMrwA2dKzOzkcdqqSiccTLW6GuDi2UXUeFdnu50JplGX
yxiWw3WNALamdulkBocxEMeHz3nI227B/dN5RLtpG+z2Qpb9r5Pj/ovy/GxNrELIEyTqeKLTzW9x
LwLrXBO+2gNQxRGjrboWeQn4XQp4xKcGmfyrlRCpG2ercNqrJoLc8uOs/Mb15s/f5SmMjELDYjUo
5DfDQp6hLF7G+ob/LP454Nfo6Br28oQbI2J65rxjcOvSL4RbYaaCw/cyiePssK9/1VCeYpQT6a0R
vLg33c9uY0bZ9tUHwtOjzE8XqT8Z5eXqAZ+Nm8drzTCnPoVSMdC5byWlhSi/yPCXjoup84rTCtAb
8wM9ZlNVc9BcFtWkNMcHYr3WMLgyLZxzzx46mZjVbWXVlAf680ReBopYoqjHco4ZCquLVElO29Go
rfBaG12WjzwSmEjqtIw0K56CnwggMXjh3peCsmcaGK+K3KjAkP273W7enQETxwwBcZvE/PJ33a/O
5LQPUCIZF0NYBzm1yYytEv2HGMo+X9p2vCjfHvqvGfxrP8U1uYR7PYAfRTeR3sM/ismN1hTO8tGf
I5VIIhzbTgOmRbkEkZgC1e+7XMeRF7XQZ22o/9ep/NhBQ9SS6x8RJ045NvDddWvDbfHEnWXS7d1B
w6Of+4g4ON6CAmbB7e4U1/0zsQBO5g81rQSnFsX/mlVNwZSUxl/NrEj8UAt3EKfnqtOf/w41Ai4i
dytX6PjQm3BYcz2twXUIp5d8R6QkKztvcrLPWYxQr2bXG18HkaaG83r6OoSKiKf6tBaD+sh2lxJh
3+mXJIa2j4+YiR5XA8Czvzog05mmysFsEGdaJY9EAwvYLsWXQfXWycmqD4CmjUraYnDvx/l+1yd6
5XRNRHBikelVhRsKuWw5LZZKAxbvHRJdVHwqdTKgJiXvVw+BY06Jh/fpD29/t9jTzYv3VVNFIzM4
rTJlh5FJ7WsZRW5DwXPxbyurCpZoH+8d+J53TxEXR+t5/a5pyAbC7M69CcxzHkXZ4tgBuq/V0+O3
sV258K8VE4hB9aHkCRbzHk9Mv4+952BDZON++GXTIrJHItwXVE9+Y5Kd0J4s2wWsY823svuWw9mq
l5ucm/+RznFxVWbGjxWi8g50JIQEy0DHnEkGdLWeqNsMMf2IF2UOi7nUt61wCAHEnWPmsOkPgEFC
GbpwlZM++yKcDDEDDX0tdfbeUgaqJWOkXaDnMibN2ZJXPVya6Edlg+xaOlq/TCSPRcFY7OktqcNG
ayJ+1ZnVDOZ+5uYa4YNwt9zLNHvy8i1RtXgXm06nAmYDOnmb35yBCjayV+yXS/mYRbzl55zy86/L
RiTtk9S3K6YXLtXcWEFkjot5bQySuBejCKAjPLUgmLuNarmZKYzuaG7zdhWM5CgoB/1MsL8oYzA0
QlAFj8dBvBt4z2yjoN/dbBsOcKPSH/nXf3WTD/gkeofK4KHgz5UAqE9sLMqui54N/66+q7MW2tls
Mn5z0NIIM0ULf4XGKMLcVshpaoiw9iSTV0ccwPxGU9ZDPG+mou16kTkZYq9yzr19T7kRVxVOtblQ
s0b+4rEOSs3QVBD00XhBFtHo8024Jx3GKBakKSfLYSqlQPUlxyT/6U6TzlM1T9ZnleRtHP6aViKe
FGYRBfofbYUtDh4G0bmNAem58ZwuN1UggcWm2Bzr6hGGRYsODEzKrEl5NJkaiAnlTRvqJaJn7IrP
uvW2N1zn9xqtoNcGNETRHXXTrQq8N0UnETrlCvqswYbzzLvR5S1kbDyYK/fuklQynii0r+IUltpu
pL8BrO/naZuxxEn5ffHpJk17a4M609fu7AwPi5gbdkQTRtCfdjmguNhaDCWYC6CODE6QatizTx3O
pXpJRiPeGfRvKsamD12dDAYg9bl0OMhqW8aq8PNMN+RvfoK7LkM5T0XVxWjhH7oBE35Batll0hTQ
YbIdLNc7SZp4G7EVeV5qP1qb8RMBYCF/2E3uZ3eFGAF3kVTjwfLW+ATTNK2oFpMajVnnMRVF5KNj
xX97XQp2xiCbweaR70C03OwXMMBlFiJ8SX5WRxuApdovtDrEKUWKd8RsDcs0PKbpzTR/z2F6Cn0O
0MLmqskCgdwvnwwJbd7mLDrQ/L9ZIzfu/TkJkHiW54V2oy1g0tJFpIVBHk3uGUTCe1VwxbJdfta/
TUuHRf8uamlAujxpgz46zJQuCz209L+AoD7Kgk5DVkaiI3cewHjdJgq9/TE5P3SShp0bXd0NxzqH
MTrebqcMtAmVxa50UK0Xubn3HGGsy95C7KpM7SzTkHkq+Gw8UOJLGjP32szcZjSsUakRXrq+XtVA
3bSzfb6yMWXLUzD5Ai+wFWyaUZV+WDFMk3V3gonQAOCgqhLKOoKVmRS5foncz1wRK7Ju2NYG9Vmf
J67q8L6N4HMQ7CbTWArMsQU2f8A9QoQrx14Ejd0Z9KxMHuPT0yu/uMRA7ri48F1jD+92vWjEPmGA
4XCUt0bWDS1gVkvMqfcKpEdWT8szqTdYJX/tuoHbFyWVSsDOEA60yCJ2FF+uyKHu2tj8ftPSUuAQ
LiAi5u4W2e862PmJUFmeBmH+pb3znPV/u+Gsm1MiLa/FDKagAghxeSXZp0BiZF5huGmAx0kBy0Qv
s9nK9R59ckwyPfny+V7f6bBddwX+yVZ/tP5THmU6ztXMTW6YWZZa4GL7hawq4dhZsDNb/NQWDj1y
EQSPawIjCXM1C/BpSdnHhEv8TGvvb17G2dVqddKNkKF/mQR42nREh06A9FdO9r08+gs/ubzybWoY
SYGkg5TNsLowA1nJ+8ugS+pyUepsAR9jBrvV2+c97CoapL+Wr3DcsSQk758z+fpgtnPdtMg4w2+X
/eva22mCoqNfUOgBwlOCoxg9HWLr8pq6rRQRucOm8s/3BjnfKGrOtaGMu+gY3WwOgN8jvMbPe5Io
nVA51pgpa/tiiIBZ9EL4GWJXUDoqpeHowFGEf/vaHwOqxLFhbrpJuVqz5g9rNicaW8Q4CteS+dRS
c4w1R9RApeTUwfXz5D0a5RQB5nCEGYNDRd79GgxVIpwDMceE9mvG/5KdruDbnLjDiETdTPmKMbW4
ItGdVC5mVocb60G7hIOGoEApolfXkBtsjbguWvd8jXIDdfr1AOmQLILD6fWQ9M7rI/8fEjAj+xTk
J37AqR1Qecdd+tSZTwt7MGeWXfQNwZUz0o8PWGiSyVFnzRcT98IacqROFrweVfjIJ/r4Xh4ZgxZa
wtHMjwh3M9z3YcM43pI4xPHq+Ek6B2sJCWURuihPE+vr6EhbsiNoimvfKK+5e7WuE+CVfPJP+Pa8
us28J8dFrNWaNoWY3V3IqoDV4Q3N/qyDor/JcgCFMbu5mra87TlKqOHL3wSDoDiiX6s+uLPIc/+S
3woqkuRCVPk6hB3j2GMH3XijydGFfJzAH/EGsWSRjzf6WufSXOmiOAyc6sJNyEfToHPGtfUMNxx0
wP8S4y2IN8WA2H9rYRjMmqMH8uI6/0ofKb3An+VIxX2XZwt6l6E8GvTxJbBaOJz1In2l0d3my1SR
xFml+penlP4Ero13kieemZ7qI8+VhaLi1nZeKOKJf8UuMEjdrTBhnQTW9b16m0sxH8IbMBW3KFj6
az0fLGUGNFnzjxJhePxZw8JIJvNhnJKCLz7b5ZLl+H37lRUCOQIPWFdyzQPtKEbbt9HUQXGF4Wu1
FASqNSDWZeJoIGIFirHLu+Lo6NBSteu8JZgPAxN8BZbGzpQSxJVXHWRRwzsoVnENEEARz4mi0jMn
3imQpfw/1y2SNFRKklCsMb2+Ee9toRvmpfkTEnWP08Xglbm95my3yTDYqjWvZfT0XJreERaD3gQt
zL0RdGqyasjc3sXdtXdjJhuIuQMQlM5gAo8y05oZYhZWfuesyJhLi9BM4pCCCt233PZ0u/fTT51C
ccTJaGa/mOhLkZbJ0GTcE2BnntOk34MdIj/mGHCmIDeXptjsn2it3f3HhJm6JfU+1E58YV54OZ/2
PNTh1tHMYLVFVEdJz62LwVMyhZOUlQiAXY3/fg43RLvVoGrJpJrLyIQoek7T09T+ZgMVIaxuBWGL
zyXDFpE2frj56NWoydgFXXfdiiJjEVQBbMgtN7JscWSt36OU7gIeTaTYBgRTiQUJuth682FF2UEH
WEbj977y/K2k0u+YkZEl94zWaUQBkpfJVohlXb5BawYc7IAimBykU8T+zHXg7fSEfP76p6oCaRfi
xQCYPYTTPtNHBv8VcduDng/VP9UjeUN9dHou8AepwKJjqH58p/E07+snqV62ZvbnD7b+vH66Csw4
uuIIcdyaSGH/a5xBKuqCAVVHdzpzZBUjDZwoKezL0gCrHThK/XfBbR/Cv/NTGzqvbLHI+/Um8NUV
YwXxbnirTpGEKJJHFf4c1kx+w8g0Xg39lH9I7HfK5RNZA9/V18Tq2sZ3UNOGLomTC47gkVUgbm5O
7AJjxrCu4PJrJvrhlXky6QTbr2iiigdwxraIZjrALU4XG7yLU8pEh8dEmszdv+4YyKuiAEq76i9E
derf9h1i3LMm3afRWe0GaVt1+dax7uZRM6mVzOxzFzG2Hw9i6NmG6ZpqBvTH2I988QQuEsseXNpH
4UF8NAJMEobQ1L5hIBXM6kpKohMTukhcuxyikCxMfY+qDi1a1zK2YenK/luoaa4wOkCzQrJXhdGu
XjwP/4VbizleNVa1G5thGrCvPyABy4ia3drC9QNNAVObm+dLVODMGWSbpbIOA1SVY/FeLcDLHS2H
i8Q943zYRF8dORGr6tgJiTlxAgKQg1LSYoU5xuhNeKWFiwfk1R4Yeymhjt2ZVDQ17VVnj3LVNAYQ
zhCgPxAcvLqz2w71db42sqcCPqJxycgRS2b1Tx7PC0+yK/oVRx35YXvr5DibaydjJyaj3jUU6+QQ
CYcL93hAMJsa/rrVeyx2klZv4vDm/2CdPIvJZoiAQObhZHDqtbCljwg5MN7YPntgwawtc9xxT+vs
F0UduOXszjZvj5WUQFvc5D8zGD4Jvr0cb0jtMhIcNEmfEIBNtH6QcP2VnqSXx0rJx65dKOIEi6mc
zzKj+bNQ89oj9XLDjux8E5bLziUAK8jsnhUUPPfHZb9atLVI5hwlUai62xWcishxnBrKxv9bLSLo
t16GiYMMCdndxSIEIaDr4HFKgZ3iJ9xC9wl7Fr7qG7/C4Ahfg83VibaRJz17rR9uLk5T+ZvgreqO
1Dvn4lf9JqbkHmApGbcWIl1RYwdt6Sryf9SeExZd+vriM3J5pg+LS25p1h7N2xzB96Sm961cpde3
TOuPKLDM/BaXe3A8N/1vCZThjjNEYeJhnmhL+9fDHX1GBrZKUJO4rItsx1vZgF2gD1dWDPRSdJDX
ZtxF/NNUFbWGlTPRTJAhwzV2CYp/djNzcO0p6E+MhgO5C4jkfouUQcPiwSwTxjt1xv/57Le1gnYS
9LHf/8ghxWikVcZR6AsZu6TLkQmq/v9rW9wJTCnITxQJVS5r6kEw0kCXUbY58YUzmDX2fRMpOKcG
SzrHpz4o2gD+GyaMyOVTc4MPBGupJSjhx85+PVB6xhbKlPoZZdQ/JCBRIUJ+wDGwv93w9lmxjg6d
Kp6kVWxWgvNlSelsT+R+URHEHYqE9LLcT+gzWsm9vFbgKHya9jXUKiXmeUC+hL4BHbh/BT+c7Xrq
Mxbxtc/BXmVq6ycB8WrHBzNa++Lo3aQoCXtxAmLkcLnFKsXF2DGz2kkXJb1NnHQzKf5U+B79dcGp
Q6yWfAf/I7+t+EWfeIKfrxC26RcrSwG4neq79fLTEo3mtacfuD9/8HWkxKo7OPN5SVPazeBPj1L+
qmpBTgRl5Y6BS+AAbP2eY9N9lglBvj9i9BVfFdwLjFAZkvbwKMgLlxBkDpl1htbUUwHjHbjf5hUh
LzGVbkKmM6ltsfCURVHF9Ik9QlkXgWuw9L0yyXzMI/tsH2Feeio0hvJu0xHfsHG+fF+0mUMIIjf2
8B8O026tI1C+6UOcsNuigzX26Vuo38wd7bEIlzcJFe0pCppwqrldDw+mMWOlFCrEbloaSDKV7n8U
DJvTt88Zz01vwrRoL/OquktuHdJpFdiNaCVp+DmnUXY86pjE13IDLmtcCkCmsiXpLWqO2alxQBpK
Wr91Kh8zJyvbgbkTfB1iP6DNwm4cp7nQ8SkS18czLuF6sa05NYzHC1LV5JwVn2XS1+hQluV+ywZh
deRlkHSH+TobNrf2FqgHPpg+7Lvla/9MdoLwRquR5yYAoL86w5yM0q6QOJuTvR1NPaROG7E8bHBR
L7xUOFUrtl6uHSpbH7VhTofxZG/ECoQCaeKanMVTLYdLpzr5oCUyAu15WBhsmXQlOzQpQNdgOhTt
WSt4zheGZWqeHaiR4fCXpeTeuXux+WM278Qey2Ae97JV74c/gEOIF8dp4VCI5pB1LLmTBxK/Ta3i
QF5QmhWuUwe19BK4ExQuOkAzHEVavYdN3ddHeO4tjFaeGt6zTaKU/J/nH9bKLIaxEncW2OjS9Gbv
Cenx43FSFyUAY31OXCYa0nnI4sHhXt+b0KOBiADH8c4DgC3whJkYR7MNUqo9LpjSvx5IBGEBROfV
AX1s2d1PFUAFSd7NglH7y5UYqXWrY8yeJkC1Ml2/o7dch3qhsKhdcrjGn5somtB/DzElqisFE3Ox
ZJq2gFsYOsJK7saEfjt/FtFW45/vbSwsBXHlcgzgnJ+AMqXxR6pUdv1zo4ierK9wvyMq8hxTf9+y
kfDMIL0Oyz4CXLxm3xTiGS/yHSg+iSyJ6GFLl2QYoVVuXXi26ZXTlgAg4qJssnj0ZuVIjcA7C9LO
GlDHWEgVJ785bPfvPKRUbKOngK0injC2Cl1SB9H7oDBKHpRneli9Kl69C4r99CXOxyPXw5YEFHyI
zTf/NiXzvyoi4gKvoaCKxwjX+sQ2QfWV/wkFKY6pIZzrh/Ey7MENOgNLa9CT0Vapzb227bG1JcXa
n1uyMgafbwXd1EczSydrq4YUVTHRbynjWbl3BM/7nnX/NV3vTcGu/cousuTH5O/ETHyBCWEK22Ez
gdlKMj8M/nizlMns6YBoKvpQcf5He/bBRi+hcjoQZhMpjCVcqep4d5lUl9SeawtJnanFUS3FtPGg
vMuF7hgqxrzLpOwpCOAny8c2awcIrigSu+MzC7vZntThWyJ1sPg9hMrny9MHeoCil6fgCyiPJ/bF
hDf7uqZVCWC5KNhxl7kizjyMMmk5/f1S3t7Q6eu2YyHNwJ/O8FdPWa+P7IvBTWSDQCxNS6BjrO7d
LqkQ0XRWCTuLMwMWLCOJn1+Ma8H9JIs9Ng9nPYR0AZm5bV5Ud8TsDvZGAHaRydhfb1bX575xvBRC
/KfV5DCn4sCVNaZXmbNQRTLUYSKGIfi7Bj/VCEGg2MguZMBGQE1erZyxfFMU9pdN6igE7tRCUa7C
N1EfzO3RIJbmqA1Xp/kQrmdKPAgP/TNxWfo5QwuFPCUx0dsxbhxRUEw3zTkXXK3yraLPdWYC6f3U
BOVdclCKdIeFiH/5NRnETXOSuv+16mvD9RHqV1yk+H6EyqORHClAdmQ/jKf+TfSmSxGi3VDoPAzS
5LGbWnB3ZHqxi/CuEt4+7r2Ya7Z65lEbEyxQp7iyVo3Ysbc1PO8YdxP8JgE1WDB+cRAkI4HrPYw2
hjJpHR1bIiQfcpi/+i/DODrMWh+sff6KUdMDB/BP5rxL5KIzIvFZs48RDwbudKCXhoSptyfsUHiH
G4dsGY34O/IIb7NOPLMAkSoyilz4RzcegBUfbhntI/ET8U2+xnmKbU2IDUBhhsOrUaosfPErm040
u9D0FcZ0GTgjzsHGLMpFvj1iIwB/24nozEQ84yxAMn8NcK1hGytBQ1gSquJoZy6UE3QqsMlVpIYd
U+7wEDOPJuDxrY5IZWfAapGCfWI8cFFSyxYlFyqvxQwa+nVM8ZnCLdGsBNv+6gSP5xqTVIOKS6tA
EcvB3OHr2PvPIenya0HwLbslHqShF7afcmz2vixJGVzCArqtHDwjmctHebZfZsth3BcEsi2njXw/
DPiZz0NxhDWj8vY5M3csQY9G2FnlIl8XSSeVEICcTLcXYAlSw3gE5SoD2q4jefs0ugTg9VWgCRcT
MN8ijjJGY8Ys9qousUEPh1BpUgaMgjMcwLiqS1X1J3gV9kfEKpMLlaRi1ZTKk7pI4ABy7XtEW7P0
LuGW/7U8j8c8KNacd2+XUIUt46t7bLI9WKvj0Xb9p8aa7SuWqcbPTgZR/MXceduEU3euLk6vfQXK
jMOWEQHR5f/IcXBVOKmkHpcZc741UqxX/+OcTrG+A/JsWuPFewSxoQTI2rAPF5OTtSA4l+9vG7h5
TuW722qpDGOkGrT1OogTlsoSwZl7Jx8ZnWNvvvNySjh1oOneH+R7vPkjNr0ChurOmw8uiricoFcA
ZJGPoA78P7ANhwTonmzydFqTOKh27K1ENjTuqSVM66dg1KX3oYGPlh7qVYi5Q4K+daEYWOHWcnBV
E2YVnSxDXBdlnPRipsmpirkCp6JqECl79kF4pSbkGM6YxdbOI0yI7twpvrlRdAJr1Rq90lDYW69T
67PqKD/+WuNgYp0tPF+KHqgTuMLh4AgHSqtQ1R6DJ/pfXh+e13Ju6ZzexnViPVeT9pfwkzrGRo24
u9jGzqjZmEIhfejpz34pqYQ7uVUTZ6VQDYJqps0mGI5yqbP823C3gNjdPHLZ8aClrVHQ+KUa+x79
yqspUyVksvxAQwFdEN4ft9UmWdp4fyzgy4W5pYxGuPpew2e3pyGpR1TbEJKnAA29qaR8gSj5HU8p
mAfn4si26Fuf0BESDRk38MI1d7H6p7rofAwwX2qA8e2hlHNP1g1dOHHY8rVHSbmXX2oHdc8dxaGO
9L9uMlzWK4+hrtw8kSr7K7LYkKntnK5mXP4YSBi6QpaongmFetP89T0m7SZFERfHZ52x/B30iLbd
CXtUt1sW+fuQyI/mw10NwyHAXl4Ws8puaHeoVAralXQXKqqOyx8/hG3VfnOeZiLvGpBxO4K+dL1x
3zGcEMvuXekLrMT8HsmjdD5WSAt6kdEOVOnSVhPoQMAesv5W3PglLjp14YNj537Xt0+W6l8x/8yp
ftKohz3f4tkzG0X5zC+iNrH3arjzNGm1zfNVe9sm2Xus3pp5wXJt2g4jka4nipXnCDyf6dHuY/4P
nntcoBwXecYGUaVdl1WO0h8KhnreB+4qHntNZPVSp2KMTFkSMiYGum2VjxA/jGlFbGXy4/DA/0An
famOs8kbu4czz3qVhgK8LRLihG7p6v8ZnUHNdHC1XlKsVIuw25oDKZyYfxsMM3r4wQ/mH7/39t5p
N6TEgNeqbhz7TMyycwb2KcpQ2hkwKTLpHkABrevYm8AO4cYDZsh//XiZz/NeVHbJ1RbfSeiWmBso
IfqY0TTagbnts0iWaZhtRnYyzOzv4vTFuH3KvyXNzMQMeXPtVWflCyafJ7RLuR7m3qQNCg5mN+Ys
ePm5oZdTeIHx/BZXlUMXIX6k8BT861Ke7VMlbQGwgEf4VdSK5f0p9kLSntlEQlgwBHDdlFEPJp5U
YfCV6OYncfW7NQDtc05pwDw5R2qIvhUAmE706WNtp1CS1XyeACsoGDNv7u3SVmlJqh/pvHU6bL0V
t9D+SwJcAyDijhzoRrMi2l3dN+73fiS0gq+/BTL3ygbLYaqppSBlfXB4mYwZMXRZVXmSfMCeBJVv
iaMTEMdYVz6lpjCA6tBU97LJ6Cw/1Vr6GyiFRAcwyc07u+JMs/npjbIu61zhz6B8gViqEHmgpyl+
NNhM8wTchKUX8SqvB8I2DncWy1kWg9cIdCeM701n9dA55KNqwS3f0HWYACTXIxIH1tPPNt+aEQrd
vrdL6LdtC7X7aKDlErMVAHRdA+TZORoEpYQPs2Nz//pBhvBUcxZNoq7QPunM6RafP+WVAyVVCRjz
JFGQU9UrTaDBEYAv4/Sa7J6iyhRcbmguxpQ67IlyT3TYCOmTzOlMVvn66indpgIui6peRQBDT53G
SWFm4iX4e/q3jAsKtvby/r2Uq2g2QlHQT9weVMnkiNdx4HSZGY+VhAD/DL9wnFJmh+xg8vUznZFG
SQBSULYBdzwhvb/0VZvRHbtG4b9b5EzUcjp5O53FG9P3LVgHQ3h3yJBNK9H7ib34GMA7uv5XgEjC
FrsH6/ySNVPTNvIYR9LwpxlYfmprvB2tMmSUfEkxDSBdYP+tL6AJImM90OJgoScMkfZqJI/1FQ+r
SJj8oEoriHBaz+vB3G8okrXEnmOmraDREIuczw/w44Q6TGb5CNYEqW0c0TuU3e0mvYCqns6LJRRU
T1A9AnQm7pz+hPSZ8v2z7rBbj5vIq0UrCCUXRmVg3Bz/ebCorOANF5DJSekrf0CdJ9wMfjCm03ko
/tEfteoj5ggyaqmMOxvJBUZwpiPvNj76xhG/unXoLyYb23HQlwh6IDnd2io0trAngG+bTCDh070z
L1QWGtN6h+AVUfx63qkmEx2cfhdUCPxy2FE/pS0bW9pZffaan1i6SIUMX7wfN8DmwGAs6tE68n/x
oY056Gz2RQjcml5HCSu2XiSAohMz47IrMFiIbsOjOcfWtMzIcwuR9iWebjq5JiOG7s+v8mwUkkju
jUdGT3rF+Rg9OgalFHz05WhJXdUDonQoK86fH7qO0gTRdnN3ebwh/TbWxMzVqoqjNGDl1NzySMb1
37xXDrghFFb9i2PmEwMxnihQXK2xDEG5W3fzyQ+qCut8M9ZXdt3+sKTzOphXIpdMpKPErqbsKvMs
FsCCqWcR27ZGeh8t9wCUBelSDZTlaTcJldbKDzkpTg4IJ9j4Zq3+piO66AcKqchaW0ZrhvNhb+Zh
IgEtXFyEyetStz8VkBeG9FSjthMhEvtqZAUrtC6mqXn9LOnATOz93Yccmy/DgvC1dQnsP7b+OL4v
ojEVkyufSVhoP7qNVORo3H3IiZ0L+CN6sz+iXfCDnWL3+uZRkLDq2TWPjIWZ0ATQhIRmy5Yqkl33
jItG3zhKrHj/VHP7Swh/8251SeH1Z94j3WTAUYYnac6Ebyx7np7FQ7DgRAIgvsbfxREh7olFOSKx
asQza0kluj/ViJqY8o7N9W9fNNll4nEKy/KJnxHsV3syrtsKSgwGH3J3fARVUZGWCcgluO0hvqeY
yZLIPNdtN6eea4Xj/avX1T45amMFkiJvuber7E91miUxCjeNTJy5jrvvMB+KShhxmeOM8yXVL10O
CTRupHE2SESBV2IYvtn75nAPrynYxE4BsdP5pw9sXdmeW/4Gq7v3x3qjUEVH4cKiguWkp6gjukj+
KXD/YLze0ZlqCDGYsFaQiH+U85q6i6q3SJoh+rUP7nQLzseFQMIUiQ2cVdTdePhOx2e+28tityKL
rcwFGnDyWMMuhnvcqLgCnob+kMldy4Z7iRaLDVRai9tZk162Yj74P0USUGJGDqydvVjNfqfQYXCr
FXpGgoi/zGFJbmWIDY8hxhDKmvs/rNWUFlUtyY4iMe4sMmsj/c5sugcXdYytC+CvjEhtPHkZc0QQ
mpUqyCBT56BfFFpEVSMxOnnprPGAxC1CboWUFBvwRIdlBvc+ZJ8Gnsg0rz3N3+dHqWC7Az276Q50
7cfdKsrNZk4ZDxU/H2fKCiW0+3crZfsXmRpv/2w+S5wPpUgrqAYXrasbAY9G8/co5hb0YYBwLh15
0a2s4D71ICmoq488JWkvDmnjaUvZmSqfRt+69oMoBh24+NhcG/9WDkWnulwVAtje824vXGO/0EAg
SIZBbC+12K3Eey0I/1fr2SgfAkEgAiGCJYyEc9gFwEh5irfM2dxVF2+U7pxGZbrXyio6IPobg0RB
7nby4L8IB8kjqylj9q3evP2vyRGl9kFIY3rt6tIoEoORZXoqd9UoCV+cfMHChK94c2TozyTVCEMG
tPGMke8VUnsMQGn3HLd1z3I08XWSZoEzxJqlDdlzuymS50vt+9EVyIS78RvbzO4rmJ+cLGLmqK8m
PUf2NpjQgM0EjBjnpi7BeBjU7z08nJ1fVdvZvTc9OrCfqH6cWUTVgsMGdFd0B2ueCjN/hV2i8RAJ
M3JNnGGhMuHdu5iJI9a0jyHVgJnxz8rrIDRhJB3vIJDZsxC+e7KBpYXibSOa0U+f7WaqUfnzcwqk
XOQ/YCyUa+iyf0H53vQ1w48ZxnC9sPQvtZDkUhzzwcD7iJAfBUreg2COGEZ+7CSHoEXJZSe7vpNi
EUaOaG/uC2MvoFgtB7wQIuvLQUYp7DT4z30tDLQ922AOqJ3svK9A/FAXMaWOI1SMUKHMotbdXdNt
0R26xp/UAsfPTqGAkv02AKlDGGsXMtATCV7mGJmlCzBpDmfQ2dMJT+uVv/gyBBv6Bme2+sDOZYZJ
ZXuZPBkNZ/nEFW1/vBXbD7IA3byEPVKWzM5Bzzf/lh9m2wufujQJVWRjl5w+zP6J4C7g5UznvZE0
ErmUyWiMqkw+hzMRBeYLWagcBlfiiqRa+klrGY40qgx0SG5us9lecZjGemqM7O/nG/lsbwAE1zCP
B05k6xpEUqmZxOO0TpLZR4ZdZKWJKKbDrYIQhVVqksPFzRQ90wwxpwE4fsvaZyBsomunQhMENHow
oCZHURDHJaQbQK5UQpv08kra0K1zqDazkbs7YKjgLVNrucHFq8J8gwPsTt/rBWclB3Lmr3rhcdjG
0k02C+tLqHxZPph/9sBgHQwZD7IZ/Xmt2HRXGBIX2K7Ubi16y0/zRWGAdIMPUiLsLIIAmfrivbvT
AroA5yq9YzRbQlIVvsuDn1ksqxr4oeRPD/dChUhxiX7P9H5sJA6nLV9G/C1Uep4ZknmXBmM0W+QJ
YQVqnHGhrgYwsO6ltOZ+JQ3sBwoSTKKuCTb0dsoVlnYNWW5zWNNwfmXDkXJym8KkFvBBBILt9974
gN7VoEWXPXx1ZG2vw5s+NEfgKqqD/gJWuG3FOMM8MQAjdf9ToBibg9WIF86pGhxRWPxqcJogMSZH
ZYK10PZ9As4YPmAGpiHgBcL9JBbG91UhHWp2ioivi7kR5CxaTUrdGtVOr4v5nlyTnEJ6Urk1WBp+
PchrcEs61eJFSPH98O8i+BDqqOWMqU4wYwUDrS9nJ2a/N55mpjrsuzuFasNqUzPs4XB8julluU5K
yk4xHUNqXIwdhB0/hJBuhWeZ70FTDBRZssf228f3LSjHrjJg5RxIx66b9TO7zwtcHcQh6B34zVqi
zqGf7yeFrR06q67Rgp9jzeKGUDv1XQAWEHSBFcqS+TP//YuOYv7ZPldAVqSYKM/yzyOXCCjx9LcD
en3DJhA3MgQyv4zEGsrS+dvTlTB3xzf3WzR5WaUJsN0p7vcRtG4vk7ks8ZhJLwuocv26A6OkDqcA
KPMWw2xFDOOzSPm9fB5Fy5v7qY3IV2kZZuiTXnZdnllhDB4AWdcVQWFqSP/PyK9l7xC7K6JnWVLH
9DCBgcyHMiLDPvcm0etjj1ckx7grYhjWUc2O2Ek30rkc463kJkmoK2J7KaajwQ6xdbZj7McRn6H5
G9PvFhnEqvH8nHF9H/a32PHxKfSzZCuje0pc/twHveNnyfUx2aRBV35WMslyBwoUUVvA25J7fTRF
+HoPWbig1hWS3Ajwg3YX8va1AXWLW7ydMAnGos1blANN+Z+YmyKcMrddbA9cIceUJq7A+5/+gQVe
1EISHhgNgQeAJqZy6Yni1hLHJRqR23TfR74IpMa5xWOLiRl1OEqJVIAy0q55o0vtswad6x2kGsvu
TrutnJsqUh8VoNCoRwi0OuVPoYsbQ3ExZoR+1QH3E1IrQLnqG26EEPqLua+wP+hQdvEKiEEqsFPT
USZFscg01wwJef5I2GordRlMZGxoGUbgrSBJcLG6Xoz6vmiodFOHDzM3egL+q1klNZeuEd4YKnkI
v2RGb8lRz69NdZIVLv/UvaRnqpVlz9XOt/a/V2IHEOIZ4wpig8WvaWJ6n0ybYaNb1r5Iat14fQRB
ICL+27u4Vt3JrhmLw/Icoda7FNTvju/kNvBn9qfLjbDy7M3bes2YEPUrP9qhDohDPBjdxO6UpuI5
TzW2r5axG9XPXEbpRpwkb1yfSPaFhMwv0M83hS2fgYjm5nDjSdt50NK9PVwmoy0JmZJjfp4Wx2+w
hTeO8hxL+vGdRv3GBq0NVxVCgAgyFv5J0eACSlsLU/Dj8ppm8NxavrqJPWKd+b7J51dPVUpH/N71
NhAjkKOdebNvHT1xaQwgWJnLoI7Fm9clz6fS8uvA1A155q2wnUvhdDlGJouB+R+wn7c3e1GHlzd2
NOQblER8iRU3epmfhOkHwL+XhTqB97Q/Yr72qGA/dXQ3sqD9od2lP75jcoDO+zWZaYW5cENPR4/E
ELErRBxTSYI9aO6ilg2DG86WQOCDr7tMJXed8BCiA/YxEn2hCxB3jh3n5ZTszTAL9lERLuCmK1Fn
fzsE2GVU0yB1g29UbkQG+YO7nYDIXbNUzDOqblZf66EckMDcssojhJwvCXobImgMjX+VnglkVhpD
g9FGQu9oM7ODoft8a32mYRRzVQXfO09+71FjOM07Shoy0Ppt7gSzMXCm3bcam2fIlkGVn9L0PT+m
+RdU/14e68iJmKMDWCXnyOgNTv50ZxQhg2XKaHrc89QLUj16zw/1HSjtxZyGFkb3wqyMceD4S+GJ
UJRYQSIuR5s5gSBGiLspbDjULPJrIYUzkCM1bisAsgla18v/q6sgt3T7EWvHhAG7xhW3Z+1EFFsd
m2mkdBPBJnDu3pb0Czo8DtKfakY2//IIdEhITlPIYkRgLefN7mIk4uigEKHnb255tYidZOr0Dw34
WZBbK0bmDpUYqA8NjYR6Vk5GHT8bmMRoqHexuzHsjbdabpTlTSY5+fPk2jZpevGDrTFZteQ+ow6m
X+q6HErVu2KC+skLKIkGZJY1+JLkq9lCnp9RyQuvg4FNIk97nMdTpXY2xYfHk+VfS8lmPNGWFXyT
IGpE1lMSbePEWa7X/y8Tn/cAi9s+M32fL/OY+pl6TFRJibw66xoccBzDIqNCLTnGgw1fZ8fV01/W
8yDHp8Ag4Sd9NeGctDH3IrFYAIYpi/NYY5lRyy8ibZvR9YTxT5iG05BCyij19vsOSrp0aaX8G8rI
BfJkZqxJOTgKtNYhU0FBCJ4TCFUWSnzRmg2z4W+bDQCf1vhEFm1mj4VFycw2/z4fVcs1euGRbpNS
uOoujMrEQWARIpj2SEjpe/Kdk/J9aocx9/m73AZDlrl/eABYyIcI2cxcNtFqWLKMw3D3zQ1xo8s8
PbAUV+qwlJ4c0SL7fsfN/v1ZXXeNkEXS8yaWw4MM/QVn/axUz3Am6oYsU9neHSFCi53m5ypPIMeO
Biwmfy6zNnKwBGjE46658EbV5EwGZ0sJuyvP6UmLixSJNej70lhEWLRu/mdY2ijz/8mlP8AWe1Ig
hZQnKBVIgg+ZAdCMHVYwbAvBkgxMBFG8mlJQGhu1t/4kYHgtMdwSZwVXhiqicxAS6GukI5cj/XYX
3pswabhJUgpOlKmqDUC+xX1b0KfSC0TMyYsIu+EQDrXFrrIcjqm8Rt4qmYNvLkpAQwu4RsK0viX3
A6hHruTvEt8Xvm2hKLcIrLvoVvdWFUtw+ADevrqZMIY2BanixsBd3hLejhiO1GA7s+RknOg7UZ2U
Fw5ZScCl6ogEqtwYERHVtD6sfkBI2QGVaY5Z13PlPhK+jhPfzYGpn6va5xYWzNXenIZneKE+/TU2
CQeHuEZldSHR7ipDPa1oK5meskLP37XA+uAexQGeeMrBZfW0UQwNN2E+Sj+GFECULK/olLAJS62j
iqO6bZCslhYznp7hJMuCjY8jGKcLW/tqwLUbyqUCYdPFybKrz61XyURuaQg2gAGsYy1ob97F4jPN
OJy+W7ycqAGGn5HmvGG62/T+JxwcOy6a/rhgbWwD6gRRhkV7jX4NHFiYUdOalc14jMCVOTzRr4wa
W01nLuCncLmLuM0lPYI7krjmbBiAgZPWtjcAthU6N3PaEyWC1TirSjj7JiqEx5vzD6jiq+nfQtMY
CLdIwzDf2e4YvrQDJpN+pcEEONPmLIgyn+soLpJzVqu04hgfiWW2sRE8JIVQL3NC0LimH4cUxYUW
+ZmaWqlB+FSu1KWwdT0E5ScG/Hsrbn96CsJnGCYNri+hFM9/+W/6nObgRCxm8EB+iEUCNWlZnqtY
e79XDBb0G/ihUB4H9JWnrKrCXi69JXFgU9wIwsVk6C3ULUIot3CHompQbchQf+IqWLPXydzq0oWP
33wbDP8MN7kUxEIxGuEzC92XfdXmtrdcpaAtNLlVJXSgYykJq2jFLCXVWD8H3j9pH+67HbHn728o
n6RLyV+smE49O1oVESCPxxaxN9CJiJQ2WiKQGM6zrkBiV/O16l3qdJgylTwmw6wyaFSD9pmRFmIt
Xe67nER9Xn3zTsIJtR7xy2gp2ETxpaRRgWCBEwW+Ffa0J84oN4eN/wb1qQTHaBocvSr8OGYsR8ui
EBj2Li+gHbcwlqor8W/077LLFxaGzM8oMWA/WyTCVmCi6EDUs4ygPeLq+Muo5vthYGaSZH02KqXi
PXNLldYQeVhvyYdFIvvIMmtXcfNmsN3UIlQpQ2FdARZidjByMYeHizN0161lBLHkHjEu1xn3ZZmX
bmnp9zscps+eXVWdeEmk1LqT2SstD3ynXIJKuYEgTdsgglHOpWH36VdDMv8rgOb2KKks87OYyA2x
XHYBMqny0bzrDur9t6FGBHb9i/tWjWSsezrmz3j9Awy3jWlsfG1vlN42oOq1gQUwwpITKfQdM4/7
WEHVnI6rtLAVhfkvx/UZANNi+IyG9hFKU1lnVajXXJCIBvoCj9xI3V96cqWQL0T+ZepZqFdJDI+X
e12ekfjBLvRnDMybJ4AQmuFPnAk/9DLRL1fq56zJfJd3lkPhehKRVuBW26NoNn1AkQzlwGOCSptz
XrCtHKVvvU4bC53t8Z6zX++SjWiuIYpJ5f6De4kAc8QWNGr6IavkEQBH0mz+qRBVCAEJDWHg3JjG
lo3ltGc7LrLWnTqY+zdkGdxxuSbhVPP82sI0DudxguU4B2R/KoEnxSw3/raOtUKDAAdgacOmm4JS
d2CfA1K5q9JXCvZpoqCWpHoVJS0t79Wl7r7RLRKZ/OV/TJBBLtCKqCQslH1tM8pOuMaGntRoNxSX
LvwjiNEXpouSKS0ksyOm58PzXY8eU74TEPYwJiwc08I1yC8eInGwBTX0h+x03cyYPwr8HiowHElM
j9Wsdt3wsB4x//CGeTF10iiZf0LX1wXbG7m6emkcmOVqwoMWoRq0ZqlN72G7aYzOa2cTEivereku
fx29y70f1w/UaH2Jp0k21Y3g3DkubuzUyW39DB+8YmQ/PPlt50C+pSvOTM2alBBQHQr/onDErhm2
B73SFIghjUWc/4SLb+jNpMqqYXRnA1BPMUpEh8A8izzBMRHXF03KgXMj9kPFoYZrGwTFnVbpCkR4
XPGisV0wN7wgPOIIv5SuuQ6RRJw9bMmYlAlovsM7L83Ljx30JhV6lIKsXsQ/jQPh0DEwZrLnEpV0
FvbDGIGem1I2wxhmc2pqjECBPGaq9ylNQrXbjslTPvi0a/WYEbHL0JKjc4zgT3NnwGexzyxUrVyv
ZddC8HU+x3Q4CyG0eStDwUK61eOk3Sx36Z7Focvxb6FJ7YkVwtJjf873rmUe58uKvIvB5NGg78WU
qBdyeU+zl3E8g2X3tE/FwTLYXr1y7m1JcysSVEOQjB41QRgCYuzVF+Rg3h8nkwIjzUz7MXZhtO+o
uft/dwE2YeWlYXapfeAYaIQHzRt/cSzDykjSgOhWDyHlB1fG00NpoeX9SvBmb6fa3qYQMTq91aAb
gYT2x9lOXYJsUxw0pGCsPtRNWcm/v15d6btzdkFCLeaBoj4/yM/RCEyrwmHhGPKjxZGNgUVkndjo
c03GV854g8Y11fRsJRiGRB2FN6iNIkGpzU9Q9gTFriZnTLkMYVqPzDfkyQ5YIf301jEi//Wh1cRm
bsxbHMi2dpMt0C5VZffBx6k3FRQh929u0icDQgjEcwsrkb04gc7KK16A6gCv8lnq6cGFFjXyeicy
2Hm703DxCsGSQuwJOs3CbUg8lJSbX9kD+l6BxLlHRfE6vUO65awlWDaBeqmHldTRdcKtrxw9XeAf
jS1a1dZTa89YYbRrWHFAyrgGZE4ZfHytsOZ+GOPZZBEplQefupg/bX6z8zOUqKN5xFpnEurxMZ6F
lDLUTaXy3VVwGRvOs/yDOsFuaN8b5R4gdwK9G3l5IfNpvnVmevtqRYrldpMRaPiQS/odk4MUX9mB
h3opR9qoZUZbp+CMCx8WBVUSucleEZgIXafUuWeoQMFZBq4r/tET+3QujcXIV/MGhUFsG+2PPbBC
6XRwRUACPqiF3eqjfAc+urL5jbpgyFOPLqQiUvgqRgNl1MT/bvbLiQLxe8pw6x2V751BB49uCL5U
qavgMCQueHObvkB9FV2FAM6eIi4hV19bueu05UYDkUp9/mzBYZiq+u21utFG9b59UkJ9UQbe71lC
qbTvO8iFUXqlVR8b7LEvFkB2PR+J9/prE+GfR8d2PbzlGTMhmmdIIZyHSqLCE5tl7tMYu6u398vm
BCO4B+ds3QAjyudzbTC0qvrwA6IVwzaSHdGnm3Pn5KJEiHpMY42etxU1Zjf6qwA7xTz4AQikDc7+
ErlEwoyINXVhpFeKA/y+xg5eO3fA26ZmPUv1ABTMb1pLPjMaCghJHdhmdvLlC4wU3kVmlR4F9IHN
12cSiPYvV+ZGE0d8aGIhxg0n2AAef5LsaC3FB1nqXCcTTlgktqMdDx2cKhBifoUZ7jl4idyhkbzo
Ao7XbVSmzAa5EaKyzu221Ko/iyZLbthtVXyUq9VzWiUFhg59TcPL8Z6mPv5490kzeKkf0RLNTYYb
AWKBQzTevjBia7cPV7FxP79wAfNCqrJJaFAoESDGOMcKcyT8oJFPNdsG+TTx3MBIha9OIjZ70Mu+
U5Loh/pa+CQCIof/t8F4R+4DNAi5TI6Tmf9EX9RxTTWckoKhu97v2rMR/PsMzdQQlKvsE0SMDxDD
UVkqtRvMXAdSrKgSZl7YMCcJt2PJX+8bLnFQf3fd9Ing5ej0wec6qOQ20shnmrVJUVdipGB+xb8B
5V8vE/KoEPBA1L463aXiaKa397jO9v43OdyS4zkgHsGga3x4GokStuM4v/QIMMPE3YWvMpaN8yzO
hf+8W78UOcJK+3AfZkMOy2EHHPj7s2I3o8ePlWYBhBYaJ1pVABpOPTHbcmqUgGieA4Jvaq0a9sPr
sboFVSxsL2Rv1MW65TLUXgYJiOzZiWE8m5Ara3eDdsRV61ie5TTDdNNC9IIcOP/xUYickY0GXZe0
p+WyCBPOm9r3YNMShmuu03bmTjDhnrLMYlSFUSgnzRaHErE3ks5ivbjqBDU5Y3LZYyyFKSMxtdQz
PrwfVubXFUx2T2tmO2w7Bi5Tle9vBkNDDrGidImx0JqzrgZBfm/jpaA8vfsHH9Au785df1MM48uK
KDxaSpCeAEy6WBEhbemmjYy9UZFWhAbID9vEI6BdiT6597i3KxbNpOC631x5YmQdP/cbDQ5cGYFq
c30gAViuj/TjgI0XILahvmF0wW35ThFrSfjm7aD+GXHNc6hJ11Jzt+WSAKviYiJoECASW2g3z6a2
5NcnrMq6HvOq7Hlm5HAvEw7xTFjuXOurMP4qvupu9056bqVDral8MSp9NtyWQHZvRwa5fg70MJsB
GYLxlrSf6h+I209HbmEfDF+bVhpK9ipNifE2TNQJsiXsh4qaPppiH+4nh74lY17EE4ntc05mKoYX
Og2W23slV5iXNVx6UcDFMnPaYYxk9yoK5rfPJMVwojzorsSpuCTBgBOcdTen5QLC5uomwACDXUTH
wgP0NFS9q+9Oh6L0n+U4Y7QjnYKUaCjOxI4F8IWL6Tjy+ovOtRHuutX9H3x++02j/ZcY9t3saxVb
w8oYRgpJIOqyBOUzNAIcjl92DQ2ikW8FWF5joX8J33xzEUOS4ZIU+NQEMHR1EVhIlv/bDW31b0Dp
PJi5i0AXlE25lFYgsbOxcBjx0E/1UA+n1UIm26qy3eKNKtcG1FarfMrabVW+wnYJfb+MXqpBE+bc
WQI/AZWaQoDV0rq7PhF7Z7LJnyQBOtvouD2YrZLGaAwxtXrNmivrLq4eMDlssJgxe1SMKHNs+uVW
N0ycEqcGFffF5FdlG7Rs7hl9YZT2STJUqdRoUE1DIdyqwMNkLi4dJoQtjNcTRE7RhpgMIjsr58fc
7PREd9j/7c950UwVmd5ug2XVzQaVfKNJ5HCHGHA9gXsKrfbiQQSPei8v0dSKNuYJ0NH6x1HHUFG9
iEdiSRJ0AJRUdUMnt6I5obsQ9IsR9+PNnTpcObhYxW6ahfYyug7WAC5yUr1rmmQsQSsB11QlX5kY
F2y5J3ld4nMHM0Hv+HcbxFNgWydMjHc+9Rp3ONJXDrudz90csGJ6PK095l3NZxeG1cDVRIt2EyuW
ycoxLDvFXRL2r1Pnso7HRtokZO1BLUED8FIHzaDIKTmWhfCF0/zXq2TyS7lDbb4CbJhDfOarx0gK
daoHoo2qKpxHs/YaRvEFTNzQu4szgaoFPRGxv0IsF4ABIIVq4Z0VgpQeO4qyaiTv+LbIscOa1iSq
JsqT6kiyZri7vX2jCprgyp//pBVzJPBiUTp1lwUGVxReKDQR6wrm3SIn5yOUgIl9sPg3J7X5C8mq
vyQFWRVT7NMDaguLWqLCNuxxhjR9TY4m/cJXI2DTGLsL6yIZK4fXCYO+EHTgzcDBffJPo51mPQO5
7UDlR68bk/znBV9mC2U+E2wTYzuGuek79peEfxXWR/57ijC9e7CjnRVhmy4G+/nt7E7HZhrFmz7p
8K9Y/wLMy9M6L04zcqRW2OR1mYFt7h/pe5o8ut+JPHnGa6Ig44UmAvQb19hqgMA8WW5qWxep+GH1
gJy7BPgLPKcIgAkJzPG8HStlKVLwA4+820PaDYaUr3DXUT/NiUlINJi1444sihgszncJxbYGdjZx
G3pXGIGvQQVbXl5wU8TDssJ+NTfMGS29u2HMH4c12KXxSiz/nAvIffkRnv9U+d4o18njYYNEdFqC
3/Wq6pRuwTxtenVAtoTiWj1tlN8qvXOLhjRMSphH8gk7vlwl4XXOFm+6FAwxvv6xxQzQ9c7a6Uom
9X2lrfY20jyCa81vugSh64b4YV9LRGPAdibEogkLB3Bm3ll01VO5PG+wbyUAIeFRbFpkwn6sEjM+
llwEVXRHh0t2BeMxoW4ybSGLgriZdO/eB03RikGNX+O6c/OauSVKdnYGPF3oqxiKaMOTNdm9LhLF
o0lDMuCeANubqgUjQxcgnq+hYIOeCNcVj1ip4WoRt0MYH2jbUlng0aH9yr5uREPruP446a1mfPRc
XY/+S8KrZASoT73Um3whdFWFld8ttmeJwSueahHM0pt3i3BM+NGxOWrGowX5ZtUKnOU5zHxQc/nO
/0wm271LbxfwJ8yDVznG/tSU0KV6Ip6oC/T1wn20e7xmM/R/8+GPk7BJvejFe9jvhs7ZLsF4S5mx
fXCHfq244jsBHu+tQTTfXlmZz/+z+ZvYGaVgnqrm3dIoW+ekluO1AAvi+mSQ3xqtcZWPMsuX7yhb
eF85YRdvCxhbe3yhoHORKrZ2lyRlsoOyT5M9iGxOWF47kEMWWYZG6fO9bCCHeVV82aWoAZ5V+3Ng
EBOwFpXO1/MMFTRAWRfCrTuyed9I3youYo/TdY3qHLvObELnZLsy+3vevXG0WFbxZ9FYkZWzGvU0
eMHL/xNFFsQ1OyJxqmg7os5k3ub49NlEa5T849tBUicfn2yyd3dWhP+qIBak4GQNr6LAOBJumvJa
tZsiiwYDCmIaQQEzh3Ph8znMIVZUfF6xFlOKzbyvza1OBlzxORxm6SutG+sy/SYlBzsq8gGsRO4N
I7BZs/MMmrLGc3owbBgUhuXhDkCShrLwBvpacOLQvGaO5UQzNAeTMZwq7gx4ph/jchlaV/TpAer7
U2alJ3hjTy5P52PzgFF4Z2NsFRvaTAon01uPATe+dkh/HrLoX2uI3OkPxbdre17vWIe5QfjyXD+k
Vtaoie6KMHZNO1u3yR4i06ulBRtpinQyb2vtgyKOJ2lb97opxH6YUaw6iFVeDcoWj8hnZWPrYFRP
bK1vdDe7FHhmz2CJRXxR+gN4I53SPzIseWxA3Xm4hE89tlzuT8tIyqIceV6cQ76Q0UdjVaqEoZxV
1PPLgQP30QoqdzUoxz3RCb1lM1s26KQp2HxryIkTdXFCzOSGsmG53Hj9PfmKmuBZRuNWOd/nbvdH
DLOEgdx0p6UYC86pDcm5WQfHMphayv3bNk5oJrwOzfEFvwYf4mpWGfYEW5hg1Ko2AxntxGtjefAH
eKu2IRhahUI2SlG7v46ZL9JjNdJo6u1pxMPiEKC3kkWvmuJ7VTDBHmiseITCuYVUf1RiK1Z9cP4e
NBaJueCbXU6kdN2222M46XZDY0UMVfM/g8xa5+YFOsdQEOKjStRq6NZ3ZKqhOVsqrztIOo+dte9J
y6OQlMfx9enDK6GhcpAX4XibOLzUSnZMAsL3jCkdflXB2sU+vTphfaaqQa7UHtMQJCkTo7mexETo
DyMYT9TEiEhuG8NcBdPS9z6Q0Hy9kHvqBxO2IfvmWyQMBR1Xvbl+uV/SGVEee/QLlo6zjL1FQOfg
kjPar/4ZIDeOm4Y7hhHXRbS8V6SvfiXyL7X9PMv74QN/1xis7zBizsUMocg4IyCc1We7DVRD9Ynp
SiqIAlGRv9jQfQz1FNiwXd6mo/8djjoDQhw+zTgvjuIgxCWbX3zky9b8M0OLBd2f0DyqyiLlNQHG
4EnFBiAFKZp/bxib1/58ikHH4cngTJtPjap/EmWwJ1G5dGdFyFSjaaP8HJNEFQfUw7Q2p3RfsEUX
r+gHNmLsn29bG2aTyo7GM2BDVzW0YNfGeEButnyvsl9g+N8yMzE1pm6ji6f2Y5bObdQFNseY9vDN
CE7+CAApgoVUoDny8wkMSxvt0gGeTjgE6j/8vX1idM57ACB6+jV/VuPXoQBU6xjIyHsJ6N5QdAdm
RMJQScfiVK9sB4kkKEXFNImJ6ak2LCdezTl02wO3/NqlesJijDhWlzX7AqEpYYxynsREUHvJIyDZ
uDsgZEBQyW+MBhxQlc6Tg8l8Bc19jRDZuT0qeLNBgjPZHO3wRB6NTFekK0fSBxE0+BQmpDqijwbe
xScxP5CgHynBq/BN76BgIrB10DtG+a5dUF0henemq++kfx5Z+wvSnP+lyB+0uhKoH1X/3SsrdpH3
48xNEVyHNTlupFyh6kbOkUd3OP5kaYBJUqmDW7r52U4doLoogRopaOzULZ4hPHb0IxWAZIdfJAz2
vgCZkx5IrP/oavq/y3AdY8XE+Rpf7sQ1QZe3G49nTnZrZhqTrQ+6I4K92e9rt9iD+OcsaS4zRPRs
OmCP0P70m5qCcz/0rMwvClGTKNHPj0/5KjMOLKPUbHSyWIdKUWE1KvPl1ROlRB4KO9mRN0KO/dzN
+IToSA4sa+hLdkWEoNS/NDzsGzvheoYRuQu+cevLGOM7/s/5WzZm4ycVy8r19FXHV2QY1u71rPSx
tdVHJE5Fg87r4KOewwmOSNrR+5ouXUcqAv+dWAxQwGneE3isfciNebosFOxeE+osp2K5vjR91cQS
jfyR36ENDuQusrQ0uePZj/MtjbqcFobvrAU5Tb8ESZyeCQlCEMLiWSTqOtuFXoE48UvJDAl1++3p
kinNH56HHZ3YlVLgpsfqcHDGGzP7CfBMmGk2aI437DeiP5MHzeAkv6cB466LIEs550OEozy8JTip
P+IqpQyJ4oqHXjsYO0CMHJ+KjBzcwlm50e/n1kZjgK5MwysCRkauwGrqpdPB9Iaz9lERLPDfloOh
PIrakZmh+aJDXL8W1VoWuBQbqhSkDQjueeRmZgFXVz+HgDcMlKCd2xzZyX5jWlzBEn9oOsxseZpo
9NCFIPCWli+lF3cxjBAdzl4cIR6DcfOHMFIsdZmeSyNGTyyg4R2ImlpznKQxHySWd8X8fDQZcmmG
RYeBV4uKncsZfTJRdnAAtFujwkNPlhTCRNxRrFQvQavvV5poaM9d+1lasZTfxzFRy4emdHvArr6+
ZliF9L6m+JiV2p1nrzaNI7lCeazYT0+X0Ds1lVukvAE95NWfwVRXRzxohjmPmaxgE7iAslTBxxEk
eIUVszH+iY4LwoeXX82xvk0FqAGuQDsCtcHI2QabaZHJMl1SIUeh/RP5A2Mqc1wJYhW4JSwdkDeb
mx987A5IzWfOwuSCS1wGwTQag6axHOyjf5TNOccUrLt0YILSs835BHwYJRQeJgCvbXgKYzhbUvSO
xc4JhyF975gDsnliDORDH6qtmcTQfbbKy60IdIxkiiXDf8UbF/hEebh0ZSGv7QLQxNN1jnglEN62
YPpaRjGRvZWWqIShjQrwWTkePx4KgM3fpvzplr1Jm5oQ9p8Y06goyRdkYF3iPOBdfS7rx4VSGEpy
Edug+XeXy7zVSglWzVVAq7rNi9vndq5OXFagh4lLbidWYIraK7n9qwWcHW9LOf9z8M/axhSItsgO
YkzgJHlklyiGa+xNNN4xGKCaBt5q/n0xQdJRqlVh+aIpHYKqCKxy16aQJlQAYhLZ7brnHwEB0/tt
zsGEdDb7tiT9L93yCo76V7FENgWQxyr1MRDLIMr+Et7CEs03EnwIsPuYaWtcXydFHYuxOI1rZpjo
IDZYkAluE9eqlowLWKIVrKqNVXVLtYK0TbwZOfd81h6DDsAnHRktFK3mkrht8jV1+rurqmXynC6P
vQo2BDDi3AqdIlmTxogGOtcz6YTNh12RoB1CFdjK4qwUD1nMNIk6i+0l26czywlDIhuwN29X86XC
L2DvqE15sNOeOZDmnGFWTcKWvxTSf5Dq1FQYe3XivPnvm2s9m/yePriRyf6nJFGbeVdgxu92XZ94
Ex6h8Jn3Pncx+mY1Hsg3mFreAwWNopVwttQk7vN7RZHu1YwNqktRvgn+BbUAG6mxnb+9uDaKtR1Y
mbPt6yxsXbRFPqwqH7sBl8hlMfAbwiMmBJNjKD0Am+3iqTtZUrT7qegKM4gNnzS89azpuxTtkEdo
ahViBluftyJDqlmuV3lQ1Mcu8ePcH2ZDbwnZKf94hRpEzhv8qnlqVW0EtfWIVaPpSUudulCgUxWe
vS1J50rYCFJ2WltTQ10gEL17+jT30VPOfG/YmjY+Zy0eft6Klg3V0EjmhMV4NTLYKDz/EH9vqT4p
eukc9E5wJZAS8h9Qdo0WuiaOoIndS1qrCJQSXe2OkfDpVBoExB2H0yZhqAfbVcEWFxsz/q0Lff8d
8uREhyywFLAUhJsV8QS9Q5uYykvrv+ZyVcNJvxXAHw5nrMWXFp3Kan8ZUqnzVgi8L+wc2/NZSFSs
NOMrXg2+Q0NoMFC1Nw9YZTPbTDCPO0Yul5kIpgEhAdKJl/XzCCX93Ca/Kj6HROKvt91YR3bFAgZZ
/bMj3hbRYiIj/H/wdf+NwArCQhd42dtoLybPt9bqMhLsTuo4FtOYaqfuhGg67ZO9dAqgbTtzoTUK
GAB5ey3YP9GSyo/o/0X7tMMY5SThj6DM4p/+dNGLabFr6VYpMFWQUEIZ8Yclfg0+smaeAzRNoyuK
q+G3ScZfXiSxhchuJPhk3OCp0sp4PPHrU0560Yrc8rPK8KAS+NkMkP85FP0sTN4+iHLQ8GdGyNy1
LFpoyVS4DRFcgtWQTPLAlnJiEU24GC9MKGi5EsnhFAUj6YRFUAii4UItcHt2YW4yFsCB5Fwr3sWK
LNVGNcQ0RuZwa8Bz7BsALVdiuC3p1YV6V73T29iMT0h8PeQCaMT038SrMi3/RSso4HLv4hT853FB
H0oJLl+23BN3kWWevg+Of6AKSqeE01203up7o7dVOA0IJmH74PiRRerUVLnW25Zh1RLQ+iKZC6Xz
GoUVzYvMZpFWlixviCfAxF5s/QekJN6sja36hsoy1/Vvzwewa/Mn25ZbiF3gyaXXduxJyq4SoaBb
4s9WX/dtBCRRWmtd0VTFEPAw2+7bd2Kaxvk7mg93CEAZIrjyP7oDXnzBNjsq77DKJPUZOWdZqLUz
LckjFEwl1A1Ee72ODQQ4htpgwagVYN40MOLGK9zQcrzF1KPDPWa59uYsCYOKQSfvR3aSFHGwT3pc
d40fEDJEISnxF9wr5niTUJbKhA7yZf9OCh4xAGTZoe47uihVNF8Aasz4vBMkeKW9QFZQn7dSRtsx
If7ngZBaRLPE1deMD2hyqzl7WIBV8wXSDuyqEVDUKFlV2KRLdyoyty7pJxQUAmVaz5PmK0t3rNv5
YjJ4o8337/z9zYO7dV9eWO5NOxjjXavVQUGJQ7lsu8BYvt+EQ6SWCkM3oXBWTO8gnzwjfFmx83O5
aztbr8X0Wyhu5pFRnWfRjxGVvhaM3jrOeM0W0XLYIgyITUzhcSMgrGw09f92QnEqt7osGJkIPpOi
A/7PQ5fuUOOtShopEoGjU/WDGhFeixzhzbhBgD5ysGZFiaoTAVVQdqRaBXzJPRTm5Sd3onbTtaio
AqdGHZmuOOrMeNIRerL6h28iKrBgJEa9dyoln4EY+ZXKLHoHa8C8/LS28Nehw78zYH7GJFVvlBh/
Y/B057LN0/f2o21EhPaLm+I3yl+IV5QZsFZT8owlJz2p/fiH7dfVndNlXyIyPa2ERUkymCEwNuAU
SUn33NJkNL/faLHmwlO/ZoFk68KhIm1a8fcMDXC9e0pLLlOsRAjgOYn+W/dtOwjPjU//8V9pSg7W
hT7+7EW2wgDjIrZEYZzlZOnlUAaq2ZSIeOFJkMk5+2IDD0LPGGizmcVWbhYuTOVtHgmf/aIRZwqj
6RzYHx5PBWwstIC1Q5KxuX/KRBU37rCrPM9jNvqzzXYpGj9+YtOMxE1JaXjQNNxn+jVCt9mxB2Em
Qs8nDN2IRQaVmBr/cSp6lze2ojGbZtWGfQJDAaPuASDtsWg+tWGDkjqMmrjxeIeIKF1fF3EEZ86V
rVHy8fxBKMprjr8UBqb3WSI5TTdVa0QQg/XQ/Y48AzkFTE5JiK9sA3p6lWlij2wsI1gcjhJ1inXT
qlMxAZ/PZbkj58zFK7GNrYHEBOwQFxCzIOb7pCAbngI4gPEGQcHsdeyv8wccaSxbxNVfoxaYbGww
Oup9oSH3wJAmdngp8PM5yDrfktEjbyzk2M+en+oS4Vnp6T0y+iVNV88HVIEN5Jkh6egkPUOCjPuS
Fg5cHpvVQi586PeuI5GbS76GfKHkIuKpYmIYUJFy0s7YE/LmSYiP4oRjFYk1hB/SvGRjX56iwf37
h4g4Vi7Gz89IKpJFMZlhevRG8mOi18xwonHkClQ5k0vzaEmZpsMOg0SU8tpq+mwIPEyNrUsf4Is7
Mf0j/KPXkxO44amNhfxDX/TYFn7r8bziQTm2NG4nQtQh0pkQsRtbqRI97UWmlGAKI09+b1s8rVd4
CI79/Xfld6uiAn74V/Gkc2p8t/0aTS0ZEDvpmODH8AJLm/yzcTttn7bp9Lc195vHJkaNaebtSs+S
Gp9ya57+Aeb5oHMS8g6HzrEcQzoCKhXB1iqf8T6rKPTK/JhNB1uwEFRCrww8Xgaw5OabO7xnuI9r
aq9fkRoQOEtYOebLw3nYmfS2qYQVwM/LIYnysP/eEH4ClNmqKqUj7WQdz6zY2v6pg9Ds5rIemwRt
ugb4ee9ngj1HTU06sOOe53Oqw2b9kuqRWYt86wRGozdzN5CxQlTge0CM2PQYQZi+0Jgptmc7BkX5
XINlacIvu519D0LcXWoOgvQYTo/oZCgZ0gsdixCRhw5F6UcN0cIoK/9c14i/1UgugtXiGyhPnvxv
6erwZzT8thFxSGUE/vbfaUBrVOryETCm9mITNHXyPAyZxIaQ8rTtYjf5IZEMIaVzieFdGQb4UY27
9vvCDKMNwngqCYN8tLETJN00kNp9mwmntHltd/yC4Bp1lMbmii9QKDJsNTc8gAXVAxPboMxiluVF
atZYpOyBdCVgMLKnigLatvh+SYmpVZ2b4nz8YBGo+eOPoQGZgIh1wqd9UdhvekHyDqGMMx6dPQQ4
mcVIy+B2HLzyp0pDrxgzqdzCQfrQ4MT80RQMw3Ped4uI0sA/CzMzp7Bl2L6u/zryxM4JyDqZKOH6
Juml6pAMfK2bGza7j7UC+/MhYMEOTp3cLp0n1jgWTu+Cq2S+hgkIJzvAfBx/1rN0ix5wAfcbLQGV
1W5T+uFYEEOdZ9Jxeq5BW7k7o9ZGxM1FsJ/lcLMtdDNVFu1EYASip+384tGs4yT31A2wJLOvsk4u
s3/ccmoFngdbRCoQQD3dFLfgrFRums2ZsqUkduz9hW814NC4TTsJ3JAIGVqOHfcVQPZDLXUIWJao
+JLSWwdOttMu7d7v15wHIYZYP/Wm0Jth/K2s6gkJj52pwbuAdf8umiNRxhbZ7lZqhgIlSrIDZQea
Gjaum8VffDNv84q04aI8teZytFLufmNuKCNrXyHidZwDIvfouO1sfYRQDkPuMdNEXWmtvPxCQQCX
kec3l/8BtXgHsfUr6vt19lv/kdj8OA/OJ3/9ltN6oC8MpVU5fpdCpSgEXA17Fcszp1pxx1NHwsBq
VK3eSMYps8t8qvPua+tmJ5L8RienAt514F5YGivxs7sB1VRIZVFTGl7vLxl0ICkfVdPyHE5eWYzl
URyGg8+t2u8KqrzpgKK8wBHbpixZvVOWjh5zIjeSoOq50FP/wB30HHCpYwWeW67FK1f1MnfcBLFV
VlAiSZS0B7a4fexUiHKv9iaiBKFe41op+5R1oMNkeIiC0J0m8XP5FBnm9lMhga9Qv+yhmUXh5nfv
FC1Ns5X74SHq+9/OTS9cIkfNpUwKOVIQ2c6jHAQaOomdM41VySl1CC5JQGhel03nCrqanmrxCrLJ
no9eNE2WOGDZ4ue5VhcjpiT6R+En2Kjc+nRHLDa5pJOHO4akLgYslh+dn7JVas02aOUIn64Uig6D
rOmAqGgplnz4xNbh6qSIKgLqlFxmVBQEYOD8RG+MjrdncUn8QUmTho14Hvh3QqhRy7OvvHU6iqxb
6Fse8lFivoEq0zZuxfnEEDiwbaz/DW4BZskXsBwqSTW//myD1G/AeOmK6jGUH96/ozqoGGtWMlRE
R1Q+5KsjKOVM1SspdYqvLqKuDnML/EDJlP9OhHwMQvBjlsYU/OdjCsonILIEYkB4V+SPnjUs44Ss
ZhZiqY3echZykJSSk+AVOvM/1+63mHrK2lSqUeME8nmSzymr/4tMpOz1j/7MpkyGFYZdoAwclj4u
9C8OEs3i6hRY5S7xY4S0bA7QAVTEceGK01lOk+bahIogqZduS3NeZPUyqdCeeLwdSHVGR5YAR3kv
Cme5YVLsFhCWdSW4qUo3FfG3i4hvzUgTDrOJDgovJaRjKS7hjeKwzaIbBzrxKZuXjzrxUkQW4/4l
uV9IpvqxROfcKuElU6cw71T+3UPywzOpX316wo5FhbHXU73YBDWo+JGBjnoF2v06TS7eC4grWFv6
XHoUKtIILwpkYwcOetXnO/vag0TPznr31C0snkCvOJDD8f0kervzFeQPlrKFvYR6luA0CZmnHpPf
qyDGhVzwut1xxFSWKoid7aip9JKaiSiIsi+aBzVBn46QLuKKGdUTHTa/RCCf8MasOYYVtDcqo0Nt
SgqwUDZB/Z5oRe5U2b+Kx8EYynx8DKIcjZXDafjahIFOF6uD7wC/w6MmydXrA1VB2n4GgEv+DEx1
0Zdw/S4cQXo4oWdn4W813vgt9s3lugBX0SfbxtgurEXEfEotLQLmdKBO788IfKSO+NX/PDVoY6xU
F/lJh3eQ7tarSYEm2gUOd7jmjM1IDZ+cpbYH+qKm9HpAUtyMS6C58bBgaEfA3v2JvGpYPob58C4v
8Niy040ltusdUSyqNZHXyMCih3d+LKfj+i4pDBqkzVSLS9j3DmjLC94AUa5vMRGs47aAwTL0kplc
Pf0SEZNHsKnhktRRtFN8Eb1kFDKdfMGx7BVasKizrvuA9qeJF4fNSyEeGiek4x4+ub76ICbVL+x0
i3ha3b3hxJv08CV8AJVOQpCusmUtGW0WJ3fqzi09/qakumhlKstpO2spQbkbhzM4JdyMxRl8LCEJ
y4cFtBCRonRuG7QI0JPBRJbkSSr8V2hDO01oBh1IDwgKu2XHknCk9x0Ml4LpguXoLsVVwWel8/ir
c95fYNuoMhi/PHQhn9QMTk5QJkipTV7cNJa5lHoptvrRrvHvRKHflr+hcT0quD3sfVlqJBthroAN
tt5pwNK5zh3DlAW8/dyOnRgZ8FQCU4p5N7K70uxabWcO9okqz5z4g9px4r7+DQ0ODO+l8ToSnrFu
Ot5nPNfUyufH9Uym/d/LE/Ah/gRelLKMj3aOFLS4wOPuAunnQaL6pIzNQnpZiJ7wfDaysA7nDLaH
6B3yxqfNvSJ66xlo0pscgcZJwA9Tsy5Xg7taJZPSRbllYvNqZjLqiKddslhyEvB77MbGd6QkQ75W
uSCknNJ8TzGNtrecYpF0Fri9KdirQcIcXs+kCk7TaL8fsErv+Vw2n15uNATeWaqysifgqkoNH8qE
Nuoh67p4qESDC36rJ0VQub+cLZS8pNKhhRTK0wwiUqQALvMm2Rj5xcpgYDTIw49uKOtnesoBEGK8
abnzCNiOhC/VNIJfyo2ogULaISXHSBTMY1Ey/eEHcM1+YWEI3Ys4Lr++GWUtMh5eZxa5XCMgZexX
XF4XUYGyhKPnQjp6R45Quxh/gPe8oeH65LUfigkVczIOb7a04vLYCbjuXpDiCaih4G0+dnRJMwqY
uDhv/ynhV7M/+0Qrtq3ejAIMLLqg5iPxxF5n56T1+csVUSETF09KqWua6LPV73fOHgxRfRPgbKIP
eRUbC9qTY636IWexMaRmZYyq4rFOX2hpUlvsWn5+s7zYARcwYYgBw4/bH0pcqMLYo9Ch1Gi6H/WY
1RsL5guQHK8YOuQiJRIkyxXoD84j7yK+C0fzBj4fp4YMkeIU1GsFigzk+YqLvPVe1iwWbTcVICpf
IF/bKDKqS+F6KjytVvBleXD7l4Fuz9OmEBup2lKcSUzO7SaPPiXt59e2PFcBx+RukiSaUn89oLOG
qfDVRLXB8QQDQ9Sj31upEG3iPDQ8+pMKirc7VKSUP0FXHT6vxF0DqM8UIhZm9oP4g0//yY4cykSZ
58di1S/BKQIpDTfPsWAfd2y5lUwbmkGmCtFEJZeXEcS9DIEV02lZFqL+5xP1zXnf4+aDzS7nxbkM
LWF4/nTmT2p9kmH4D2xUWTRIeqKRDA6J0b8+q5ggx77hx9HMtVKSm2KnOok6hPnoD7iy0zn1nKAP
Z0DjU1fzqw01UZIYPoDAKbWlMHO1e1H+t0tfQ0DsQX4qxDlTxkbLCMuvLDo9WWXV1BmcrV35IDcA
ScslnGJSycKBWGk62+CDAJ9LBEUxDPKzmqHPSwqusmFmyxZJDSqaO8eOWo7pOVPQ94vqrOV3LdqS
cMrVwtDAO7VLnK3hRDQLd3uDtmwgWccmoh5AAGImDrDsUMffS2SofoEzwwBpwtdfCtn8/wdmTAd1
CxpAmKGPGR5G/Dr40fnZ1bDyWwv9tXhd4QoyVJm8L7AoMnaxzc56lJ5l+80qG6qKf2Ll+Y6+lkeg
ntpNDIo+uCURStb3K8Y3Urjw9FyxOypH5VQgFuz9fv4LdkAFfMopzz/bB8t8H8rbSFi3BKVI377w
lNOUBmikIhXwuV21ahSXncTKYQbDHjzUh/sRZB70fVNr+zq7a0GrR5howCVwPeK4bjnqs+Fjz60v
J2EUOAp9xLDxAwxzHuZh5PD4+bHkqFkYiurAVIbGNokOe2hZ3OcLQwhGBrWKHPrpdQQWPRnp6Y/f
yI1pIV62uyT1YaSvMLDikDGgG9VTKNZA70fPIeDT4C2XoNxFkQRgc84UHdUTWSZ36izE0XMt3m29
BX1ILm2bJdNdBbxT8J9a4Jq10dACELGeR8sPeifS+WLI4HqxhGj2DB1cI6XBKR+nvCdZMVUcUK6e
mfOrkJgxrC1HG88f1C2Ghkb05UwntCg7OACGzrt5EOhRV44Xw0BGb8bB4M/JkZR1zDjE13fM/bWF
CooDU03Klp8P2gLCxczcSETw6GjiNES0lQw34UH1t5Voh44P+UJNPlFUwvE/cmrO6+o9yt+2ECE6
oPsLa1RhlnabegY1SfLVGoGscXvu6t5duzzDuLZbMS0rRnTxoQOFWaY5yJyGyC9FXT6KhS9ehNKq
MwIsAAze/E4E8NZSPkD45X2sgnb9rCXa5KMih+h48kJIq9rQIIvWsCno7h0Lkhims5sM9Tr0hh7J
fx3W5IHT1xL78Wc2aSHJxVSUHCEI14t8yQvCFTnB6yYj3hwR2zfVsp+SqG3iugI+jnpVGCdpjXIB
4W5V5xi0c6laUg7ppvAJk/6OTcyM3FQim8f3QDoDBFfcJ4JFZErj99ORSPnKEDMrmsSJcO2XOieH
nfzidu1LCnYRXHT/2QRzvOhtRtGUGMLjRmH3tdcvmWllFcAwJQdUszpHVNnZU+0AEWnISF9Dk7ff
92ZV7Vb6sJw0KkQCUHEpPWwHbYAPU6LD/QzDAxZCNTAbNW7im/ufjZLAtp2J6gwAA/Q59AXrwSlp
4f6rst8p6QZHWx9PGo410Lz+BrGUQr8GlDetX1iRwxfKhWo89BrS1ckzUsC/w8BPs3kz4Dtnx4kA
gJCXf35jERQD8Xzn/ihal1Hpv9hQtoaoFT0uRhVRbRJ3EZiYDPGeJ9DWQ1dGHFn3BT2l2Q0m3DfQ
YgcnhMU27nR/WLklMlZ0IUWlclo2yHV7Rg3tbufiPkgOEazJduN14HRbjT/6FbF2ZCap7aghev7t
9pzhfvRkCbGCjfyLa86dlpjYbYFQGblZRnlt6Cb8YiFwXKEvm4XFCNKiks5/iGDhUCSS7JE7/MRP
Uj1wA4yrbqgz3vWvCSgajgalgj4VDVEpq5yE9ziFGkzPGZWJBkejGihgqzc57dcMcJY+itdgbLCZ
BSiNVd5NFMgQBBzPSPU9Wrs5YXQfwiH/bPThz4AyZESLdsycZG59O0RxNgNdbEOPhgmcHmOx19Ar
zliVpTT4ltXEGvU7ONmFKJBH16Fjod3H1486l1iT/BIR+1Z2WEFfTz6qKmczLbCszNu37LwSYjbH
mS3GHdsMZWbZeEVH12BVd+q/yVVQIfx1QvQqj/pXSCLlJpFjbMWF+6Fwl5OnOLvLNdlglDwwF/MW
EXzzMDVhJXU5m6qrKW+WGgU+OH7/2s19OruOFAbsUWguc2fLszY2pgbB7zMj+2YqyVZM1l7keSmL
PyS+Xt4urx52IfECtfDal/lun7G4wEuICOJi9ideGHBNL0Upr5Jh0FcGuNR7XZQ1dde37rdQ9KcE
zlEZDk5KVEXdwJtrSlQ6xJLdMEPbS/p2No8OUiqsxBw4bC5AyZ3AMKnEvTGBe7CXxEmzVkISK1pp
A+Mk45Q8Beiok94YOq4AhKcBihpLQCrjaHiXdu8pZl7IGT2WZdFxLmkP5GRff7cZsTXgZMoAVn1f
QlHmy3QFLJXpR0qsSCi6PZFFxpkNXy2ph401hJjrqCiTSUSR93emG+55OAVY3Hle7+yH/pybp9EZ
N7TnrgoBe5n2X4E23TYw6GKRTZzT/+LOGFQS/gbhZ9ghxULhZF3+3nwn00QJxACIowd3dFCSV0H3
RxswrDUoJPdeCxhmAOBHuzzZa+vnWclFTo4bwHYE0nflxm8P9ew0Vi/cQL/Apz9QfEL12oNrpEsw
0nOQP/QajWGdn0R3/EaN8vqLxcJTELTdDBJVUsjqH1eE0Ux6EqpCObBlKmLMz21bdVWrAlmchHvK
Utt9bdmg92iGi1z7PqXIgDqHNnVoxoH0BTb/erMODZi0i3fbmoIJYf1ZBMBR5T8Bp4U3F7PkWiiL
PEJFj/4j5eyXA2RC0AZwxsQVacK7HNlLQ2AemSoDNvSaWLe4VAMSm//wnrHzBjofzrpLpTU8Bw+5
DpUOk+kJbsY5Lds7n/TNssTZzaDo1vHuyJ3pkWEgL5Q6SuMdS5eTzEf+Cc2Xw1lN/n9LJGEgduSE
nhNJzHKCkVFMHBGlmmGSxVYaUcOv8mtG1tn8/WFEz2Dje8CyMGLwDoZvNUf28ZsQLkxe1zmFvQRK
4TAefr4h6oB2hdTwDktQtX0iOgOAo8HSRlPVlLGJFd55kSbwrnxSucNweN0MFSfgc74bL6eWP5uX
LjMJRHsksK1gWx5h+DRPsPmxkqljA1T7iFIlTd9OwC1ypyDYF/QtLv18hx/1H8wJDD1hDNWUGKSX
YmAtnu8mP7eOemGUgqFgeBQv4HnCtGEXMjBKX/WXHWqscNbNEKtdTVyNE2+1as1VIklp28M8ViYB
SCNDSOCpP5N7w9AUgR78vU6OVQDcBm9WAWZrEj0jOQdt7HOKUig0Zh6aWmxsf+G07yYJMiS7gS3Z
RJrzuWGA13cqAK3T1b3lIi0ZI+vuTw7ORClhdZNZv3JlevNHIJUDP/nVLHomaVMmu3LUzo2NLlrV
NKhf70FbKigkGCjl7sCRec8h2KyQgaffZHqcdXTtFPNb0+q/ZxjZ1znKf5B4LJFIpw6in4oUA9ta
BaR4PGKsGQwU720zT3w+Q4D68XtXK/0NRFpam34HjdRePCsR0ySXK816tb/2Of/Vc20CMo2v9Ble
nv3y6V99OVgDDNmPoA/UF7uVjU88zu+sq88ihG75v2p7QqbI8d6fFvlrkpsaY/3Ix436m3NGEG/m
ZT9YsuZtpRwnn0A+2zg567M5qSBnwK+18tkwn+JbzPTEURfbkQW9BK1PHq/28mJ6gAU49Abgng5q
aOkj+iJY5piUT3WuqfkHB7uZqBXXIJnOhuvNjN22sATSk4FB4MiG1sZdneMVZZtrVPNoPyTuegR3
EgzgR0uD2+C/KX2tJ2CNYQDL0F6NUDuJEJzm/XfTeEhCfa+6LWP0s0NZaqwEy/zsKaSgXLtmNALd
q6etULJNbq13QtYE0HFHX6D7wJ+ajLOH38BowqLNHHPyoTmmOXeD6v4oGOj5GeoY/QeJaEUdSfvO
Te9ciosfk4XWffWvhmHeSHF8qi6jjm1CHy5bsOu8KEZSf/XI2EwksPxoNaARw991wYML1gBEgFNp
n9j/f2pPXQ+koCpz+JpRotfKn/X5odU+ioNmn6krG2HGzhrxiucewiTOgoJr0dMEC3IcXdjOdnUV
Yepp3KF9u12CdC4++AVETnfA+VjHuqJo2WV3b60cmskR0T5ofg/hcmAIAMYoQkKc0yo07xnp036T
F017+AOM2YHTSiB1DL5SwmoRByX/wEte5co+ZAM9ep2pnfhj5LctI/Qde8Yjve7RnoegdEGcmWC+
qST5DFZYolPyb9FAgygJEpYu7JB7ZyxrmbVcuO5+1pdztYkGwYmZY6lpdW/i2juCHL7dP3LHEW4d
ZKB5qeN3GYc8fo0KTDpXnfSLaCWX3bwEx1MIcYgwlb9bYbC6mTGOYk2CjXTWimYQApz2mvOxfLLm
o6kRHjZQMzx8tRZ4f+WTaTHv8x0692YkR6gG8xYHJhfDqivWx446bAuocoYMaPEegEfPuzzRKDuU
twdJl6U5P+sM8uenZNEvn9LQhRJFjffr7rQ5kZT3jitm5RIXKxfaGxoUOSLvOJdud6Fr011bUQR6
pgDhWrCfSD4ZV0BIIl86oAmAz/QXXwHoD8BaGil6izbdqKCR02fGczTfEAaz2SjFlM6kAxSTMbGt
TMkiN5/bI9mYJK4b4yYgAE6M3eMvHhjEElbIhngDGr12guDt24Sc5hr2gbiMo3VzWlQgsRZ5YDaw
l5yq5crX0SkX34BPmysZkPJfi118l9d29Kg6zE84b56nOYG5zj0yEuAT+vZRfEQ4iuLcO1tvCPCp
y6NGfTTZtnj+fydfifEBj9wy0x4L9ZscqqC9ByYFIUWcucGNQlEghsDXyQ1JgmoNL27ioOZ8RryD
MAvvV4txc3NUniiCof40qzqLKUIleE9G6gMIXHv87wvsX1Z/9nCzBoPeuQgvDdjUjeQJdvj4d/Ba
ECV52GwDqAEeWxIOgvvhgLflE7ud7dnUDPPHLTg8HnjN6ERW4UN3NP8S5zeuNlRo7duHt18S4Br5
IPeucSLE+dyiaiEtGI1ky8EeGubeYr1cxz96Q76dkF7TefK0pqshzG2D0vO9aYYrmDay8HPQkdHE
pdevFG/DyCkHOAUwhAHd8n8aQ8zTewKZchcYe0GquZN+CIHNcudnGXYjX0bvvpzOIb+YZ4631TKQ
pWyBEeFrBK4/Zj4ME+9QBDxA3OwRZ59M3/f06rMJb/0sL4MG+UKqxhA40ptYzdyyTyo6H9r+nhry
HevRvQZ4nZdOTOEXa7S3rGE8CMiCuSKh2BDmZ9yXPUX/eKdxiIzsfRCjaq0AhU1YoqcfjH7EcTgg
5k2EnnBemHR/h8uQ2ZRwA/QYzYdEN6oJwr8EysTttq26AHNnCKCMgP0IbwDr+OTibZ8WhGn/65vN
mMIRCIsvHvnLEbaW59eNJhTwDG/qcCG5hN6rX3mqYGEsxjKi3eTpZWO3kTbB5UTPEl+3VU/Pr959
kMmf6TwfZP+BJhhoqLF1vkWJ4daVls0f7RJnTzRKQvHPEzPkgLrydiFSK6mMReZlNRuLDgIITk1f
IGVYlAOepDIwHt1N9bXZfja3yL/Q0o1+NXDMwJonaXDI0hSFuSNbZ9XopcAEcQnh8F2oHpsAyiTQ
/ayLixk8RtSuIQxiZ1p4AI0iK0Qr+nb0kBFWul9nezyocdPFay+dwUXKPF89SZU93cAIj8q09iPP
Rvf/PU00qIQdqQonyj4dy85qEhvT0NJe4kp3VDdvUJCV0aIPUkl2yPYq4cvp6380yJThcFOcNDMT
0E3u3PY5gwivPEhaKJcpASshOAXRJyeLVR0XU4GZsO867kVPj4yTneLldzLzOwuFIh9H9vn5i3FZ
ThpQsG3JCg0/LDKpN3pUAxfNujhqbFf6D4IbKjRKvAATrb0Q4I7nK03M++oxBLjpo0rwV3hCzZQO
ZnxgQdeztp3r7Bdz90LKETqrtSbKbXU9D0pm5oACUOfnC1hprcqgyKZiOqg9dVbExkb5Ieyq5+f4
vK2y7kW3fA3xbq7jCz/03g5Cs0pd9V4FAK9ihNK6yZYgt18uzrFjS3ZsIXA+Pf+44ef3VreNp6Yl
I0fkw65R6ILrF/ZKX8F4/BWj240NAACc5s5ghoHKKha0fkYuDmRLeg0+SKeSGAkCzIOSk8Uq75m0
D1chDdXOcafUPmmO512DkQwhplVOzZAHPx3ZfiOKQuvZo/+1zdW+7ekSXzCfUux4gvR6SRnHL/T3
B6kBW3mtbjMcC8SBDDZIZ0/r5H+vNrRoOyVpcDke7vzSKjZ2VcFlR8WXU8Hc0S1B/VRRasJme/gv
vcz7/NB3AdNDMNWu0YiHmHKvThMYQb+IDwjC+46R3SMpCRhTRTENVoY6nI3Jx1CU0e+JXW0FJ55+
yonXjYFCV8q9xJ3R2JVr/AjVCaw2vP5GX4bQEhb6rMmgAbaMKoJ0FyCFbnPQl+CnzkExtrt1Isb9
nE6MBSpUI/ZYj6lHlSdc0hOYN4TjqT1U03IJfbcVVbmyWQH255b3mhMnZDseRd9V0MJV80qMg/lY
vmFb6B9jLzQQXiktnpgyvs/ow8ErtanyjeNuUPWpytgZ573UVLE1eIFBnwhAE+dKQNkeGA8Eao9O
F+q6xOAQCvphKAuiJ4S6p6ZBIAsJlKsiggHLdLhiGn2+ytk1tm8zdIXNUI7Mf/jqO9XqE/+jrJAK
8V4FnOXmFkR0u62DV+rV/rjkGLtr//2k35RQJ0Pa9Fvd52J+j34ircmZJ3dVLljA664NkH381TvR
pDSw7X1NzzgxVVLB5nTfMTnVbUfsp/Lx/de53kORNr4dzNgqIDQFDZoH5mx8iA+WpiiPLcx+K9T8
WZNFOdpO+iT2gPOYvbaLklKMaj3qNJUPi6Nv2O66Yvgb3ora3hMru4uN1xJ3b0Bo24YxyOZUC7Pd
twd2d6QeGZsjhIabKXhSJYeFhUph/+b6ikbnLeeiptIGoRmJS6QNrn7jajD3YKTJIgiI6k0daQtE
uAmFrpXLq6I9YFX8UzwwlUrSLMJRD2I1PMgZEd4vJIFPYKPQ4kYX7P29rM/P2GpYsiUUzCZ4par7
QpOncr5rRIYiU7I+dijXQUY9FJaSjVx/cW3kajr48jcXLuP0CMLg/YsBmppmVWKIfbxfEBz5pxRd
CRbBOEEI3j8DcsO+aOo9z6bY/j6v7cvtIJHb2mtG7sF1TQyzgX+MhIc+Y7lGbWH3X6xGgdaGJLoW
Qfz4VQzkYUNY9ws0ezbb3rEyg9yitJhvlQZ7lUVrN+Gt96cqUUVte2YhoKURfEMjUF4TNT1rUG33
ppFATCkAiIsVIpF++hgz9NGM8qgdw5IQdmvb00qMrMmQx2hvy+BB4LTpj1ehT/XtWRXvoNzh9H4E
UtObUP+4mjqThVUpKMXPDdS1ewea925TxJc4fVBwJaAsbfPcSg3X/cGD+5rWouuWNNuayGf+nAzK
QnsqTWf+WeeeVWB62X7XPaCJrzlbbywlfMz2ouNP6gzrFAyfTlWivPbgt2O1yBqsfQh0Yibpv40l
IwygQJxc9cw8sSjMiKnRTYykwwFQGMF8gzewJ6P+UAUBYevBN4KP2ANZsyMT9Ly1Inf1JOK9Ljg4
ffc0P+y1iN2JTWiIoML75NU54A1VOMCvn0C+SNJH+XrJ7b5wCz2NUU8ybp0VCjroOih6EZyzcAxy
3pOTNHnJLKNR/rQnMwQWQ16mMGR+kic3zEgMK7BMZhLgS4eCiB7Sl5ZypdtmgnOgSy2CjBQXMsSA
OPn+EEVRCz+dSawXPy4t9cdSKqvf9CYpYsWG735zU7DgW2RmClaM7FU9NI96VxvlHf8aPLAWHtyT
EssyEi11DUnLcv2kmCJmdDOV3easDXUC8u3EwCCTpxhszKQDE4j7i4ukPnsSKWIKKOkEIZzFR2Jb
oZQ71vUl6Nvk5O3R0YZ1KD7aVe2Zt6St4XIa3Hf349FPh5UzaAH+xW5nTfWC55Mi3RTjTHcKzE03
Yzul4BZ0WfGUSukUMIi7MRDEEAJjcHQ3ELL+g/ohwAE74veyTTlLhV1Z8hjLNJhTb3el+vEstcek
90isMQdmQRSBoiNdqR+NARDXXtR4j60PZWOH2cteivebC2l/q6pXo0oS6CNXCXblDJVFDTrlaWFU
LZmP8uMiiSF0EWkk3qGl52CS8Iwv13yes/TEXYZs0l3YpGbMj6E/kWhUdRd6bcdqbzUoeXoYTCzd
0RnQ1hBxbspzKT94HWexy1v3np6H+R6JW8kTRdu+UmK0oLvO/8F9ZBAS9NMN6qoznIEHgUV3vVC8
+hz52lx1szMHZf6AljPIq+jENoFvQ2N7jb4w6xafABQ77hRn14OPFM89w8c3luYKrZeOlZg4h301
6Tm6p2Bi/gZEEVA/61PZAIQREvQ2zAoj5b2kpixI/vr7zp/nc3XtqPaUdHYEylsFhQvhdFyxaFxP
rO5sBOICO8xMPw1tQSQ7xIcNTgbBrFd5akI1Nio4CIMFAIV/XdEUUFwhdvJAJeIJJ+Fed8rxFTsB
HYyLejMLpaUb09shd8lmHumfshiEpUt9WGBxTOV6KX4Lg1JUQXfMyqqHjFAxspaCObK41QgQTmdw
BcV3esXZUIpUg6TYksZFBvUTykBlSosLMd6COGc7JEEoJWvF6hMtYcwjmZ4/RJNVMiOYYHgMXpUG
nh2LVilWzcOywoRH23XTvZlGSWd2jqElcYTFQpVTcOCkdK02WrUqbALlj7TKI/WSQ2KqNHNROGFo
5mUaNp1uqt0rnKdDHsEGc1BWnP+1TTw8D5BO4pG5z7cwkLmVuzJCX3UrXu656J/1oh617wZtAiLM
gU97vgELpOtq6KD6P1/lSPgQxLjlUcFlyQgMDi/bFXYmSyi8wWDx1Zzlsc4lh8rwSNa/n6PWmKkp
V6zbtSDQzFgol3ofWbO8AhOI/rIEVu0glAopMrF5IvdY4jOMNw3PBduXerJpk1tnjNbO5pQBmtqf
vx3m9vAzEaLN+iQN+blRryEkqHOFXelIzLTu0uwlU1+WUpTRrE1w305Up3S9ZrqdgjzV7EXfmhQR
lD1SCElZ9/SEGj/Te3AzJhbEXLWFNNEVGJzIxe/m737qPU611+YZIigFu5tHyFrb05ak4BIaKLCJ
33Xu09F3ryIqd2LDkAGGs7sGdZo0fUr4fCSAWmiYFcImMm/8W4ZRROKuSzapKcA7qZ0g6cOyZOUh
FqhOnAg6bZQIazPtXGvVggJFcM5YpU4ewU8fbcKs79IqVruGWWHgpou37Bm6Kw5Pv5eGXJ08VVK1
xF+qpFSKM7BCiELUKOLwk5xYsjRHYKOYPQI41fCn4U10iamKnxA7fmmsCvGoGREVhGiwrfmzyGNF
daIyfi6mIm3ENlGbblFMGYL1qjob2hqA7HF7E0r+9+oRNsHWctVKvG1pAg39mdQdDmhoQlkXahzg
SHMYpxLM/CKqyf3jJZedlEYzI1WYkyXfBamP0b3psyceFzQrekGJrLF3R6s4m4RLjk75WuWOkszX
jcIpdBi0w2MAUG1Y8m0ql1fKeOrS9khAkiKVnPxH6Pv67bCvtf+dVAc/Sz5CWcOe0fEGnYMzfJoR
UcQsSavd0IYYDGv6gkzEQS4J39ps8mVlfA7YIFnaO70eeiptRWKLkMhkgXXoant71peth5C2sXku
i0FNSKbUY5UrXie4SIgjI3d7Z6rlzjNz1iIuWgpdTmWP3XAjpTXh+3WOtdLkaUd91LbU4fU2+nCw
Cnc2MMHaeJSOlljmrGuXUhUVDAhKdrQhOTQFcHtf/jaq8Q8F5O3fbHDpkAuiAREgtaMQat5bJrAe
4YaKLx0WYrxj6SAriNwyD00IcCpXPCK5vVsBOUJSdui2vovtR7qJAwGamzaBePijywEM248Q564o
+TzHUSOiTtFLPs8srYmqDOFrAp3Y5qeoQW+0N37ycYRzmHjdgzdo/sKRFffzNEqwSWehdQbBHdDq
vhTZnzDxLovyalsLIUHC039Ovm5f8PMROzU7Kpd9PSJe1AnerhPFSoURMRjJnriE7T13ZZA0wHXG
fmlR4Q1ing/96KtvhZKnUUCdM6i8UtAne6UnUlRif9rqktzCHEn2fMldWrz9/2k8EmNm6bllNDVC
dijvYSs6ytVsHJ2357R7SQD3oZZ0gDl5tyJRzuNWlB+oZTi5e7BFqUhZvKcBf+hlSZlWzNoPyT+j
EvpnNChMlRuIgmlqpXZF/3snvs6kolRp/hhzz7qF8T8WJ1773C3LXzY8XzfQv0XfOJE2hBXUoKe/
KOqUpNOpJWuXZD7/XuEu/prbOVH3EV0e3dhg/juQ6soCu8Ggr1JbrGt8t1+w1R0IR0YhKGfrSgZ7
RbfGbnEE1mnsmeECdF7mvX7KX7t1anWLF4MOLUMHVUQoVW47RCf++s8PACV0U0l5Mtk4fBG+TTHq
L1z8E3AQqI+dUuCMNQg0y+GB1oEK1ZFV1axb5F58UyiNFYp6ydP55R+BQhKW3/gQO43orz6jmnEa
AaHYLd/Naxhtcy01vZF6n5CW/FkOtoGr6qtMNY1TZgjgeEOC1uHPxHoqEaWf+JK5kCKEo9Sf3Fx8
O/VUtHWQrX2koh//ONWddZXAYLxB1qE3ftYFYHeeUWuVwnrj3D5C0YoE3/jKVHaQBsb+WBoL6kXs
8hCf11WjuEWar9LBAZs9e2VPGj7LQ39YC073FDar/zy5ic/4umJo2hDD4borThmASm+3NySCt0y6
OT4ARkUhaAe6k4XoGsqsIpjdfsdBqXrLW4K2MMn8qlkbty95HkOQyr+/kEU26Kmdczbe+5QP8biR
jFBk+ohYGEcJ3VZrx1nfFEiHmsnMOAn36fkq2/PC23YLP9mAyAiaCNU+flsEr9+wV8B63ayPlcfi
N8qsuNswMKlLAQerNyBs7Tzg5k8dFDcRej3X+eY0dLmnsPLQ0H48m8WlqoJfwdNO1TTxvWHI1erZ
rgD/zpqXflHnsvC6f9htWWexYZe1TOdL6SKZkAA5liaqyHh/3uPjWGPCe8LGQzHStRkjZa5SVy6v
k6OeGN5RkZ3PiOC/8y/pkoIVyRg0XMUVfm5jAcRVuIROhC+LfjCstIEXd5c4FUgYuS6SSUx2Miuw
iVn7xBa6PW2KlTdgHt6HNM54LnAzPbE/1f/0P5JdG62fBjo5WZ/6v9D3HXBfhGdvAc/2snDy1mTO
1CEaRP6tgZQb876RYz0dzWRWrbgjvQJviJTvUdv7bTUx0xEHGW8OLWyVzedkk19MaYmB9tMV8R2U
z/zfUs5REaHREvpPkklI7Xf6XxwzO1ru95COG1c1uVzjM7ExEwr8GzA+yzZ188XBC54itlhjyzGi
9nWUWCrryiNJXjOcwZ3emkUFVI8mo+/jeZWBfXJqujwqz8D6WU/7IJt/o3eA1/XuICJL8oE/Gx0x
g+ljvWseoPmcpcwbgOQRo3GHNe06FtxU7/1liArRoUrOF3NJBEFZxXXEQ+ld5cU4eHMdGSLQN9Yo
1pRMc9Nk52KwQ1iKncS3yyhMXRt51bzAr1Y99wIl76jlgg+c4qI/S7Lf/8v3wAw9lgWWuPYjsQ/n
XYkflKoAcHFQA8OpyZplH0rJh3mFnKB1Crt+2DVQ4SXz5xZsNyZHNgmLpjIqW9SKnGn7zJjlnBQI
B1lXuB02qsl2lUJi3KTG4qS22/+MvM0J3Qd363VuhuYdludkPhofwW1UEKFYxA1PIWvufnXPz59E
5xgyYQRooxreId68w+xN1Z/gQ9+zz/AcxSd9NVDKTEpKbHQ6J34i0dDdjAC4dNoG5eQ0k9WkSM5B
uL9KOH1J6uDXP0j57yjm4bfAwl4D90yR3FHeJ5Ebm5rUmSNqedg9TnuqCy37pQqu4rCFdNNlaRkN
+dusdaRZINr2L9NZ/2b3Oxh90/DQ4MF5PKH0JDar0I+H6Uq/JS9uUsAuA66unPY/QYw+t9/nvg5S
zQtKTOXO8ltwIWVfR7Y4YQcVPntpXR/C/XfqMeNl0TfI5z4lc3Wp13imxDFHCtjwTBUJBqP5/a3s
lpCjznkCXs/ABBShXs3eMVg4EroiiLM79rwB9nb7lDkwaIkyFJPMKvAESebA/Lve1ZMfKvuVvRdZ
Bd6chYaFEXmww2fZSCT5eLRqLNSaItfV9JG9GYMtEJspeBwF60C4+OMjOSye4dRWrcuRoLl8Oqb/
/cLLFu8xAqJBShupus45qTworhFqdXhH0ZOT9cd1/bEB6xe1P8qpnt5895G/IJBWI2AsiBxJmE5j
5wTV9e3jWsd52bQJ6N62mujnZd8YFhaxT6/5wA9XaIV3Mo5rmYzie3+YCJgu9X8RLS1Vw9T8SR77
Leb78p7cUr9tYvrZQErfKUcnXYMhgGaJjldpPDXESzx57jndqVvxoBpVlu03ZdFfuowVhi6QXI00
4QyZBTHs1jOdOqdC9Brdfiz/o0NusFUQcSEA07R80IqgiygZwkQ1qPRHZ5vBju3F3obK3WGeT9XG
wA09pgZgVTACKM2DnIdh++KYAkqHdgnqlXszGb7qKbuwk/ZwqKAi12mjWlD+w/aN/b5NaVQkXru5
qB7TZc2dyw9uTeVcgigb6FHW3nTEm5Gb7be+nIjXqZZPFPk4fRjlpE5FPVratcuwr/h//K5//hZ6
3IHu5chunc5EVSfIMPr9QuDvoCWQeki6TBIKpcMeSY1Z/4b9jlAFaS/6jMp3hxRVsDfMozt1gltO
Vff0Cu7zepqxvwRIMxwEsq+VkIkaWqmQ71vU4hmL7hEKKd0ltHsXVijNmir3rdcXTVRwfKLrKir2
aRb2LLGZ9qX49X8h/dIjKGDIKMh1cuhTQH3ZaMd6XavVCktS3w7tvKUEpnFo3O1GZ7rA6VI3UN7M
tbXQcHfEP/YzV0SvbEqIJsRNs3yVop9CO1+y27EhLPTXDpeEAXz/4HAwbf0UCfETtZSDZDNfT0Df
iHgLRwfYuaJFFmIfZSqh1shanJV7QHirThP7VXh3vSBT4cK0KZQ8NpHeCdPCunn2jYrkeiOA7ScX
NaaGBEN5p/wLmpY/3R13jBDigbpAm2JrB3ufSW/3DAP4PPkaCxZ+0XJK8V0626DDD6nnPZiPeGRU
6n1ASkLqMXaRe2eGfE1+K5yikMduYgQ0rcz/ZqTc5JMG0qs46nao2SvxXdF1ES0mFLwrlsmGx5tq
wjyC53MWlgRdB1rh8uBF59cbqA/Mje6cc0oKpKB0vpfjN2CyrNVLT4aZyliV8CYta175aZP35uPR
ZBj8tCTTolWKdfuiS94NaN2LPN/A0y68XOzcDT0JOKCER5Tq/RJ4afEJieSWnC/XY8wOQ/xXiVRl
FbfDOYXb/Xm5AB5ibemOWGn2+y7We0Q3bdUk1LdfC6YtzBiP93i0EMeoQNp6uMuq81q19eGCHx1G
4oCkPVyj4IJIV6xTiZZxglfOW1Fngau2rkDeruwxFmJra9SV4Zkk+mzBwDm7J3oAdX+u+nowCvsO
e9FTb88vpx4u6sHo/74+KXk8M1QGgoygiWFk4uRHaHgE8mG1+/3ouJEvIH1jj770lh8Qqf6xjYpb
qV66TNEpYJ76XojB6LSuV7HtfJyJJh7fSYJbJ7YqK758V7sV7lpWvuCqRlYvMQu4o0aFJQvWCAea
zKg7eK2hWrI9XyCWB2RbveGPrBDy7Cn8cCGSYOODx07Okzs8HsiIngW9nyCzA3wzoATATas6tns4
Yn456YPu2oXqDBdTAjCmahdqgN5uoadI0IfQY8EZLGmUCoExS6/e2vCjiDJcChPbvmJH7cO8cAUt
Mzm4k5/y6pAQzJQaaYSZw+Qa8ogBtjXgOEA6w6wKfNF0cS0B0zKHq7B4y7fSntkX8y7IjjPc/x/m
iSgKyYrtLKsWPKQMnuPv8bWFHCm/b55UnY01MiCwDtx9bZK5xfdw93ZupJ6QkTu7mBQg80K+y2RW
6V6I1xx37KUxPil7JbG2/Uph7v/bMxZstc529KTC/OIGO59BKFRW16Zk1WH0tVSSWpwyV9SPVji1
ZZK14jZfb7hzcdWj/3QP823WLp0y034ybOeB2PeXOQcAHzhnZ/l+TQWaMHUCGaY+Wm8BSE+cafqw
64oq4Xb12Mtn5vLA/470vqz1HPn+YvB507wMXsea91OGqdvos4dt8f1xeqSzjRlB+OAh/k36bU3T
J4HyWQgFGDrGqtIc+xIGr5D2weysoOwlnl9A4XKfIYK3Fb4MFK9pgMr0X6QcMndYgkjGIu85IKcT
GbJpRI0aNIQ9D9F2+kONVhleRAhQ35EUW7T0icjDfS53/NeTLIu0z04oAzN7CFeLcLa2o9C75Ii/
OeChJoGNgZG9nhT+WaWa6sd2rN/LkMkk9Voo8vTeEpq9i+bGFKrcOP5OZo0RrjiRE9js0md3jlyx
yYB0Dk9vZvoRQyJn/2AwxEcWKRFxTt+OpqPsix2D/jKiyrlXQMv1hbG7lGaBA4p8UyK8QGyYkmtX
8cWp1G5252K59hS0AlQEMxSeawqlm81QbZVZUaDewmmuWSgGNTR6PVmNnxlkammd5Vu/TNjHXi3u
HEiKcs8LSBZ9IMCSrYVhJ90j+AwvXWhA92L1OhSiiy8NCeTh0jjpCHY8QzYEVl1T1EKkKDK1j39+
3IevVLlQ0GUQzUxp+0xOlKH4GfQ80P7IJ/rgCIz4KEhLs//tAiFz4Oy1v7fDbLxtd8vczKtaf5Ko
YLR0/FhawAqE6eitd6CwrHSuaeXXZZt5ygI6/12prOLJDeDs0pb/CI7ZeVHjBX0sVAsMaPzAizcu
6Qdm6+ssoxqkIfyjKeO+OVbue+2+ddoDrpSZah3mqWoMhoo8cflr7bjRmbKi09VdMtPi0e//TYoQ
oggdaJUmZ4CWqv/c55ptVjHdiWD/Lkus0xe675960X0hvpe5L11lySIad0447T1HWC6BbM7IHhYh
X3fR2r5FOuQexWejH6jJKW2ozOQyYyOMaN9l5F3qu1Lva+OZ2xu/yN0WuDQtusL/lRN6Iy/V+9Zl
k6UXYmggZz6CNOXSpk/pUbXYaW8ScNaA0iAkopm9I0es/54zkXVXx88nq8mkCJeOcVHU9eTUd4wO
+Z/XTDoDvN+5v5MmkQIZqf7za/VREaDc5XUY7mf9ppIzi/tdAQutkHL3PTdM64RGzd7owwR3S3gi
WGi2J/7UR9LJbu+s2g7hLTlEfJC8f/eEsBVP/myG71A9oCEpGUkJSMNaxP+Blwn8eQqfgnfmROmd
CC9sm6OLKc/lu1abNyY7Fs9R/LzyePR+nzvkaZ9z7gAPH9on4agu8Th19LQaW980volyjsGCu61n
dLJPC5xeNecKA1DtZ97IY5aPMUjokkIFpyn1X132U4iNG8EOcqSPq4SWgmenjPhx0/3kxJrQqB1F
x3P5x6DMZnbNbEHv0QT7ErhRWiGRru1bhZCDzmCmSlfcjqoqzcX59HpnxA8QmRKKS4ZzQLlhZx5b
2wO+TbEgAVbnHEb+KuSUKPY2Ke/InkicwFKmbcFJCuszxjFaL4gmq/Pz2OktRUxEfOUO1Dh2hNSe
+N7PpIJ07mAh212NciWx9vfjiL/K5MRA2MMkATXbL3GxEe+3/kas5T0TYolUNsUa/pw8oJyUc8zq
SwSxVpR6VlBcAmYIQ8qmDK0HtjqLRAzIs+Sr25o55kIbJQb3kZMAhhYQofHoUl4hkOnVfRL6Z5Fz
gZnKdnptK5Mh8EY04jZtQfuqe9Yp/VFfhzq/eaVuaio6ZRaRjRqrx3lRREcXAtDXBHOT5ZkWYNo+
BZmV1SRod+htTL9Ax9j4rq2l9KC2nl0dncajTfAAcOewwow6GR5HzCfp+vHuzP5AuigUIzg8FIkK
mPuLlOwypt4OK3RG29gmLSohSt9nUEw5rMpEsV/ctfW9fuJZEdYOLyFHqVpUnchvRaXfWcO6vm6B
w6+jvQDSDj+qYPlGPcEwY0jnh8gGdWSNWMM5Jw8x3Qtw51ua4xxU/rsl1IHYj0/ChDuOxtfICzZU
NGji5yf/zpw5j+S/3DU4sb5JX7CJdePUie6XxemTsVstnLsxglC6kRGlyIU/luOoqFIEP5vgubHl
iFYwnWDOj5Z9EVMMaxxtdABTgU4GmvV9/QwMeUWFEJvieYatr3UemIVIB3XYvyhJ7q/LksBXo2tH
cSkiWGgj1I7WCgwXEB2IHmNNHTr3/uqM/zfysKDBl9yvJDRWRH+fcGiVM3rbIaTY1SqpmgCEv3FH
xt0ZrPMmPBokRFr6f1TVaRa0ZUysFI93vmQFTjmOrHjmbat3DUP9z+dv5tephEKGsB3tyymsO+u7
hV+EKk8moJhyO/0lyihWLd0T7eqI/n28mYX6mv072Pdz7zO+lQR+o1jCE26gT4tSxUBvGKI+luRI
ziO/aAq3/ndMiwtdw9z70ynUhh95Qd13kXLjjoCkGSMs09+X1m8ONFtgr75n4DKqzYzStBEeNQtN
EG+eZDLBcDLdWtg8XXbTH19zVnY+zgytzrVPd2E17335lDhPjpuHO+jzbCO4Oh1+ov4RDvel4WAm
iZkzUTqepTAmquLJ2Pyg9FZhYSGdytZIzMjOLdcv8GUVdOS9qfWkdzCBCaLzSjv1XIVEncEtsKRZ
J2MMAQEc/u0r4WKua0p68okmIXwFd28a1YspZNA0aXrQs3nkEwp8YT2l5AeXx3S/ai9zi/kqEies
mKPWPFMZitHr4l9Bvjj3Mi/yTbFzHPStiufwF2JqXKH78bsqHJwG2DSrS6KOPEsUqM2T7VpsQNDn
hXxks3F/gFSM89TLwJzdAQEwK7RE8eaOm8xUjZU8ArOyk7VDjhiYxxA4QO7rTWyUJGspXX96T27T
KyWgbDmMAWGFeAs0DtrVsP2JgfKZghqv4aQZfHBi8ShIgOaISc477fx24F2LTBe3+YWzq1iuPQIs
N+ZA2BBx/VmQ3nd4sW2KQjZKG6NZlRopT6UdUAnh0fKGyKV8W0/7n4+XC+g2lCA9ZDfEDnERu99H
S1ap9wgJmHrxrx78Jx3viqzZpAuOt2U4/PAfEJNQmhled5KcJ7uDm61s3ablyg/A+c6yCS3Z+9f9
ZGcVbHi1C1H/vHw+9FVZqWemPH2nRgzqaW4WMKa+M+VCx0BGUg/EfYh9znNTSUSw8KzEk31LveRe
s7BX+U5+CD1vCIrK7jf2GS9h7bax7tn2SWbqriiKU8jHr7aj8kfswNS1e/Yt0SKuCWvgYZj0Cn77
64/8ynf8zKYYnBLJqjUDnkuQy4SE4ApTd6UQWEm6QQNlOioMe26//4Ih0Z8ZGrR6STQ0ZItmFw9f
IbP0ReTt+oO44Ix+kxT+TrLRkQu+27tmctecz9ePVOiyuGIJoGZ+d5SDJLY+0l6FQTDuyYI9b5br
tKg6+Hza+DLTBAT53jhwqf4OhxFkAVnDtv9iIYXEpFxClG6/vU+AnenEuf4VrmzB5RpvsfMB4FzT
3emMoaxEhT685V0QFykhWUq3Jxg5jGuqvMocqlNlyfo3vNvsuFCmaiCOxzVkoPn0tHdh9tful4Jg
8P1arJIO5sbzj9PMNB7x6xmqY71MzkljPLFe2D/ubi9qaYglslnnsmeXNlU0HkfOfij/8/xvV66y
Tpqe+Rs61l19CTUaVe4i8IZ4Zm47skKhH7iWy22OoS18i0vPcQ2sCQDpJaIsnOE3SqR78ebLSrjg
VGx7h8IFCwSzUA0uRP+x0NhqO+PDYk1JMJRjkXftz4iAGBA4wcRG44CG+BDiSgOX1uAF75SjE/by
Gso9afEylMrugot+eukqW4KKsvqgAHkeLVolQBONpjHov2g1mXwKKCkVMb0Zp4C2CbolspQ/ash2
k2QKfedlcx8UT7vfUpBrEoJCQXR05HjPHBHsZTJf955hyQzoGYyMNjSM0ZwQeULJ7yHMaFRnhVFH
6jquAHREIgbZ99MEldIrzorTGnr8IuDSLbG+ET3HI9uCVNlmmRZNwULpQ42WpT75WU64VWxxdL+D
A6xCLfnLZwZyUS1xshXTHIGz8JmGnctpyVHMYdSwC1A8FGIc+3wV/dgcxbVs+xns/FJC8gBO21GH
RnKAsRQAgVoGQfTPzCvLoxyHPD+/r3gsCfg+p0PgFahtafk5TD4qdFzgxes2PvzoHk02XkabE+di
xo90b3jZ4ZYOk3neffbOBVLBd+qIGH5QabJEOm7ANSea42fK/sAampmjMKF1P0Ir1g2uInkIEiPY
0rMl0bCdWgWz6jIPYMY3dQyFXhC79j3pFfy6v1eOaCmCkrC/8MWDLeaJKIavRjOmhZINgBrB9DKu
wu+QHurE3F/0tLtc4xahPJR7lWfTW5gW4M2hGSV40SojmRVg/Uc6sBsax8nQl/2+QOnS/Kz4FQDM
8B/IrwZgf+RiWot5oIwofTVIYzNB2ewT7RtDYnJJyGKG9K3XLQx4ynI46jBetSaKe+Zh1mYZZQ8o
bP5vG0MImFM8mtLHEzz92bv1956TrugTYSTYdAj3cf8tsWsaI0ELeCL7/vBr36Sfsfzzbi7Sx509
ez4O1GCt/JfDjYe0wkYKpdQ0TaywX8JfwedU0KovFUWHvpKbigRI2q5hz6jxhXZyd5yvtRyNoYww
oNz+/bJw28Xkg3hkhMVHqK8KIpCXoiQMMk39OQoHKexgIbfQ0EIg2EJtqOVPYm2SRqST7n24QVdI
TG4ckEIvlQ1diabIFYn6vO7LgMrpzkQygqgaiXLkgwOEEFiC7Ufx99P1PAVB+mIaCrEBM+wzIcKn
WXJ3a/bDt3pKk7MLPoyM10lsfHRhXkG+Cymiv8f6/+Q5j3j1quz5GxZBSPAEBRNQH9oISIuXcddG
O1sQ7FhpSpIW6CY9hh5LO9JafLt9lWAt5Laye9uZqVYQT7FGTgUl/R/AsTaS7DsGOcPBdtISnMtl
KJyEOa0jPCkg0n8H3dt0FOTktygpKszuG93UpM+Ml0EdpSn1BW1yk53lPoKLh6eV0ABiYuhX7CHE
tS4bRcXIi03723p/btqLWRoW9awywMYV92cilI9ugyPBs/GIe55dlEXDKurTKNSY9t5t2vHLp7qa
V4t5rg9mbcQDQH6TVdVw+CCqQbc8B3gr1KroV96l9H/ebXhJChO2REW79FHB6SsfdY+xfh6PG/6u
+sU14gBEQlEsuywwF00AETDc4wsHa1Vqy/OpqbeOqUlybRMAwtZkDQZCSL2q1F4qUxH+eKDSjSga
4EbGak2tsC1cuXDV0B2Apf3gVCdOn3bxjz4rGj2JVGMXI1aCtnM+sT+ZEe1A75VrewyGAQ1PCTgD
da9Fw7ilhLUYbvmw78uGJ3bvlQ82RjlMQIqe2OVYghzgZZwzmxKAK/B3dUUEQsQ8tnsM9nLvFfqv
ZkMqtiMBNGjioAx0uqiNeJMEIDc/h4Dnt/ChewMl4oPxoQRDOh3a9bvhUQaS7tSsyP7T/a1nIrnt
DddssPXX1P2ibhf+/lPptxncSLHi2Yh+MKviIUYvJtZj1Sxh3W5K+jbquOKQzVZ/7rea6Q4Uvouq
nX8fkTXkfhP15iIi0M3U1587m9fwgjI9SLXO2uA2KBNfMyCrzJdEloUxGoof/aeM+MCSaF5lDBAS
sldwNRHFJJrDtjv8WzUyYK8MY4535kS3VNOcnaTN2AxYru1aqHlWg11kmKp/U1xSyH7rV2JM21mc
KpNSow1xBlIzrBgAibeqfpR5jhJOfO6iUtPZHed6/M1rJ+aqmCpiHDc4SRlro+/4dO3zadB22c3d
8SUcSq33fMRce8UfS2/rgzRtjBat7RqvSc0nw58RsO34qZXrGgr/n8OLw+6/N2vonKHNeGnkBafe
tLIAlbvgP7f0aZZVuMVsfJfimSFGlxVdPmO0t2r2sjknhfEVlwnsKMQCttRiggNl/nBsbN4V2g4V
MUUqP4H6RVXxf4xpWPEAVaaohViU+RlTyUDt9ch9am6pSVatw/8aU2I9QSy/flhYxFO+M0asXmLd
jVI+jiyGty5Ns5gRYN8EMtQBL7ZuMdycc+zFRDNv/73cu1vQhmz7AYPvbKNF0Z1fDqLFedDADoOt
uJOcVfgp9Fw1UOGv3639CNAKHIloItfLG43fSbCY8jeeJe9GA3CGJOUmkbXvwbEM53OcME2jJNhI
a+qBEKjaP0mv7YslFyKK0Wvg4s6hdOwkrM3LI6dQoBLAcqa4eqwoRjX13yfoZU/DKvEJ4xduzCHv
TFyAnBJLJcYk+VJnaahUf6nUxtKLZrIRnzGOUC2mgFL2b6lLn//EmMOMH8t7j8P5eJs0/o/4ce9X
m5lWBwVbzcbyQRuSF1i9mJO+VoQI46Afr9ACU7DP1d41gGS/sNniayBxiZg8GpOaH1QO3yf8E0zp
FOFPl/9/VGegfBi3cCH74yD1+Y6OLASWusaPDV+0MZp9iRXzS+9MnZUrXdeEfUl0rOk9mt2/0cg5
6uDkIOtAWQpZ+Jvg5OqfyW7zrpOTIYmzlba1WjALw3K/bdSzQoVS7tsLY3nA3lDg+oDASU3LWrf7
Uk6JvGOexjijQCMdR+gBvfqurK0yY2TdPNUm0hZongadc9MpRKXJtlkL5CKQ37U7Rson75k1vPLZ
orA8cHK4h0imD7WeDjxADI8V3pCu9E0eupaIecRNECfzaxOvrP1KrZqgbnUsGIXynLf5aAQgeKIp
qzJZuJ5O6eFlqYDKpmf+mQjqypdGa+xLdzp5/P46BeTLSmrdp3fi6NaTHwlxhmClKYgvxHrAkW9J
QWQd91/YaGbgPCExBIPANK72hSIb7bSoQKz0+IUoXIpIT/+yBT7O39NW67du1z1R+k0aThy51bZ4
CfE8S0umisS2WTCgXjIWsNtJTVdSxr3nPQU6SdCvhyIkkmPBJlwV5wu/HJQeCtKQ/J+XTWlh9OCy
EHCd2bz44jFFt9WNeRQP4jrzPzVhJkN1Vq+pNSnzd5W9F21jWtPUNZhE4ebiKhRT6T+cvHhTP28j
x8WJy7sXoj3n6DI2GTo38yxl/ybnnx4coqGsTHdfuN1Jux4O8V7ezXrI6+VkdpLEw3xD9Ue/n1Ra
5lRjTKxmqJi+5mWGsdv3acvQ+AX+KEz09RZFU2UCUaoqXT2YVxA/vMXVWVsimI9kze6NzLVkpMjz
JZTumwUcmKeOTKw7hueYu/s/QfsMayxo2KW1N/5Njm8n4SG9l7elWSKyyi5ImERxcuk9nWt2HgKg
FEB2/cu19XNBybm5ZoMIqUxVF21rD5s/ka6elhNyH56cqgGdXc/KxejbMnYyiSF4xEUv7jfYjqqN
/ZyrYQw3/vM88i5NtTpNV4KQRnFjxgRZE0e2/A4DB/lPr3kh9V4JPdNulzG8DgHWV34N0zZpDNlm
X9wD1m2ZO93WrTCSUiZcy5nSCIjqb32K4vhu8uptOlGuKItIJDrewjh61cE2olr3DSf9xXuC5ZIB
iPhBRdpB3lWxnap04UvMxKy/cv/bvZIp8ILZ+aXGhKI467aQEQ70W7sc0GucD7rehCje/ZAi7nm4
X9jo3/8hPRojluZAtvTaj3B0J6ojwlG2ksSrIAHkQ0G8ZNrZL8i2ZdyAUVF9tpMRXe8IM/6CyLgc
VQgIkp2pA/UafRTE/OenMcDPdr2Yu2xDCiPibiwirtjqE97rI1sHy1j7DWBmby6h5c3bViwmjA0P
oGjNZgm6L9xpal8ukAdf5vmCa7mFOdwnzJr6nz8Qn7Qp2s6nW5j0xiNzBOLapLtGEQOioLV1QMAo
Np0t9TbksLC65kO+aXw0gsWSOamH5jw0IC9jKta9bTC8KA4U8+i7TKUy6tTD5nwQRXRrhCq/2WKt
paaEU13R4KrJbszvOeomJDQKJp8VF3KWveJeB9WgYl0ehcFTGEIWU8fuMWZ3nJ/Alhd32Nyrlouz
vMy+F4O3s9qIwoazotBtC6vOQzuiC3SVRC8H/4ByVYenhS7cK9BkiKej+Pp8BEISxWiLaNwjQK+X
q77V6xhcDarTyKE9IC/widUPFo+3tw8EOG5LRTj4hj4dIqlhUaHUkixh6UV825c4ZlZB1aTwA0i1
i7RdMk533VXBFKQThrrM///ndeJkNR8g5n89BpV5Mq8ci6XaV9BVzbGV8zihH/VoTnPXNbBLJgox
ptpbJccl6CWWsFTTHkatHzHxKyUzCkaCBukv3cu72ukT2v6NJTn67zLkhDUTcS2WpXYpqDA+phof
rAYrYpOIpZxX1B6HU74kz3oKZ4R74YWvHigX5LtqPKFwu/1gbly6MlZpeGkXoIklvuO36LyjQvwX
QA1v1QMWWyAI6zuYgJSuDpj67/+5p69JGx+mBAb1XRqqIQ4xi8vKzrb1oII2Wjb4CaQhYCAE3Xtk
dmKPU225mxH++Pfcmy5KNNJ/1kdJ2k+W4a3JWk2B/iFPZg5dLC6pxBPldEIc/+qgWRYa2Tsi1Vso
TJCix5+MP7dxtzsbsMhRhx4tLADDClT3Tz1SV2dXMHhrZV52t9R2EyVH1NzU03pMnpnhzoQoVV8N
la9ZvnKOnCB3lLuyUcgEG8QCsaAp1dWwgzeZaPXA0nFXO2RFy/trGckFnflchuh7/StVlV2T7lPf
aoUEy5xqzNIlggJwI76tHB89ouQo7kyAQkH4tyhoA3DVGifQhgZVxrT+xUV4wqsrTxq4xo+B/AUu
a+4opC0MpvxwWzvYUk3ck213t185hyfAISSmA2reJxQXaEbqLzncxEHXwMzrW77C20/sCLGPGsaq
OubbGjONaOnBjsckpRfiM4+5FdJHM25/By79FUgW1KxU6W+k8NJ8PCANYVaAlQvN7rdPHmLLT3HU
HCNOQ9qpgTLQMPsdQxBcu7A9HQnz1JDZF7xDeebM/9Yx7yKleYNWfLBv2NeNLEmEV+pzXFct4Ho+
gAOlVyMdJAkvOm7GAuIsV00fDcxDGkRmWMouej3ugtttZlU3uS0jroD6/yl4mYi2rr+xAXrtu67D
7YjFPC4xaei7xaAfNiOJlrswa3dPHiwg6YoX6IgFBGH9oVZvtc4YJX6mHll3ZKwEzcXRDdQD01Sq
tcKmlrkmn3FncfswYcJMOmghgvwq1N678eeMPbrTuXPzVq9xUwfBUwSO04XhvRv35rvpfegwG4Mj
SkJ2CN61dE1sDZmJc38GnFcuEhP9g+pOEjFzlaOcLsnkOsWFyFXw+CHR0kBUrLlodL7qdDN6u20w
Xg8YVBQJ9rmAuEElY4yRA/0gPgFHnMcRWJGEz+GmmHY2e17OQ/WnmxT8Io/+KeGLyqQM63+Js8kN
FIdMnXX1Dd9fQv5063vanLSnZk68j99KLN6K+yLap2K/2WaorwxrqumdBzpu8VWWzEZa4YTidLkm
Re7B8irEtYXydspzisMk70HIuV8rKDHG8PToCmyPS+EMAaNMrbxEegNxTF1uOXUFFhxWXC2cTrE5
IZRyK4ibrSoRw7YgO6Wt+868O4RkohJfuq8L7biGJeQaGpMEDrMNr9Y2/4LBd3A3FDV5TroUItbl
Mfz4FQ1aCgI+WtNDLkOWAABIDybcJI0kS1r4c47FALuhoKrlQfqcgB7mBP8sax3LGjVxuCt0EPod
2OUApgExd7KlC1tmDSIcQAc/7q3sOtue2RFzzWvxQI1cm6Ux5A45mm8bshwVJFkDtNqJc/DZyPRn
0jh7L7h8Ot7XdN95YdvXuXDuo3EmNKr9FK+IeaX/MA/7zKjvA4EP+9aJzmXDMW6GPmBu21qsPFpD
eclm/Pl0ms1X8m2a+f6aITuOwrx6sUnxgkRtamAvQtGa+/kiTKhfTbzDsbt9P5ip011MOj7tCUZM
OmFtWCFz4SprS72wXEh9eYl+NT15WPQZ+iYJwcDFFJlJldDQjvc4DcmRZ6aDnOsb8727qyhmolfp
8bHfJRpBO1ttf9FxdQ559buOAO8chYviXiy6UfY+JyE2h1OI8jjKtkT9q4VD6LBIyTbT/CDQVf8V
nAo21MoOxefiWa+nPFozMfn736zNbGhoHOSEF7kGfvtd3XiJ9UznZf6HIRvjxdxhYWswiFyEiL3p
ipTURyDxrmtpIRQJvsl6arpOqlXAhnBiMfMNHDNbODPm7zP5CVU86WC8E+NIPUQN0fKVSLnsoi6C
F96koT3Yx0qGrRihpmvmQXIO2CwHTJvlX0il/HcjJaoMX+dJSRqcswFIwZ6ZEDJj2MlWzbJWph1f
tAs7WApplo6iF1FZKj/7d7ojy3RFa/STP7NMR7M6Bl2v00+JWfYs5S6DpDyEFsjf+2+vp2IITG/g
6i4EuEZJE8zCzhHKYzNiCA3Atde6ZX6U6A49J39rGiqU8+s/5Nz7U/mQO9/W0+SOZwDi/BCJQaXj
v/jeFembjPuC2VvoXGTtZA4WftLvhsb/Ey9aFvRDm1352JiWKK/FUF4l7m8PGmtb16oZy84DDA/y
kY86lhE0xk7Dnv7E1HDOHIwyPZQSOn7iEylcbWs2txZO/Li41X8wvIyZ702CEhqKLWAScVKRe+f7
U8gCBAW6LKP+rcEH2udMcrl9YuniBp0caxbOJSwdTZtLDXVcMBKvsAVfTYKQWiZDZx6Ofb+/Rv/H
P5ESzXyyNVG0wVegatBIvAs0YHwNxDJQ6mJiH2kgY64fyJW1a8KjgoQ+fC3I8amzpG0kyKrLczYr
qb2ATtcQE4nWrs+ecFG/mmWxCTAIjQbiR31sK/F2bUz60GUPycwKwNzCa3Galb8w04i7YtO5BxRE
rr7+mEPt6lpfeJ81yjBCr/u8IAO7sjz3QJFuSE8r7fZd57VUO+pbOI81F1mYgYCG8YkYGh0j7AU3
bYqdrbG+q/wCfHrIdbY4hWcVASwSWxGA+RSOp9uQIvwzK3OR9/Iyh+HOvMbr2Ftuwx2CeRHe+LMM
2J+3b22EcaTuNkTM4uml05FGrcDmQJyLxmsh2qci5oUwClN9sG44KdRtT4SE7GUkPyymm4sAybaL
SVlJQXQkUxPtrbfo+yzwLZIKQySqAuhjBPvqYSfym1Q4WUOaDoHvSvCSGnb0T4KblJPq/dRKev4g
+/fyVazUuKpgAVk60JVgKCUqe5/pqAOni/a1276B0lkPflszN2qnH5kTwvS2KIG3JFdwDYDbSIKA
2MZpJEOTOBLNJwD7oL98v/qIt0lnOAt/N6daLsX4EuswsOUfpImJdR1BnscahTX0hAMWF0JMfeXN
udhj0JUHiAmSIZbuccPWrC58Gb6s3tA91WFB9dWputcSG9apArwODdQ/CkJdC2A2XjcSjgQ12FYI
jMCbqO4Rfo7TdgKcVIrA57eEmnDnVXZD3LOOrPCDiQ7AA7J7Ag/4lVgQpHDWIGHyEdsF36LWPzIq
04Z8pHukwfSWfihrFMMdZZqu1osjEuCQE4y2uL4vCu7bYX5Ani5gXMwy0yNfUyxF5/nSbzKXR5dN
RvjhHfQptfbZQ4CNkUyM38hR9zjbF2t4rzTKT+Zjz9b8hRJt/LKnGaKpNaZWYA0JVgHl1ICKuPjJ
mqGipnYWFBvAulSznuDnlR+aoQpA+BRzJd0W3Niho659mABnyiMBdBWkrNavFADZL7TOaykD1SQR
+wln/nhA4I1etZhJtDJV7XH2zQyzLtx05OvmWpAEhoxiBTW3DlqGUdlFxEGMprJK38Eh0llq1jqm
AeJ+iB9/oJQjPhMhWlJ0MZxbXowsf9xuXLN1HLUWjZTjE6C96LZutWHuy2jP20BHE4G+asiF4lEF
u/linqfRvL/R7f0wLc33bdav5IZ1CQvy7Nif50v5naCRVvi3AuKXRyhdFgBdf1MRoQYzhJIxlCkK
q012AohpWmyC998Y1vjBtd5IURYcvlQC+yFANGUZEdYdCN1zE7IDKt2lgWPe7p1t1BX748M5vYGO
lv+GccG8sE0PP0aiU++uQ3vbFeGePYgqcj03ZZL1hU40kPI30ktfs9g10+IP+dm/0wsMXN9DoP8V
HIFPXn8lylOGDnig+gMEMq3ZdkSt0zRHStAGeLvU2YEyDtukk7LfAtL0dx8iqjtuy/d9ioin9itl
A/bxS4oQi8JaJzzItyfWSn5g7MmYuD6MguzgRZn6iPy9JK2DTj+VnsoeWmCmvPOqujNy9v0NJns4
NB6Ai22MkKgnan+DK+UdwoAD/PZ0ygSstEPx/Y5nphHiQEaKJy9z8NBpAkXIH7iXXe5kWjbr1AJo
0vr4MPuk8PxArnHk2tkPlRygFIBdVI/n6yerXt5Trkw0kflTvXFyw98dmZbwpP3ItM1Yy2LESRtJ
UP383CvM8NYo4LSVW04F12d7eIhlP6hTnOExA1jWWlMZH/KL7eRKKWgqUm7kCDPb7blYvtP/dUB4
vM2hW/2C0MI4YtaUQ/4uulIxPIUU/d0GoP5at9X1frXMUzpW56ub941xJjqFZRDFvwm/qGtyoppq
0/Pp7lHCHDLwmUVZ1fVgnj55juKXlpKa112C0pd1ib//tPVeiIo1Kw47EQ9o2S2qsPX1P9PsoPlQ
OKv+uKKvIvyBQSw37gYEXmVnAArRGLqFVyw4uXQtXm2l2nq+QC90MgsmmzTmrKW4ZCyomiAmUA9q
I/0Q0S4hw3KN4KPud690fd7zYOQx6fi6epyZ0FqUJ8H765Gb/2S1RuY3WstssVGHc4Fp8/bjFZkA
RHKDXPlWgAe0IwcFh5KysL/n773utK91TrUICXtTcm3QYdskRRKzKz0dpJqaPZq3/kapRxcNysHW
yNapqi2X0dZHgf/UySLoGxd0PghQVVkLmNP1pNlCX7UWRx8aCSvi7qkcHVTPuX3PSZnTWU3csoRm
DJCPpj8jVOLFJCepyjFMWhK8KNEPHHJJEc4d4yTC5ECZ7OhqQezPVCSs0esGn+2vdEwV1fv5oN4/
HUIicf698IrFzthWoSXOuPYLcW+jyvdzoNwDBqexeF0Iwvh/XcDs9ArIxexJwg6cUF68jZjKp63L
vP/dbBYZ8slq3kBVBeqEcoFrEoXHJipBMTF5iJAPviOwQN/bGD28F/9FcdWux9cm/NPFRz+iUiaF
t9odVv3z30VWBCCY8HMeghwVUJFlNg5yI33bG1pm0E8ZnfLV+nGevSYaEyZV3neU8FTQUXe7T1LZ
fRWtf+u4WCXcN/dCLUUT/JKaqiFwtOxH0/PO+MGiq6q60pHkz6x5nxOiOCwOF2WbnO5zZPerTFsS
qi+5dvnl3YuaGqEG32sidPpdWobcUyQXkV2qnTt0/zlfVd5yF4fyxEH/lJ79uFeBbMAQTKcWo7mt
hzuw4D5tH7dv5jmAHjFlrDgr1l/u46sl9/KQuzlC9n2Zq+8/H8RbWLWyDQfOnsD8plMChJDgh4Fp
649kNpDnF3Fhlp6L6VtP84CBOhS/3OVAAWyotWEVZBjSWYs2rt/Thxqv1I4ATLAy89hcTDqB2JP6
JHsfWlufo4mTMWc11Aq/yYDfcZixc6hBk5uABBl849zi/Lq9CJagt41Q/Aehaw3OdbDX51qh8pCZ
OtWGtwuqwwCIAURNicjvaxAhce+ib6ZX77ZIerzXsWdjCwOlq0Ln6XiazNu1YsCW3aiIzTppA1I2
tvK4zLoYtYUJZnJdP16EVSxl+E5woJPd5xyq8vnJ2ctAZnsLxO+I2o2ykcqyEveZwM+EMawgbxYY
gJHPguqxyx9FX/UuPW2JFQKW7xXdyCCpHrwuVtjFj2rQ+HtWUb3zSMUmcXXdh+ZN/bimYYwDMqIm
aCYdUB/0l4d5ecHKmSRu+ZdAtKpDAr3L4HGSku5n7PwdX/qdZMpPn4OlXHw4bQfirOyisPLycZEU
5/vDWkpP7Q5z/SwBCAg/uaNC+E6XQesl3HVwL3nltANSzy3hfPo7D7YKB3x6JhawcGwP+DL5ajIc
br1B26lKHo0zhq+SVQqlIEw7qxPV1hGx0afMAX9M0qjmhLO2kZATMvbZN+k2LKSNli3kzxUnZ9fS
qeeA+e9HthJnHM3yUIvAAWuis8o55NEGSirq7MJUafdBxAnB5lbZNmt56uk41paeh903nwsBZdmQ
xREMzmoJx1pxCIlskIVH6gHl8LEkQx7edSeoheQWaV0vxClY34d5HKAaDaP4PC9vPqSNpKujbd4h
xNGsf1jkiOgSv/ObL1uiAh3HOIdokKZiP7U1ousVAyJaNhTWsOOiFnuwTh+0B9r8GxcbAd24wLVQ
NYNWYj/QYWq7chMFvuegnM56ylOFUF3z3acYUI1JDbqXXkqXgPYkC7IjouHilyUGkdzei23P6I1F
mC/B6VMfrv2s92PKTlmgIf3Of/JdTunMJFti34doILM4D7uuTzr5O9Uo6SUnhmVBQsQ5u6fRhN9E
lMFWVp8rJT/oZzCIsbtp1LSR6tBX9Ntt3XYRspvVxgnX15AohF21knQRpQU76L+PK/adyClO5fPi
5AAgJ0rGaFulI6QBNknSEB6F7unDEbICuT62OA3BDbp+T6xlvMYjX3BK9ZhEBBwEnK8U/3XG9TpA
ggqmLmNOX5ODkRYH2QtYdmMxnM3a4KKVwlmsKyct8EgA9wsiCTyAeGg8tb8qCs+K7FKF2YdWVsvw
0FMWhwMiu27z3RdHbM5I/lEuamUVbddvnmJvzRa/K+8ccrDYjZJv3BLPVckUMlcypKn1E6zozK8S
OcYU8WDcUE+3muiHyR0zhm1wSQyYOD6pr7pCxFPC05aobe542W0MaiNwWkEfNntRs/I9sCJUX8oV
pjkoC3l1BE1ZWASP5iw+J7KHTYFWoPDklGc7vyLcTFAkV3vIHqeXN4xTGTqB6bEvOfy1cRhbA95Z
eeEqu02DydvrjfAp+4+IonaH0G/pU3Ihj1GhGihxP32R669hcFi0YxSzKlzEl6Vp/8zxWEAOjmfO
FpkipshvK4JDhok41/8uZjHez17KeFoxt/bEP39SEF+aR+A7RDNpLXVxkUohU6w9bIQgDB7T/bW/
Zbq/f28O6n5uYLRsNItC0xgF8WcBk6Z2AkAL56rcf3DZ58tsDMiwmAxZQzkmOrWG74zAiItYndri
uRtjoZw1MxBa0Bk8dXH/qBbtJ+yRRnkMqtJ2qdO/De+/H8gQm9mYNB34rVBsjvFYYJOSxhfVYn3R
sDps7ocFjfr1WBL4v7YmRBOyZZI0EDrqrqSVJEoHzscu0C/Y0ZMB3QUk8lGBpfNQIGT8GHcsxg0C
rduxYHLIrlOZx7YfT6Myf+141fH9evC1mMM2p+ZBI93WVgwaaNu9vX8srUURXVT7gDtN7FeVTzXq
u4GZUYl75Nuv7YJ6Bw4pkOMeLq1b17Oy1v5f21Pcq7eBeX/YZp1bTVPwy18MWV/1HK+fbAe1LPfO
B8RxpRFxqJ75CIWq8JcjrgOcmjSzFCOoChIgpRAfUqZxC13tH+0ChoB5O+tzqeohHogLgNUu37+5
qcSPmRTKVA62JiwG/JFUxAPTr7ow2W3JD85IMNWay+0gf9R79VWjKieEXemvbJdVbaZPrcI2a5Tm
XMW6y4y+CO2WUS96UoOhkUKYA8odNwbx4kTV9T0p3f+1Mn4EmoaMjTujkFeXyaQ8KHjEN6BlNgBn
s3BVLqSIt4BJG+mal4246NdAaklUsd+7eDjFrU9CpbhZ84QkAmUQ3wj8QGXygMv0SzEiHmVQ1R7q
Nxb5JSaF3ULJxH1NfcXrG5YyhkQJ3bpuTrhTXdRMxzm94GtuatDGgdLccshxVVoXHaACrMjvvfxF
oSbEMfUEqhnq7r3anZKYop0pLDY+lEdZ8XqLlBnPzCe1B+6xMpQa7YRUfzgBnpzw/8TDWpUC6CWz
/y33YtfKn5YYlNKnsQXjwAEr6PD51IezKXapYM1HV4rrU/6Z8hxorJWaQzJmCKYgCsIE3E6ZaDqB
s+1ErhORsCvxvo1sU685Aep0AxgdcZjjCw7Ab72IW/8RQdIwQRFRPVkS8BYC3UXeSq8EP0lqQNWr
fbe27avnhWEUhVzpXeLTE/myYLN84r9WXVBiij0GOPIDv1Nu5732D9znNJtE8zXMYbLjIlsfP53f
M42bnLwnMiaVbi/LeRqVGhUkgV3QiSPRqcJk5k0jC9qFccIGLyhYpwXnkA9e2cr7vfXFZG9eIdSX
vXTyn6Nkf3RgYsAzhJjWkpWkTPKWP8Vm3eq3EE2TBai3+Iuv1DAZAtkKQPwGnwURfeZ2UA5r11KQ
b397JkBaBrHLjXS7lzoJiCDrjnAjI/bVcYNEM4EV1EQWeE27L25ZHWwlja20jHl4bYb4k4jufSQm
hyIWiRQOGHskiI80DVUkp5ERuPTsA+FNwQvGqfbxEEMhe68Ix2y8r4QsrJzN3I1KyMBh4EJWI2kH
uRLKqvAcv1Wej5s7+cRU7FyKVJcv0qgAuVt1ZJtk18u34Sp4yk6WZBPCDw1jqKTRFZMJEzsUdL2U
bVg7j3k30vNhaBYdq3AuJLfs9h/UhS3EUVqolcVusG+n5ca4gpBJ79CkqWClkLGuwNzPKuTj4NlA
/DL2WQCGFcyn7guXwOhICklk43uSWZ2HUS+Hl9ZCFwQNn2TgW0E3EyKRBl+c4AOlFXB9eb8dKnVT
tUVmSzXo095V8vFh6e2JVBgl5G1UGk8FCEmXY/q0CrWIWlFpy1z6AFjXx61wkXSnSO+55LWAVr0H
rZjoy9jj3O6qB8VyR3JFm37f+dRio9ysAWaEdDAnHZ7X327fhdcm6NpCfShvLx9SX4qtzrnnHcQy
aThVHmp+uWFVtzy1yCr5LtnZHNfhbIzZmFOFZpOBxVZ7I+hXvmrRzPI/Nu+q6oSPbAo+UjjilDgR
iIWZZB6pyV4M4pFKUDKLWov5UgzfaIrUQpgTCB9dfEi56RRsAw/HYyFL+2Bt8aySXXDHetIOoffM
2iB2nh9YnrBISeswkNk2Kd/MJss3+TSr9wp9+RfcmGeXiUHe7gGzvOkQ6hcljZ3d+szUusFMzIE+
UTK/tvrOScr/UkxONVlr0ViURQlbtTYYbeJNKfdBBVSrdiHwr/u7bmO000xIBiQnEPLBBXBGSf1L
pTWjSDQlYol6uwUQ+Cuj95zuQMo6H8fQ0NSvce3cUUezC58WPSfBobATfKwYO41mLo4gyOvBGM86
A6TzxcmL6IcmgJcAKdx1rSyACpmrp4XgesqXILYAqFCDWxjAFnSLRZIM8oCtNWdgwGrrRzSpL+ir
6cQ2S926eqLWC64QHYXJ1Ns7a+LTvfzZMYVQqvrkDDelCfS/gxUb+zxkjuGwayPpc7wq+aHaDUFG
SWNuE8JTh8Iz+hukt24qoVlnvbzeNuXcHJGzG2lMpyUhZ+QLH0EdotkznbavSFMa9o8TVGc6sQf8
/WYYve/hcNofj94EJ491IE2Pwu7X+Uob/HoPnRHdY/V8m7NowGjRn91XCvpTROevxzNsVRfItDY8
t1EI2MXpL1ikQX6OjYVqg7gWWyOBMkqTGEOGWQUZBCx89k7b6hkSCkfQuaSpXPI4ITVoLGR3A7m2
UHQ0zW9fHqDnhCcLNBwucowQCW2uSQp0QJ73ztRA1NUBEONvp/k0El/wjn5IRX5duz1VWl4XWx74
+SqD1P2rbbnCXHNaUI4qJJ6dWiKdLKQMc3bjCD0e/U57uxlb3m5/tGRHMqNfViG7kLsahXd1Zeh0
Vksy7UgZZGCvTyBxsOggKPiSB2w00XhepRPe4Z9cKvD/DFVoxfOVym+B3itqa4E5opDKd/UtBp0d
T8XSAaT7EO+qF4XFBKFSjnCKDZIZ85jUxb4YNHv1a0K7F0Ei85nEbYvypx/iT596Wz/Ai7ih1nw6
tj3xCcbUqG0TFtNsejAKzm2a4oyMqZVA8TbKyViqKYmHCL7Ma1kSWolwEROUCFyRTqEbtE6ts7wg
sJCf6rOp4MnDmASmqAUccekUcjA/TTPS0XBMzEnX4H3KEBQp0QNl3NolUpxyagah7aM8xbWPM/70
Sr/hP+COgh0nYVQDozqlrVP2FVWDy9t253H0oDrZSXdTqX0kajqq4DnTTjVt6RPfRE8riu1vgILe
arfbxT+/PRsa5iBZBw+3mEPW7LhnQ15iIpNqjNEI3dZ74nYLMN7Pcek9EnnsmGZuH61ka8hjE48P
iK5SeRFd7jQ5vH97fhwxa8jbf72nnCdQHZ+sSLyoja5gz/xZS/PwAQlemZddLIX2hHY29rLF/71i
gLxf2st3g/+aBB6rGaHW0CgDL79a40PIzTx/ArKJ9J7IG1bekYNz926Xvmby+U/BJr4CCkufRsgl
A0TP0u7cHd0m1NVxPLYllkpl+WfSxkhGrC52KbF/UEWtzXLVriy8nquY23du+8klZRzDlqeoAM2a
3FCFGA516e/SmHj3wuVmdsMAWZTxDzPAhoBXyT3xqbMeRC+3wDcs/CR1DwBMAYJw7WaQFgHRJvCE
UIQB+KK8FNx7ZnKe/B/H4Mv80nOz2vp2IqZoS+GhlvOmurFm+q9VG/k261xKtI6572wiJjdFS7bM
xguFDouYGvJNLyt7oyRAvJbaeyV4FvIXFLQO5aSATEn28KN4dYmH1zsuy3UdNSR/F4SosfEuYl04
mpH4EixtQRGgYwsINXjLwuwvA54pKhLasBCOKWj2cme09vYe2X6HjMP/Zr5N4oUIo59pNUC2y9Mt
wpn6xlpSQeVGY547vQievN46UnIhttxzb1arS1QAqtf3Icm8FL7GHicvh1T7MfBEn3GlbShY/y4M
jc4HEVzj9ot4RJ4q3x9M5QPh1eG/xOyxxRDtYtGYDj0QJVtywKVi6XDYc9uy8Od1tiNBR6Rz6LpJ
WS0HOCTHQEVmsAyE4vNGVodeGI0eMFe2jqAad2HE/0L797SAXXnsQBavvZxnwd6VBuvHkaxeshiw
AhRxyey4ICLVf6qkECRjI4qbz78v3gMh9B+AyeRP/FkK+0d40xfCSRc4XXQg8F961DdNIxn2MH60
TMnqENJqG80jnS5KcNyVlctRh8C9kBUsCz2MQvyIrYFMgrg4izDmCaMG3PtZzTvKcyK6Q14/XhiH
nWGjVNLYsQN2mE6Hvb6xojSC6XDu7zAmj58CtdbkzMzRZeOHhprJC6IXqYZvYf/Dnh30aBKrkbOV
5NVWKxz8O3JbSPqTIhT686/xN246F/I+t7ilS0JpXUdvcp+LoWbFaMIcMh6+kt6Y8CZkprQtQrpd
Fn6cwQOZVNKtUn5H3Ek/MOyx6H3fVtTbpgIvXRxYzRkW6Bp3Uw3jhB5WGBxEHyODywsGDqq4Ebs5
EbCCkXTt3YsbjupTvZdRrU1a5vdZnBiMsHD6VOnYRaG33OoHM1GEKZkqrBg84AWnEDURfHCHpp7Q
nXS/f1sbGgRya3HHbZaskWjBWjuiqYo9f9037MQLj8Pot42Q/w0V61xSbuAFwcgL+jIK0wqfiAmX
/vYgMFYj8e1MHaSMDm1+Fj6N2l2ehFz3BoEsdyRKBY21jOU93a7qnis6WtkWyJYlyxEOVksUqJBa
5CI8sPmg3gGI01dmoPm+Mlf397COhVKNTJLEqN6s8UrdjYa/+4E5DdwuQD/BjG2d7LuddQH6POEd
JraODYV+lR5oZohsdiUl3Nk3xOFH+1XOHppT1OAb4+AF3Wsa/FyGGd/1iHo8eoKSSA9oR9E771PO
ik9ZsThlUnT7e1rB1SQ5mxsGuPpY4bsIHIMxzsgmxTmazk+6iKn/plZwfEwMDCQbrl+BgBV7IJ+E
96RDEHyNcgcWPxhBoS6XfW2A+VO/uP/napCqsW2DSnm14v7gcR5ZR+xWO56rcOu3SwlyeUO/Ylzp
PmWNHQHTOXaT7uv9xfKgu/bCcak1OYPphnA5fC3bdzGYdPfvEGLS5pYhiFl9dNBA8QsXQqhKKMjH
5OA2jEZRu8YSSm+whb7DREAYR2vTxIgZJHQaZ/tf2XTfXkJf8j11jkwbNVCrR3JI6fnryOvFKn2T
VC2tADjQsWoBTfdyKKBKCjSsZHUzReSk7tqXVnlE260aEyRrRYQmlNBVCCdgbKnmd0agDd7mYJWR
y9B5mhkOzLgb9LrvBsNIBoAPljZn5uwqnIxymU3PEX9I7x01M2+46Z7ZLzJQgQy7vB532DLvzFNu
bjC6LpcU/CUnN2CQ8zxVGndQeNDinsUCzKsKkNR29yXxye+lqHiCNOykS7wtQxWyF86CzBtCtJVm
duNUHMGZWwLX8tnblCZYNKwT7gCFxvDCOXkjObly1mnQEP6hP2AbyTyC1KfZN3y2N8LuW51Bh9lZ
RWHkcjQWLs+dgPzPgpdVol55uK7a6a/h0GB5nc4GuqOqKEKgrix7OrH0ER9GuXNBO6G+4r8ejmzO
DRvPYsR2+5Rg4+rFBYKym0A4R2Ys8K71SIt/IVyPk+ESi3QSkC56mZkv0kc9/BvEn6QHM0yie9Io
5cbo3/ccq8bFnDVjOec/4GEQyBR+egW8s9mdRzNvGbeyiTRH7eGaMYnQ7dpGotpfbS5fpctlrg8g
qxU6hoif71oUU+v4U+pkXUI8aF4PiX5HCXgwWH4XYxEmb8wtxzj4uXTP42VlqMeNclLTIwrRwaFb
e2IS/lO6DfQZWoGv/grDVHbK+mkMBJkXB+U0wrB6PnMLusv7uW6cHclh7bzWwsDjnjFAmwxup4/4
RD0vpJ9kLEjYWYo+BkmaC2tAub/4bw+uZ+E0ooKgVOSpSu2sH2oHtaScxYhICpiW/Ba1G0vu+sla
IAyOHQ1bHkuWpuAaKAomzbsV+VqzgT5UjnBkhUoVEX0kIIPD2JfCRg5bcEn/ujaeZvWzPKl4dplA
GADoJ4Dv0F0tJD3Gw9JOJaut7ZUY+32iDdkouk912BNwEmeMWky9e63XHGZdxXcI9cyfl5mHWUA8
yR6VQEO7x0PL4UMghwOY1m6snELaFSnaRfAFw5hisxnGdlzll4ycvyUrPPnkvYnDDTr4DBtblUNG
HZR9QEV9NM9/62K7mLnWIytQ8TnQMqvwCPLZBebXgCtpOTWmJkJrqAzOPGrTXbOPZwzJ18WaHXDA
7DdHMP6oIDcjfvi1waxoZytSsMoFl7xy1qXRjeiWrTNx7UAb23mCpkG+7VsZeyvUow6BK6K5eM+I
ERGk6rH/S43NUpheiE6fmQ7QxlvX9IRKjgZBT/2CQpsFaJAjDSaz2ImC0/ZN5svwmsy4Fpa4UMQe
vlS9RLe83ZMavsW3+gNpyEPgi3UzrgRmktWIkG43X7qZf7Ji0CNCRjtKiEm6yIY2QhnBtUq3tb4L
I54/wVTTRI2w9yv7j1R8dxXERSrFqmdpVKPzHMWlFzNPPfiT5GiXT8lkpWWK97je28O5H6WD//bE
e+kqU0PdGjCeF93qOhycdSyiwTIv6uvf4TUCy3YuuXYCHu8a95fjHIu6ksZ9vnxHixpGiJjGvdqJ
ZvAE5IdZRZ8fdmn/DHoCV3C/OTEopP/cognrMfRzog7Q/z1USBiZHyjnNeG7rK+Qd6rLEf4ROAWa
wQX8kVP2vpPQmep2EWXAjpfoSchLP4bNv1TZ2q2+4nR4+G3u/+PhVxobLfCs1IWH0SIS6fp0biTI
lVqdSO0O1+TFQZXfc4xymMmcKyNwrjzSrQN3J88jtAJid33v52ZkdqiJEBh2ExGLBGKr1VC5aMHj
tDUggb48WPkKbBBhNxH3HNiKn3ZMIzSGNcC3OZQGNRi/oek0tGfzC3S8ffH0Ovb2U4bDdPTscA4S
x8V3HED56PM3LPxJkX4DFUt0B7z5ls6mxGMbrlBrL8chOrQLxM8vYzlQLA6zZ04A9MMoJQThTICt
63uLair1XPqsLlk1BVRDZbRuCqppWY3oAtZIpREjGz3RrU5cVvDpohv/obReZzTb4WUqf08n07eA
8ovRcwwdgtclQYLOgrlRzkGo53/sFru0DMGEwHrIgXLY1NfQUD+UyOnJThNb9x6UK1b4HHtRIe88
Pid1RUX0PZjlSeC++DXCmh1Vi0Kmew76uoE348ch/MXm15tfSFrREC0KsNyVs/Buc/gj/yNSXXfl
qPK2/fG556wlgvpLAbvnK09C5khbgHpNTsRB+obJsujJ7f87J1WekhOUEYuW7SUO7KhJUC9/rORy
olq8t9PRaS38TtRj1HT2eQq/2xZc6pKuvWEE9XnqVqq7HUutVv6ub11ZgGjBQL9/Bwo3z0XfrWl9
Nw57+0RqT3Rm1+nPXAbfcQ76w9moJD3KpUW4v4meD7T5tcm+oOTsG3ZdQPJ6mvFiYOOMfyBaNHrv
yJ4nophuWDoVdOOBHGMAj1wcc5ggBW29Sn3y2U6nlR69/M+DJduzeMvcdWUUQH7zv6Buyf7GR1C+
P3b9ytxoADU19X5XUPsSvpOYolm0uVxNf4QZng3mFzwSB1dhx63HqnMN+HBlSNN8bnF1/zDahtwR
86QRO6h9q0tgG4FSFsRJr2tMLaopDrKQjmCVeF0PL/yRhAYHSnr6kDb4f2wUpf7TeMiCkcC2Hfsi
D65NlNpJyQgWcJR14obZFfORROvGDgcP0XOeV67giabCmWY30iB+1uz6T3+XxUf2XJ0E2sZ6JPkJ
emS4CvMNh8QWBKvRsAwwNpfvHuBbBr5kpVt/PKeUF3a5ICaiCEyJ2NsA+hMfuDxRzCgrGsO6Y4PK
VfeimJ/9OUG8i+0Ji5SumCCifeCmSLwBh8H2oSHQ7hA/IXzgOoBaxZEGjrdqOiqNAOOyA6Sj6Pkj
V+5Mj3p8mI6YgrP4u2NHeUqUXYpMsjO22wBzcZSgK+emS9I7QrSltaJhyw/V1ZZHX0vKjndcs7Pn
l5Vo6zPYOhp1rGq7yibkp51I6gB8vlk8WZk3lB0fCjp492ZznJBnK28VR7VH5FrTU+LF2VSh3juM
mqIHpD0O5nS7/nVy7/qulVurlb7Ivlhco1IdOePa5Jo++BggC7Bt3rK4byblMQgB2F5qniSe8LBM
RsFbvaXiXBnJz8qrlO/c+hbQXXCL7MbyCWyAfs9eLv9PDxGggc9WqXLY/mVV7lYvK6LDKiOPvZWr
B/nM272z/rOXO+JzqtK5+3oHEiBxDRZ2sZHMYqFCyAJvAB1XSbZLY/0vnM8SwfHy/m+jm1OBSlUN
KCEetIlkbbLjad1k5Pgj9IhkbYasLaLUChamqdHrDqnEhHtgm2L8ehVu2GrpB0XGrj80LwUu99IV
clYMifY2lopRQvv+Y90l+ICLow7QUtZvpJdfn3ana3QfXw+iOOENlFlDDfivIM3RRLwmdHnkM0dv
lGsAWL+WYf4cwsrRKOh6+7w0sq8UBsS2tgm+42s1eH/jHz7Mfg0v/zH9slDGz062QH8tA4BjcGoM
QFIKCyTxFy2QWTncgy5mBSsE2uzkp36nl4w+wqPezTWhMEZJbFpEr/vBQMID/mGLVJF9tuZEmlwc
AMVFCgdxb1zUSMnZB+H3oM5DYlf35qodTrZlIQrnAJavsLQGA2GrlvZzPTrQ5n1Ydm3zDvHPtZis
Sp4aXzDDVuiciXg9aeG3R1J6dfc+v6EXO6b9rIQuwHHCG1ZXCQ0JukGu2KxUvVBTrB5/TlDLPUCQ
mspz1jCvm8Fqnlqz14mBeaIwQxAJ1xUMfv3UkaKlCRh+u01qHoIpRcF37SccaVY57KXG3SRbE8Tm
Na4vybupF7qmEKhPZrrzNk8omDiEkgaa4ykFlX7sASLry5JRmBZNgrPpINuQbWczwkyxDXmbFVMi
eDX0G7+AgGarmPM5NwjSogeNV8j+xK/YVhb5ZJTBSd/Ex8PCpaK4uQGLcPNokLwLF/ji9ORsnEoP
zInrKPDICVy9hRrcB0+W1qEIldQfaSTkMjy4X0VBxIvMo24lRZVgpii2jhsWyQm0F23OMr4fKHja
etleBZnSADQ2ZMJViSfulvkIbedsLmLRC/BtmIMcNCYnHMkvl7WaPSPDFGpy/jGD5y6h49Z7MUOH
3AkktRELoNcfAyMN2xp7mrh53iTT9hYiR+fBXFEhuo2H5Uc4U3OYMBmTomKR92U0iHFaNAvboo3j
+FSID9Mt8GfJqI3sWoOFpmY5E1FXZIflU869V8vJU1IFqk1kDWP3SMZE/pXWrIaUf4Ix5Ts/5kvC
nINEsVLQABr5D0VD5rsyrSjTiCVpYhavh7D+jt1ozBwhhHEm7LEtIdPUfXD6IHZyQyRWydqdbdtS
waONixDYFr0QGO3W+NdhtFpiDsqvo7KRTdMdPub1pzpYFoW76oY77BCw5werWUApGaUHCW5syUT/
CoQI4AR7KirzC3LYCAezHBa8vgf9z66XyxY+yYowlddSCXRxyDNdtrgZ/74GNuRGrFbGEOwVhUwe
wEOzn+Lu+yYiUOM8y1J9DNxnkJDFt7BP4queTLWnYsYyTrKBbRO2As7pi1ovNNppP43QTJpFdYSe
VaSqbsAiPJ/98OArN+2niMl8VnjSi5cPXJ+2NNhYKCr6YjicqAZX2e/RJ8rpHbG3Ds4e3SdLjE43
V8fxJS9VXQyrOu1qUziPUO1F89nwnwdkDcqCXMDeesxoSfcJWwQBDk9IJDwAkGdTUPd+MaCnq5re
ax5uS55gMvH115Jy9JXRqrCm+pdMu0YbDZ1hA05DKhw9f8c2BTBAcayzeazEfsZmeKw17cN2rker
fjqV4/ZhyC+yRFYvF7/YbyTHUPfk+B1J6pEgbY3EM9YMiSGs0eqEoWcFK1R9fYDiZWBEulomcPJn
P2EC+YAP4wVEZIR9mWa75EHAsh/7TtRl7zi9ST4bx1/Q95N871GtSSHLDQcaZQTXUl7DhKeR9xSq
aiz2FI0qkvdxdEj+38GS2bhX+N1TZ6+kjNWk/eyeZ7C0dXYriFth5vhDqQGvlXDX4lbtTtAOiTCD
vqcPkiuV2vBzbIatENOor/LUD/2AR+uO/BqS7UJ2j5lT48L10Q/dMABQg3zXbOZFEiUwuo8IUUnK
SkNMIGv5C8gc01aYIrjAy2D3R29X/skdG4WMPB1G/rFrVsuHFE3hG/V+luSR5CWMx0AezVGYQyFl
zOUpo74Dgwq4wvezmraoyCJO5DLAsZ6jkzZYn4A0ZmG0VIQ6D/lrU5KPvxmRW1HiNsTQrDcIo+1h
yKf9kUgk1yr7VyY2F8L5XojMT28qNxjTiPy7aBM0tvSdhGrjO51BS7qWOYRtvqviIHs5A/qJy1Ek
TEXFaVoOLcmL0nCdm3xhMgwhpCvCKpQj+UIsoCDM2ESXsxX/IpIx4IaHZ57w4iXXfRJMuY29Kcqh
SSF422X5IDhTfrzIFozVCzBBaQcEtUuBFMIbH+wUsxU6RNrlpfiwh5vtgEHur4fqAp/kCzDoRWz5
ut8Bh6EJJ1obiF2kNi+oFZ05h6d14istHdK9jJZ+fG2+CpxR4CADlXt0pTzdERrFq0K4h5qt2hrE
s81UGe7zXsbQ1t8mVbRLjqU/yDPj/d50TXmKsc3ZvVfzmQTlVhUg7aXJ0rXoSc/W0XWtFhyLPT1p
cOrwk2xsGOK6XYsubomE9581nab5lSMk/MoCsUsEw5Hnr/eeDiXO3lrYswymUJ00tZ0zHPLHi837
WnQtD9j2nrmMTShYXWXeyZR14/uXSNuf0WrEkMpXoh4NuT5CJRXbtEjQcdk6DsyJb7sutvSacc5w
QK7UrtB30SvmVg3eQjKh23xe7+qo8I8l6k7Jnj0uAeHttYLHyqPkRF7d5z7pyudONXXdC73ks1MB
FRv93y5boCd2xf6w2vlHBNVszVnTqHqjM95h2oseaZL+euF7z0r7MBaqNc8dE1h380jRClekfyAt
5IjlnW2ivLoaKjeheMRyDPHEGvREEKGo8Hhyon4u7FQ6fZuXai6q+4Yuvgks7mHkf2AvTCgFtqh5
cIdO6db2QZR/mBMeypLfaRl2hpE4obpKTh/TarC5iwmygv56uBfv5LdVwHpLY6hzFLy87fRdM2s0
ofPpsvvWggdpDHSDU1e6Mn/0MdBmuntXrQiDxRBDezz2JzfufCE8DhZhg1R/8eJM7PN/39Vc2s/Q
zVJukp5/fYZaLMzlMTV81ZCEfWG9kESLblp2OE5Bk9iYqWHPgMfp9fE2SBpRnJZcNoos2HBKKxh7
CJpc/fKsilElIIwWp4OmelCTipReD1DnsbSkKJxAImq/8Kb1WMMRN+3FzD3ETY7HzPihFAXosDkw
2oXm3d4EASD+Jq0S2dKsw++3wTLgbKRfZ9GhYk+7Qj9/Nw7OwGA5CDYeAfdtEMjRRWK2FNQHtHoY
DJcKrEGHkweey1wgp6EHtLHoA80co6zgwgPQdPg0lw+3z5W8aPGL+RDXy5fhSN3fViERIu4mhiiQ
IYjXM/tkS47DvR59HMHUuP2U4YObwJkkxPHn0p+uNwDyS6GCV1VgfwyaWc3KfoFB0wUK9/SQuOav
KabAOVvKbi+gpSQmV4+3oYjjRXdQOBVNK/1+xPoJvLZU+eyPASlY2nHv2pG//Ipy8q/+IGlXNDU5
JWswkl6LtB/RM7S56k6iqOFo7qYfeo+ZlHrspnxCpLIhg7L1n38xmPFSB96zyIwOrolOSI0YSSRU
zdTTZEDLB7VQd5ovvzbiHqAszkIWLwhJi8GmsjfULOodl2nx8omYFDO5K9OjiVG6LMrUTy+E1LMY
5JCuR1oLRRgL8VRhPlbTYdoAsaqyZ0DIbGr5z8iMJl7B/GPBXzCPKWkMUROrysouNfPNXLUxnKlW
rWHSyo+Es3HAb0M8KZMEEsuJESI593i+zhnqZNlMhhbmSV/vL1IZxydc1BEvt7Qnkhwz59OkOia5
oEy2fWUK6ucSPj53N9TLINpo/f11kKwqB9Fw7fcHOAiY01bNP8m4kxXjlcbIHAx0M0yM5A/BHuwJ
dodgLaRRp4zLmI86XXkNxvmIWWINbAGs3TIHNfQyy1gQrciVQy8A/15e+dZB/d4ZmA6HPrliQ6O1
sdJwwqKpjKPKVd3+vhCyO9rsfCc+WKnQBEgMbs8/P/1IysL2tC7eT14pxlRg5E5kYno7t5uf7McU
m6fuSvNcSXI/JDexnq8P8YWitwzXcpubSl8RCRn6bA4WKmTuw+FzsD5Ws7dki6EQk/9/q031TqPn
Wv03CO4ay2xf0rIQaGkGhFStcvnphUxF+obrS7Db9QqC7HHSU7AAS94RBRGa8jKEVNYQeoO3Tfob
hdL6ZymjiEYUb7/obvtGTCrSlLIS1crmpJe8qzYbei51oSrBVlnf6oTEhgzgvKlhwTb4ovSvZA55
Y6umAyLE4WLJ3XGTv3Ailq7emuTHO7WuUuOm7/VwVFCv9XsyM11ehlb0IsqjaIchcIOLnhKtVTH4
hDIwxpeysXG54eecIyF7kXjmuy7LZullFa/OdWaeoAg/lenMfl1nYStOkkvPibRNd0/z8HWJ+hCO
v7MF1QgtHpEnkrJbZQ3e5oB3rDy+gNq5sYqcDZA1NgKq3OpjNxCjsPRUhHWGFTYJXXZiKcmxrGqd
gokDG8dzckmfPC9SnMJNF2tUWAEmo62nhPWPetzOrhapr4RifnHfJ96kkuqP7jOzh77/aOeDL0f5
UtpIUNBn+me0YTauIBlWuXd4AyM4agys9VlGIrPqrsZCjpUV23I6rm2oYgDxAEV1jp+gvajYI7EA
mJAirB6jgDOMdJ1buG304c8Gachy4S5hDvzk2fU+EMYbRFYbWK5IiuM3KgrinAqgomgbonij/3wo
w5ml4naO1yMUmcGDvJPD9RknN6ePogkxocMav5u5GMRo07uph718NJYwO/hcMf/3YknPFSu96j/f
fy6qzZxAv8zKzlIRnSMh3rG4D8x99h6V4ovcF6fwgDejD1WOK3Ig+YzaNzPhovcIt+bZ6No34Q0g
9F+lkFUI4xTW4QDeqRzvEtQHrT5OBexhhk9BMXY4xHQRKCItu8LxsvVGxgsVKNuD4RXoz2Lih3Fr
dFR6fBaFKnpJNXhmtuVNgNCJJVm7oFqAWj7hbW/Uq18VDMvmNux5o3QLJ0cDHXO6RO0CkrwzeMLs
WRnjbmFf9z6Bm00tatDDZ9ympy4BaTdNteXkLMBo2RYGEX1s357qDjAnBjrHZOk5h2I4yUy240/c
iNiOTEIp24JqJ1vLzsjHuC06k/SD48+LMFE/wenw1nJiSeJ37jKZHz74xnMpqM6+7r3NrPZF2tA9
Fv+xgABWF2gmh7dwH7eNbSXwWkzWi0dXD+mMMBy6G3sL3nRyT13uDaN/IscjYJeuc1xM22hAKVro
25VNuHDauMzw3k+BnbE9ni3mIi4In2ilN2wGgi/mhLlGBzRD4kLFSsYLIfz33E6L1fObQsbuMnNE
cxduukAh/GfOa71dJGyc1IzbMc0fCJZxcJ918QzxIbcjOBl+zvVhr3dwMUqU0Gf7u+xDGdlqAnY7
j4NNhm5kdFqoCu4OSBgyG+QwoEYyAMaUCzj1MnbROR+tK7iv32KBoO32ho3pU/jY6r12AXW12wHQ
DtjHP8tPoKvf5s57i6w5lMdPl/C2x7boJT3lFZA9lmhevLeHT8wVIz+jcFRwHiUGyxe7xh56y6IE
15D6ss4D3AdAeU2Jtdid2Qm6sBekPuao+5bKBe/EMdTmz6UAT+r3esQ/vnJTJq/OMOHRraR19ItJ
lfERu2ZVVEhyqi33PYio+gxdpW6wJodKlQ1yeFEpdkwzWFby4Mz0Mgb++6KFiVsUAY1ik0PQ58J2
inQk3sZfgMZFBRdZ8WkvWGKJHqp9bHdtxE9ZGQO8Lhk+jy3SjxgvFWW8gr+3bCujVqWLFd05GYyW
yh0cJ3TMcpWicwCVt6+GLDdSYrjpDfdC9ury0AYqNAH5YxzOE1Z17IOUE0Ai70RHdw/bgIWPWRVA
/By3lzKowXdTbvx2ZrH9Bn71eUyBGbHKNPbq2EVizCXKOpjF0USYXoXPHY2PsATCDk41qb8/bLK4
QEhdTrmY26hIhGbMcPxBPQ9f44gJ+39Ju00TBP/ifINBWLokNe7SMMhZp4QlGBxIdjFqGkmQEdPE
9Ngw0aLw6QyY7yj0QQAvmVr/k0dRDm5nOoJI+F2sDkkfeBo6TxRaVka28K5dWx3QyVWFgYt7Kc9U
FKTvKjvredJhBghpWLnfIhhDpU+7D50x0oB7+Pb3nzpEDThGQfNjIUbIzNI0cw62jV09omj8+xcj
0sQ1LHYQtrRwUbIE3IJ86p5Ck2mJUW1SwXy830Um0scUlb1AsfgFVVCNgL1HkmXnNW7lkzY8AqBx
zv+yDyjsdsvlR45zktZTRlJ30E3//oD/fomjBjBeGsRV60Cl7JgXWOa0p+HOYtZdpK2x1CWvXhg/
D8qgfy3rrNL384ceIrHLFACkaPKWbcKV4EWoekj0jeG97NFJge/Cky/a1DuyIAtfbX0grNThAZR2
bZUAWRmq8o1j2QV33aNLRkRvQ4Y8qVoVZUAK0NdYfoamya5LTLOg46AfMkB8UNg9JpiC9/iQxEYD
Ksrv1XWVR5MiNtVtScNTFHHKLrRsjY7gNNeXcOHViXVPUnmCOxZPmSrhnery1JDlYWwIKm2LZmVG
MkP058Rp0zS2NZcf3OHj5ySj1nUC7FfzPsmZjUmyQPtfYIh79jTLNUFnli3xcU04BCYPPiOQqYx1
XgLqfp6/SJRN6DZQUmjGSZ0pvVBbGv9OFi+3LmQ9H2MwZjnoWAYm8yh6S7/oljYfwNnz8yyaz2C9
BF2eK1zNTgFMLEHJ3F0IwLBKiPlzTSaxeL84fkjWJ/uHn87u8lCgiGnvIoqHcolaQ0Frl+d4jKNO
Qm13INaackfY0IEjx9jyFcu7lk6DLzVydhSQiQm1D+QBNtmzVG/dnqu1l78oIEyRlZ37u626Le+n
3D6FaaI6JEHJ5LjzdOlRTgPicYkm8BEn+voUuEfsIa4VzxIkG9Bom8JUnwbPEeFj0jHPBKSkzu6s
kpB5ibssV6kPVpoUMAIBhWgo4Sh/SYooyLO6dwQ3n327O3JFGLAomS5/2s8p2FD8mLR1KUatacGj
9h+SL8Tg6m4hkWngMSaz5NXoDhfyajSPcHSdidoBv5o316aY5NFGYswIqltPhEqHukZp+MScAYez
d1KHJkSs19WVwaovUtZbhQYI+o2tF4wRg19ZD4T1ubXyZ1HSQu8uz+dswTloVl6bUgWuvK2qkBzS
IkgWdQi8lCBxfdHHfHcX44fzFRna1D1J/Por/a7lAaJ2hVl3b7CUPAPBUiVQSGiYiKHnHslzWp5N
+v+xvlZPubwe12P/HpvNtYUs9mAM8gOLFREZafsUw7b19mDJbNKS17q9sFKhQjbN9FHzssq4paGL
9RFTdhrUc24Tf3Jswkx5qvtYtvvCnB9J2wqgQ8ThjBHl6YY+fzxgUhA4htMui5OhEh7dF7Oqt48u
milyhZTlqFvFYPSO0dTde8hJzPp8Lk7G5ZtXlZWHAr/RaYFTl8o3UnsKVjaFc+LJVQup3YkpvLgY
mGtmMNBXF7KAGMdNjiMe7o1wTtTmOpzDF7nAJOj5blgtf5JTBQFf9LsnaTuqrSfQIDwgTuZRML6M
uUEGyZ7/uEW5o1+RGMsDmpilQP/9SttlmXU3u9DrWkUgJGWVYWYQtLFV2v2zfvxpb9Y5sENrJzPi
0EkhKMw5q1WAUx8C7/HFOkkKIVYP3mzWJ2l8KYJWsqjIb+ExHmYmzga+4qg+l/Ls/waS0wMBNFzM
Gm+mtJVVKnJKPIFghFJxXOiNQnHVWRPLcpW9erAFVFycfCF6E0V6bH7gjWAVf57A6iTZnproqyso
ZMI2tDZ2g+A+kzC5uuw8gtmVtjTpGWD2MTmzW56KHvS7Ptr+t9kLWKO9IbtuH2sy7k0el9x2DhZV
5xuVL8Hr9R5luBOckfYlewjIZi5693p1FrqxBAdIa0xaYMzMutkpNE3LGLwX6gtil/vlLA/0RLm5
uavT9QJnMMUJrYqHX56EsaRjZpQW85DWlp0WtgG3DuSei8mrYRzGnGk9gv/cxMi0mbEiWLbNJY1V
5S2Em/0MSmUNeirD+ZYkXzs2c4f2v7RRlYFKXJcj/q2JBZQTA3+nIkzxNVxYp75avr2zprH/Z8dd
LsHVmMoXMpJqVaiKFb5KLreHxpI86ysqm1/inoYL/b3AJXhexUyzDpPpLPHQX1E1TGNpdr4uUyvS
pdPfQMJZ4Te7qLF70fP8dIdM4xIY4qNll9P4pzyGRACIKD7YFQ1Cp86Kc36CHdXvXb5J+MtXcIao
h9l6s1ecdFYX1gcFBOgzcvT63HYY79gupOYSjVUu45/4q0xsAwKvtJK9XaJ6mu/jfx1TxpCMjU6m
lMuD+PvcoL/U93R8IcECUZ3scK8wIc1kV+a2Hyy+c4t4owwVmfvIW5U1j2TnGpVs+3DMA6uPwPhu
bxPz5AjBXn9Gjprw7oQfWzojqMY8UbzXIJE2neoy0xGou9FLGj/FCJjxyAyMgXcYHnTDrB75hMlu
/HLWTIUBQn5r/5SuPC6+CRbkSlmHyJHO5nu8QJo9Qw3xXa9FQF9BkIFhzkLs6voS5sAqtJTdiXKv
Z+rtcqeR8Q0Lb6Y339MKo24zjHjqL7QAVhXimoBQ0ZfsFdbsUiZSSkGLKhnFTaTQXMeMy2mfq63R
mCTj4AquRUbzP/BMpgEYZFg3QZaqavWI0FTuo1NJbrbE4VhC5e6E0Mgd5BuVhmDUoywX0kE24Rli
lPSRlzhGbXbBPq3+UBIVp3Z1RU4fpRphVcEQ7A4+qazikIDn2zuGYRm/1RAbXI+LW+1XH65nAxJ8
q7YPF0QJWJt/wRJ87/Q64/asx90HOthw0M42m5f9rIHWFeuK2dnP/x5+L46noJWN9TkWNyYpDWGU
EvAVzXs8Mo09/3xcMPE71xXIHjC/8hDWHfQzZXQP7thGppSQjDiZhBIL4bWn6NNHaZ+0ghAw37No
Abv0ed7xQ0NtuIY20B/n8DQcF6lAidXOgUD5OTYWL4I5AunXJqFU1VMa/ffKNH9OOfG4jC0tx8Sr
LCsr+Dq+AEC+USIDQ4+CvLqxJZC1ciG2/GYQ4To8vmYDHq3SZ5ngnNQMzyENvMTOUfgkbncdH/kv
hAJn9iFJbpatR4zzmZPmdO6egr5qdm7nu5vgkIt/JIWOMYscKQtYWihKqFtvg5epScZ1jFIBrw9M
qHO9NuEnCv7zeubCaDBlakp01tC90mDdRTrRYzPWieo56chIJLcm6PkWfrtibsbsPqoBVVdHqSZo
LO72lkafNEeU2k3r2DxPMvsdz779/A+fFDoyJFlEUnzXjogp1xRKQCKYXRepmaPs1bvqauHCGGZP
9ziL3sK6yUw6M4GNSOIsJ/of+AzsT8m2jB4/bMwo65kPwVxUyVLeTKJMGyx8g0l3hdogqLpOHGWN
1NtwH8nFtMx1Fxom4317bpfhyW/4vVAWI+D+YALA6sX4DRSXw0mkmVQTlqhaBS2HKbEJtvdYCEVd
zmevBU+xUBcSmcmZ4GlsapCFdh2jgwW4RMWyNpygjKUsq7zw4Ynn6oURIF4/5NVidWR0divyRl/t
4Mckh74sFYnJqC+XXslFgGrjVOMr4yEuX51yvGT1S+Utdy0Q3TCOhEZPirv6YFZ6mMdpIek43Gkq
mIBxMmeSzPjbH3Ov6w8tIFva+GwYZgIoO8hOrh9KGrg6Y/wRfMWNdmTKHU4MIGvKfqqNdvxfYf4j
82v0G2sLxLQl6yz0aZ7ieX2uQ7Kn1CKMJ681fdPYBOsLbfKFnOVsbxgl0bV98ZJPAAdh+0o7PHoR
NwC9KXY13W6qeuuAEemDSN0n9hvnrsE4oWcOa30mDqemcKABmdQ12JiywuI8S7eQYQ4ia+eFUVL7
tqX9SJYovalbrmMreVKXmLxy5dZT7dMUrMb8Ak75Psmh50YMuqkyk0FF/NHO6gqbA6qMzk5y/P8+
XJ0s+D/wdS6Smcr/2cx/jhbi99cCdVJrkg0bPECBDz04cCm3DTpUboQCKQPOL16EkZydJU1EIBQ6
nuBIpjA/uZ3YMJjeNA24cQfCCWAYGYU5BWwk/wweHMCp9gBNr1U4rJxXNyjXcQcTN2uVMLG7jqog
MFMd92Dkjq0uPrds2kFQRceZJArCqYYKiT1KdNv5EgP1n6uQjt5XCIiS/exFkTJtyv5YbfLCh9aD
Ul5q5x0/gSQrppG9MVGIldDhAKPqgg3kHyNgR+PFu7E/tV/PRmGrEVX1qCLGVP+dsavZzLjhFczK
7oHWBBliytiISw2K/ort6bapR//0+9d9FyVg4x+nkcybqhn+T/z/pqwfDxQaXb10x2X1Mm+GPU31
s+K8S23gfeZJQCs8jm8R2jxJKk357nng1XI11Z9HItaZIc8qXGHreaVd1UMKAwt22vpsex0TiQPk
GW0ZnbBzc6shBbhSyW5CmShba25magBJrgIFxMU0eWW/mvSmoJVYLnZZeM62S/+93YunmUg46bLX
krr6tUlVJgQGTE7pN4dv18me3hWajbWblf8ozUNwAde2rFsNiTxBOjSKMaLcsnStN6zuTvlAKIJg
xXZmXUuL93lKigrP58+/HRJk0oA0/Kdds+wNn0DYqSFdJPYEwtYxmhvSR+kgqagXbm3EVR/g1btN
JgKVqnfRzN7yf0mCx35R02ieClZIXTQJV9YYrCXs+DRVTJYuwoxqDaXSiuyG1eRXtDSOXdHhiNe4
Cq6C8kBlTdyvRDPgUIY/LtigboUQuZ8RfOmCITXRqWBlO/1qsOvg8+X5CUGjL5nduwrUHfjkglMZ
3Dc3aNwptTRKFiNlZc48oAXL503edNWup+4exB3RK5tx275hEtjTN00K14u8iJcMhOTlUGxwgNh+
59U/YKdhfB8DKi5D5wZhhO4ZOFGfDqUq02M8xNjhY1yn6t+taQtSxGbN1GjaJrvfK8SKsYTiHiLe
YbchxKlWJIVXF/EuI/gb8PHU9gMgFvKJ0FRg6odwQQM/IP134lHo54XjFTpGI7osPybpaqlw+6Zo
yGuYs4VWBLJcFKOJ6VM15jy7gIVfYxFFSoDnLJl4PlNibdqcvs+f+VwKDiRPMBDf1xQqg9WDi3kx
MyyHD/DlbRsJv+wqdRA6o4dAVex3ZYaO3Gdh4etnk2chKdvNj6vsSOApT3LHe9xhH9VzYgeD6oXL
CYBf12QdtfD6oDUvrQBUTZcmkW3gj4Xjqrvq6MeHQBb2npD/wl829dM8K/B3VDgEMS5RCDrXgy1Y
0pNHoTFyv+od2sf/v8FPNsWKGK7kAYlOzPJ1VUARPrGddvolceQ8SNUU5Wiej9SAOPv7KnypPRX5
/xwIxc1N4z2NdbbeQxHZg+21B3dS7aghuCRetf7FGdJDjD9V/7NJ1cykPza5UbfU3NsPtc/MWo7Q
U+CUV0v4MTAb9rzmZVra4BqQtsDfwv3qqVRMcMJuGdLmhNMaSQ8uXAHC/UyEMGeJX1Mpn0AHSyE4
Pzltbsqe52IANaElOwqU/UTyAI9y6JCb/LPHDrnzbkRtBwEZEEquh68EusdiLVRi29LXbHeFyWcU
HLBnxMhxQcKXiULKy34smB03alPpBq2LviQGVJpI85hsfjGFDkStDGrgK72ctFYMNtFnnXigNuYU
kpfRmF4eJO+8JIMaYCAIuB2rqd90qccGJTnkFyUUglML+ThKStnQ5OHzwq+uW7i/u1HicLjzuX46
b+9Jlvp92ZBvs/ulkayLb7VbcImspQkTV06kd5C0a1u6IYsqGHjc3xYYN8vs6o6GGYP3kYmFkbaP
76M27UV72GJ59HEZG4MIDvtfRAOJKCSy8uvjZa4tuU+rjr6knYyKt1rScQRy91KNqr3pQhRzX6Mw
2spid+T5AXobOLUEB1B+GM7Ct7+po9i/jU7niA7EW7xe
`protect end_protected

