

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
g7azmhtm6FcP7uNFjuXJjN8Z6yccOPk3SSjzvKB27peFKmnPmQmov5+YTGwYqqN9LpdyiUExk8K6
vPnJqontvQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MFrqn2K0Cr7TmQ5al162oDGiY83d+AkTWOgFyXPYrTNznygR/tx44RAp24ytphNK9p6shs2EFMg/
Qqz0l8DCWiVEoJ/T8vMpnAn7Y+poGVGS1qAR3qE2njrl81VcGBZJeFaWIudhfr/DLTuuf2T/dWDU
YpelM3KbfYNPPiPy8PU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FZca5XZouG+/BYoQ8qrJTmnJanku4IprIWRkO6VciHehE5WehR0wsZJhfKlqLEeY1oTPA4bXaxmY
NjYkrop4EOwW8t47/hj2kFLI1OKUAE/TAhCGg/aNSOViUbB3dUomG/y+TBuDt9L6g0Arj1vb/5Pt
IChc5ZdEfRr1lJMTpFfP+5qmEH6lePPdzgPZATPB4Zrj0P6EyiEsU1FKBuAKd9iYNGiLCxVomaz0
3/RwK2Nl+/l4mc7PJt5Hso+4s1qHb4s2wD+OgbIwdH26ZkEnKVFpaLiuWQKu9uhDLGnsBMPf7XDE
p29f+mrvP9Zi/3nonA2aBKrTwR7XuH+ZYoakxA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jP68OjlYJglq3zpmKrXOhq7Sex8XNW8fQKp4hUNmuw06OOoKhQASNTnjtyVjAIk/VXb64ViBu1ds
cNMJybDSWBhnChfJq4h9PNybShGJXxSm3NDOo5wUHKf10Eti3fSotB9rVks+tNdTEZo4O97kgfdD
G1FNOqlsYcQiShEGLLiEQ2yYtgJBxJ+jc8mFjIEfPhAYy1ElrvtFEpnhkNS2LfE7xdWOQdO/XoKK
ibeY08pgncTI3pvO6TMbXushf0AX2S7hgfk8ysZrT+0gktqFrJnyR6oljS6VVPLtRNW2vo/cC8XQ
Bzvwwt4cpSo5KLS4XxB6qClZipItck2AUEdIbQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o7jAZIoXlFbFtDYmtXhfRBlb07dhBb6Wp03mlT4T0FXtvccSHWhWZgc+VUNwt6TohLihOwvSipPP
XVXpGL4pUVYNdQBCVpFzhMkt6jhyUgsF5t10yI5Of6YEfQrDHigceoBukM3+/zJHPprrPQE6FUvC
wXSGhBCXnHJs1R+n4l0714w8/WftPQhlD9QGQp1qT2VARQXUKBRxcRjxe9TcLfs0P4xnN7uHu0R6
JTmV+MHmhGpetSZGx+B2Wa1MQofUPURqwE70IwBoUhdXH8+39DT5I6x2+wMY6RcVATnhNd2BCgPd
RzAhwfrcqRiU9aB+eNNdFR8ve9M2nGMmV2JxZg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Cl1Dz+fZIDYEIQuUd0pSg+5jknmtX/JERd+yOZ2SRaVra/4pU/eCTjEXMzhz4VFGYB6dgUxMsGBk
nL2WNdn/uaSPpi6mNF0UHQvZik4pUkYPrnRbFveVqW8i1t95SG0RW96uD19206lWrp5U1lqc4fH7
sfKHi8ZpU3MAg0DOO0E=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Qqp76m2aV9ue8Qai7QUavb+lhRYdu/txrnwYLzwTe0vS0S2OD1vxr8VeIT3bF/ZuXlTGm4S/UCSF
bgOPp7VqEOeGNfsSPK+VpQ+foQMENCQYccwKquBDSg/sLjpPK9uuoGLBLxjw2OwsRzplVFXiPcRN
LYK1/FmCP7RJBNgmhh/ti99a+WSl6i2YIIRGocNplQlG8FXq8ZTTHd/x2Gtdf/zGvJOy/fNsos6S
Oq9yJ0rMmbGeWbri5c04gZM08pUmXBsivgOHm2IVEZZFM4SBqrsi0xa52hs2kelc3iKJcWiTvU3X
0fJP9qNFuIjXBPPZvEYwhVtIh6DwiIC2viSscQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967856)
`protect data_block
XpVvygUlf+E2sQx3D/s3JmPbLunAglSuMdiX6YqSeQL+KaT2T53TYbSD1XYoYm1kTBymEKfIWuj5
3W6rB3Or5dlDEUtEN4PO2JcSDvDz+iWho/gZgyBHWAE20b1QOiUPUqdT9YAlnrfewjbUb6ah/vL7
RdGg1B5nLvtlttZi3dTpze4SNpnb7iv8Fb+ZnXhT+H7GvEP7D+WP3qOMNg/Hr+9N8L13Y++OhFDw
5vgY3G2d0m7asZ95oFlWKvPuK1WrKhCmeL8iJWewEWIXybTgLBFtMWXIcpak3SW2KB2cSIa7FxX5
yZw39+ruuy6U1ohtiG57U0n/C89YoIxHJbb3Y9jmVXLePxpR5puHD8fM/2xU89xJX7InLA5svicD
Vc/V2i8xuDQMtHfidYQwr1PGke9/x7nZmlT7irQFYQSAPc4KXatLJkAYEO1OF182eC3Xfft2nNYU
oBUai0X220NHcnk/SZFpxlMx978UZGohnf+PlJ46qlaMoF/MKeSj/gWo4bOBqIglbjCQHTSyeRGT
8Ib7FiuFR6xWjUoiBAfPaD20f/r81XwRgypEx2Rjty6D32oyYpZJc9nqmiEAL7X6MuQA4faUkWXn
mb4D+jBOH+3V1l29C7RWLPnrN/Las2Zav/LOSVodHPHKpYyeyeREk32C4FKRuYdUEUieYFKB/lX2
QTtENZKok0DK+o+IAl5Gm00PjVFSBl4LF+AJpAhwNVFzya4XPAc+xNKt6TlIMmyd2meS5HO1tFuN
Bj4cbybyggfydytCk9HCsNfNDCjaf/qvTYqeajcnFuxBh/Ruhc/i1a3SHGElmDoH0uXhnbLjRhwv
9Fjaj6cbDiQj29NXqsCScR6wF2fB9atc+kWp4X1YyA7huOTYN/52xwStcTfvsEya/OQW01Z00CWv
eQ9yqnzAFz9OqkCW7qDWqSzs+D2bsBzAQemFacQmJn8HJfWWliB/d7rI8RfdDACthrtaivf472Tg
Phu68zFGZS41NwTX+Phie9fSJwKpbC0meG95BXqPkR1d5pSme/N6lPDVaefw8wycGGQOKxaDTeTa
QmjSaR+BhaWXeZZHB6DpJKqp9LaN1cvD9ZNgDVf8KH6V9w/1XLE5EcRroZ+Cpe+LYj5G50aLYg5/
W64/ACONHI/GRL3NECpN8mlg1Vcuv55RC0cUGJokbP3n1XzzI3hZktLhZ2FNPhr115HMd2zrLJL/
gsMqCx3YgWKtWB50lG6wPGZxkcGRLuDiaBQa8URRWTkBzs9/ssl86mg/KDzzGboTemUTPV2Bb932
dgqnVZ6DdzCCQLnWt2uTOXPeIgdWSswTcoNKhvopjcqKRyHMVNecVXX6AAmFOOK8zdO972h93NdV
04kziYuOddOkS/6VblpxFeh+lSho0XglYR/AKzu3mWH/C//7vx/DskrcQ00/hC02P7mIZs149gJJ
4Px7W8asSDw4uJ+OuQvHPAE0e6xvlnQPp8kj7tUcsr47R1imCnjMTNZcpuiUJQgofzOBzCdtak78
onwqrfTMrv1jf975fo2JpH37UWJ9H+IRQXdN262qR+mUd/UG2ceWTQgtJ08D9ro2/nQ/gYhPX4gy
kHeZ1D+DwEzgGLh0b5HUL3QpYzOupgvR/N1MVC5nQyM6KbDMDymBNzZu4eGSV/4HK0jzBMCpdj77
WviPN+eqbNPZMmLb0auk/rtOW46aXKZeWYb0fWXvyx8DHCTAb8n73VOSH5RjTaBNjg95dp02KAFY
APgjkB1CLmTW3guW7a6N7bpWEzkKS+YfpCIoNX/wyIdy/DNNLhlW1lU7sDm+hDxtjyj1sn/Clz25
Bi+bqSCq0dlPM96GeghMBmcDBraGGUViezSRFs1waKLCje81cq8/Rxn5ml5JMWUUoOpoQ9kP0rmH
g1OQgnF6n7ZTs2v3u1hkZBSbTFx7wrzr1M0Cn1l+ZVjrfWUFRJmologXSpIxgefUNg8HLXaaSZJL
FzynWV0uTvhffCtXU2hTmLI2coxsEmx3AGSUn7ntNO+C+N+bu0qsuXYGKOQeWImrdc76y9uhTmpe
RPuAYAyz/z9HeJDj/pnj0h2LsnYQpF4Lkyz7e1x2V0IbO6Cv6bjA4Hj1K9z936KKT523a2t3EZZa
mQkJvXpc6GDFJ2ajSQkPMx38tHtIFqz42dm4o2cxBh4QysJNIt/lRQS0ULY1awpd8U8/eFCsqBtq
fOxcLUPbNcRjvFv/4kW6MmG+5qtEgDgr7NdjKWfWNXe+sCjcYL/ax+uUUTqyFC9PR+OEsaHK99gf
5w+dWoWGBZzrFlPpJCoUvDqVjgNIOSE22sWFp1/skWxXeKshU5AnV5USXJwaXZPCzKItb5xzVP7c
0gnlxdvcTA17beZYi+tLH8Kh/qOO4hoL0uG1brwKvoVRkCycOLFZerQqqglSfJIbtPvL5+x5trJ5
ujT7bJckixytr6PHf36DJU1IQcH4gZz43byIwYoawiHWWWcp5G/WfCkNPKvIjls4c4Z/IC2t3uXD
21ei0abk9Fw9nLed6hsgvJHJfylZ5Kmyla5Fug8ySZu8S2f8/ZBn5vJqK0nJjgfPSvR7MQPeeKW1
5ygD0fXiymIgHyrABx1igM0BU7eI8rVWkPWHioqLfoyqEg2OX9Z+daFkA9Eeoxpnp6LMnjzxieDQ
VgDLFa+LIIG2MYJqj3AteY+i5WuoOEUQDx/FGNNI/tkDcq1nZzrRQw8TM0EmvH0OM9lVzUGx4Rgw
VwCOxVC3BXoP9A3Pf9PtkOYNlmQs9qR109ABd3PFs6BferXd/8LuvlJUTn/gfC2Z892KJgHF5kup
Kg8fF+5Gcj4gKJVHvswo8I3oiSFY8XBJgarhb8MdYkYJvWiaTtT/VbAPANiDXcTwi/1V+9kJ9AUx
agkDCzcL7mjLpO54DHObG1Q0gGMG8aFTd+c5HbRWCQ9E7WHFo1DxfP1Q9gRy/VnvxRA8QR9RSJtE
XdDCzmjYhr1saQdD4zAnu42xyEqIP9bzT1MRDepfBrHX31lEqOZvhEuwHbabKAhxhBFm0Su5jGYc
idGgeUBLtVLBRetnlj8/DD1ikODhrN5AXdieqthbPBGkibF+Tn1iTnb725TWzQ5oDf50gpIFtoFF
Pj7Zo6pxW+dq/SrI+bDhtJUlEU3Le6KvpWhZb4+vNIPsKvUuTCnm7I9hlZhW1YN3UZn14ZIWENuE
SWYhoRmMlYytzjympGIVoGVbNn2x8EU8sHbDdZxnmz2HqZlvBbP8HzxSHY8BFMvAdWbObAX/PcPN
8lqGySwJ8p/RVz3rvNiuKmojhAEk3VcFLt6go2PBXRW+so9/8D07zWqi5urW4SLSDWVteIeodnEc
rHNpJW9NCUg1ULgQkbf4m0fYdSbobk62GBJdkUNTfWi2dVMnYAl6a836aV/ovE5GlwVeneLylMjf
tg3vefTHdBY6+MmNoGTi+CR9q630kcvB0TbOfqVCM8bnD6wOuSzMEziZsU8rvsCXzIBwjcu5/YFH
5XeJmqYoi2E2XPUo00trSwYe7D5e0J70JM66PTy5THB3+CzApG+Gdx9v2Ki1ZVOmaZYny7io6NFA
oOGCMF/Uy1HUUWzBIzTuc04MZbE2sAUYRpB6i+aFcmNib94XH2sdIkqvs9ABT5EQYldDEMZONFIU
iny+OC1r1FfjZExgP94QKCfqFBwID6SeGmKUfzVKQb3N0eG5eTBxsIgdoJg99S61+hSxma0pxC1U
Sw9fTA/QI80XPp2E9OVE/nJ8b8TAOlY5bKUM13DOdHlA9m1TqkK9MWWlWb5aRHIoy83U/6a0FWJ7
guIVQQNb1ddbvQFB0lgvVuFjIZS63FIETpKZTY2oWDoiKIETae+rzWNSb9FC/H4Sx3yQ3mrzlB/Z
+yiiw0PjwxNBnuAR/lYNnUUWrownXlQizaBk0d0MkqTqsmhzu4+Pr1SBzG6GQYoF0Jv+GY43FpFC
x5V9O0jwrEmha3Yzg96Fs9SS3bOA8TK4cFXHwzh2bxpwSB1sOdWnak8krrhoKSNPjQjAmZqTHu9v
uaoFA8glKhaDp4BptPnrMSlxIegmfKV5t5pFxWwmhvJHUfq7U8/PXJWEEFMIvyGPlXmZ9bV6DyRJ
tRvLIXmYDiU3XbWTwWFc3vSWF38aPVXXp7R9APnG1ZFJyrle4rxuI4i3xVvw1GY+la/pScXCKsXz
X7PX8X9tpZ7sR0BW9uc0ocmO9YIly4JqZyFE7dcILJ9GbmFtTTQnE4vstayh4XeZVAjzYsmAZ5C+
qw+JVF9quhSlVQB7eReOZ/xL93PXfR24ZWKwUR4iH8OiP2LUqvJgGEMxmnRJeXUTNpZ+egkB+upA
XgqFtw4oyfQ9pqbjDHrlAS1nTa33P5aN9HidTw5Zr0m+iGa1173sch5sh4fX9Y1SVZuHMrH5rJQ7
740tVKiU+dV6+0P4nsEpUCQxn2PNrEtFeQwFF9CDmk/+zd0JrzPEFXGvjvAFPksPp12CJ5K4L9ig
T9lFJ64l1nZS/GpQqyLJca530/IqqKmKwtFrxhF382m92NpJ3scVTjfQQUpvXTvkyrteivnNwTAp
0g0HMNaMnjfZkW0r1ph8FkPHmK3y54RsekmOY2PnmIkoPKNokZfTXqucpv0y7jhgRObL5ia5OSmR
eEXrWflq4x0V+7KtWE/RgUVz66uUeFKYr/nUharQoD2+EeHnbzX5ZCx3FsHpwWG4Wh2f0n6dP24N
YS25x0MOgYcWlvWsB6C/VWvDh4+MBqridqt2xu0N0Lc131892K3How6WQfHL8Fayh0kb03UQwdDd
NVZjKlqH6ZKU2M0BASO3d+EQHA9nnYbYrDyU6ts7iVirwOl6pT4d96OD6Wq7Bh7bi1wzgGKgfZBx
JIx5u/DfiMo72HhfxJ0kBCbSprLJ9pTfc6FoshtSMx7+zznoWRgrwEDHfmoUkq6nc/BLiS8vwMXR
Qnrjl4uz/WD4J2J1wM84tcJpy6DF2MOKYofo95G2oA7OUC8ea2r/fQ9QRMS5o15nToAPHP8Rj32W
oa8tzrVMZQiw6YQrhksH4xMq97jbEP9adNFg+TYE+BOKUkPtxRpttgHW3rhYpvqpbpSOb8Oy+4g4
aFp7XwcVCopVvekiKgAlu0AzbfcUQZc8mTNu9aURo8s3rg2608TPuBtFK0mcle4TFXP1jolUhOQq
dyV4Bgqs6tvXY+xMKqmCf2JLNz8rVupwWO49XwS2tie9kGfhnYVW4KxvcDY++O2fDQFD/+8J7/2K
XQ7cPa+Hx61jkhIiQPaQEYJQjjKw2AFgxDLmVaseXKwr8a6Jbu5cyp4iUzF788cy9oI/rrBqwt89
qhe+/AF5xJG3v9CafddqkJmWp3ARq57vBnDnM/PI3xwOYgJWND4w2ralSFiirJxW7Tf80Ju/1slK
VKEMmBq+wS5oN8utH8VjqFV7qiiaAEHFuDTzVqfk/hMcqbLhwsWQLrbKpNxQiWfDwrbLrN+4qZJD
DkIQ1Wkf0HJKl0cnQDmGT74QylbXojWgxx+WyHR0XeJMVQcmLUDi3bw4la7QqQ12ny6mky48H8Gy
frKgK3cdhrFu6Vvu44Tmu9pJoLO/usA38CaAmw5tSMvXgWbsgMdxsFmBeHevnn+557JsjZqp9g0U
XBU8+ZTmQWhhIwzA/q1AgxEXTUXvfmj7imXEX2iMTDnFKldlhOWwXYbAO0Eb3D5zJz73sCCKptXE
5cEKJCac/y0XByqtZmJQD3dnGPweJfXLbC0W30fEe8/Q2dc+/myawDNKsgBnpg7kS8ON0N/MAnYy
mXjGVlaPA+UsHw/9nbcE6QdFJDNoYJHS4i/uohMHTbAVXXffNjyoIYQ74Sree6glVdyuziYUW2Fn
4gI4WY7x2m/hsx+iC1keu2dnKtiYBqmhRLDbyf9RDp2sjXocPTj/Zspk1nm3LF9b0YReINioSYeS
ToawAeGYIS6SyVhwKwRCjh2d1Y7sg6eBWQ6TvPl7Rg50TMe12rAH2LKdjUjmOliuraweCEPof0hD
DuzT3s+z7dnFbMy6O/82qVaHvts3Kfw6pcixTsQmJEjpdmjKtQgGmdO0/n30o71f2hX6WMBG/GEg
Q6CTXGTcyVsq3+k8/Sv65AVwcylQBsXcW6zR5UrumvZZwckKn0jGFrEUtnF59j9wujBjTpgrwQ7R
JKSL4D/SG6xhJS3vNMAUNeV0j+oUfDJUZ16M9q1Igq6qdtrInsihxTVDoOMoWQlidbxkxAmVMFmw
0oJvOQ4a79UJj2kZTH3jKZIp4VIQdnOF0Hiwc+Exu3o+sWp6L8dKd5TXnGBUgbrlTKe+7aJa11GZ
a6DFDa+C6ON3SKia5GyIDqcKnZfoIn6N2GabDz+CaIqaBHWjhjEmtZ48MMVN0hTJlymCpVMhBBj5
NtimcWiasjdsnSBFbBnfP/YUGf+SENkFwed2vrAW2CjC7QBTahGqmxKGUHhgUjpUaLFcUrkJ3QlH
QhxmdepSiKCjM3edfI8KLrbOUHxsChlFoHsvvc1Mn112F/MzVRg4ezC9VsKTGUv4XX1t0MAzlIwk
le5Z2tn5NvSYdSHy+e/Yyx0ImU6WZiwm+aPdKzBTOdPDadxAr/rJ7zWLZ6pCgxvHdPknSa89TI9w
ugJRs5rI7reDS0r/3PEANg8riMYwbStPOzyEELbEY6jkuDCzLrNOHgW/3qY9dIQy4imGOmlfxMFU
NXWogsiVgarrsOM9yevTz7Zqs+Lutm0bohq0u7nAI/SS3djGbAEs1uerJx41ARruZDL2KqW81umR
pYB7d5IQd3SsBb21TjVzkpo+upsMEuxgpCjBGdoMZbThbFNDAUEfQCiHEUiyT8Tkpo8CpjHv3MWZ
ItONHBPcUYTjr2wIOFffxKGRJ7RUwO/wiBIJCSd7R+xiiqe8/wqYUvG8anK0IM6XDBHVAkEp9ayb
6jYshPRwBwDOmEFPZ8D2dkm2A6SiC5xzoAZ1rztXbWPMS1BZdl1BbifBY29Db0K854jwVkyJDNND
Uk6XR4SHRMUGK94TPTJ9hHiLQ0MxeIlFu2XINh0SlbxsrmM0keqJshcBtRgzbF3vjXYXO4k1tp22
YdabeH8mfpwEcPtHzccuzOICy34j4I+zucUQesa94NUAsw+OkLYNGJnaHEDgXzvYiUPIorqtUJEI
tmCWQkIMVWZynftHOPWfQs7rK6blE6TP62kbz5GiX6AZiJ3os4IfS0FystL8+HBNA7lGKZuIKlQh
2dzqp06Dak1cJbkwV6eOWLWSUSTRiB41nJmGZYc/BfX7ynROji6/vAMEMauW8DrpHrylOnH9yPEI
jvrqoL2BlmIkJEN+9l4uRIJ9BzOffdhWJlmCVe2ifquWAaqeWga8eMgIHIOkiyyFm9m4R69edM9q
phmrPUDYegKdaGk5B2AwQcZKcuL0lqYAXcNbSBhR8A0y+739IY84FexXi1doze9vuDM1Mfvewrrq
RSd3W+RPtauUEOFwV7HXsOE3dIsK740fFsYcJiToepAI+FJy29EaKV9keSkb4r4WXyboFFVZb9GY
vVHWeEIurSJ7SQqHY9dsypvGNSxSLQWgP1DmrdXuKrtAHwm7bo8hm7mbsDQWnHt0LYN/TnceKJSL
xUe8inRRZn34OT2V2eyq8gBlNKGPEDgdiidF0Gxu0EiiGVAX19wzbG6YPR93Djr7Y6H6PC8kwtUs
elCh56yWMKMjlhlMIndD37z3arpjHL1yFNdV3LWoYzZu/jP9zclF4NZjJg2AyzqtouaH+G07FLSm
w/bEgdYGQCVAqJ3q7loG+einpt1a6nRMAb9K0/+t4R50M3Xai5HiEH2x0G86+FzzwQB3GLVefj9x
nKqJjLue/dTtBNQ0zcE1YQyt+r2EKUJA59BzQOvwavbZ/7XR3mvu7+JgLeer/c7O3BjzAyuubx+D
Ir/OrQCn0GfHF/yBNfE4JEzkzG0vZdhJRtZM9lgbDbTp9K0ZLqBQlnKfQ7ifEwANMkDL5tLUj334
rtSq/WCQW80cwi5iyRBMDDwlWYyNs+0yNcq7U43FvRcIGjg2/aUx9OD47A0wcyipi3dZT1MXyRHm
PFK+3IFvFStV7JMIGeTJgBezDVG9atrRLaJ9PpQMkLXHVKGPPltTieNsI29B7QFy+qsFWwPE/LEg
8ZbYLLEH88A5/ubQQhUDvnSUK9IVnI2TGMFIGxT+KV/Ma1yTKsiQQnMYTJletgm0E6dALWeggBUC
yqFGZhdl8xNscYchPQGvJef8RC2JUzEOOKL70M33Tk3aJ0pHTFY/gj4lA5HCwrx2aGdFO25hKuRr
91vaOWSwSuK8/pa6eNsA0SPCb27JxEaRp3Dj4V3OpRzfoZnfTiJPkE1S7m7anc1GoPg1u6iRuw0L
PgzEJI9MVsai/iTbpyfKp1y4per89wpes0ep5TIUk5w7AjZaaema/k3yWKoITZrmjrbEMPUMeR25
VJnmOTv0OxPcsr9O2kg3g0rLACW0B3Isqx6p7qvaoDIYCudOysVfeoQMYcoUhIv7bKlpjmqjfqXD
1oPOR+DeeZNNLe5eovhD4pc9eIjdZOXklCd+NE8pTWGasso6XXcypfYBbE+tA019KEYg43Wqg+RB
cBXjqwyjwWNfwMa6EhGgGH3S1BUki9NOmr3e7KzIa+rJYOt3f1RNwBI0f42P9kmd8FGPoqvtzOpR
f8JH9sdVsfBkIWnYRSvV86UNtN6m8d7LTDq9QojacAiRCqRTsNIs5pxLxqEtTw3z2xVr8IqXMbw9
8ES5dYopo+ufM8qDdALYPC7iAr4KxvxHwt9Wmy4uprx0lILK73SBLuTNNkLBU8pcQhNqR0iY1AVs
JV1Q1YBTNr4CQH6UC+GVyisS3AvyIkL0vn25MXcHnIlkF3HhvupvjN7/pRvK/8pq9h8aQfXiXLHD
+83iSQY/QbX9/v4ZkM/dvm7Q/GNLY6KmW7bTib32oD2eP8CetOVwOG6LFwTURqQTtb0y4SEQJZ0h
pKr5BYmDRaSdr2ye1Ebybl6REqFlh7ODOmt/k8Bw2cSR7277Xx62maCbcyEKHiqFsUGt4fuvztWT
9sHiwNVmj/cLfWSdc5DQN5ERga5M2thRO0g7pXJiZSUMZIfT8O7EPKNd0vJG19TIFtdH1WQWV9bf
43snhQUP3SbWaa8UIwxIh/wE2G5OBtxyjb2521dY7lsiOnDt5W8HnRFz5NcU3k8wN8OAZxg0v6v9
D4mtv1/faWLpthH99dQDeDeJ9I0/2KqXAgBGEjWCqu69ts1COxje5p9ysx4lDXsIL3nv4AKDC0aG
Vth2aSHW4uS6B1vVXhXjydt6Telgp0sWNOtx+b2wjy0nmJOHnYBoaAKqq1U7bmyOcUWJE+Sgnm2q
ibO9K+RwouH0tNzgc7lQy51pIiFPNFQkR/8aoMFUyjvx1J+lJKv1/kFc2oDARSl3S21AIErweRro
dQiVUZrfBCfxExd5llmT9XOIVSU0VhHKaSoKlX1RMFe6ADRxHQCT9JnI9NBeG7pix9FlHqMba/6p
lSSs2PqKWM+T++GEz3donvcp/FZnPrHGc267InfNQU3RWuzcONwmKXwXzNh+2A7u1eOayFwKm6bG
G5gWAEOmo+PydAGBweZYumvVODff1fFWmJuk9DtGse/PsMHJpZ8DTILnuf6d4cIHMysYum/ce+PN
N1+fTCP0anGtzd1gC7PfHZBTmifEG2MT0dOG20B9DMtrH5k0A6y/6LBSSIfP7anRoRycKRRvXYBN
/u7X+8mInjw+6SS5GP1L42VjmkR+WgfUnL3cZihnqS1MJOVOXcFVkDgXXKAjzcHReBgG/zNSPVyY
WNdswuhMTyCLRVBwzTopYZ9Nb49lfXmjt6moGfoOfhLA82TykbIcAEzt7iqwdjVJQ7vUdCwybZFf
AUMnmegsIJcJvp9vW4cfedfrbWb7w/RYmGIldS3cX70TylPSNFx7cCdACBe8Uf/2qHkUaGI7CRn4
bWxs+dQYp57rjAjwkMj8pNfT3XTYVkoUMV8tjN+9vCV9oZbIWkCD5O/qavR/hcvrM/hJdfL3jp0g
hO66FOXpt0ap5wYXDykBxiHr20hi8cUs0JwdLVJpRSQbe5csPRsgfnY2b67Z0NPyUcLWNejUjPDU
H8GZ5hEwvjFetQYSoN2c8FbMpg79vz4SOKgzwArY1NJgoXosIneE9WAWvZ+qMMQhGkShW6F7jTpp
DMKRM2vV5GETK0EDjUkJh6sDDlJe+7qdJBhyppmag2099QiqHXhfpF/BSkA8miY5TqWQItazNnnw
6zp9E5ix3YvDChFsSuzP4yoQDJwYj2Stk0vrlmmqQjPlgqkvbNEH7D030D/pVn8+d/GpBXEl7nS8
XSXSTRCAP1Du+D/GNuWdfPXcYppFId9nui3k2hsuV8F/hQjKeurCH11+CjIPirUoMfNT1dEXy0KC
Xc92yxw7b5yTtt+rwG6/NCNDBkQsCYWQLYHViRvcRG6abUolXnZ9h8l1WaWTveeWmp7/5P8guNfn
7aJqE7SH+2zhiSG2GmYGilQIcHEmafM4JOQWRzw5dhIQrDfFpvWm9Edi9o8tgu5Ww9RbYTJulP+S
i7jYZwyhC7qtzy1TiBjaruxHzX3yLt4jAdvQiodfArfE8Z8K8aqAgblh7wvo1Tu/5Csuu4cP6f25
RaL3SPxG2OADCPKXI1hboI1wRralwe8b0PBI1is/8kl8b1iKV5260B1NRKYmdtM9xe/ACcImOah0
fcAEQ7fsEdhRVbzi319SNRzeIXaWMFEw27cyWcAng9KzuXews7ibrd+bPKzqMtp4O0nJnMx6NR+Q
F8LeKF7W7ClqgR4/sGn5Ethw0xRwMvYYtovCN1KlbeE0UTUFffLjrwsnwAvVdlRZ0cUxMguBuABf
ACcs8wFv4+MPpWjMrYiE0E+6gL9BjNUzN7MOthoS83FrkC5GKnaVcUAuDvtvzfmJirAVdfI08XlK
t4OtkqQGe/bUzcRNCg2Eeo88Yf+qXRZDBBGKxPiRzIV9LGhZz4MKffo7wYhFq8UiGKKuQdX0T5uN
A7VphLLqbido4z048kDLPDD+97ieiBJFfI09+CAur9j0YPeCBHrwZLu2qVbu+g27rG3xCy4tQ6iA
8Mnp5+9k1cgjf9b+bW7e2Vh6cd2WJI2x7TrUTQf2/+uIYHdaEayZC4gowoIXwE08ppHwJTllAxQD
XxU77HDs2aMJEBwif+qB0juTkD/TCjl+Y5RolHf8o3n9U4yrbs9UhoiY7AoCz3Srtns9KYxSdExx
DbHls3KE9D1WRMQRmsNTCR2DMLMcJZYMF/fF7O9J01QpXQeGz2oOyNtB8yIcac/VeNnRe87KSACW
WCUjxd09GDtXIIUHuffrddfBv3KN4ejlogjj1d8t2nia0gwHZN7l7o6HdJXmkms9TXPGXHmvVigq
6fC34skR9Jqk5kaFHrwwCPELBv/1QBExLAoK8RLKjKtbVSIqcugRvWCEFiEN3tQygSts5AMTNXnF
OvPXMLOF6b3iPx09rripelElZ43jWuvyl5OEuyoVY62i8IcqKR23bkfqGidvTXT3uLKYsXQIfQ1m
zqLD4TdX3FWNrfkUxP8pneXXjP2hzfhYTZ3XmaO/EtE9gI3BL7fhmjgoJOnCO2gkastVxXsJJ5rm
p1/AdxAHxvswiIuxXacaZu+bAphNKRHKFxBZXxKWJwZDstUef3nj1rwsxWI7QoRoPuTjyhMAh1J5
fi6ECRT9ScvbeKX8Ym86Vq02mdcbPdTby1WO3sVhnCNHfob4ZVtk67E5n0dN6EeXCHUQkqSYqULo
tTclGTLJWa/BrmVYgFRycCDP9Wseahnlg4IaNkGUvG/RW1QTEqUYFQSkLxWuBKzQwCTTFCecg5bV
ZWEDkvBVkJ3roasmjl7D+zrajRwVKozn82jYUPdxK+flN9OIPvRnQ2po1nYrGzEF1QZU9fQaELdp
aS6TbGfauNsmVE7J0EEyEqbAHe7f2DtrEmiDo6+HTm6BOjxxqA8GfOXebi7G98MKrDMdiHR9EL1C
mEAtPUCe6z9bI5ZT/L+Er/U2XLBpaRZvbGse5ZUcIz6iV9iBGBjc9TwLdRGoMYm71mlCccaTGyWp
yFSA0HIFroIuk0OuHApiTOteL6ql60vRSwCkxOQ2yy/ZVHqhSE6+sxtCvDbZCuWOnkZNHsfntT9q
Fv+TWTD7dNQGBuFkgUhF5DwWfmVbeRxaKbTvyYtGV6nBS5srhvlUXowH+kRaKJMzXbp3xzBCMu4v
3J9d5qNndZJKK7qsshuafSdEscit5c4vvkOpg2vC3TTX8TiNkrNngW065pqTReN2DFGO+Wi2FRb+
tvZo3y1So/MFaeJYtUp+3NSh3iS5B4SJFhDY5jjw2O5jr3zVzOlVire9YgLrGvCWOf0gVAgHEQYH
NQ+aQxxJ/yU6Kd8jdpPcTNAvB4dDRjEF/CaFNhI0TunER54iDhjFC4fCg0gh+FMaZjtPEXO8l4h4
tyXDp4g8SCE2+sUQe9XdaNXTOvJs/W+FbJVexzgmeGuVObMn3RjNaTodV3r67LecS+CbUI//Oslv
RjK98l8BaoVLXxUDY7eDKrWZVDfXBePZNZcMw+iz0G+36FO+ckxymKMKn/Dbq6oBNGMcPOgD9gkJ
7iF1ymjaJITKyLHB4cNTiRReBb88BMDM2yfVOJeP1khfKppEbdhEQlUTw545zocTU30D/QPzeDtD
6gRRxG2xnU+Cs9KFgcTZjwVDyIpzn3glGGuKELJrEJj0a97PuCptPugGBxn7AURSEn3LvMTqEZeq
iO0ILL1gYzZ01CAr61Soo8ZqpvhQpvuks2eNFVcLgjdNRcUj7fvlbNVvPLwZ/sw+Zxd2I3Q1aVEI
oMbgwSj+6wJuXIIWt1mWYO1z54Xgv4wuETlHYXaGcklXplQMxSoLXkZk2csuNxMsWJUk4IWvfqbN
W+ePlHQyorsp1yilXQpXiTRQL0Z7c7N9lSeNRa37ZmJdf7LYXI7vVYhP7phD5XKCTEpGTc2juPg7
35rHLh9D5PSgU9BOQjSvxZ2tCQww9bSYAqA3lkbPY84hbz14mJxIfH6Q2nPhYw5zh5+32v+Oq8gG
uQaNqQWaYl8FRUnpVnhjGdTZJJ0Qwtv2FdYNzkiWT4iAoKqdrGgpVjGB7fOgctwa+mnIWpzBwlid
uPEXjsihh0jiRXon84fpnCSn7eiJixQTfPU+T7cxLr1Radh4KctTvR1yCuSMP2uNojiz/x5Q85sD
ahjoEh+vdvVlEuLE3twfWF05749Tr07mMd9QWSs+5X+Alr7AdbVNlOUdmGJSpANBzijqchhhWvKW
VSYSpK+w+34CLE5O363+1g7TR9S8tdwdshJzbHsvL/m6ccMxrnPFmUMTNLjswwTrcZP+FPNuRJFc
/txZRIjmsJMWbuqjJQk4tpQa3YZvvljdYVW4JbzPJITzjlORT18XK5cKXwY99Jti/LJ7LIlLMnXb
BeLkwLXYX7G8xnyamkP19Opj586c1omi69Nguu3ut8HRh1dEODjNTW2xUpPAuSs3R9zwZni2mNnL
OlVqSqe91keFT5sMtOFFYKB70XpFNPLCD5+Bcv427KOFf5EWAZpHMck7xDqg5ur2yxneZ4N1O3rp
vqK6K17ix27IEYTuPSsLF514Kgg63oC8Te95bzF5CHaWcVcK7m7sxVoi8akhWFj294XzWqP3trxS
3R6SGhKLcIZLLs9+E+b+H0vhJ6E5ikNjSQCZNiIkbnXdqeisPYb1y7vcICgAMfeS9HYQkARG4h3K
rvfn10VGbDQAjGXrG3sTa5AtxqhBT7UCF9m1dvjfB3xmCRQkoJwPlZbv8oTTAofgiPpOcqmfZc2p
D4HL8ZMPZc8ZijR3p0iqU0BoKC33orVzfHb4yN7yDG88W1cY8R+vFPyuvj84lgLFdGIUywvoC2er
9b1eyTCRWDM5A+XgrXs1S7FnXtW9W+6wVwm1NC84yr+2od4RSIqXuPGpnu7zAQ8Oo1zJn4EtkRBQ
LmR0KZa3UR2oWQ8hHmzHSHv2qTy0s1tjvbIIPFBRMtEHz1YMQNAvb/N3tIyAwecfhgEFGl9kbhYl
mtGN0g9NG2whYruXiLnzw3tJ9lqDg7o1ReG7bYgR2OkiPi+SUIn67GWMidgTAipDqK3PNgU3MeeQ
aQ5XrzfzqdnVG0OoBy3F701M4rPVuZ2CeRh3nAKGGYtYzPtaJo8TI5nzgtDgzesC5nqCiuTm906d
ypmmp3PX6wLC5FBJAxamp/G/iWe9WKmzGkiMcIorUukEe8Emplmb0at/tR4ewj2iGpPQyfWMjhBe
Q7BgCwF51vUMx+Znd43ugAITJ18RS17zm10NuR/5K8jwW0kVpQ5cEygJn9NFAXHqisE1dAtMqrGq
Ezbeof+DkCPE2lvJFb+HVikvKo45YBi8XW2S8ouCkwsTmnBIoDO0L/SndiwuAjE0XtT4ffFd7f/J
YtsDJ/e0D6raIz2kZQj0AkjwgstkEz9FI0nT2FrBpsKOE6fD8kCaEvkH5hKr0TfUWCKsn01dWwJy
6HJ/kaxukrgf3Rg6yQdF4UFYhfJj/MS/Gj2iVNYTdv0YwEzFKYmscCz4J2FTACQwNR2tMxcX3DLa
8Bk6577VSdwMeSH3bGZ9R71jRMl670a/r+6/ViNJ/H54EcYsZMXJjVqvkWwDO70FJL//a+TbWdNa
HjCKqE/Fhv7ZHfZGgwaew5r1n9b8XlW8sh7mLwjooUD8nOTM6LXwNlYoQtMzgO6pl/BYu4h9vSxr
anQcBf2kENXEtpoyCVS4y6enQfB7umxp2Jgi3/v1x6kYsFZxd6x6K38EhkivN3zbElaMwAN6n24o
IMtnsVPfOi1JAroH0q2ff4d5XqM7pg1mvP9itSsko4F52WQ85jjSjeiXhAw2idlmCnotB9T8IxZ6
uvhmvoXX4x4fjtXFA+XFdSCLoWWMkrT8KW27HYFB7StshyBb2GCVYsdnrg6L3mRUhhNCjrnOwEEP
HD9hYosYx8cuVNTMfghMvE+A6g0GEBSnPpACPvwP7r2s9CrFZwptyS3whv3AxFsW+PQcw4Ogmn72
qwgdzqLzPc/AFrXN69ZclnGyqnn+fxwnEbqovK9ZKJd4yXjgd/qEnM2rtZLuy2my8qwRLC2euUmr
CnmcONeMZDN0cgU3ZkrMnZCPNz4JRiYBGD/FBWUobb26CORGoq07FuknwWVgFbkLq8FKA/lDDbzh
Ow7oh8VGe54Pd4HvqJnz+jYs42LXExDSOep9wMuSTntpdmMuCoJ7brGGf01xC/F/v6htU/fjbNpl
Soqdkx5GbnhjhwRSR2C040SBj5+wOQusZzN/V7TpFMQWLGg2EEo6IySYNNZjcJQs9CUiIDCybSBp
u1d01yv9MgkrVRW786axO/HCHZ0IxBmFpAaPSr1+C09q3uBbuTGV9YPocj5tS/JqfSMzGE3B2ZJC
McFkW4LS7wOnqOf2bQBMN54IiQg+8BTWOLn7b6LAtOBwTL/ADP3PvBppmqHNpf7YYGKmkOmH0MHt
lolxqPD/VJ6Uv/QL6+5WY8u3fPTpCeRU7FPsksjaCU2eX93Tv7JyhHyqZwKfzrnjcfcUyAQRe3rj
PFR+yvpXJnQR0MdD7+P6b+0MuiguVO1uf7ZzcYgU4PnlJ3mEWmDZnzz2sJ1+SM4QB1pZPFVcfJPC
L7YYDO4Q0yUzn1N0RkDUmmuFYk4jRkqASH4cZa++XeN1R4Dhnmv+85vwuaR0D3PDvHGKow9V8iZ5
gNsfOxNMsd8sqqM9VMOJviTO4HhrJby4ZS4jereNuawyTI7vtbSNyj7uDNT4Molo3bHAcSCMbCm1
MQ6ECruNVKwD75hdBjgvyQ235JSllYOtIDtH1y2xLvJqVbrLTGkKcbECRkV9N0eZ4Z10c+KHBNE0
/rI3pZDU6y6c0uPFOQ8OMWoJMcJpUCp3s7rfQJaFBxfnyuNBUNtSAlfShoOYVIvii7pf3YWTYXuR
BZpuWpFku563cAjLF0jkYnuOndAOpfUD55aeaRBLZoq68SwcnDWrBeQlmDkUKIk2XM7ZkWvoPpJz
DY9Cf9GnXHfbiz3C9XZdNa/cXpKmEFDlvwo7WuyR6xkTTOPvy5DthuIJ7O3bN+a7CcKGFsWV5/Bp
NA18fJy1RUu7fkyfHTUdxyaFeZNPOLgpFUO/LTBZksN/oZXwvhUNv8tjmZwIhmgmJb2tMl0Dw2la
Ntaz1WnKqw21N70Z4xFJWNfI/iY8lxkojULoxDAfbImjSiPe2S8fceYXNcZ4VxcPYbKn2/1m+0Yg
9+DtTBEIxTpRpm8u3sjFmGn54XsROrzOqwzYnzGVsWme2clTZ8ZsJPq8OD9ytVd5+cw37z0zsU7/
W4SQQISGsv+ZX327gIW2Pl1xDybXn3S3pxKq6sw5BsferHJyg9+Dms2k7u+kJosrqNGD40NbQ7kC
NDtFkWoybx5bZA2EWjiV3WTdP9rwk5GgkNXH5ScFvZ4ldH1iIuiIGpX8jjLONIXyYvDjD5MzUGig
nfbnITizpJSzkrbptWN418DBrR6vWq4+ar+zDzRB5zkAheBKV6idTsn/53288AwQPVj5c/2Sua9p
ZirnL/Hi+4Sh/2581ldMeybzu52g4uy1hIS9oz5Uihd+kJ6rRnKGugWEqVjSzNdqZUrA9cU2CST1
ERS0m27NOvrYVNeiMldQTYoM6MoUmaZiRp/CIS87JoIG4tUpWN+aiyoAnuLVJtF8OlFAnTfx8Z82
1SbZGs4eeRG+W4LNFuZFruo+OcQNjht9I9nkt6QQjftR8GwZwNpxStfKbDUjOCbzpiisTlmGjZ9X
qsBbrFadRiM2N1yWYI5pR4Nfra+IUc4eeVGn0ntxLao8dS3I19+OVoS6MfGkXjJTumlTkYdzM36Y
5Gok2Y39O+DaUuO3D2HXsnfGmKFfSkdZx5frEMNN8HKzP+9mAzsg3fTMdBgKDUL/RDavjtZQs3pH
yKkuHHQTXMjKmrwTsXQd0yqoRqTNrrFvjFi9ab3b9YJHCVV4Y8Dq1WHSZQCf+tykSaVlVt1QQ0x1
cTSzujFHvinhSWRGxrzowzaRd9Ge7ZGL3/qBsC/QEI1dp1/RFuHWaSuO97CY2FUCK0PD+YYqM3yI
H3nqrASVOkuOQ2vQrQjkWUnh2EXh7qloF7/vFAbS9r41kDHgizVg3TtjBW+3v3P4Za8svf1lR6gr
Vvy6s28FJFFWmG3iXaxRT94S1Y2y/6Wy0IJJr54tfV4Ba8tyIPrGwUANduKz4wu2FyEHIBnSX1Cb
8g3lAlSf9WpwpP1sJ4jiAdDjfbp2wpHLoI6YN5cKEWPI0Ue1PtlxOnd+iz59C9Y/tHjYQa+8ghcH
Nl3HrZR2osdFEYD8vSsWdR2OB+begSxeUOvLj9F8q6wUmRARdM7N79C8chFXQhoeOtKpsocBVlRr
NtLxZqXutp6P8LoeQ8fvY//La4+q8R6lZc0xo784OJsI6s+c+Xv4X/dqd2b9uEKLi31/IURxn6Q1
vy5zjvMmxN3SDRVhoRPngOvB5Q0cdrMpy/+SQioETMuVvK2yfbfYGjjMudQ3JwufM/8ykdm+HFF1
TH3uVjM2JTOsR2H2/fzlSelpEXEMExisLmv9hj/vRlL+TMitlK7kySVVTROuZxXhyhwD/fcTa1MF
fYtVblHCYghpAhuQK8PuYG0UJMJNLrHglRgIHnKAXo2ImwMoYuDHHb0x6/q3zHZkW5hB5p9K8jZV
9dndPL2bH+ADu2mPZYIIjuTpDkDGXMSJzzRX/Pe6NidhNFQLjQ3nDFL+KhSrGcCBhIJDSfyoiZVe
XvjkdtGepYoDg8XibyTLmINs+Vxlwgsgmttv3x1oHVT292ASvm4EkxLLmUReXCP6MEpRtAs/awQi
06vbSmWf9YPSOtGJJw1jH7mwrZpnRd1JDsww7B4zoeinAw8XZuw/FTSGrg0+jM0ZWXjSF7dqa47I
J3Gub9dDTz1ZhyOt2eZDvGVkiv12qxS38+c+lbIzPvr7/F4XqQPcH0L139HbqnkvGSrSvl/Y6SuT
YThXDJmsmNe/AfP2ghHdsklddoxjqgR1aOI2mfISc0sv1Vt8eiZ2kN/HQsic8kPjiI3JCON8yFQ2
KczVapdKreQ4g+iWwBlJnETyrzR8/TBg0BaFz62a0sOo6BIoXTVuh7TKJcXT+mgv6ey82DdAz+0F
TMqAWTWtILrXS2nC0JBFoUJRjQlVLxJVEpS2VQ71NPAIXar9IsNgQKrb9+aA5SWRF7cG/qiaLhpF
pYC2jV9o+pw46LsbJ8p6UxffHv5dvtlYlSf2ucIZ/SF11FUlzpSJf0aRtarJiTWq/bigiANIuupR
7guYUhBRsMu23AYI5el04A3V9vbafE6dePTnTvGscCuvfIlDBPPcesguFbgOmnYbVPEyubhuLqAs
xayXwSjIVtdRwY3fqHwi7wg6XFGDODzURjniqlwmHbD9A/bJQSi5EH3VxmfQRwrEU1TcmX9JO3cY
mSyUgXwlefkpXGKXt6qJf/7h4NSHgzUK/GapC07bxtGFHHDycm/lvESLCgoLrWzr4LBs6bKtrQzD
t/PcesU6Wt1d8i/u73gM0W/TPK3XLmMIzwwjHv1cTRWj6FmmGZUAxqeF5OsHwC0ImTHIUKF6qqvM
BTL7CljXDQLpOjEEgm6rx5HywRqv7UouDe4IDaUxLTZKKNe3BBztNuqdEbfuibWMa993wGD8G/Ht
X0qRNok0BC0DTHIORQXlZY5S0kpUCeYvOysmYe1srwlE66GfRyyVqDx4rylVRQYLI3t5dnkO09Cw
3VWDa1t9VKw0xsHKhUYZb9XhPasmHSSdA/MQ43MlgiWnn01RYs8YgG3Y8SqsY22u9THZluA6K3cr
nQrDQNquaz6WbDK2OnwFI80/KA5ozq8Z9k0CVQSiDT6f9XUgWvlCJKQsWb9vfezcodY3zmreyI5f
GWG8UTiLmpuvxnxn92bOPKMgpR0YgrIOlwwy7A1amPyLDCSCog/JBzFfS7/fJ/AB1R3O0mVSDhsz
kJVT2nE1C4f7hl+PCjoMaJtGi3XGTFj+b248GHtlRTUKdhKNeHfg/vh2pHhz0Jcs7Wl0zJCzsEzG
922WxFbNua+5230+nNnUpluvSeIbuOIsipZWdCfTGoYKQ4i7+qA5gFdqEbrWkHVNXppcI5fz8JGy
sea+gtNBYq5fanm4T08Zid6Qz25ci/rU2dQmk0XYuiiat28OuaMQZ4jB/oaml45oPAzd5Zb1Oc4J
KH8eT8BAGpxb7sl7p7NKskIHjO5y8rAekL8qtB0eKnsWgroNLE92qHETeCdj0QXwPYGtXW7q4ctj
o6A9LvGsCoqvj1n9N5MCb8DfFVqjTVdfpaUf9P7O7/0raHvaUez1ollrWwi7kc3wh3fiw10QKeHZ
NZ+qFrzd3m1L7PSpbtVluUtznntpduyHbOSTIohYbWk9apL+/x+wZ6QyimQNzAyqnDpJ4Rq4ZW+K
Go883MLBzsTsHrku8qp9c9sadZcPEznFYhNTfQPG8kyKHNF3tVM5FT5/RUpI1M4lQHg0kHezMlPY
bxeMoqEiV/A5q5TCW+THv4ABEqi0sC+2z9AMOK+Ae9HDjkspadwNgeGG2DZUInLEAaTr4YWI7GYp
Cazz41mWgPDGIjirHGsjtwXF+qecgedHwIpSyKX+j/5xZsdiKCQODGlGyvyFCOy78Bmyg8X2gi27
6+7raDCLRgZFOQHESa/97b9qi1uLuEL50kOodXifMO9BKILV/7Y/+oV1CvD8MdpUxoJj/8t8deDf
lLQV11FnKUXWuCtm+W/C+8YTVdvHQwBHg+L9gk6Rh+CB/XE91Aqk2okML0V2rYdpsEgquPv30uNW
1AFp26GI6OmNYWaP3d1fF9Wc/V0GKGGueWtvRMKTawK/f5bR1z57dhppAWlrU5oQFYKTXHqPojbo
OUdww8NtIMz7XiLMEaOF9In7/JIDjgg8MsNmW9RN34eviCLKvG3oUk3pkYeP6XvGiAUy8Q0ay9k5
L83BJS1xN/aks1OkKWYUrnzVvYZsrv1//PI2oVNEXMJ/nHzOAh291In8uJfwRgjZP2drvngcIZ4A
wtR7UT6qORziRLXGfRF/uK2rpFMhukIFEz100SISEYiDq4Th8zXNwe9VO4IlS9JbTMYqPjltiAbY
rbNLz6C271dt+sjxXZF3D7SJjDpcTi9SXaYrmTQ7W0uQ/XbPkEXEvsHHhRSeNoX9572qhOxvLkh3
LQcjUh9AKRWiRq9OxLKhI53eUT16HRL/b8GUP3wSbgI3+/aq99BPs8Mg8R8f5kOWBFWqpkb0CxJ2
qQ+JCBrLEUs0+n1j4kTqJ7v4TagOtH3+e72m6YZYC2vxsKKq3eYR7yVeiJToQow0/Cp/huQe0j5j
66mSlVsjT62jdscoKGUF8udxGXQfqI/mUloMY12iPQgGAeqwbMFi03mAkjSiBA/zzXqbn1SiDzed
IzmASpeI8LKFKeLI0yEE88qDNZ6gOwiR9q55YHfGww89y6GvVQ0td4+s9ttz46SpMEy9R54p40TO
UfBSKPT9wvDERuKkk5KTyqrvl1CK4dzd0znVz+JNIp9KO7YJxmw87O36y9RlRWRL/WW6ztEOJDv7
UWtDrgP+9OPXAOE51JuZe171QuysVmRNuBPtih1F2nKKdWlog5gJSvEdljCA1XaTzcxrresQ5WQv
PJTvB5RVfViaJlW9DlxazxQcVCThlkzQ9JT2OabjrxFTFvfEWzn2uR9qdaWtN/KBv0Uvq1rpze5S
GySpVFhxBPdsixVlo9VmYFC21AZkctbJKUBqoewOwffG5I2TiHA3kFj6cdlCGik+G5csA+cZTuvW
cXC2ZdxK46U7JzyeAvW/ZwL5eM15c/zBN4ZjD9a1I72TmVWA+abbEmMWoZmsGNv7ogAbXV76u49S
YxaDd9s1RnMD8l7OLkTUuH7NhPKgmkxu990E+6u7pS283F8j5ZLZZ64MP+qXHUdVtMurQhVFdmn4
P4X0m4/O/WzXUcR99Rsl/ycKbthIjeQiE3HHXjEuW3geGG6yhJsUbCquwdhLh4CTic4+A/ZchSfV
u5hioAl2uTaumltMmNxGkIr/N4sepWJTF3mAOh8vbukz85ytVgr5Z3UHNvRh1PI8V9NbIcVl8d6E
Cr3nobwzpeyzTdNjjNcONtLyKrE6/iKVTMDH4Lixd/C2OrtlPyfHi3nDToahdEehdGuS+Dw5BGIZ
43bZgetJcui7LxNzfcRKJVeCVZl6+kGRNr1SAbSPXClNjEzym/r8qBBCQEvicXm+gjxtDw8eXkt/
kUdu0yIBV9CFPJFXO1MJBcR/btwxSWDEUJbRpHRttYMbmeIkstSMQA/YPqZDJPIGcR37jGP3eWr7
7olStcBzP807dJlg6zH9sUQcqarkCwJL7pUgVYDnLSEHG9/JG/adyx4KA1sOFk1fKNUd8CwJ71Sr
8MzZbtT4i0P+ITqEDgDZkBF1/nCWNtaOD2I6aHNF0GkHPv3+ne1rJeeS+aqPqasesOmdL5k56csu
Njt9qnrceZOgTtehzTBayMBLHGJ113nsqi2NIb91eTaPPdtgSv6TSj9VlhhjkZpEG6Y5/WcTlolq
sSmNyMgZgWPf9nhsyXuXyXtpYeRpV9SC+o7i6RsDWP7qsUG0/9YHb57mANpLeTuWDNrS4FLpFC6e
Bc5KDK9Xjm8CDQfAqtYcfJz/GNUNi0IP/v7JcscddNEK902jUynU1kjn6w7HlWYm0UAJ3celekaS
09ExgVY88sm8Tv/4JlLgcyzHNsX3PiHIA5uXAjRS2wpKJ/f4nf31LHHUQu0NMsXfwFSLUMU1Qh8q
zZDFj8YxuEgF1p1KJoCFb6xUVrV2nwtTfS8SZdVuSs8gWwLFyn90ca4ErZrQDs+7Jq9VUK7+As2s
3vgp9SKHHhC+2HxS3f5exRLwxyfHXkAbEo307Txso2bHL58q06OUcduqSxLRQ3338BDGzKh6FCQj
8wVp3pvehtol5L523TbPco0Uc69i7oidj4RpwOT5O1DVaelFaWO38RUgJ3qOok7qlhq6H2zYZTLh
HMqEG7AOJt8MPofLYD2lLfXr53uUrIxiUnrIjcg9K2ZZ0D6pMn0q/9M5oZm2XgpBMR5pMTyutF30
uklh1QDUcjK0RAHe0SJU+/ZbcWCtJxOtNwqF+Q2joA7dduwwKHg5ZvMna3BezPUoyR0L1aYN6uwT
/2DJclURmoomKSWOLv+bEYlIEme8999UxrKKfj5CrMwingMRTa0e3hwyVFLTlXQPjOEBxkitYKj7
LPAGCaTmHq3Wg6pWBARudTglGwvRJ9kLazfGfAIiO/3QrWodBogQsr336jdZSZmS4roR2kyhzv2f
RWHTD+D2aGRGECQMkK52EYPTMjn80dune5jKm/FDfAF/kMTYnfzP3Fr8uscmjxJ1/5zMJsXl5l2U
edqAX8iVvNcnvqFeTGpWa9MoMNqmfx5QVLszh9XL5hbYVtlBPJSP3tOoT5bbmaA0sEmQzJAcY6QJ
5F451TxvPDuBVgTJfPDs4ZCQbAemFgL6+aS0ZpvZKFfohTi6Obmb6LcjSXQzU3d/+Fal5D3JcB7U
NFcECWCfSL9tYksLFeG2c4tO+Fx3hTiywaD+WTavhasF/PTcTQqCUeBOCgFly2B2oQudGhTtF6iU
ijCLrV0aGymXOhklUk3FmEeT1pLeZKq3gKvrXZSEdNcjVJ1uQ2jo/jqcLNLF32ZQrVy5EBmA6mS8
Y+9HrFZY5IeLMV+gXULIJb9UpMMpvT27JakAxLz0gu938H2ys1jNuiZplFy6KBBjxrXUsKTGKhy/
4SVysBzS5gYKjB2MhZB2MeK/iEPNUWZP30kjz/4tVwwEghWXs76rt27S62w2YgThLNWDmTsiw0qQ
pYBO3qC/wE05BEtIsiF6H3k913eY8orR4hJexED+VfI9EMDB6uteH+dmMIAkYkDvpHra/OmatRHk
6nmm7gS7l6wKoeRr4SmZB5wHEv4g1egfkzTwR1+TVxOBfgjPum1wwR/ZU0bcDS2j8FIqJo5PYlsf
7Kg6t8MRmwglcKJ6Ubb1W5mRlm0SgNlwJH1jxeFVmgeySFBS4OFcIOrD3d659GTLmc9aqW2W96b5
/T+J2CUq+QsKGUbHvHrY1Oz2Dc6s5qtAlAlnlcOZMFh0sk7/84zTGjT4Rk9QM/G6XZGMTtBTJN9k
s47PAtj9bCAg5QUn5AwpfTmHzcPEu/RYLx8ekKcLVsHtAyw2maIfeqqbFxZwBdMIByOM9vVQXTkV
wLBru+fPaKLTGfnd+BTcMlrkFruo/RbnXZ2QP+IzRQXD8A3JQGVg2JFtOMoE0sB8Jlz1PFnbbOZ5
AYLv4gxbb217j992F/Ces/P0OEphCfctwhPqEYCQuXyhZo9wITsdIcH6OKz8Diwu8oXVrap1dIM+
iVKGwdJGyKn0gP787N/2cPCgfjnZnIoDZ3ufR0w0B0qXOTOcnUCzyuTgxTX3p+2kDXyd6HnltOSq
PYLmSqOr1fcB836jkt+NlckTrZDkAfdIV/58c3l0HqAMntLx1Iq7pcuZ+L22waOJfl4vaUkffdAp
hQDXSnHJ1aovRo94B+QfZ1p0SBwW9/8tVhHvNVH6XXbcTkDm81ZBVg2lda3a49bkCnyoGxYarXbe
2y3O/VOXrpJzhfkZ2pco1y2lZvo6ZAfG/R70ZKUJzH3YA8n7E9EqGKE010XzWtVg220he1QY8Y+E
TtR0YbSrNl4ju4GVrBNHRAxKr6hxKkNL2bkgkxnLljcOIKWModZT86Qsu7xafNyj7o1XMpdObSaq
YcChFIBuQR50Epai+FIQQcgcXuVkGZKaQ4mPOVv2IBslBRKcMW4enH+T037okF1+jZN1d/QqmVLc
+NtvGoI/6JrkX820tcUwQLMR5zGmZ0jo/evvvcjLTmSyxEvuR4SYcTfP7ZrkQ8ovpu5w+7I/zXak
QExdzBDOw7XTybX8BVvxAXt9HImam33E1EUtOyL7fLWAnk3WktgwPa/6YaY9/MbxTMLhty+jTlas
5PP+HJIMTr86vKlDIaVmcAZx880jIa5lyb2h1N32IpKaPQI2zWurKDMOfhHjM+4g+NiuMN/DZjgO
LXqC+86B9zk8ytEsJduSF9dEgQM8mM+ZazVKlG+F1L420jE3IKIr9R5UlBZUw3gSKDfrjERsDnOs
SJtBkCceM5NyTfxbnwMkatBKAVFmw18+1HAo8DzAhT7N2ZaTsMSSuGlQJNRGuG0jjTfLfdqmbem7
5yJENP348YXOkItqc295aAfHnAkcnCEyyXBqfn9zZAiGFkZjRS1728fzKEkL0xcZvTTb5LJU5y0C
MwNiQ9s5DsO19k/CP6Uja9wNLOO37yuVFOclCeD0Ds/AHebI5i2kO5AZ0Jv2Xkr2Mmbe1Sf4Uavf
FDSaweUxmfD/aI/5XZi1KFukacOm8UOw0I3VgHhWMbhUMQAvMnCJJeMQIZxmte4Wwz73rLH/KOS7
iWyZ+YPMKuoxCbrlvXsV5ROAZQhdPlrHlWHKqlYC6+CiLvSAp6x93dvEx9B4vG+3smZD5/pC4bKz
PN+aKG8XJ2UGOkUsS5T2Z+sDnzC84/0sK8S9+g84ftkrRHufXNwNtsyIg4IT7YT7/X7O8vUKTTTX
t+p7KW0tRzhDV3m3tkGx95VV/df0wBbW+vmYTcpsLzig3XwXtdoAIRjGxfCdLf//LpjTJXiK5jDo
aiWeDVmXqrJ0HlDk3NUxno2Zt6bFwxgqxNvJ7Ylt8oG5ASLio2/AmnjA1ghFSVyareUiFn2VJy2J
aTCorvKWl0dq6Ng8eis0kgQkLLqmIttVHE3X8jh550lRYp9KnFyG7+SpvWPSW8saFLAIGL9uZf97
BWWI4qw1gY76wpAw2b68NR6tOl0JCqJeTfF8OrkQ3ZPgNanvFScJe7freZfNWZCFFVKQJPjqhcmN
QAV6BAIwE0iBs868JPX67apAqKmxmKZ2URhG6Ri2btAGtqK0jwYAPWhFlxrJxBAflE3cBTh0mJuc
V4y+ZT/rjuq6kab1Ie+m2XNgQ+T/v2Thl0v1ET7zONkPi0H9lzlzl5+HxiHiyWM1LpEYjZE0PXrH
puROVbw72JmPeO+ScNXaVRRQ5NsKKvS4881Lr2egnFdt7lz2UZmgO5RPqZApLlegW9AbCSQRjAyx
nGyY8a4T9E4g0K8IwbCgCmxAgPJQmmGfnRMKUcfbKYPodjE6khaFZqVqmwRZHD3OlYBhyzBiLBpl
dnxc1lxMHIES/TeIT2aowA6Gcaxt8mZY+M8fwkaSOiqsQF5tzVBVV54Gog11XNxOq2061IevEWL3
BHVj8sMtYRiOFzrTvAiF1XOrUR2ojxw5IjlIkKkAv3YY62d5o415Zk7kuCP/bOEoYppWgqW3WLiF
IWU/iViBnkCH4vRQoFbtPtGsrwJxvEVVocHI4/xewvFMMyO4xyrJVaywE3qi2ytpBrlEP2pXvRFi
R/nI80YdDPQhHf9N7S1iW5iXDBcxQFZSzcOs8rwxPwtXLWUeeu/wC9pJq+1jmQR68YPbmVG0Vgd/
EhIUT1WhZw/oahGXrm+MAaM28Vpg6l+iW2C4rCAzSLvOnHR+AVCC3tPN9C74XD7Wm4uBqFNihL0W
YMuGfEYPVM+CZqMax31jbtOrd9h4iP3l3+P9Dgixt7rb0aBKqUU0J40CSumditOW6biONwrI1Sjb
Gje43Qu6Bkdu3UolwK0/j6+bas9ZufdsxtQT8CJ+r9I2hgS2tf8XLSb9AMiHQxqbmzPo7pIXVW1Y
wY2V/HPKNnFpq3yjitxrzNMkYrbBu/LwmOhdHon3D/2kI4HXdug2xxOlpKYtDVyXiMogg0KL7E5v
a33rzFYjjGDKcV4TnGeje7JxMYypwixvfLo/oJ++N6nqGkHeZTtrTUZncWZIz/7zdWRNyr0D9Nb2
lXajXUS7G388V75X70zQRPQjcm7mr8CIGH9sPWgUMo4ao6aCW9sDnz5oluLaFrtJkSZdPJu8C6D4
yq87p5CZZ88ovdIJvDcfst6vnBfp6TIy2JnQq2gxxaco2OISlTUqJkn0NVHRLJC+NUp90qvOGvCS
oablxd0kBIFTB4vFD48JS7Wm+Hifm8MmRjpJfRgVwjCYPeAoyAREs5J5GIjL85HQRsDyIpy/YsSP
X5fqQU75wyxdoFjol/f7ekWkTKvP7ToIT5OCIDXzpKhL0a2Nc4QsdvARwPZ0lWby+/IZ5+m2eHFj
XHZNj7yGSRsEjUq8Sp/Q3vcchJNfl4iUq3T/SyThgsT6FqK1lXzqD315M8ldLkX8d+hdl1h4jCbU
SOljTi55SMUu14iWXCsVXt49+6j7U17b/o7G44lbs7h3seSEjUYsGgZEmoK5nrUhA8GCs0EpViCq
TTAMarbmsR+hgy160kImZ3AorRxWyUx4JUhM55vAH68aKMkxbkH0VdWXn62kDsxZU9cVhhwZrrWe
G4S2JUST39B6AuqDnsmAxq/geBdDgkCOmiaBmMzMdzDTxbV/vtz40J9Dzlc4I09MBHQxTZ0xHnEO
YdUv4vkQTPOHoLxGg9wp9oMmO2Mt8ydJChnPyQPv4y3+g1fHVp07FhOp8Xu19tHhFKgbYDgmghWp
716CpbrH/6Ag8gAzfEtaH+FfZl4Lf82wqzEPrQzpUKOteo5o2fb+0mZb4BT8okFaFTZdtXKJey0M
2vvNx3FJHcctHQDeGM5Zj5ksvgAT5upZXLVE0SIgaEqLYoQ+zQXFyNK90WaE3aNbbdb3EJLEEkOX
63lvLln1lK9SZX1BuRj6DhxVbp3QCj/PFXgD4lAzhFAFIftWxD9KetDclw1wzwPDby4NshnyIXp9
e9VtahdjPd9SaMsogH2yLvc1Slqx75nDq4TfI3KymeXC+IXTw3UG7ZgRosuE1aXWjv7iEBq+o+B8
YKAdkTdaL3V5/2nYNX8i1E2OLTupfen01D0WBp4sL+aEE7Mu9Kll07hPx5lCLkmh1CAT6mj1uJ+r
ogUozLMNFs0t/9LPz2ON4n6xwr98hPDshLI/0++qwY8xvxDY6G4NFdyrAji2apOqbWi6VTUC107w
Uoi2a/oP2fkQB18WJOqs/OTWsLAThMVtrw4X1QJMDak54yFAkIyiAPnmEkncFMmMDAgczNv8LSsi
Nde46fVbnurc61bJUZonxP0tt2kFVTWY6GcKt4YpcNTaVICBuk1Tq5TGg9ztsFLq+70+QT5qgdwu
QCywEyaKNqHPFxycDKqtnWnkbvYtb/K3xp+inBZ6qLPoDGicaZpgGuJi1weqND7jBptVSIJXDQtf
YyLdYrz8VS1okySbzd/I0MqilZkfMkeoOG9cBzhbjuyKphAkNntJFooNFB3mnSyhRo5KlKgGUg6W
3sYcWoPJjymSLkW7j/GqjX0J79KedpHa3renX2AQkdux1TERI/Hqx/n4OYB5KtY6z5TVnME5st3R
gAqUIYvpuI5klRwICNYAAigdRi1t+jXJp5s+O7D9aRmLGNBAStxp3SrL0QqNxaZyH7uuRfzx7/0O
/NF70ZQnpw8DfVeBo/AxFqi/Iv5BfZvlA6h19phaDjHA1LBdtXCyYXqp36oNPhICDloSyn0nqJ6C
eaQcfwAM1/79Oim+9ZEYlT3khFZ9KS1XxVTmnb/4h6HeZUUL/bI+Zv9zb+B9oca5k5vgrO2/vaHB
5TAojqhc6DtQ0AzMAKs0ZRMKAS6StsXs4HBrEwObiGmJ+JE6FTDKXyfkollMaUK3Q36POTjDu+pS
I4sIqsgqvEU3XIxXur2LJAmX4pDOnQ8TV+eiu4p4bTbsM8n0uMd++DN4GM2u3BOz9nLuOTpUQF7t
ONC18Tge5IPBA1GOBM3QUeTZN590CVk5Pya0r8jZA38/BaMG74hiTmMrcIHd8e54thGbjpAp2kwg
WQg2RlyVaK1ZH5bxC2hPN05BUwf1Tm6oRHfeTNKzKcaD2jc2VDznhuRCKWifjLjlckWYPFYTP509
vlmHv01TOIrzVGjB/rOkDJR/RhNb+vojcoW2rGRdT0vNZcDfH/r8YxiasVrCumHyU7cT4xgPTAf1
S2ad+KerPAI4pKYCVfwq3M2PG5aSlUzhBzIWQXDgWeZ3n2mIOfSEi9GQlZiGRbMaqNmhc3sXKErz
3beRWjskr53E3gT6UlZXSZ/i+nZTps6ASgWjmLuDt7Y99SHa5x2B4mVhLHUwKYiDrZNx1VMSicCs
2uv4F1RDWdvgZimi1xG93buLM65TLKQmdqaRpzSa6pO31s/tDnjCjIDLC5r4gCgglXdX1AaXzog8
GrgZBrZLB8v2hW+DdUknnvzTfaQi7FWUqpUNdeLZQypBvRrsWXQruVNM+H5ZPCGgDTQAR3FCf+a5
nMHEFyjiIXXYm+/ec1wonWXD4s7jW1i5iS3ixd4dEV3EZlMXXV38+aKnYev2TRMim/wW4/cJsMIf
ux6UiObqb7+HN2ta8YHHJVOM8KkISzCZqC75iH2Uq4S22ip91FncBqZzUAfVL0AN0idbQAHk8nfo
IuLM9Tg5l5nipzV0wUCT2J8l7mSx8d9wK4Agw7jJX1tvWmDFUaBrUkHV3IcYDJNeKyrU0n2PCLGi
kb//mOamClM2kzo9VypY2itfZYrGS9n3voliDlHsF9fnI+GMuBp8vbf75k4RYJOS9DfjwbGfsEU+
6fdkxd+oEgEPGIV//HKSuSzp0IlbXoHbrSgWJYRnafjhGx/IHWo6IM97q3Lze2M8gDkKCsIT95JY
tA9tRgms2rSaeTLkO9irOtpTqJBRSJABfAxOqi1fDBcmUtFg8oCxHuUUszLSXEpbiJX+zMifCtI6
p/YEolqDJnu59kK1pljoBD5UPUM2oazL37wP84SNp2l2uEX/ZTnL2vWwTMJbfJz3GVLIupxtFEFB
YdA78wo+roDGhLne3YlSYzuXhpchIHP020KJK8ptjCjun3XHU/Dhsjcj+4Jwha5byAskbcjYWZBV
ixkjs5RbJeaxmk7GuS34ksRxdfUtccTKsuDDKlSUtQcknwLbCv/CHr8Eihq5tJpos/eakD21B4Mf
9LPFE+/SQrdAFuI+0RxCAdF0fS+xVLhOGheGIpPimpWrOmnVQ0nhDcA1LebklNufpA+rH1GDqeac
T6FHPOksDpPF8j7TFlZW03rjfLxF1sZGPZGFZE1fCG8Xyg2zdogVqNsQUk8rG0E1GbGsgnlSoVyf
JvHkf427A08Y3gdCcioqdhWc775/wsUkPXYSwU1yDffFtvFnebMR1fow7X2V3rOu2/0BKd+21QvO
hOMkJSnMmlqkBw/apWUBDgwkZuUnCXg9BpRHatxJPZpw73PSnJKFG20Wk63iRvSvxOYU92+txu4u
IU0ZvhH8aqvcgbwsvTr8E5s+QwwhBSoZ9BAhbhaYDhztbQNvQNcLkl4+pb4GH73aLBVU0LiO9dCM
jR+1tKYq9IBRU5kNo/zhdwmsawXwVS4r+4K09UNmnj2TSR2oz+pPi59XrXWu6+8yXbJKdjD98DUv
0LIqUpqK4vp/+BoxBKwH59efOoMRB8eF9xa3gWfBgWq3SEqtyAjUHLuHzVzNYt7o29L7yRvN4AhQ
M1ne2bJKgIEosOO6EQOLYb1rOjYBUY3vvZ1WVf4RTkjB+ktltVeHDBRDSj6r9KfrdggkD2f4+no3
WasKY6Q5r89wKfZb1AnS/Qvc5QLvYW6sIwZfd3tnUCwCibnapUiTgxtniMokplDNqIHpDnJCklHb
bBsHZBshDPzgKdrWSE0ojb3dd2pyQLWYe6HJTzdT+OZJpVz3XRcVX9vGXKmVx0jRJL7scze4slmo
Zy/6rRY0RpkEGn/8GQK+wH2HE5asdYfzNgLJ7pcM5DCLrlloPU4m8DE281n3z210GO2/ed4thCfz
Sh9hOr0h35gQvUEWXDVf1mRYODTaDTZDDI6KnKijnKM2iXLKQlJl6jVZSj+JflsxMIPYwTbfRv9h
XgLN2BIESmG9BoN0OUmBzrOOlbRQViXM+BKaACF5vFA5w77PiQd9bXPQJub+AhzW1uJearesScsX
TqDw0CSVrtMs+6iRbHkKh0rCS57qMQ3PZwfFitg4ZL44pxE+etf7hTD6AI6meCy3wPlgDerd9vdY
vTiv875wkp7DB+e69qxx9ZcODDfzsEdkpb0K89VOyKYK1bOh3BP4Ct2GqvjOjIbdCskRId/sQpJv
xpA7z8docm4W9P9PMrunOqA4mg+wPJhPwP/MZRqH1DVxk8tY2ztjGlONhqGb6gl6okjvZkGyReSs
AQNUB2azrHnU2yJv5YZiuEQQ1bD9nfd2lq3AMq0fvqnrIy7zEh70/2JXRv8RCKq6di8vXGCFYJJs
vhHnGw/sgtZ5cCVeCNvHrGY1F35vmIg2nRK1yNFiJBipseeQh3yGWmh2oy0eUs89ci9uaik93WIB
hwpXbsso9DBWR5vIRPra/3W8XEyZHnUUhDvDahxG3sMeiQofzsWiHoSJWB4O/DbfllSdpds4jEZ6
7CPsloRmH8i3gSrR3+iis6y0NEOyPl7M0qyWLviXz9vy4b1dWaz2EimjQprfBaxoCpownDzyfCux
c65EEGmYQSISF4lYn1WWlXP1G/MybQst8pYF/YBUbq6asWy040ISzQP7oVSeIiiwQEchWVGPa0Ce
E40q4Cz8WtJcbZqwrZuyB1LZ81Tg77s/VBjK1HvL1dtnhVCNZfDOSTdkkUKqbW5m13si7XTP/QoI
SpBDnkWwUIe/bN6OxgdfzmWffrQQv3pDHweLmph1QxUIQ+SeuxT4fvcA4J+uuqKScoAA6X269XMj
R82+IsTEpIyVMVtNxVrJJg+h3uQ9oFlD+NQWGRbdjRxFO3r2ZruAQWMg+QUToAdCvyOqQg0ziG3O
3i3v5q8K9dMJHns9/bQ1NOVlvybJWR+s2xg5BsO6WJ2wydmS6zeklbUL/pFq0EUWtEGtgsq1Inro
CgbDrgBMyJ5S6jMFGJKFM02DLIoKz6BGJuh5xU3sxLoJtQyZKpK1+xO3yadDqKb6TKo9kzbkSAFk
+dCYEfaT2oQOlPjAbA4ol1U4bDxUINZJ9eRBi9dQ+Crlb25oux/k88ca/0mCkIgXnLMY4tgqJTZF
EmhJ+HqewT3TrqX4h/Gee+VSViuw8juVGUXnN6UJ4OGsQ+vrOhDkDPAFk6lpE6xHrYh6bSF9rpPi
2PvO+qrvAEqxtWYSZv28TJoBEkJAInzdM+0k2XrWR3rYrdh7u4sVPUzu5UJLpzA36oKZ73+mkOxf
neJmDdMKhzaPRJicBMpXvM98XMvOSggYNFGAbVjVzZKqJn7Vf20DsAzuYfpnHK3gRttwZZ2aN22l
7vtpr1ajapCpG5Z50JjuxRo92iOR8evq0JhLYiDhpXNMioNGeRTxPewWjCy0Dyishp5PWPGwf8eK
NMnuBzAojmizMFC1cMLgc3Px628uH17QM1/p3JTOXZrUQXz5FYhe0+9siSCtwj9iMyRC0cgLIyQg
NLtn7r3nLMVSwFwJUAZ5gvLRV/K9FZBnuTnNSa0c5jf6xtp97PpZBQMhMDcHk1APZXno1SC8Umg6
7YFnkROTdLoiKyhJ196N5h8Rxhx2ybtmJtIvJEG9EgUZ18uCgYScahtr5/IUjbGe9qV1zrl2W2wS
15/a/6ZOYS3ZP2xZGK8AqdmSa4WC6F95Ut6ubsFsdejGKFBhMjNGdSPdjtWGN4Mqj4FhI0OYwcPi
9CANh6ZVIhQPr9nBm3lAF/i78tEUPVbFSZDT8v1LsVoOWvLefyCvsnWeJ+gwJRYuZXP0DjbmIZPC
De4NP0T1tC2zIuMVjkpaRTxv/PY3otQbFf1A+DpoptQtJzWgYURK6fYkZ5nPmQ2/bhP6t0wZzPSs
Pc9MfopMpjEdF17gf0Jon9OjQz5xdfj20XIbOMx1ul9WQNlL6yist9u5yn1gx7lI+Gac2zV1q1G3
aQz7huObS7R2fj8O/J7x3kjc/e/RXBN3wP6LmgXXW+a/IZVzxkIcHJw4h1Ag1Y/+2msQ8h6yqd4P
kXnP7Ry+U0fKVMFrnJReMTb2MKo+YjT75se0lFmbxc4xMsK1lAlNG4yTTBCnwKoBWj91jz8WyTir
R+68No7A8SOHZACHRtFWccP+GKszjOteBh3m88+luQRbgQL1Si63/useHUngR7UO5VjjoUXidUKk
lgbCWRDKItPO92fdejmS0lQl2tmLag4uzgX1lcTCB+SpmWyzAnS1YUdpP4ZP3krfujAyL0gg3Suj
2v3NtXEwz/25dz68jcyl2EFr5UPVVBiRzn6lPAq4wgzKtVWGOYxmap6pVriVru0qQxjY/lSi4EuA
jikK6I9mz8g8z7MjIpm9p2UfCqlalKRMu5FbQgWIE43zDXl8lzyWjBV1BCfYfIzYkMB47UJwML6e
hrPn3w1y6V9z3KDpk/jTfxIvHf/s0TsTV6fET0hEBkZ6v0lInJVdfUyRDl0Eh5G1fZsA+n1dUKE1
7ZpfmRG38bn/RfDX5hvmBgpeWbsm9S6NyHFUMCM39Wf0FWfn6tFT+RT2N7dL9aQB2K0SAC0Q5hjT
wsfwq5NAzlWmuxeN+WjjZfjBa4zBQdjG3Qf9QiBG0V6r/p9rKz8sFF4o2nFpcl2x6G+gCGwK3InJ
zHmYVULtMWT5xJZkA0d17qGsiA1FuvdArpyTk5mrjGpTVgKkYww2iVXXg8rXl2ozPqCs8HuS/8tw
gEhuqaSKg/sl6sfRbEav+JDiWKbpWj+Cty6XmR8bl9q7HOl29DI49vZPCT/IGqrmEvUOEpD3Go2/
D08DQIAx0IOzwv7H0EVzoivs/75MvktO+e9fAiGlEWZ9E7nLboZF5Q4ZbMXo1O7rQJk7U55f4MtT
ptchAGGdMQJxjQdaWQjKQs4HIGfQwZbeGKsss/dHi3V6hbbmtiv1J12dHUj3ZfW8DqvzrwxxRHTS
8PNYRWURiyOtsMYQBZQu2jW6Vj38lKs1l4N8FwYAWyfvOL/V1PiC2GbItTk5IOKTACc+IekvITof
9x5sWyytXOUnfqG5TO0+yNg/xqSyNGlxXqbPC1v3+/OirZTkmYvTtA40fyIjcWiAx5dbqnJz/g49
P6gC57GDkHA9dsJWSLKTForsYejY1yiRg/B8F8atSJ+k8B/LfjSpeW7JgA1666saT2rdV7RUvJQ0
58X4/M1PoHVdb425Mw4IGz1TntpGLQAvicKTnfd4gzc1ppu6JR64gRKsQQrVabiS6KbdgD+TCSxr
+EP1yrwDen9UdpxRTGhkKFuqiKoX3NN34nh5UdO1+sWZqDDjmDpYRXOPO/y4YoJl1d/Pg0qPO1fz
2G2FQO3PY1DyEklUWcUQopqDZJvytTnGvF3q19AL4PM2EUlPJ7Tq1QN9+yzmd1ODAIv5B3P85uwS
G64FJevnawvulwT6TKI9WjXiM5QnZYu43586oAjmNZIr8rDeilEA38VObarJ4oufZFZbWVQWLGeT
65FiyHpCmKD+n95ygGntI/qjm420yt0ORfLGdLNHh3P03o7h5p6ZxW3WEjP70QdVNkmg6LVZJ1ql
zuLV/WfhNPLe5rsbvrjq1khTLke80AW8CpveOQeIQRD5HYzwYRDoRNuQkGVsieS6X/Qw9flygBiK
Xx3AvWdVT41Jor6O7gQ/rhAHD30uXahWmG/JhXZ1Z/s+Q8dpHYp+Kkl4ObC7iW/qT32VvxWemebh
Ge+6h3F+X1REvtJrdYbpaNUinwg7sfv1OMBLhGNnetFYWhU0hij5p1KEdkXVdyMks57PFvvMhRnK
/+jdCCqt0ibnlwQnATp7SbYL0hZtMQ9qjq3pbwhjJQ2JMQxWJzQN784DcioHLrLoqbgTJ7+Q/Oi6
yBlkOkxQ9Wa3WytHb5IQuyQ7BchdLGIiXQ4tPO3gtIZcDtxLntGKxe2P870M0gLeSfE+Vd5HQPAw
s07MtZy5f7/QwBwmPFrkNacmJXHZO2Q1XDRK8MElAU6OIpakg2UuGSrW3LnPCuoJtVqVji/KzSwW
jIzF/Ijn0/vXHazggnO2PF2JTJWj/jP1bEfvEBv4TgFpD3R7y8bUyblSuJfbp7OFCQ3+o5D41xVX
sve/u6ZIBmes7UAlCnbQbCDMUW2aDu/ze0IvFUYJ3I5Nor/Czw8IzKX9gP3S1/yrs4CTkkNcLLLA
+tsUU1mhy+II4lTL9GzXxbE1flPCkTS/TN6YpmStdBgEmC8esrHaxUi9ZuGb0jk9E59bBlga0+u0
OYWJjrs5ZIBlT6Xrlom7ibbl8c5NYhBPa2EYD/b+qJFioqeebTN9716Sopn7x/Brt2CnC9QT+xfE
tMileEm/oi0ISCWrCGLgItsqponhMnJAimb2ADDFzddFe4erqeSqc1VURUHx34XJJILFaVUqBPQn
L/fCBUljWM+Adav63KbRo118LxdHfyW3xXG6xGiyNe0oB1O4NfTMWkL00q78eBHSAFlI4uEF/NH5
UsAExmitUO7tfn2oTfaxn1iHHHadsPI1x96DaowyHFC9inIU8O+F0+EO5oyAzVKhFDMqyLgRs9UT
bGNq73RXiIIVUFvUwLSNTmrkZbIuwtyGCzzgzZ+ZK4R3RjyUolvb9Uq5Msk1nrXPR/EMuha+XBEQ
Qkka4RBoVmxHhOKoBvk14Co9FVrrYyEcM3piFiJl4p20F6OU3vJXkWFVG1lNU8vruXjVMY5+zMMS
IxmjAdsQoMoL2X9oWqxgsJjGXZkyau9qfHSpyOlj3HYguYSXNkYiCWOZjDykqKN1YCWv7viFMgTf
/ynijxs5oa6Ak/Y8IMOeRcSzVDgH6A8CKDsPlSXb8hMakgdkKZOgZ3DSEL42aK8LQ/Qw45T/g4/m
OQyT6UaC3B7rBYivhXDVxiQ9yQH8MUblrE0Wg5VtzdYNe6oafofEv6d84bKj4fhB3yjZvbEbiVce
5SZxcxLQ25gtxI+9T/nIIkI0uPVdoMU8ufg+1pq/bAUsoeyXTjXc3dX53Dg8xOq35TiMzCHDKk0U
awv4Y5Bt28x7ZiAL54+H7NJvMa++/LSnO7qfHk6C4HX1rsBiK4pqQQx3S/Xe7eHnYRL98qqW+A8q
j/vPqrvyjfFSDQIq3ZXDDsSU9aiD157a1acdv3pq9OaZiOctHLFlfhBhnkIloxrqYwyf1/dYi+PP
100frc6OL4nmWN6/b8zJiquEWL4bA2Vs2QBFGshkrIJXuYPdVYNBrf/mc9OzaUgDG5FU7M8BAnLM
GHmXNfE6x+AiZQUxYUbTcycunObPYtZNyPCSPorFDGmhbxX+t/Sl+OQEtgawHrFc9WAO3RCx7dqH
PmmFw02ZhEQm7r3dTfh7RJ5aBVRFMFKtTOuUtiGkPQxmFTNmEZR3Kz0r9i3CAYvNba+8WN0LMLbB
a6c7C/nj77Ip2LXK9j52OhXR5aF2uraflSntz3yPropC8JL2447Ewldxlzq5xvtDsazdseHYnyIr
/pegNHEoQdQdAOeDAcodrBvzS/NYS3lNJZyxCa9m35evPBDPzXR34LgCQfuOQuuHI0qCLhNzcQMO
XMxP1XgGFaROADmAhbfjUv04yERX9GMk0tXjQtHzQ7E0bBDaysfZl1PFSJ/Q3S1sHEc9R5Qd+HSR
IplWD6iru6AmC/lU+PwCfzIShSZTiW5n7ZxIlSl2mRR2rxxJK7ZKul8dAi6C23kFRqNCNkrik3Er
O5gL7QJZGPCgigDQCQNmAp3XrO5Oj09L8HclAdpMzHOSzG4/AXGr0hI2xIPxOOvyYHmVBOBv5jcw
q8jktNT0Z8bicTLldVAhC4Z+pYPjAV9suzy75aEayQyUT9aaEDPpDoFRpwkbYU2WhMxXwaofebmc
cx4TOV8SBu84l8aD0gncUU8Nyps5C6VPConkAG7DrO2vPkdT+SUrXFN//Oci0RmPHbXU4iXMBQR4
/dNpTT2w6FWfUI3Ze325Mx6HId0Vd0VTCAoaHZeSci58C+roEKIv/+j2NscwrYIudr4ki24mVz85
E8iHut6w9kXCnLqvGO86v8qoYk8sALh3ur9AOXnOFOyr0R/AAY9aUEBVNyaOTo2w2JQp6vQ3ZkfC
dFfgDUUZ5ZWnhPDjOZ9jaiDqnf4P1I1caEFAmuvOOs3m3rd3l/nHLAoBRnt5cCu4C3zicTv7eCkt
KVDhxHPpSTiG8K4B9RQ0i4BjJPCwxii+bU/7A6YITJcnMf8a4jig4JFkYIfZJd9w6m9nT8ry0QnB
b1/CfwEj9ccQMNqjBWbNxY+1bIbaYxP2aVuFZGjk4PbaUUtOJaI4BemcyRnyj6TQqSMxayevRrrm
gz3LgKFk9Vnge8d9dzazemfLewXCdDfV51PqqbuFO+915orkYVRLnclDBvkqNhFAi9HWsacmLRd6
uNK65wLt9d02PTVicE/+3aZ3JkAX1Zuw5dB46UFiFZXq3ohljRymCY5HtDIE4SKG3Bl8t2KwiYCP
ei8ctusCHv0Tc+XOK5/jD7OOYRdKlm35DfdzUa4vC9WFXf6bqyjTykLPc9vdq+QbsHcA8J3m7z0n
pb/TPSSbZ6d0ZcMCV+oJF3XGXma0SLarFfgAKoxGZ3kdYboIEf897zNRFG9l9cAONhm136QO/wnY
/sWCk4Tz6WpZGWzfGl19ibOmVw5Qq4bDiBYLi2dMafGRpUTpc7CBUE5hNAw+N4iGcJGdkwXRZwcB
NrkI/i6ivOm3K+GujuiVAr0MYt5L13wcrlqehHzeSw+0/Y1d5VnsUSThPi6JOFqIcyvLFVEBkwjA
HlN2+DOA2/8S6QVYhOJrAt/glmxba0hoPNFXpXrIwRL9MxtPsOWdJ1si4NA9jrlajehbMCLle2jp
U8LtZ1iF01UFzKC1FglhQ/J8WKJpAMsh1HMRHoE11tbX8bo2IdsP/LrufmLbpvxynsj785tm3MeL
liNLrL2t02/NbBOllAvYttDp0ouJ2VQRUdCue0/rtnAG+WdFkL79AuctYiHqKxjUXHSRlUuUSDyk
0Tado15yBBiDFmaRM2eYXQXDA0l87rbDYu+7vRxfNpu37Z1IvFW3hLLuC/YP9EnPqzAOEjXYTdTU
r/ezaLDW7lCKV2rgD2TQZsUvd+GfXyEESW0qBlXRKB0DIzaKsR/htgDA43xihj9hegtEGKYe49K3
xnlxNwfp1RYbHaq6zltJ10i4rg2ktIy52cgxEO/Omih02gBlta+KXasnn2fk7dC6E6bp8oxYSQ9h
8zVD3IcjF/XaUxt63kvAr41znPd3w8JunKlmY90FjQ1ZXvhq/q6O51k1B/DmJfBfRGNO1dbxtpBu
BuagvUP5majrojODnc4JHQlSfTcO2oJsbuQ7Ju6BiNsiCaHz+JP1DR4lebAyE+kSCTd/s21r1sJm
gTmlEDYaODwd5SW0sMy0CfW2Uy7LIAALyY48Hw4McSkpOltGcq0Mxv3/5AkYyhpYOT+yFWthldGm
58o9/Klg1BJchz7E7ecIMiLQbTGQwfjKzqRNXwdxqU2wJV4PenY6fIyYHwBomPWKn+QML8mLeS0l
bbfEGQPqvUiDNq5Cu1DXVYFxIzP0pEfLw0qhJNOwZ6JrBrQhB9INIMC/Gr0eMoGbNHDfSxH/whOW
Wk70PBN09629+ft4EAhHmGyKSin/dTT+UfANVkBFZjPmfZ+hBEo7sDAM+oPERD1Dlgkv3yoZ2ohk
W4yD/EYRoOE2haxc+YWAsR9PdozC4wcfqZZHlKpw4Ik20O0hE/+vLNO6GS+PJ8u3SyGTSvJNELyX
4Al/SFQUowkbkQMORZYYDEyL5+VPIoE+krx9HwybkBYQTxV3qy9J4YNlI6A7VHUecGRqK9MVOJrI
ub65+e6AwtkbgT+Wdea48yAidr27IoQEX69vZG4IT3OjQm4ebZRrkxIMNgsyVuW+AjR1c2ZVqq8/
t9Pa8awLkB/b87mUtNdSBvFb1O+Qaf2sTvz+PmyxSfIMkwZy1tsEycCVueTzm+TPwLCxDEQBsm6h
nSPYEp7WUubmxLyLiRW9Lw0LpsTE8Ufx5oGrMayGAwCShenrGJ+0nuy6I3DAXdn+GE4QQqrXsMN7
EWP4DlzbEkC482+vq48U8xAuztEqlorKj4OpAqqgw8eedC4Jx8AwrLZDrnOJjeh59sOIEvpAzCX7
2cKl0SmSX/7f37otlSZuRAy2gka5fRs7KGmMGNRgQkAeSXY17e5pU6DQLbhJMDwQAynquJv6KhYa
u7Cgg0EVGZXAzHfav3kSg+v68SaIQiGLTwFyMv0NTtxL6wjSnIpFl5tOAFtNkuD7nv/vC2roAHMZ
BYyqh1ingfS2NoscxkukI1HSo+CDCbv3d/UbAkkw/2S2JbT4xKLZfcgxnKwPohpivgwBdb5OHyLF
50n7aHj9y6sDwTQBLCJlINnVHRxUga20vJTqp6ljxgts7TySoSESUBUlhWazOMQzIZYNXjQoElup
lcdQyR1qu/vs0vrbr8h98iJ/6twwZ5C/zxc3QgzGGUr6suntsfTbcoNeiyECUhy0niYaw7Fdgbyk
nzhuTogkM/V9LsyP2p+z8xrXBligu1ptd7GKSLeS4fJFYCNnXhvPTkCk8CRwJyf62lAJBZt/xcXI
dkI3idFPxrCEawIsa4haIkqnAm5g7rLOeY+71lco15jW6qeSj+hBkkrBLp6QdDflvrLJwF5OL9OR
8o5FRObCk2724MNkCT4MkSzseHSeLud0JFAmTOPGsY5ynkSo3D/hb6it33qILx5d6qbrPRJmxUoi
RvjQD+JtvwrFiDl6Ulj0hULdn0Ezj/7d16Vb0jtx+J2X1PxPRa36Ssypm+7KP7Sa3GHdi3JiL4v/
wZFkn6xf1FWSV8xZO2VkzVe/4DnpV19bhu0C/pVA89zoXpWNPMhnFUzOQpd6sPkbHHEEBQwLXgas
qNEWhyQ/qvT9+7Aq8cZD5RBdeXu5uLooEJRPWY1hg29LT0E+IT4BFVrDQo4ojyTAt508rg5gTjAP
yBmw7P/DPtmCzQJ5GlSt7iW+f5NLaDlH9TC16VtBmsSIslKDxNgDN2z9cW5DlD5+epjFsEYiCqsN
XkAJ6sEJXPZyych5J3WZN5Nt+Ggau+wCgYnBcFj6zLsq5tTcq5GRPKqwqGNh3mFLZKZHZEigP0hT
rQIObv6fPzCHbrAyPHcKMxah0SInbALnRUfmmlaqhVTl3NTtL5nais75XFD8+Jb+fNIYQrMbkDOT
yne6UC4L2zvfQt0obClBR+rKSKaWyQ9iLoNNaajuVc6ImjPygsd+ppJVkfb587Cc/S2UX+G+U+fV
aUKM7/j6XoZvUZNjUKpI1ozh6HxAWnc+wNYBx7879w0kSsFGDu1K5aMHhBeV+uK+3Nj7kSG0EQoW
kEShLD5MkilwbU8RJHJ2GSD6ynDsiGTk4diJG2wCjXOyHKZfl3RjbHuvYEpp250x4KcniFMCGcrH
vdQC6vBzbNIExhBBmhtJTFTsA/CazrfupB8O2qrl8F0xi915eoG107tXMhN+c3xyxZFHKUkmUQ3O
3QYMfyKs9/+41iUJZhOuwjseqKvpNmyvb9BHrjwZNiosMmm3YP9ppXpcN0DiwI8MjMPdCZ2I3bQZ
i3F+Qx6MhPhXcfSjPamb2xnqPjhyWN87F/v2/wnV2pxfntYcpWHJOXlKWPY3jSyzSR+oXBBAtWmn
44ERQYi3mdNK6Q4hhyuWIVFvIuJYe75ker3cBvQ397QfS+c5IL+tWCSnE/9vEqsdXF8sRDLrxJlL
V4mBjotLZMIg42iFlE8ItdH6C4/aKVzKoJ0wgvjNqKuvV0gwqsmtsHjj03yhyI7MGfQu3Y84hCGS
LfCpWkp2FoR/PfU/CJLm1FPfrD0rlHHJyB2Ksb58Drhu6GI6tLNIb0DV+G+uGsGZ62jFkq2c/NBQ
I8chNvgNTKlY2PJakcSpgQA7Fn4w4SZbPNcREQ/By0265Vwg/vK1UFvVqmCCtlKmNLH8nm7cHhbd
NHN7cofGfIk1KLmCsAYSIzmm2aPv6eerACyUc1EMc8pOiAw1KYZ8J/eZ5Lr89h6VqOh6b3haaaQr
8ttaISMJZpBWqRILwHQXL2tPqGQ7c1X0qttBGMjJttpnUc3zBJAe1i/+CIuK9M+AAuCwOe5m2H1W
2rE5X8OyGsDLo4G5RgnKcujWcPTznMJi94hK1zHDVgOpGF+xa1j0ctneDu/fM5vvld3g3TJMsbOB
uL4ZBkQjr+MeAaDWj83JBmSPNshjAU8vWqK8fjqZlyUMaBAhllWEFvc2bKxUODkyYiobvI1zGbK3
Osg00EiTCcy9ZdEJc82T2DxSSefWzCOItwhYHmOwLjB1C5R/XgEqsXQnfE89mijuyOYmQy50fZjv
7hcMBTzqS5mE/Pviqr3ueFlXZvSIMaH1EpLootcTnKXBcwb6Zoajy+binPfLqE3i8Ku6wrbDNOvw
/CnNGivwZH/VOHhDHYJYFOzfDtIrD5JN5vEmA1Ec+BX3MYasLRgpe72phpzG1P6gp2yOa3GpCttQ
fpd6Fv5lKTrnL1skwGXWLsC5au0hO1F8A4bJIaFPRyRFDV7rD27RbO6aN+TiZ1efSYir2KfphSBv
Kmk7j8KGSjkjcU7QXXORCukl8LWWSa5PzolLAlifEy8pTk0L+3ZXZ4JsGBeyTDTD6CGAVYgeYOd6
hLDdvnjN9GIakEN+kPMcMpKTye5XRDTy+nisgR/WQLAtMX556B/+mAtOOFpmCuz2vS3fjrg26kCt
KolrbtJapPEW5ITRecElwK+XIg4BFf7YYkLjYmhk2tQ+G4Zq+TffUkAaBrW7RkYjl3dSk6NknzDM
y4Lk54ncC4/rXf/cT0UgnK5uyNmVHrmZPpy6c7bmjLI5F5a8dyM7WJmllxn7+wQqKoNdHLFe6LfR
pUOUDgrCUpXh63ypTVTiMMNjjj9KyyBjgtiCidCQDJ8kLpHGTsS43pGj9ZHviXev6+PiVTeECJid
4zSm3jRPifd7JCLoCcCVR1WMUzDAiV0iX0tZhplAihANyOJSwouPhIPqRT5acHXoYcXKaAFOVP0Q
PtpCdzOYOtx2sWzVzjXGQWrffGNVGc2qmIZmEf5ETheYPYmeYu3aS6QqKP9u8LhS6gHyuDOgAopE
FKE8Sdo5OiSD45A+cv6V0lEo9JrYWzpWxlwTA3CzymXJULkQqViSaBTXJDdKH6A5IIU9hvQWfvvn
Jngp+wP93ZMXeDynXI6ZJ1/mXw/nDDuF9FqvvTaYSVwQtNQV5npcW0LTqK6Kx6KPxE6wpWuz8kR8
c0MmPf46hc+U3zGaezgyqxx7mb8EG3R7WzSoulqnKJQmVlFtZjJ99rHFqNWmzM3rFUEoOGlMJsNq
hOfetIllXq30+ZJ+5S97ha+y7CjtNtwsJCLlFlS7PUhMMdKl1T8WLGwDeCf78+Za7BpVaJSF7TCG
um1kclyZ3R2Z4huPgIeK8UVLvTSkk3RJGtRaUdIg+0Gyp8Tz/eVrbtbYHKa2OrAiyyBQgb46QxbD
iAySiNV9/N4YIUop1Wbhfj9nVCUuo6JuBq9vaBmpitHgJbDf6ljtcYg/NgWxXh+Dj9Vg65zxo6SY
Eyf7shtjG+yvXFizXETQArOaxJE6S/kOO10pd5orREnV8JyZ1hIXhgx5ynw9NUx2QLhRbLody4+J
bw36mRobW97HKQupMKdKVCRDkxbXt/z4xCVVv5hqei2GD6ks3cQFQ27ko050Sul5nD1hrjXHQyFS
Vc4+qexfTHKWin7fI0rddcZwe+Uq3Bvv/Pmd2622a8SMhULW60cqs1vAoFVBiQLufm3gbzncVHRN
u5fx+fx7zG7uzBtXAPrFPS8t85ZUCaZeaCELIVFmTOaA5HmNnM8MFEa8PUxWy/PbJHXeZArfSK16
CdU2vbqOTXWAlaB1xXTxDeNqVOY6mQ//DNwIUqit73bsZ/i25yiPs10Rg2Gc6wOgOPvOeNYbLXTT
3g2v6ExNsIi/PxU/jJWuHH3bZRfUxut3piaOxxXI/H3Wo28dvMc2LWMHOXrHG+yXYjkJJqZ5QNX1
210djbVG11pu1f52FvpTvf1RvxnHpVO+Jb0ZtXBgU8HyiXlNSOtBLldYVRgUD8iQktxv2NDH5Ezz
fCSmqhv1YpQKTfeTb9qTum54watlFFzqit/JnXa21HRBLjBUfWl3BOixtvctkkSziLNj4HqUsqxN
exUoEr63vbaqRAJnVq6+0WtqW3BwClCf+DM/Utz3SmMO46SxXvcGuvGV3zJ8PQMhUD0XGMm4D2tA
zf53N1lSV+RUGo44r9HGNSVxyP4rbj+si3FopS9G/Q5JBOwTa++Y3Oa/5EZyOP6kq3AsGjJOzoP5
vKp20OVk7qFcIu/6wGB2sLgMbvb0JiRgXW0MMffw04sztytw+LccL5rrbk0uyv1cHJnkIrHyGFOR
C5YwrtM3jOENSW3jKAIcuZPgJhZFJdnuQ66tbjSF8JEtdtVUYP1IS9QbfuDSQL2zI5PZ7qWxCzkR
ZZ+xB1cVctHNGrY8PDDmZZzZJWaxTojNRnrWo9lvO5SP6xLUe6N4wu/R3ixyInn3hNIltiAjn0Ou
Fyogk0oiocukmUgzM+nFqvm1S/XB4l5dN+fKypFZh3yBIPgyeUPFcjyD7Rl0LsNnnsvD+t7B7AIs
awLA3MDxzHXaUyQor/xUzZMWxGz2GiI1x6OhZdsVwR0+BmQPi9wgeShJq6E2vJRIyWiH1YY2vj+c
i2klQEgNpWkRcgRyAvf430DPxzI9nbEoxN20Uu5g2sm3a/yd8wWRZH7BXLwtvTszVh4K0Y2r3pjf
S9n1zLgKNGzRNIoNYLl+ndkPuti3hD2GLv7+3mUqwVTDrwS2iKjW5vrG9q1WMNSRQ1pFQOqBW/Kj
2swLrEJ+5Bw3OI0IUuHFafGEcaX3EhrwvnLJxTmSgmvObeV7ZMQJrQ6tAdKoT2iWZLElfRYBxtv5
T1ywdYkwZ946FNY4fftwaE3YZDKxgLdP+s+gVJNJ2/SxifSrYqAwhkHlnZ0cNLWDS3RX2iZZOTYe
cMTlEJ/+J4SEsJBftXvclfEFL6DErC7jpBAHPAwpB3yf+eYDxih+yZY/3ulGyOy/Il9t3v8N8lj4
s0KkLXMGakXRCanTIcCPn7YGurACxeHcZ2XDuMraqwl5jI0k4S+juh+0S+R9t8iEHYweMp2sQ83x
kE+jeGYt8l8//AJ7NQn++GtiRJ9ZDP80s23TEvUgCWjCj87AqNG+6JItVqh7zZR+oQThEzkXngyG
LEMWlN88nRvLLpWPqO1jPuLDSDbbYkhDn1iKxONroAJyZ0Fwet7RKePzEnp/uGit9hoPbMvG/jw+
TMKxX5bprNu8T+qRvsaoO12GJJOLs4XHI/P970lNGO++bD8npIrWbOVpw1IvtssjZsP+/UUYuQyk
itr/g8w/Mv+vxo7XjBhTqsyhKGtkh3y0Oq7geJQdZqlfC1+/BSVq916o5paUjssrP0IpaGXIxQHi
xslhk24f8lbXEvy+aZzS/ElKHzldlFdlJUXvsMO7taXjo+gUjVOWN9VYhdF/6oSLiGB9y0yO9kyI
BgtWgy+L/qIu3YQIFCAp/CJIIoV+P/HUsLnu3/hZHcCQHLzADcWk2Vn48LXw+Zy19pRe0tnrrh2C
75BvmA+Vx2Klcn/5rlgpIUrhXo4sOzQPdGJFXCOo0ouHZlOJj0LrIUSc1M4jXYiE7p4ZR4b60JbC
fZcms27a3BWQ83iwiw2oJCbrjGrGgCFKG3li5ggUIaxZn1wUpizavBYljndHB7mdKAWtHGVGcofm
l4PiSf+AhdMpJ95Kcb3J0EZdN8taLyHGMuuKBOrK5GlAX8CLCICN3MTenDGVO+PetZiGc7Lh9lAl
3eMVCGZ097rDJq04Ysj1u0ksQous21Oknt3u1gT3s5Lxde7ftVBbkfs7MUX5pJelOPtwXfUrSCuQ
GrjUa9aM/CVSYJF6VV74Y/pKOUVm9tOfGRZdReY/m56IdTCvsQ86ewh+ContjKbvOXQzXglfIl4I
WSc5BpTEXvIZXbKok6hd8cgqpcd07uAdbMRso+D2Y6ECD+SQUgyQztAO5uRXb4m+JMDFUGganJ/L
f829HPWcpSn6YsA3lROAaIWRbrI6tZsORl4SFzPoZEZnfZCwOlT/UkEm5ITEg4Q8npe9VIZonTRn
xp7vE9gvNebbUMXVBpQ7PfFPmoJu2kPzY2rpZO4i+M1ERqtn53Zjo6SBSM6gj3mRKmtAY9XvRCmw
9fbcgeoX0vF218gqgor8nJjRznS2b9f5EJXbsDUb8ThWNSa2J/A9FFi5cVlGnFNPygNaypN0Oj0O
FdjxUxGh0x+PVeiEOneo5kUYReHwUA6UCPQ7X4DPf1JJZc8pFNeFAwPuJQfG+9NmT1knI6YblBr2
+CbznLep+IgrRLUuGDSPLF1vq18QTKkvTiG5tpmbGPFsbK/4+fGFd56lONFhyFLOG4uRm9Xl58Ap
dol9JvuCd7cFj6qyRmK9o2q2Y4G6IWaMEH3AguEX1EtVwHXWsSAJeX1KgmJUI4xkSeTFqEPIqb0w
bBgHyGK6XEN9CI9/CpXEy/kvwklE7WOenYKETJ2S+0idD0tAGjIUVY4GT60ukKEBd4Ziv32uGgTZ
MEEW/v+5JtR2fKjrG6zuhJu94rdNzOOFuWMRwuYLX/Y6Em6ImxiSQgqXXtnQiQdwdlz/hu1Uay95
y1akMSmK/D9n2+SGpTEk+lQQ7h2Ir3Qm9BA9+WSkqvGrzS/5866fES9se5ZOLI5ZNRLtApRlbgVD
+OWtTqOiZK+y14JQkWdLC5UCdA97gPjV00NnZ6SkXkSwkYNt0r64hSaRCLN/g6v7JcqpBRPim8uG
Fha6IAuZtKAJG5oHbvL/AB43nQI/WYE/CbO35FMT9IimA2M6/EwOe5XyUfdKHfz8o7ePJj+eRDiB
aciTFuSApLSrbNLzruCCh5Qugc2OTLU/mYwYwLkPtkxFbqKN2JAf/ZtdHayl3nRTNsYWkyLRiX6p
dkbCy7yweIkJmawl0W3YaFOk3Fkv8ULoUd9Amvkmf0H4jAj5Ptc4MnDX4doIzBmxyUIS6HSYMQqc
0RDp92clkiQEY9OVtGSroxHZg0KUyhGqgFy0EB2Ej2igc41LeZAV9e+UMLvAMfI4ujNXxVcbwC7F
3/feiz0vQJoB5kT1V8lXL8N5kI5Uwwxm+L+SRnI48tLnYToWyvcyDI1SDRQIIPM8E6AvoauDXURk
SXJykUszypjsFO5eeBd4uiyA/c5iLFqbtGDd8cmSZg7Yq4ny77ubawBUN+hxTq0wsGAtHsiaLCiI
EpDZpWw/+DX8dk18K51X8IKb89h5m/l7+JXSl/ZLE3wI5YkK+Oe4RkKnEeByh+f6oNobKxZpGoga
pl3HZoGWFJsKmtpy6iKrZy2wybrkPz+uQIlkN15Hy/QgT+VTlyFI6OwNWnLuVVNzktIq6JrjPp1/
MinXOroqHpF6Y/y8g//QQ+kWKu9gcV72rBsyTpnwH9QJ+eccWqRlxuFmQUOLqPY99xTi2rGWkF79
c1aJwKbeFH09uaigEqlV9aKW2pi33JOHRdu2vFcd9aabBT006Q9a+pLyjsA6NoRCi9lDblHria2E
p8cEuQJ/7yUaCUnlqM6kwN6kV4J8ikwtuAyTgtWj0YhBRRQgvTPs91BEw9qE4j/rYhFUwSsAzl1l
zv1kAGhcPt9GoV8nd3b9z2+zZsrpz+9Ka4dLOyy6pikOy1eU6bRkcW8AxDTR/a7DeQJJa63yZEzI
ZKYKClke7XOF+4ujr/FYeVZ387jDpWM/SxnSSWhhWFVnwm9OXqyyNKnnMcSCNRU8wLB472aeUWf+
f4W1sftF7egYpLlOQe69d/EZyhjC/M0Qr0f+NE4UrPBxzj2ydq/sFETpFDdL+F7Mb6uIDXieZ0ly
L+bwv4x4wkO7DG8dArCFHXaUSMYSkvVJioADM5MG6VzruhE4O4fmpZGm53f2C8NsujSF238Urouv
jL6oUiElawnngA6gg+p/IRSN1fN6IEG1XfDxaCkjkySgviyx/RftOBrkqGZGfqpDSit8MhjcK4dF
hHbSIFS7Gz9Heqx78l4FvnsFOwmtWoAsrK49nCmZjZTyCbDyPIGvG/sHwNIRFGRLQ75gGNQttw+K
eXU+nCbHpw4Vw1asLU6ajbuFT5mD/Au96KsN/6ikuRDqmtDlKMbn6SvkI1FN6c6/7VGCKmmVOjm/
4GyeJW93wvYp0+l44c8F8nBiSmfB8AJQkMlqfJ8EwMNy8Nahgz5OkVlvVgh1wCabCiXi8I76AaYh
8mAL++ZzEq2zVCWm4er2S65hd05qkCH4UxWAz3rvRktRHCwQseO6pvzW21XsyGCSAgI/RiSfdXhT
iDYbLFAz0qvuZ+3iRO11WBtHKjToa5GZr5n8P4vqbMjdivecR2rZ2FBN+UvSzpCoyr+3GCrfBr1C
OPzCstu/A2nnSXuietNZZfrMtg8ArqScZmV2AKjbmzuLG2IDBO24deS0tpu0Gy72j2k0pX+bbS8/
Sr9xitnTF1R1zGP9peohdYSUQmVYww81jrToumeS/SfvwZ+HZYTvuoBVji3dfVigLoW0yM7RnWFF
F7n635o4T3boZBKItNhcz8TZBSrZ5Zvz4y1Ky2quiLkLFdkZTpqHvdSK/cNFAyxu6l0PgZTvo8Q+
PrTxjDgzfJSWtNip2HjDq9A0tMIuA7PK4J759kEdE8aymcUlCzkPO1+KRiF5P0sXBBy2G6O9PH+m
0vcu2DAml/520ck+l6M6zzvU0lYzl6qm68q8erQ5LJNxOAvyrOQsPJ4bkc4JFfWQlZ+3TyHN8Cq8
kngm37kuQvorjtnnH2Tw9QEtVjnXjA23mNF4PGfZokuqLQfAhdiOGaCHUsgc+0NGsIwF0JKzO8jH
vFavLAKh6hWxKZ8dsB67GyFdyUfMQe+U1T6pNiWEishkCeux79w5gRW+k6BU9WIQz75LqeZKKSv2
dVxDnNmpv3irK9TSFBd6bFnhJNuCTJYBh5MupHdfiXeVBd/oYyEHzAW11qu8OlBR3GWwxdRx1BKS
t9jEGXW5Iq7soZDjaguSy8sW7CNQGNDnTR7LyD6BQM8G4lKSNDQDLYdgLBwRtV8HjNJCp+eIdqFB
28XH6bz5jaD+YtWaHUmkdmiKr47y7KW2p19GAZZMPnF/CJcX8MPE8iYBuVn0IBESYJuuMF8FkgpZ
0heDRkJN/FIBlHg7Zw2I2myb0HbelkFrelKwGQeA/fzCF2898EKtc/EbLIVomTu0xY1+tFLTVclv
5+fqE2rvh8a4U8XdkAgrd31YNgVOtpkdo/ypbYB4UiRKKIGjUSI8P2pi1X1hGI7Bv0985JSBSh8b
QNqvemDAi4mvAmP0HEtJF5mJ84OYAFIlN0Xl7jz7CrskwvS8kxlf2dIIttxIuVj/2xo9Frmjd/yY
LWtfn6PXUboTVsQ6IuHLlKKs6quCGSsYcZ0tUVToBNWePUUcCO/MWSfJn7JMcRyHcKp5x9M+mRzT
84Kz/YUdgTpV+qYtQh2+I8s2J2w3wyGocEyvQamB8yvTqiVVH04lfU/BKXD4TMQiucLnPGqPwJKK
XqRH/jvAA0UPXm+GI20qzPRqEFBi1eJlIIXYISThzXB/15zaoEPqjNNAs2+6sBNnqy0AFxaWfgFH
lvp+x7DhbM5JLegac66uvWd8wgRWjeOwT03XkwLUdY0ZhcR/QzbqgltcaGtGoDkqmKWRVMnIYahp
lv86OTFqxvUT+w1v2Vam3uRreD0lBdIAs/jL2YEc2mQWCWNw5r3sbrMWXEubavlpoiMdnrpzDtxw
M7pSSBRZJVysA/RvuKuBZvhTg8NgazBdtL1gtJc9PlYy899d8Apk3lUQobykjBEL0edUSIt+WnNv
IMkJCCwrogEhpl8Ra1oxSUidsvuUpSdh0vRqtUdOxITWd7EvLrovVZGyom7QA+tHRjrFoSY8oIUa
yXUcFBxVMTQPdoF7vTttyUl6BLr6FhNi23sOwXeQfAIFDmPjtG49udcylXgFm7CsREurw6f6o6Qa
76Us9qf9dSFXYeo65gG8JUxz2muOgl4nfKUIwVZq0ETIH3ksF4NtL1YqzY+G2dsJWW22KZo66OD4
t8MxTEe4iZYbZwNqlbOrKrUYhjcVMkALWrjsG0YrD6R3dY+hzGJW32fFJRSEPxMBP9/nGdgd17A0
Q8ydqtpVwHbfLbD6NEFeW6XMGm886aLCNr5eKZHg841fd9S8bdySC3Sz/uKjJfozZA8FtkZNWQv/
Ue1L4Pwhriz0IJKE/A9Cu4TnO50aR+2GZN1R3ETObJVH0InT7kT0sO5mLuDVu/RDhdjY9boVOjLd
eFTYS25/fqF3pSx8rajfJ33Oda2dKZpK8BglvrhghVUUlqR8+H6vUf2sjqjPIZw1CzfR8D6W8hyL
AvEWkzrRrviCN6Bn57gtfLO88XHWqP2B1ttaPzrU9iUpRybnn1T9M9gVxNSByxyLAgtVhp9l8z+f
8iRjiSVuE+4Mgpcru+aiFQoEK0oyTN2ZmzzSF532cGoRA7wXy6jhvu6hKnq5lmaPWyP7w0v/b9Mb
TVbL6afXb8Xe2zEQfK94Lu1UHRAzTqWqSF0puaAbVxPqaI9WFrXHAseFha3q2qMYhhdgx/cdCGgq
kdy5mY2k2JGy6PXq6q/ef08+jZj65G9egCjjEaAU8MoyqXuZLqmb5AP5kRYd41b45KyxEV2gP5zL
Vl3aHJEFtIsleVGLyYuSHX8n8InqRbQiR3BRMaHHzygIaoeMc0EBMST9cNm4wvwwidlSE6ozAh3C
BrvhXHs7o7yjATJZ+fS4B3VhVV4qpXilIAkWMkbaLra6bRhNuNvh4LiUEIq9xGs4TLpsy6XJCu5u
oxhPvTh65qSoLrti+PLotvL+sFZ9AXDmuMaqD1zagPJs6eK4jq5p6R8M9FEnLiURcL19HVMxQWEH
xvEoMK7bfO06GpLZtLHuCDOd07WSlReR6n+bU6rFZt3HVtt9lZJ6HnEXT4hrvjYieKHpSNQ91vRa
wjnlixCtCZxDKWoh4vemfpKaOntXvus5W2CHIcFuMLdQIlri5jM14AJPsNRzVU63g1EJSJtAMgTX
DJFsT95pdnLg1VKRSsHlHaF8HQiIO1HgxZC1eA/Tc5zmcKT+AZL4rJVpEJHaOH/nkNHT7xcS/1/Y
6NYDL/GbiLPYxr5LSypOQHTs1wC/H3tGL+paqDTMAmfLDCuZobwJgng/0uvT4eXsmcNAwZUGJvDr
xI91YlDBPtz0Vf4IzUa3QrF+lJYuEvflIR/JmeK8fAK0YoAlSKX6xOiVQjxkHcna/HoFBClECmyt
txqcyhFlAr8Z8BNTv2lPFWZei7u9sNwWLXVjs2+n1wWOwRHwA1jdZ/RAqDRmLVpBcqBiowhYN6vK
n31fNvI5yo70jrEQUFpxgke5mQ94ht4IA+cImQVELALhPNZ7bEWdblX+E5cOYWogcjAM8WS520fI
sUQMjDDoXeRhz8XgP+HPmOV18z15pHc8fnIP2h5c3qSHbAv/BEn3I8XOOtbPVaRCW2OKzW93S10/
j9UmwG8V57EuIc2aclYPj2H3k6iI0/Mlqm6Q+lkyFUhv6YAZfMR9qWrkYMqpDM9oR6e3uDgqWkkX
zduPrLlX42QlSfD48DSqVR3GAlvSBL8zk+ELgX3S4bMnzSupLyBUkLBo4nq0VtfNK7QVwDapMrQt
8exTORMdpu8eK3KoDX8tmrvwXHY20RtUsDK21TZftiBDb31cicua6+u1y+4CpclsOUond7WTzAtn
neh8UKP1s+D6E/OXMQ9PzOI4WWAbsJxMnPxYC9C20G0V8jQDdeshBdO6orRg1a6VEB3bMHQpOk4k
N41mMwgVHOoAtUGfE5AChmsue7L1FjVI6c5nKYmeYRLQuRw32g0Q7AKpK4yY0empSsmXMjo6+Sta
j+pdmJMDaKjCY7nrZnf/oqT0GTUXGyfKJWm+W+9q08iNtYiePz9AFiuFKNDLSKtEQBiztcZSzuup
HTuhplQFvkzjR+QR7GPkHA3aBBfhMW+WlpN2gAYVD8XgmRKf9lP0DNtJAo2wenMlVzcDrm9alEIV
NaGfccfkagDznGIaVCdS6YTd/ECd8qNkO4lRok42BsOzbx8dN7/WI9OZg1USWIR+DPDbhmlV3sPi
ZgEPo2j7g6xjOVUs7oZyf1zgDswkDU48wBLGjx4OL/lAy3mgTvG672b4fdVF7z6tzcBJEEp2yHUI
+m9K9r3hpVv7KgcNT8TS2j7F2TJgeznc/1vJKK2IjBhTV2w+OJ7hmKECgsMfpKXKLseqSnjFi92m
dpfdiLQIghsWh2ITHGH++OYuOxiamSXIKBwEecgpi4gKt8nH0u7DnYB5K3ouNP/tSWK9WxRcor0+
svnIgXUHoS7BihUmGRclIM3jo6114H4FOSnW5vBZ8WE8W8Qf6hjgWlwV78QGv0CNf53Zhi4B2m3Y
xMkYpa6617N6IFvEt9CJ4k/muCOhhdi6eiuC6k0P4A3XavVb8J9FeGAA0Wt/aw/4qwp5ZWkNJ3mo
eB37uCBDVZ1opGiYWxSr5ngyNitHxpHJTRCZgzZjgYvHA6SKr5yyXnWA12Qc58g1zy7uz5z3bsyv
rsy8pvpQ1To1ODmt8ewZI1uwY/SjeMbeo4594eiRH2zaZAgY1Wcf2E/QRi6D//OR1aiT0k8lenGl
OxsibtUH3j5gxTZw9z+liaHztAfpF1tX6FMFqmbphvcfB53x3eRHBciQQVa78EMTMY6WYPFJeO0b
kLJzCOgHwlOpNn0vRnPLR+xiBb+DBZ6aU9ulaDqSNNtR6eRx2MU0mhkae+6E8DktI1As64mv77Dm
vTtUY2InzEPnUWgfpyLWZCj2blE5zDZ5UgvUwWps5HnUuvb0wJfE3dgvM1y7sNGnE3l5j0yq4bMK
e95lIK+8EweFbRTjNP3tXoWQlgDktj0S5rDl/Vz7ACm/0KudG1BaRFicoTPWtC7JrLsMhR3BSQQm
hm1ps8y4sXpX4jy4TgLUTL5BsJrldHooybtHNT2vCwtEhlMWIviZawEJrLQRykSDSh7u0pN2QxDL
o1RB4/9LlRhHU29uo3RwAXIoxv4WmeVztg2BRhckrtRKWz0q08lw1VF23teOBFYAiwCo0s4a0Zrx
o6enAVAaGm3VBku6YvaEq7O0zFNmIRb4gSvj2VJScoi997sy9bqx84ckqFCOez4P3ip4WdN+tOd3
u+eqdqqHzJ9IjBx/cepHDSm+kmkQF3QYIzXrkopoDQAPtsTpAr1EFIv4eDohuLhe8vMMvYl4LfAM
+G7tXhf4FB5KiKBFfDIT2O8vWOUp3dOmBSTSbe9zDu2tg6HsHfO79yY/IbIXGN/PGhS9kQwoy9L8
mkjLT7xqzgeml2c3+w7urVXjtxaCWp8RmS2iPj2qDvRDJD67JykJwcpeBqdiMrEPQ3FSzd7YISZ+
c3r78+z222ETjj2+ZfFfdb0Cw20Cd06NWuWvmWQJnC5uVkyl8i1L0UXpEsgmfyc433VzkE7LaOHL
a5THBsm3BbN6GuznRsgSgffE0Ja2gFLbiPRpbFioz7onbPu8yBCYgvUeFCoA+NZLL5wV9IgfO3KY
7lVq8+pLSeJePWiJ9jeLjjFwFZaMDieWPMn4zsVXXdfm+NThJgC2A5JncILV2NG+FHkzyTW2kd4O
966K05/sOzyr8kOTb9JpygWEiEJDUZMC9/8e31T0/wjA5+X1X2FaL8bXcuUzljnF8dWJU1LS23Em
CGiyY2nX7YMF72N+BYX+N8GFY+UZKmkOSYmMYQTEyWjUdUAfL0txeiegMbZEU10E5RN0pnJw+LtW
OAoG2bBazMez0gtoivMGXOG4CeKsihD7z2IRHDwBI0cYSE0MrTyWenK+XbsEK4iQn1E6MFHFlaLZ
C9YktEOTlqYwE04jFrFnMWNG0DGzhK7q7kkDSy42O/op/Ygp4lJom31M+pxTGgVeyfGSD67FqDPK
XGI+aZBcN/NXaDxCw8H6Q27tG1ZOZlJf7Z+iZFT9KzfeylcDtqs5rUApygM6JHeeyVxmBcSqeKhR
trw+EH7R0ls5r1oo1Zcx/aGgTro1O9sAZ4pQWRaoJqoTNhz2xv9Gipp2adBhXqInQZD4Q4QiHQ8u
WFVHtpGdpjTRf5UsS2Un/13hSzBM25tTYVRXMMvFHYrNdC9Ia8KmCI5s3Cnz1oln4psfKTEGupjU
a84s07iJABSyx2WleHoiHZ/HNeeWuC8qHOYqB96m4RaRsBs9aXorGey39s/OrGgOyvETBu0zM8jS
5NkyHuXUGIhXXxcU2nJai+fH1/Tx0t3y3HkwJuda7tjqC+4ynt+s7njzrKx1L1Uz2AUQW2ulS51p
xv/5qzm1ENLQXZTUO848oX2Utlz7PYmV5hgGJ1axD33mAL6XUkxHH40kf41cWPiafJXs5Ye4IbBu
U5t02gZLn4oCZwq22LkCaPal5YTLbrIeIi1c37fxPhr+JL2v1UI/q+GrWNaTNsiT3uIq3yjQo9TV
6ndyDoWIT8JHsDSMuVQefxioNYeo5PyD4f4vPYqbDObq2wMlfIn1n6y6r0sNrtT8IIRSDXny7Mwf
dA1lH/f1Wk6zzkksUq9SifenfBK+BGALKD159YzaryygIo31o+7ZNBCSF8S2Dm6miIEZ/A8GraPG
8Mg+p55d8E8aHByo8gunjlRjbgw8C2wUh6Ne75pKp0QqenkhqUU62D6nMNARshrFZ9GqkYxh+7I4
G8NDjZOFIGjL4qR19O8MXTJf46gFApc1RUdqKf/ZX9Brj8d/K2RjKxQszxLLKEVUrE6qu9Mdn0Mq
TTYrC4Bp4ltZNScpCNi+WlJnpJA0G9azarVzJogPUhs6QXAMrqNaDHX4AO25rN6Wbx9WQ0rwhl5O
Am+b2LwarF7xtVZhSdZ6gG7nQTep4Tsrzft7k51U2T57NBfmWfjW7i6loelu+uk9hO9Nkyke32DI
/5NhTqGvnmE6bQ8rn6HviTHG+K8eyn3ieDvjX7EV84ysdZ/in2jKpxeL0bagsbA5dLFT26B9SeiH
vn8rhZL5gBu7SvSH/OzdAXy1qqpnE+P6XCVtEMTNc6Ey5hVlP0HTgFx85pQmc12bPaZqA2rAko81
j3uNvqZJQMXisooH+it7y4m7W3YeWdaUPS/1D+qfMuSfFEnwQIPRToZGH0F3qO3eZ8RXcQniNXsy
op/sFMBipKQmfN1Luibh4vkvlmvgc6z8kE9NcCc9hC2cj/fNKYiPu6EDwTjysOhs1e5BAYcJ1/Jh
e5LnAyA+YdCoKGdweZebd389E+9MsXX8kfMseZ0CeZYAayZHz8OC40x+2BdOaOGUZGwgwMFT0pai
IPlOPSYfTDipO0XF+h+lGarRslctBMtlL3zO9iXAAO2OhMLJxEY7tnGYUVRij7erisMVGzUxaUS4
GgHLHzkKDlqZKT6Pu3IY0YDLCWSLRGDbOK4AfPXve60C6IW+qlGaq5R6er2mV+Q3jaAAsELz1S+9
vCs09TLo19Tr4d8D83e1/wJDZfUQ5HXWTqoY7B4YHUU1VtXGvqgr6Ac5cl6H3ciS/trOHNk5z3i0
SYjjtB0vxsQvnge6fh72Z12pOLtIrMb/k16Fk9HbKghmtjEtt7LQxUmhbgEiH35YginMex/TLBsK
3cIlBWexK2oo+eBUlyMyu2XqyrEAnWfi1+BfsC3uKerEdykFsRq6o9xPMaYKzRT73tVD0aOIc0IT
r6gfQYWhIrCYNwqsoMNvcYGyEh3g08AxFaax6gEcIjA6LR4WAz8UgjN8szi1sjcEJn13r92+L3PU
xDov4tWUklZxHelCwNYZZtjp7cwdW7mQpEkVhgIzcT5z/G/EeK/HwM6Q4Ky4c0e3TCFB2tRZRQ6v
XKbu8AFShoplTFshOkdMz4O8zB3Ylvc4XZuxv49j7BuWkY2MoOh2yMaWK3SOC/MmMrug0yx7TLtB
PzVFfQwtEWftyhgVqN4TBu260YqtXtzsC2979Ui5queXutkPjZuUkmQcea2qWqaKjtCV2gFHvu/l
YkFOSwQYqnUfVf7/j1VYtavfNaba3F9xV9tcvMwJ/4eR/UzTeXgjbrHH47aQiyhRhWHIBQ6EI4Cl
8+9uTjX730NrQRsgCwZqjGgtZa/Riepb3xZwPONVs86pmUB0oAoHK0WH5R2vQtYMX2tILBOJRPaY
lxPmtC3vRXh6EQs3GGHmKvI+j2NBwi/T+xJb6UGQX8s4u9czckk2PjL+ELIM16nvk4lnK8MRu/TE
lXIBn4DpdHNDgHRUJfeZHVggWRIUMPjkwcOvArTb9DM+QiWgw2ZbD1v05yMySqZrCqr5BCKH5noE
a0JjgltU1wCAlpuju3jQSKNQ8ugJ7+6457Do1ZG0olpCFaN7aKupSqaBZjOgVYkqGP9/3DoibGUm
Z2TMFJjRb5i1LwP3bwR4GdMssZloqkIcx4PdcbhOnbKKmF70LCJaA6+g90RyXhwm9uRr76/bJc44
3GrGfsmkP07LFp/+6iH/I4IJplkkYJhQlySC3GQbHUT/rgw93ZI48oVZy0fxvf7tTXg2Lg1M6HJB
dCrjZ/tQ3uGADzbpAbZdDp+k2GO4SrXPyMo//coNnARgRe/ZsdBIi3jOA5TQ7ST/FqzYvoX6/CX/
53mcuD2Ol4UTEVByqi5KLaoUTWknYbGXBlMpbILA+Zo7ErTpL1rh5IHh/r8km8FOD1tvQbH7s0RY
W5r7uyjKUXvVEa/r5a9py21e+PYo6AaAwIGH08/s2QAV4wCu6ovK152BbxPenzoNsaH+vmj23Uek
py+qj75rZ1LMeTJcE3Q1N7JkkL0cS1a2yTtS4EAr4sLyBZ6UMislL9zDz4K8GP2oZZywSvZbrOEG
H4g6ciwQtmHuDlWVHZDfMqRLNrhrmVv5QfYaSbl1IzZBq/8TFDrcY/5A020pdxyfZRdNFtEXHGdu
bV/bLvmA+3tpz7pidsavyMIJCgyoWy0jhl0bdTtQPJm9eFmrAHi6NmLHXhH8JeduBOBDZFnCoZxJ
FJfd8ysflFOcO4o12gIhLZ3PKAImo22dI4CiwoYIlirm7l3/f4sRYb2Eu2dId0txD6tlGJrq0eR+
Muu2XCdXanSIaQ5OOlamUBHiScavcvJg788ETSiMiWMqLCPuT+b0OCo9ecedodlAhbqPxU5PyvVD
EGDEsmzQNaS5GfsAd6FxBekyrgDZ8GSvWcRHLF2hW9xrGanmYTpxckEo70jSaZPCJQJ0/2pJeXgV
tdkjgVbV1qB+y4mJ/1l+KaNNbHloGHQG4C7s1uc24U4/lY37X8HTDfw6hzuvcfn0bu9WtX34qilF
UZOGM2tic37e3RzGHAAx6NZgV4brSpLFXXqFIE32ITOXr/hNHWsoUzAIYXymWh6zETaTDuZnlRj+
rizeGXM96m415CcEi01AMshCEFluIsRS8fLZHoU9B44EoZykOa6Ty2VNeotYGmjXCCh4f3jBW6F9
3EEz069dCUBRUv7lXUpFtpke/w/w38e641nrWhwVt0fWKOKqvMzyMhwRraU6ykGlsSVWwTjgIoCh
i/cvovnUPeQ10sOYVi4xTCh7y/4w+CgVWI3oeSotoURsbFMr6/EPqPHJWaIH5fknIIangg7WGMXc
8EU+tfXCg5NjUDjcRjQ3sX7TS2MHps1UZOlo4af/fyg5L/8lFDDv1ZDB+iFAVNq+v3BUPiFIcniu
31RZrWBZDAivcyooMbVU2o2axFxgnmuVM2eLChquoGmlYiG2TlKoBXcdAILxYg55flH7hbVIemOj
3AM2v83ZlgFSKPNCWkhj8wLdn5Yl9Y6KlaD09Kx0H/8z4GPbTZY7SBZeDZB758b0wyshOH3hpA6h
r+/Oc7cgvbubCncrmtxsNTCKoDB1zkflWC191C673CzrYz4ybzUiSwbVYkD7GEgp8TrN0+FmocjH
D24lojRWtVhy9WWUGFuBjW/EojdZik45UwelF3ykbW1fBBSBBUSYdH0+f+y1eq3WRtHqPUzZQGjT
F+rUEIOfxgIBhTTzZlt/x4xEBcm+XXlVs1ZSDyhU2sPSoKDucRDtNxvKys8ZrhMu8Uko1XYffeLk
goiuHFiT3PFMIS7K2+q/ztHgFff30H3YEGCojOSP9pRmJfa/P/7eNOZGXTp3t5M8glhRqprz+hBb
81E7WnBx7O+qE5M16ZD7YCaA0qJDanNvxXOwuHiPTywcCL+Xr7qB66Z98dyKk56dj1WbUXNx7osp
XeK8kcZfCciFe3pZs8n4WtGX7Po8Pj7gwlyjl9VLHUAl14yliQoDfd/U4S+67DZgkPz749qjEj2A
MF6uZHFUVpin7rYJ39A4n09boFdHldZgILj56xv98uKMXDAN3gZ48cbGacRk4M0v2THgzVQBWgiy
2AiDuI2VDOVvxKVcArkmxg24nfHSq5qCqYVBBivDs/zIv0T/v5d7YDMIjZxIbElqT+KJ3to5mRgc
aivdbN9ab9/XK40TcoHIp2gNM5tw6gaNV2QPACKSD8WQI8pcDRexGvsKveaMXDe7eDYnYWP9wRFh
pa8qOfIn5ryt4lZSW2JDF4QxEOqbt22XQ7z6nLCm++hOGSOBun0YGX5hPUVat8Un54nRRRJC9cBy
yeIOCGd0N2dQdeeLOIxOWpeLBRsk5EN5cdirAL5BlDaltbjthJAq4YFIH+QEGCYpvz/cdkZz/FZR
zlYghkD1yxhB0AoXTlzvEcGWGKgYTHutvuvbpmI2R8x0XVOcYFt3GHdoI3m9T/PFwtvO9QC1sorK
9xXlt6xkeq8JO2Qxie63V2Pb7tEaDAGcrgRrzGVOrfCLA+W+oV79qwavsW8AcxK6T6Dwpbyfp9B6
aoRp2D1TLje/fQMYCwGdBDW6U2eAkp8E9XMRm67ooauzpdb/Ru3bfy7pPUmSOw/6tYMxuRSZRB30
qsjLXN2IyXbeAluvQupXq6gf80zz9Rt+kNl0qmoXkSk4OSYoAPn8FPEPQtxLIWPAoZurEKUTfuSK
5C9D/T9oaM74TNWL1Rkv53XoXonZnvRjVjoNwZtSVfcoUZ6/heV5IXse5t/e6vw0F/p5HkgdlRrf
6vzE+p/w9rwmOZl5HMdupRrpTfGAwqghd7lwhgG/kAiidLraktdOgTPvhlBCL6L2miFS7FAGygVf
DRger+kosFyKI8Lfp2/aNibLDUs4aU8/8XavKEgE+wC3m764ysFECoFoGSPCkXHbmq+wW2a2HEZ2
4e5rGfGPsCT2MPBazjeDVd/ztoHqYJL+DjQGIPrFuvh+wHMiI5XcsD3HDBtkObx05D3BUG5qH/PF
mCYNJ2dJJwOwvSZWBKRUFC8+/mNRFafIvGvFenfzYYFTKvLV+hAasCDZd/vINb0yaQXgOZQV3XXQ
90yao8oNPSC5h//1bZ/3H4l68XlqaapdHBy6iSC4iPkmZVucHjT1Ocgwp9M7Mi3PQG5F4UcqHGF7
eAGtZX+lvthukgFZ5PUuc5qEbEk015pf2dcWhcktOfIPGpciJR2gk3gHEG4bdf0WZiu09caSqKaY
xyqp9luk3NnwKVBuAkExV+TFMfMj08CJBXlY1Hk5rUm1Xl+mnrVQ8uHBRRaxVMvQ8cLnweMOx0Cs
u0k08j58LY7XIzMUAjxlRVvG8POU2DWEhFutB9CU0Z3VvuLukTmsCggUvbnMY1PElUNTmjhq6oXi
eA8ZrluJd8Wm+uejSI36EyfJ1RRO4kG07II5n/tkUo85w+i5RPJtsjJG38mO/X1fAf3IgwSw4+ys
LDX9xcHB41X3730m4VypTIIX8JIToJab5q+bEPaUvPbeK5RKfMxk53HNE+iCl4kr5mqo5I8nr/gP
rggv2mwMgxQXPIAr/eCkqLuIL8CnB+eTuWSaZgLR0CsIdmI3YhNvU7VDSsTuE3pfo9pETS45FP5u
niAZG78xbpYdJhnH4sXyOeavPZE53xNGHLXC7XfUZ3A9fsgT4k/yIBfRmXc332EUo5lMrutnDTOR
AycJ9r7i87qr9VVcQRYGqMifm/YRocxUWdmtjy57ityQ+F6Pddjq4jGhuWQf6iNNxhGjJVkosvy9
rKrQtYMZdL7grUL4eWPkZKUIw+1uomT0fNkB28NCp87D9WPOW7mOTvquiSiCZ+8SSFY2ofnlSqL1
7+Ou1+0xg7jFUFEdQJfryJPct1Xz4Pgi/j+8gEIX/KbdcMDbc0UkyO9gWe6MLYBjkmi8qfo+DGrP
ZmYc0duwRbjdlAM2PznRnhXBNm0vB/UK18V4Ide32z+0VvekQXGxwC9SWljgB2+A7cZuDssUuezn
y0oxOsJF39ROSyqa0WXSlXyt/Grs1NcwgJ3X/wMtbw27XNtlxHtMN/pXx1mYQiaourEYN+WbUHzU
sLFsd+mcmB0ooZb11cDYgsaIaUvWC8rgVz55J4IUALOzeoe0siVKPpyUMXS5uRycLKQDwb30r9f0
D5p6+jcxYfM1v0wJJ8QYHkIZDbp3QiO5oRoykTj4SqX/y3PSxVhVpfpwp5BFmxRza2GGkMP2Q/Xp
YcTSAij0ALpEF3MG5AdPMj9bYt3BBAtO+3gqj0rFlYbm3CF5WGJXmeyRVOGYMoQex3bTQv+HYyPJ
nkw6P4ZPg7rSJUtq1k0/Ex1BBg1fgUmkTVVMqQftcVXP71t4XIB+sS3N3j0xtO/0Mzl97MtHHDyf
il5648ErI0RPdFDv0vZPStCXGY0x7gxGnSW9zUPgJgbjXI4R/OliO9ZQel3YzRyCQiQbJ+rDF5I4
Qwr8XONEJeijJHmG4nAEZO7Ux8ABWFi5mE0BxI83xuBet1Y0l43tUdGAQ71F39WDZ00QABzFGuXP
YHKWd7AmNW1GZw734wIrGVm+Tm6GwJYCXVjqVA1yWcKd/NTZv/0OWs/MDGhQ5rj3a/DEU2hBtGoe
NjRMyvtitpZQgQm5KqlWfyerl8MoND8nQqB5QC2zieT4HXLp7JfQPB6n17cxveDpzoVWEayE7Szs
1OQJvFVhOYDqiHeO7TZY5ZYq+vpH4SteFC8a24gbs/ObxwVB+df/qLke1knXnbxnTpHrehWSy5lL
37vuFuaVlqDzuGdJ3hoJb8JM/5iJxrgXhAjr9sk3PlC+mbx9WwOj3Szqn/5yfBIaXT7Cb6Qd9Q14
wjhqd+Udyr28IcuujE39ukdLZaLVB7aYlLqlHuRUhcXy8Ai9qnlLVy3J83GbqQFIxo0YCph1JgLv
nYMkJ8mrJE3SK2b1ky9Ce6SPoosq5ANpmEVGGcRPIAt09ztnzmmckW0X6DyMuFcqcwXXBZxNXWoC
r/FS0w8YUzHdZS3bpbggP5A/BsYfIZ17AQTV+b5f86xdw/eOZ59JrOgg9DgKyy4xxi3cKRMZOclI
8bnckgJJ4yCFebzdxLoVu7FxYH9Rjx9B+ggl5Xya/CC10TrhfEHuwtoKmmW6iWPfHH2qKW+x59ga
YRnbI+Cikjw/hNbo5VBBIi1joNGhfqfKp+OJPu/ooa/qAABPYZ09Ppc8UzkBVlahcJH/AwWeVT+A
jCsQSwfsBY2FKxYGEfkrfauafOZvTZ066krol2G30RazT5iE/KFWc4TnJPC8SRwuuVfJfqa0EIEb
kzsZtMTo7KBHWFxHOzY57OHDX7QksRHYQobwtFLzBDnpMrx54+Ny/AYnmd6KdApGrD24W2QGndME
8JP9Vxz1seqqMhgynJjTPEIjb31/E/8DeTYU3IF4STtJuRP/H+qMYDzPHU0NDh16PLX91tAVb7bP
umNAKC4C9tAVfxCAXNpW8LFcSZdfbJMNdbBGRE8M+/DPj+/1vCM7xLjHNzitrmx20uYmTVtcRLh9
nmxPGysi54TWuHZdgSgPMyEAklXRbS39d9REdCMBsqV91aqdB+S09WnmIwuQ9m91Rcrlrb3XJ4Zf
wmDhS1q1WxH5uGqgpWkXvybdTEFmWaehAkmKlHqDaAypCVyncrdXs2igzsjP5/OuxIbGXagRfpiG
liUZ1ldMePNwOxX2ZQ+inKaBoph9e1L7pHbRee7qbIWerqYpfKx5VtUgbdSdNx8YZWe+9J/koRQG
6bKOrIhuvYfEQ6N4MeOYSOYiO6osSVGUt3w2jRvhthW7m6lbikOHD4zrgMmfwM6VfBGo5m0bdX9b
sZOA7DLgxAEn8nS1BVmRkyf6fhrgddkYZ8SDzHq+O1cJtCRweiFdkWpCMa0SE18ZrQk6ovt9rD9+
uj5sHcssHKlKJ8F+k52Bpqrl7GJwSmcMGIJvR2CnRR/6LUiPVDcrMlfQvNvMq6MaIgseOUCoa7Lq
xiue41lN1KAkWKXEpYw3OJ2vomg/CuUcIUtWa1EOs50VaKMv4IMjR8avaOnYtgfxjbpn/zF6rpnC
cW9aFCau/7lZ2/BK+x9OsGhyZ6L0zKVJYVAStK6idZaThndllDyTJB2oNzH2O1zWf01aK94drF1z
GGLAlPx6TrwzE/ox446SLgyMStVaLZEcRU9kwYRX3VHhBWkRy8UYRtRfsBve6lj2hYVQTYZlxYa6
jWbvWv9Xn30tH+kGV4iHWiwGm4ARZjtkur3g5Snr+RpE/+j3gI1v+8dq9jzgVh3/xEG7DTg205Gu
rCnrrDSfyW6OAN9q5yFvfHZPAZjeYW+ZsqoZsCqcojqU+Ccn/IjCBJT1sz5SVE2eNhianmUO/25Y
k5QAKskwP/wFt3LzLz+Pz0Sl04UMGwFACjR5ECOgzHUSjF7k9wW1U/wb++kiwMPYIQ2XfqmHKl2A
e9c4boJWNVeNiJPuoI2afQv9RYxiqSzUZKR3LTgxHoL3oo/oMNAGH5P1+piFwnsB9YlnyEZm/TKP
+U2BTJ85uyrY4V6zOPAKG0lKh7/dz4pyeg4B3KdsHliVV0Rlz8zkvEKcYjYN0eYJwjgZRjtq09ty
OrlVXPsYCw89q/QluxOzRg6dFuArE53YideAqd4ZU4nHZkChXWQmTHYLW2D24rUuM7Ope8cyO3nx
nZ1wMTKkjsJt4maEiyR/WTOgQHbhznELN0nXqnsmwFEtjZaDN7yBJUErKESv7DEn7maLThP2lgGH
DnSLzEUx8SrZV+9hseSxFhIyys4ULYEAlI05f+9Mu3Nd8J49yqebiH9JoCz//sUu/qvJrUJOhdF/
TMUp9c18OhX3uBZZJBLMz36u/WQfsoP2h08b/9oabkEqaHG6rsl4o2A9g26fRjMFBmK9VUhi/Lhe
ll2/ECycyM2e+uq8L2LDyvAP2ZCFF5sxSvn3JYu9sgjbvVqqlrAQiFORN+5drjx4XQa1CvvU2rul
rnHhwpta8FVnWMIJmn8vESn8vISusC9cX5fWuvFrJ8ge9yK9zfsk9O8kyiEAzx8/w9YD3adbmU3h
dyw6+4YXo1jfqQiQ7wOUgo+KVPx2NYyoiWXPUJd/k3ck3zyeMdtQp7/AZBUk4jDxG/paV6NrNOew
NyMm9BQDH02uHqNJbzub/X9eC3t6zUwvtNC81q7hEcx8317puS1CwT1G5MyC5QOjsrZGYMtuJf1Z
LB5P3Hvx8ApLVUaVAmEvxIgLW6SLPGnBtD7535wfDotxW527ZPhkdkF2EDDAkPjF1+ed5RukfTmb
tTbN+NerVEgv7iqIQvUwaejJiOQqCXljt5l5CyAhYy7IiDQL236adts55s8KeZYtpkwx8ngPxOk7
KXpMb75k9vG1X0R9R2qw9da/s6XReqMiQbpfiVrWISV6e3ptRCgjjveIFQFu222/G7WoDlvNk0II
PwtO/stO72Ln9xuoujsLllWxNekUpGv2ydXXG7rgjmD+FKdDCYDsIiczYnGKHvpjwKjdlYrInn0i
ZCvTy0wkm/qdIyum01XyAr0Baw1ePJMsmB7g/YyvhKRl9xrWyUPbHGGIsRXA5/wVPLdcusgwpONS
wboA7+FG7RpGnSiQTHKwnVv6QKy+P6x/EgKOgLMxhut9ePW5Copvq31ZoqR/mEE4OcKP7FYS7x6j
bhzMCG+ydDADurwTet57Q02XvdJxVWy3qMNdd9mNl0C7C+YIozoWDYfPWJA4+QAbtcCpxmq2q4FG
IeUegszuOf5OG54Uk8/T63EttcZUg/WcZ7QChExoYvejY06aRZ3WKEjy5PB+atsGq/trdz5MZnWc
UD973ptRXRCjK5/JmTfYPRpTTXMJZXl8JQz0+CDItHMPmf7wo8zCZgUYK4+WoIJk2G0A3nvlJmEE
JM2NkVfWesNbkOj5tXfvx4xzlx2UAJK3Aze61Bx1nfzDHwdoDJ6C9A8885yjzi1qobsIQpaCimlF
kjbDzIVgZPS96lcJNi4T6pyx8pljlVyartMJ/zeD7XAHRYm8vweReVb4N1s/7euW/O4v3JmyTwCf
K2sAEOwbkmaKz7ovZXzIwsEr5ZUdvjj0jlVNfW21rOAfGLOjeg1kcWm8bSdE0rg4fvUIkwB4OoXj
zakmtygQS2AJncLK53lqC1X4rLZUIoJ5lyrOdkOzqHCCwicnZmYVtypTt7WFXzpLlDhChQguk79s
kKKi7Zj2QBNt33fBIoCuYCA54ReJvG9u1HIcuS6/lTOfvVlTU6Tyl5dTOz35cT2oqRbV4qS9JZKL
naRHnaRT49n6287AVaIlOo0QAJRcW/WiUZrzaQVnCQHgg+TZ9MA8qGZZf5nqeIj3rt1B0dQrO3ww
15+2CsbY0ztudDaUKf8MnQtTQaKfJAbZGxZ3SnkRk9ip24ZUz/a2RYA1c2jvVN53VMKWarBBx7bX
ulSKlCN41UHNyKWZxdmsoX8o+eagm+RG2ZoEtW8S5wQgKoIYJRHclnKJTh8S0DrskLGcxnVjIqF5
7wdcwhbZ4yHEM7yhvkeh9HAOWsulzUOTbEC0hEfJkndS1HIKazdP+U93Gee5ZSM8iRurRqP8FLKs
Qzx0+yTPAIIF9XPo8Rnrftm0fLC5GEJhJC9/qwU3pHsby6wTbawk6itMAPZhbFKbsvSJbSebbQ6N
Fbewsi2pSu/J7DEVrWYMc4LsHQsDUQAn6rrZoSRj6v+fEc6uGGO/rJ0C5q5YXT85I5S4XpiSeKQp
BkmXp0L+syYezKPTLDl9nrifdVI7OWMVXZwsgbneee0kvSti+uveSBWTfFwC9a3ZrEm2VoURRr6t
o2RrX9DLM/2dq6AKRvmjD1qmBqgcERtQYCHbCH7s0Pa+boyCDo7BzN3WaOcMgkIHI7hunjRsezmo
N8x2APWA37CItXbSS4ao7ryEbc1TCdwZhsF+/iHzkBn+8fSSI4qZce5D1Ij1SQGFGOdbL7RLgd7y
UOT8+IOCRSNDbWAB4kHvJIn6Vcwvi2W8WwP1qQmLmLqTP9Z16g/rXP2dPS9cSN6Kidz8Twz7zriS
V4cE1WNmCQU5Y3QpK13aIjEuU7VgjmHG99OW9rrvIGSILeZHO7HcPdmsK+2kHLXx06vXKvP3CH5X
1h8o75eMKUvFNtdYkrMxf0xnKdhJ4daHqevewj7GFN3dbI4eXUvB1RZIZE+yL1XcE3uUdaHqA01X
Oxk0NWMd7jPxKRtQZi4QH8noavDwqNS1CF5HdwESwb2IyY5g9xSGcdvMMHdnov605OtPJBQkkRxU
pIc/2MNQ2JiYPweyQz6quZpf7Lc7y3yWHPSdy+L2f0ow2Bf/AKrgf23L2vsAEB+uN6/KrDBBP4BY
zAoz40MiY6I41HjDCLOqAdxBRisUWFMdf0bD/97q/YrJ0/fXBujWPJiqqKmIpnFP7bwlvNqZMC7H
+w/Zl4jO5NQxllQLqS2iyKjaVNGO8Bg0F7xQvuiryEgHOWfif5HaeeVC0PmvScCM3BphiYqDpfwm
WO03F/24qg6/+4qjj/j5B+U2bC6DRXS5LbHfnP1t2IFlDjb5unYQbAeXsCOEEl2wCeTxt9/ZXQjb
zRoqg8JJ4EarnEh+L3c5yqznjfEn+9IM3xqB6Vn9PoBtyVcBhEfLTVS5QVM5vx0b5sSUvmtfqYAI
fmZlmJd2uAlK2dMZidySj40z1tbdn7ZukzX7y2Jg0VH6rbg42e7XQh523TIkCtpqORLEtqScQKOl
y0cA676R9J0wAjEVKdyi8I87qYtfU5w7oqP9cpIyqMFqGAjNFNrmj7R9BuwRWOhRyGsMYu8WxNSJ
elpI7j9/J8EaY3ERzUIEDv8Yt+TojsdDEow1Z/DqTB5iY0ox8W/23Nz6SUyb8vFLaTqSLpK+K2mq
ePhYh2/HU8nYirTJtVOnk5XuM/cffjXK2yfq6HsIOIAPmuTK0NcdJRmd3FYi9UaASHNtfnNS1USU
yRQGrAWV0nfgSqg4Zdge19F+vyoIdcCSYQhpG9O7/v92Mz+pVgHznmA19tFlgiZ+ibO/DYCgjSbe
Tp6HfxuZoq4s3ttGWg6HcnYKyLbZKVGIwNysjPYNsFFXlHl9M90i9NNSJ2+bathsjC/UsoVxMoIs
CB+C/s/FhU+bU/fX2ORzOGTtAyhs6sNLQOAQXht3d2FsD3E7/zzeGkJgUJUk0v93wy7SiIrp5I6K
fQHj++GFHHCmw7mEaDIi6nCUnRiHVoC1z93b9lZYEOXO3niQjqPFDyl7cUuP4EN7ceCbNIX5lDj3
dlYkCuwQgk8pv7sduIuFCtmN4ugYGysoUvTI2yA90zjJzzHK+RE5Bb4+APONU21MgZi5kD3ueXSE
dpbwHFm3OI04kyzKVijTHrD4U4NHmotZpmt/Nv3eAuDSmfpuPnrZ5AiwyJve7iaxCy6ZRPQ3jDm7
Nbtop1llUDSHSCmQTufSDP0P28b3dhMSedG3yWmRzSbpOTAR25SLQ5zAgLQ3T/aC2RTvM2uDnSut
GJRsQdUdi7gsh66sAvb2hxdXux2gTDq28QiLd5F7UTswQBnpoY4geoaIr6oPcTc8pn+JDtyaSIcq
s9khvqKW/SssHWu7vtS4GKtrL14Ud6VFYZt8zD+WxR4zzKSnS+KgakBp+u75kGy0ahER/PD4udRM
wzLZPbUcDoBcPkyoykBTfTkyUySEUpFWvwwBCtSNvJO6nTYjUKmEBpjQncKAWrkarGP6N3Fhezmf
Afx4weL254cI/y5TiuM0Wr1bMCNgNc4PDIr+vWJpYEL0Wlolo9mc+UY7x+x9gYbYpUIr6Qv9el3w
cEpapWV8Hb1oRhGXi1w0i79xAzMmUZUrT2i59TVrzmBhuAYSs98PmdMMbu+nq8A0ZOg1m71a0lCP
cN7NkP5DLNo6ND6dpoR8x1Tf5n6Grnbhp2Dty5k/tPqHOeBELF6VTQbZe4Dp8jDNBLTukMqK3ITy
qHkA90aTa8HMWjOyLMnhJ1ZDOsdUIBW6bjVjcMzcVRAcWcSjTic9opA5m6FfOotDR48j8+YL7jau
pICow8DU2lVN+hYKTJlDOV70o1OVlg/v/G6VfuD3f+8c1frpHE+utvkpG+mlTxnL9wC7JrghdP7M
QMGWjwvfozfZpuYCGyurJECmUN+jbjAeuvaQCu/jFCXG8FMp005fm4eyaYtfD7zBB/zYtZZa2fQX
6RPqL5tW4ZqYhF9Rz7gEtg9rakdfOh2mCB80GMUr9rKBrD4yQLkAqa29astCvQRXKBVRDhJlVzuk
cKbYkPZwjg3HpCc37XqT8mx2Dyj8+9/yd9CafHfOwWFYian4WF2eQiT+nhObwpGY9MK0xsq7XbL6
EOQHtrOpCJqlZrEUs3hi7GSb+eLvkAtcNA2ZaCHTqCbJ6naODRZpok2aLKtHKlw+U8t41PCWk4R9
nytjHlEwVMH8Odb2cB8etPa7sgmDNstUpMwVUNOAY8Oa9U4WSuCacy2MGcM2BHNo65ve3AkO8A+A
OnT6xHXVJLZse86Hp22ondmk9HSWZ7wGzN+Suk2722p+cqaVLWVINvBmDxYMuZv1id3b0Qp5/qo+
KNsJDvHzSBu5VpRktHFIgOfXfnHF9v0tonTBSRUubcOOj9gIWWlMLO4DQZRTPZPh+ic5kPG2m4SJ
9B8rke6VbbwTcgxLbezURw6LcatTlQ0/6w9fBgoQCuR6lN86BPtXce9Ol1xKbpmKyMQaLw3t6/4x
WocrAtXvIgRz0YfGtqBJQtLMGuwipLhLKUpneP7y+0NiBjLrfaap5g/hCK8iqF8kqOlDeGjIi5yl
K52P3ckvLlzF6h1yqUilu9/vEs5jU6ncKqUGj4A7h3gkpYkoIJhJtb1SoPEn/c8m2tOQJ54zQoLG
lV32awXLGBbRZ4eTtxeO8G1rVVTaYEUeOiyxIShzfC/LXGY+NFsVxBxTc2Kl/Gt+pvx4CFK4gO2s
pqCYWqtxoLcT/vmMkd9hUo4L/RG7dqd4mWTnoMkDkn86aWv2XbfpvmRQ/JHwPJOg2GNqHQ1Ly9OE
l4Ej36PQNlongGxPdRoeHZxgCKibbaH0c6+vMqhtyyggskwuCzmX0bYJflou3+mJLgjyhj4NuIRp
QM1V82hIV/2UoCtoqEYo8kEbDxx/HhddJPv+Jva2/4oIe31HGhHqUfXlFybNAOQEaT0irSeyQBgQ
TNjSUlT9Tyd3ymRb+/oeEp6dc3wcvBq4/Qdb8i0tOMndlk75MI7fVm/awwzJcDLQAugfDCdJQYF8
wx8Nb8Ct7/DRzf2CRgYu50xpXay6JuPevxtMo0CuhRywfI/+eW1A6TJ0fiXzgzHSnU5zepfkGsiy
uDnbseswzYzRJeBIUmyQJvOgCykdYxxS3GfMEitMonw5jRYkVMpmNPI9znPrczgBupyp64LYwOVv
RJd4ilC2UoDyPgzAPEsLvQqDWJekpa8bgW8wLY89jKxT2/hsvMrcsck9LIjD5ftGkVzHoFzTvkiK
93HcKoKT2nYl/6QHP7w85AOvvxo+dzKbGjS724YesU9biJi9xZYTcnThsM6koX9CyIO3Du5IkeKB
XvzxgIFLoSdcpy0JNn0azHSvW4r5UaF/MapuCyzOcvRsKzBS4UPLVvtqK2vPvhltloSbEeQxt97u
1nOW7TBT3TmOrbwafh6IKGWlrjhR7rklfYi0+EBYuBD8FZklwILS314T2JAHaTELbMHwOVRLvp4D
+mNNOi/Wh07hTco3J0HlNSSnomjjplGG3/pRX2E1Lnh4J/2unvu7qfBvl1hl9WkUka9VnyyT7rlt
Uf01AbogFlh7iASXdU32KxqRaagSdDJHYsTtH4Qhv0EKi4NsqerpxUYpKi4F9IWFcz6Ns2KNZ/ki
vke60l3UE+eQqrjp7JbvkpJC6/0WflNY2HWstUqAfPwt4g+tD3/+Uh37dWinNlVm8ZvuScTRQJGh
+gQVjAPp0X6Bb4guRe7e2f9XH2L+IOLWUbbfDHVIxpUKhnZFI4JBZw8pHc6nDHsUvAqNfbuGb5+x
UuDumSC2iUVR/pWf52b3xyD3ZqA8UpQs1/r68tLB/OwSzQ7Uf40WnnFHJ9UpiB7LbO14RN9OqHaf
XgyCdh8YTJnf7ux5Ae9MUouHH5eYh09PHTO/M36VGcF6RFk+YLNmY+jJHgei/FHzN8aDdJGEF85G
/Tsy1Ijtk4nNqEC4JiC+O6/5WZ1evgioz9MH8rZ4ghfdidOj+1B+f2qErwv6OVvHU197Aubvn311
zNtwcieVrv8SK/2hYmXDBLCG/4Rjm3IWw0r8xEvNeoihr8aPksBTb5LTlip1MzK7Pc5U/tvWEh9A
FoOk1xA+FEUYK3oTxtQjaw2icwm6zzP4qqJkKWTc49KBDgyLF9dErl6zP+Yd3bEfwINc6peDLVHg
FAAWAsk1dkgyU9c4oTF9R8BwoAHTVwezioOWFNwTW0W/ICU2I6DCyR+2EQp8GWfc6V44cvwNNSBq
62QMJCf+qPX2vWMPaCtj6EYGMkS8ZPs0YBAxS6xOipmPAx5K3YiswKKfMMYL86R10vo05hAKzP+1
UI2RhwlDSWLxv0+X0s7UMQwRBA3xW9xGEw0WXHQNyqZFX6389S4qq6JWYu5cvK2Jk5TtVlHg1ncG
/1xnzWqibcf0UUb7QI1ygV3hAOuLSMvFI/o9dkdAtKjrnK3l+YFSzhsfnoze0VpQl2ucq2UoyZ9z
3kRvFNHX3ucpsrg+QpoV9jle0JCZ8hBloH/LIYFa6U2X/6Ckwn7eSuTg7iWyjX6QQ7DNgInsrXYl
27owTK9EkeXV7Eozzv4g8/dwUQCUi6n7ourpMinuM5u78JYH6Bax3DM9EH4YhuPAkajkI9nwp66Y
JU3Q8yZKHxETcatPUnONYfg854fow9aO5M2Wo/WkP/UUAstingiNcdOU9MydAnXoy6fZ7Q0ZsyD7
fvjFCIoMJDAOwso8U0HSVSJJkUJLaS/9kNfI2sT09KQImODId2CMLyE/MiU+YoPgNxI55AuIE0Bz
PFHQvEFmZ4JMSAPNDbcgNV08yCpYes1x8vDA4gjNJjB/hezF88KFQbym9lkH3uEq5WBC4z4yOoic
QJF4nJV+cUuF6KB37uha9vdVxkNPQPsxOXOWnTHtb08oASNghcjPc3X4Dd1AAuW4ItBDIsoBS+pL
f0FZ1UjBN/NYyMTfvovEnspfKCDMfhG1YjPhI/VB6nu0fN9fzgzpnqA8G9AyXMsLFdaBT0ixePd3
lGK/Zq6B0l9XDSceLC373qBs9G9iKAy0Ui6o57fuEddXBEwJ52Qyzk00jPP/1dpYpb6Dn7/HzXfD
NBLVb5T+b5lsiHwjXF3I3scZB/tvr9vOkRAcovUfgQJiuii/i0L1YWKzCGTGGV7L1pph0+suxcTY
5Eh4ejWPh5XPvAilbkxZ+vH8Gd7WumO9DiM+abWvyIaAFq/V6QgwjqDgdJeatEUtL0+OusIVBZe3
rtKcEoYlDc/LqZImYbfyPfoEthrYv+y2warWtVHOmiJ7yoZtVygPupPs4aJ+MX4hUkMbsF08cMtM
UY7jRBChE4pYBFR6KKUmDopRS+cpAH0ywUAHJKRxzx83bFSJg0J6v53jz8S57FRubhmSYVe2lU1W
k79JzZ5sL5XFxhsEyuGhul5/xijxOGLomEa2yZm7MrGsBvH5A17VYZF2uUtRlbsACoyVgIvVaRie
9cD/FrbrrzAX9rAE+zbBtraPw8JfmAWP0DxNXcFUH6cqj95TyejZWp7QHvPJODbSo+6brwuziC7n
4CSEwbzl9qynRujIoILgCqVP7MmHsjvT28Gsgd2+6PHhnW1G07xiuCHQIVgG/Y3PrV9qNRPRK0tv
fhLZuQq9G7fhFqyrp7Ea1D5NmoOwGeeLJFdiPmm0e9Fz0Tf4RIfHjcghIoOgAuWouEI4ck0xf52D
waj3Y7p2dyiQtYXig5mYvjWbBbsLGftcNHtCyNX6EeXfJzoK8Zlu6yE5imNxFOF30HWhiiHDL+RS
duwvg+xn+0BHJToC2e05La6Dw62vnUqUTOoD1cfEkZdd1KPNMTnz4ebTUDYn8hxGn8ivXTqpTTvo
UNWYpJ6lvRZdkKQKPdrRoKrvgauxOllR+7KcrlB8ddUzJgfTFx1u5gEMoDe+J+EDxedQ+PsiOMEQ
ojSIvtiXXeZAJNvrJ6JDfFoeBBHXPYi6elYs02dsvGpTfqpjaRlatnkkXx+JrC4IotCBpjJKiDmX
0OrrLk/DOm9y0uYevjoTAEG4JchPGBRu7WiTtKXCHKkBOKSiCyRXvccwTbbXQyuUoKNuAU16Zqfo
1usEPQerFkBv1a55N8i+pnIB4PcrSAK2uMEtjOGkgXNl59M756m/vWOvicIogUai6UvcKuSI3d4J
Er8QMmiq9b3kjaypXCDY6BsTpKt0B7RGilu80L0FnPgJMN+DsSuBgPmyA0WoXk4bjuamVymyaURq
CkL1j7BNZKcYJnHut19ox3/Zy5pwEk4K4sZanO+Fi/VuB8VpA6hPnTsFb3RnAQ20WzbFc2IBuOll
8K7uWkeVGJbXdX0Bz9UczxhJ0oD5JP4bqP5K3dlxc9M0vIOXXMohclkjsGdLgeeotAHpLuAhA6GU
7mLxYN7mUvgIlsjGeeXlGw5NQd/jcSiLNUg0kM8QOl4bbc0GscObUVLo2OyvF/qTeHysPtcDS1SJ
gU6NH/oFMv+vt8IoPJCjuJhKaO4qGq+QNH1vK/8QiVrcPjFQGhm8LQ9dnlx/vMEeTY4fWIZZdWPL
0KtvK6VxQQgusbZUqtVjKA9WwS+XMJUveIYgpZj9PjXkaXHwy/MoibxKWww8hek1q6LKH9SkhrI6
lsWThVxLvV5hTj8c7qAR+iL4xr/EUwbMRFDcEO1yjAa96Y+peWjPxbgxlFUFrfU0TkS7aFDKm0Oh
b0bFugT11Jm6qPRO9F3qbLN8mRUDpQKfAdi01wEZzawIpQoLDe2hQxnxTBJm96Pi6VS4JGcTF+f5
EjF1iZOHR1/h67KlSVV8R8i13WjKjydJ6zfF0io449Hs+7opjFe19sMFcsHclp/Yn8uIM95lCJFE
ReCmfXni76trPJkRq20UFzLNsErIqdXZiaDZigpoxZBLdcRSdOc1uzE+EyL7FMecXL2YayMSHRxG
SQj/AuhVUY4LHjWGr7x0BKiiUTLHJvFQ24iwR1B4lMhxBEE0yz51c2PhmRwndTWuUy9ip/GTQvuY
GRTL06miCMI4B8+h5Q1TEWHv3ZUmpCT46GjmN+177izwnByEkQkfwGoIzStNEusoMSclXmbtZ0A8
36Jp9zZSPGxMUtyvBIxsz0YgwU882+bCN6E0UXubmTo3PHQRNWczJWE//awmnxAHTGumJZ0YOgiT
uuilYwV3JqnfrdvQ2woVLOST7kzhUoxOXlULnKeGy19apYlOMax/0ywRtm/M4nFPOJbyNyBqhqY+
LdKIUt+wD5/KqgQXCsI95+EQN1+XnCVknddONvzoGdL3u3iTzMV34G5f2YfFXayQ5iVhd8HFTDIg
Z/nP7lCJ4p13zTVUsaKWSgEM8i5cYtzdsqVmdNmja5+j2CutFTVZaI2jmnYxXRdAJMfhLMqrp3T3
44DT1yW6xXW/z5bLw6sgOaQpuup6117+Foh8JPo/LApWYaStMRkqsf9RgVfXsRoOrbmVJiewLrnM
mm3HdK0UrLKuJ/foH2SUiF3KMMO4KlItTkLK4Vqg1HWjqY8hhznT5dCtNSTwYPCUc2XUhBkvK4I5
Qxbr/6fiyu1vDjVPKP5Pb6tHbhg26CNRXTemwx3r7vUROQChAps0hPXnUvcvYl9r6tXtDTSjnbWc
A87eX/0WaxS32QcXF5tsP2b44lZ7uA8IRzDeO3yw8M79+435YYykqfM4y/+GQjEW3ZSNh5m5BRqJ
nHXIHjmJA9Nr/oap2bv8MdpZ8uF9rrdq7FjpGmCssmDMTE38QPh+NfuKx8XeMDMja6lcF6MZS8wX
9ol/pBWeumTNjMMkTIOvGx+OC3IHvmn2f4Ga+837OWRuewj3WvXklV7GBEw7tOUmQjunPdX8kG7Q
bDKSm2mMnRs5YgqUH+7WPFlr3lt2zFF3TPAAC3/r7WDiixTG3Oz1mB678dCF3TGuPmffrvpEQgCx
JNKXU8RthYl5ydQmDsy9DNmDTFPzbOTbGXsY4LefJ1KHDvnWmi79o+khb1jRXszDn5jv3mLvvguX
CLP6vS7Ngb6M64p9ZjYEWVuuXbYFjM4aUfQpl0bsonu9JtUcT9lKp8W4TyYn+2bS4hW1mqCj3/db
s+xQQKFSwLUSSouEE1N8Ya3Np+3ptbn3ylLswLvIbXjb0SHa258gJpqWb9sqzZrUiGM/gcgepcC1
5Idz1kn88VZoxH8b3Y0GeaGpkjHww+QcbW3QUrFtjuKS/gMSFejcUiqAe0VZpczK8U62B+JMRTPG
sVyzt86l2s+53urOwy6AQxrTvGzumDM7EmdktJh9bZyyiJ6wqmoVh2dvsXYtEKqeILlxuCgKgqZu
R7zspsMl7a1MHsMjG9lKJn7EV+53Q4crTc7omKjzafvDCOjCTPfrqxwUtrAb6NLw3+CgzvuUNBGZ
fTZbN4l3ZehE0rLsXppM0Im0Ok0Yz/Kl7UkXG7GxxqCX1bdhZj8pKcXk5Gnejl78Re8SCU3Ur70F
UdJtd+gVcKewKOkV5Yj6fqmAlsM0Tn3ymZRY48BHjUM3iJbOLgZ+TJOg8zAJVbX/S2wHY1yKRkS2
0oJ3irQWah6nDW6N36sw04uaMkZxX8OmCVX0nysip8e65TIxq4tXmVr7r6eGS3yUOHZ2sXD0SXYv
SloEk5K8j0pzS39DtpGfbF6Yo1BeKOkNDj+Y1h4Ayc94d6Iyck5UWT/eW1EMa6o/u2jcJQTcosHl
tgXly30z4qFqJv/ykQ5R1DPpLqBr4KIxHivyDzM47d+n5oE03KTl7xFiYGMQuC6RpOw4VS/EX3Kb
0VnSuAQCRAe5Zx2ieXKzQiM5S1Smev/LWxAbG+zGDY7icL8q+vIwq+dZ/4t5iEih+vtJgrYhuXOV
DnvpGKRg0CoqNqu3kNSKEzn1K5baeIbyC5Flyy1Jud5hKta9tMFqef5jf5WXbJX7BNC54PDkGPTZ
bbyDwMD3Jg6ot+iBkJP6tUXqKcIhm9wcx0UJXn201Du24QkdspNA1By5W6OqIurA6HYvkiz8cD+b
Acfxbuni587zjKpB0qhTHUAOLtGETIh7umc3AZE+RZeYJNpF5ldwrlEoN0YLCiUQcOnyqEnPx8q7
nHldraLnGCugNwsz7Vb61RS8x3O2tdx7Tiy/jJxjvNTIe12QY2uTASyhSmBSd/H2Pd4DZCG5YGiA
vmOm/ugKqYGeRkjmKTH843RRBsoQOlGQz4VMRFS5h+YyKcVckaCRqVaqD4Ct7JoiWjVNF+Be9pEC
u7nZlu20lIpjDA3zFxefyiI0HUMywI0gKIfQXBcSMr3Dzwlc4ztGmvtN722b1qNFMQp45T2k15Nv
VQt1ZF8i/7hbefC/GGZ2/tmg1Yd7276gx7Myaqfgc0d63g5d0u4q6+hyNmjP1IFqaF9w4VIQKTzg
0ZIsecLDMyPSvNASvW0suKQcLUzBMPmHNwlKWBDIf0smjxgeAeYf7hzw2gyb72oaE9bnKUaVfKH6
ATVb96+JtXLqYG/Oxt9bRGW9ECImvhKzstXcoLm+B8ah+3AzQ6RyqRZXMtPhijlsZRKREb2eMRiR
VoJ9RBlciU8lFFVkIUcbK686FGiygMm+Q95B4SlJoyQXaFCWzv0KKH6tQsVydfQfjkpUGOTlLhad
uobfQXJ1nulW7ewFOXq9d7wB7vsEXo0Gbm7RaK71ILN7xBgKSlYdqAisKzjng+KCRZfWvvVvZ0I1
hj1vgtGx1/NwC/RO6Gw+bCspwGJ1oj8peLSniPidPvLNSObfNT4XcYNydPhgFGSXQZMkJ9LvczqU
KU8Hw7BntyvAxy3PW2MLGtxxOfdXj3mZKd/BvuCOz8zGGW4/FDGLRb458TQU8X8YcWxaHsBEkHCC
QFCv+keYWiInFbcRs5ZCGmIErAt1L9OCehW99jJXikZaX4OCOyT+4j3Ud2/BWeXoj8SjwFAkORAU
M76G71dNlKtNH8GR9lt4c/e94MqzJg5OjSEPVQcFFVPP/HbohnXESInFfqfVdLCRTUApKVhJMXTq
NZ7G3Mo2DnMcBKcVqtr9PjY/B6KUxxk9NYksPJ1dq4lAtP+smf4CIkrMCX8m1gbRWnVIoXvXl7wv
5F+EBYXBsfJnUvnRKKN0O5MOnyUn6lTCsfDTJQlK5lypZY4jirEFL0JoOAWh2VmEgKf8nPKk53wV
pX1hbwsp/KkcW4105RLi7gvcaFTtxuN5w2KXucG6K16FpjIKURyUJa5DUaW9KLAmcTneqHcj81gQ
DHqxYQ+8aIfdg2yp7XNniSuM6MSlQSGWanbd4lNt3mOhMQDaOKkxM5HMm6h4C09QEpdEtZaBnEqf
2Dq1oSAvOVmEtMHE1TfbapEC+Fag0P10AT/e+UGBehLZXiNRqGDFI5DgIIo6+8+iD3qAb1JIVtP3
j+rAlxLqBcpprkMiHf7lqp19VqpUgnH8kReKVc0wgemQ9b20TzNbvIZFOzccDPxjDNUyOyijnXsd
o55Se4U8NwfMhzTryg9W55Me4UMOBaW2WjJRS+Q2vEwi07cxUuBRBxXH3zOvCCZKRPaHO8Z+xaAa
4LKEcLLUgLe/lgUXnIxwQTuVjf45z5jTLhEhAP8uzByee//7N/I58oac72VPSOgztoRANRT3eWCM
NVA0UfKPx6WBTpYx2NK7S55OamU0mw1GtMetyMazNsKay/Bq/C7b4jDAWluBUW2BpdwlXW4THJex
OXGuqdIrNjIf4rROPGVpXkhxb7HtoouyT/7c+/5zRlXq1CPR2m0n/hh6Ldq6Taw9D3M9L5faNkDV
h9TNVwduFzC8sFh9vBCCfdxqMKn6lzm3EfXlAFYftpEEj1F0pRiypeDCCT2tdSsI/Ey8CJo/7lTc
fDpDdPsRrlwEph6+wcCxk6DHTQD+0MBELfJB0cSW2cWLyRY3gtJnUc/UZVkr6O3q40ZAEGv72khQ
IbaG+sC5hAUmDxWWRlm+dHErmGLoAfsTaWNYKMywvdo297X3eo/87Jg8XLQqCnl377TdaW5BGhWz
fUi8U1ejckAqpZSeXdIS7Lr3CWssu1PBt5GYlRMUyFUD9tLMwCGpe7UYfp5U16GVKXqq/uhM/Vsb
EYN0yBBy9M0XmwqG+vqRKCynfuho1SmSXgb+jYHKJ3bBe6eiv6+nvKocPE96DfNpYW9tLscG7tVa
3Le+EpQD/QjStGvsme5bOI5o14eJnB5oacELJwU1YBOqWHnI6M0Q/Af5wj0UxuBm9tst5PYY1ZoA
UoT08DK4lafRrs/TIABMEsQcruHbxIrSJF24xPlt4yfIgbS1FXNK8WuGl+RGueFWLM11ZuqRp2OG
QAN4+sG6cGz8iJ90CNrT3rNzRmU0OescnI+1GCtDgrW2V94x7tD58f2J2dDaVqh776sHwCsRBrlA
qhgSjSHTNetCVw90jaOp0TMwbhI5kflj4SNdsLhi+oM0N4sgF5BjU8yx0CrIGO01/tcrLfmkPTYK
QPe+C0NHG+IhzMjhUB/Z7avGW5ceCHv3Z02Ly73WmPAZEbO82i2f537whFU488ZHqrMzI4x2Gg2n
Et7Bos5ChmrkZIpStl9LLgD//aABXcdI0Kss3+8KugFAmR+B97dUFjG34U2nCog10442RL+xw+Uf
FddZS5oFUUOo+Ads1Je0qidglywB4q7gVxIp0RQpX+6Uwlp36s9onYTV6sWLrqpAxmNiw7yx4nwt
VrYKHFHlqfsKZTazdQYsgwbLmuYZjQ5U7mc7s4bIFJ6J6vNlwVHNyPSzXFF6knt2UBqbocbIb23c
UsKmGeF45D0u79H9MCSS7uduT41m5DwEvLSDbuCi0MxhsdM1CKNIhgv6xsNzfP4tSm1Zda884V6r
lmmSP7eB4Ty/PuRpaN0c/F5c55yRkP1GSBdO2u7Px1tfn8GtTck3dMJWWvt4EfgZ9uf6sjnYhqIQ
9sorfayDAt5kgwoziW3bV7cSmxAyhSUwfeXdcz4PmQqCu25pGLB/PCoh4HeWHW+ABz/2/OF7MN+0
v4YxbrS8+gGhvaNJjK2PRhuezBM7boTTPuyOwqTWTAedG05oLvcwkPRdgXXQADfVXVwgU9TA0509
DRoetNuCOxN4XG0q3A/EWjbtPLkzVp1aoYH8dgLAzIsakpNZmqUKUmHnD+NhHgEyesEaoisv6TuI
LpnC+lj77d5BpFZ66NHy9IJ6wsTiRItip8tZ/6if7EGqgLsfjC1qn9sxurEcp3Jlmc5KtKcBTL8H
zLi0PWPYETLHG5aCK1ciZQzFC3BOnozvp2FFVPB5SXy+9NGinAEEdloTd2Eh0lMvVzN3Oel2LIdf
dkRa6KilJ3PI1xuvRKoTQzwQvnKSyhWvYMOraX9p/N3b+tfpQhJZHigjO6Ni/f4f3nkmWFZG2nPg
UBOOLD92qjsHyz5Fwd7kyOsaoc7HPRLTFryMfybi5RV0RTPfT9iU3CPVxXGQY39XtiAQK/nxJsL5
GEmBt72EV8Sf6Tdw8gk7MckQkLm1YKb5tLTg1k9nx5oO+Yhm7wNI24P5d3euepS8/BNn3A1QKvHw
VI7DGKgTolKE9Z6Vw7We47S0p4qhPlOkEqn2M4NEf+5RNnCDjjJ5Vgt6bibdWgBzZ+kOoqZ79P3t
yUoipusT3CVeIdNnAvvNL9OwXHHKtPBGtXx0R7iChQhmySA8dwhIyogl+Htfn2Xj5dgJRfJlMfHw
mzHFg7cJqpPFK5D0zS84e7OVKho7QCW8QhE6YNsXf4Y8yVPhqAVZSRTsz9oL1Tc15FcZ+dRiDxEJ
THiOOxGahjjSlrSPXLWdNenREQmGsb+hzNRs5GenePNDNWqNpr8DHPpUdCeTZp7vCT1hM7zTEGsP
bG6BrzXAJrUdN+tssDs2CfRMllafgAvr8zh928wjsBN7RhU2gAgLA9400szzoQL5q02TAfbk3BpX
AwxHSQaS4Yvt3L7FIARDx8phPW4G8w8l8grUGjPxKVpcbEiQsXCBVtPuo3hVeTAac/uZEGCIFzri
WpaKkyuzbV5ERpsSAlJpf8ZkHOJfd+c5cpvDhMdLIJoIgZrx8ZRB+lw2UqdTmRa+guxm0hyjsh1c
AA8R5zpnoUYVLsjgiQundlz70hPLQr4DqkNi8+r5wOPqtZ/Eebnynh1PyNFB3vzXL2KObIlj8Glv
J9y1GTl5k2aoluRzwYhyDv0Z6yu59S5w8i7CEAdPU+9GnZ2jqFnqJ7cSsRJXTgsBJiNz7K29whGi
mbcbPYWbyYl44UTgKDeo6gDfL3K6xUaa2LoYukhrTh0+YEBjG9x+1RBuh4IyPuIUHcy4uib5nrP0
oyDjB0QT4N4HOdfxDCutFGgPWIdTDuu4O4OKTiEWfJ4WjwLuwu/p4K0JwHATsb98iJhuNsCPjixm
kipd574at8grxgBUAhxkFyOZqucSkwNqOVLwIpCsKegh4C3LzqwS2Q0RQ08bz2u01DW71dHGBeSd
55YlRk3XfTQnbBtBubb9PT5DJDPSG2OZFcLPQL/V8TiUopG733frMrdD3cXjUvVsvzNfhYDKIj75
KtJxu4lK1djR+gonO/e9b+6oiuNQ2ZfHgSLCCcvpdDWrWgxhQ3yfxo54X7RdPGZmhmQyIT2eEUO7
92wD0NHYshDLhz+5QgxTsZ3213KhxMtsSIUW/cPGoE8B7ho44451djFGD6NXtf9gIyEO3NE+mqBM
w9Kh+KRtn7cJRZAJqsB5G/asZYpVdr/5zAoKFLWRpO0NFpD1qjUd4DpupLWI8Ym86RPnPppAQSz4
LlEpzHh+oLUv9Ux5Ho2xK+7VKUE05Ei8YY48NFLbVUCBVWCmWn9ESSbx/JxGzcZBUbuqeAQRXPZX
UeVA2AfQL3gW3RaWSOF8CnI0C2Gx0aYb3xFlipoURNVhC74BFn+YAtaRxGNqOU00in/Y7qKPii79
hlq829Fiir8Rqsvu4Qr1fm7NtlIf5iCv4j9if79n0WoRacqQuZpDizm92erAyhTnZRonfv3aQm4Y
PyAC+VzmTdAD8SwVp0J4RmTzFUYQb/53chOrr4UFvqSmojbrWgMJouWKMYYx4pHkRODpaW3tbu0W
PXpq1zqQcfE7dGjINrwOHKmEhzswwKn7dn7y6+rSrMcOiYngYlEF2DSvNo2s3nynyL4pWudRFzLu
GblgIixcv8q5yu7scASXDGcALaxtEB8Ev/M0eDd8PkJl1cWRApeaxT6S2vnG6aO4kQYQeNzlFz/a
z2KBCtlS28XSnTYgZoshURJRzJeIWKlvgNheby/IKPKq4iaFOm9HnSehuIf7IrcmEgpA/O7xgmdK
A79+M2zSS5k+gl5DUj0YVmW5SgKGDNfX2x0CB5kJPVKsPKGNO1Xrceiv+q/XCZLSubGAKocpT4Fg
13YjepmZJsg+W8S0YYOfQezyVT0dJ2H5lEdX/WjigtUJzEhhMYzidGH6Ke2PLheVmLMNcamdExrC
WS6cS2JfUjAPuvZTAT8Fmi68Fhj2ojerZhpZIQxtv6Gx4lsxfxUIl/n8aAzi9GmmvItYVLuayuAH
15QP0oBzM58LP6ERs4u61ptB/asz089ossSxPzagYeUZoiANqerjX8aPH6vIjSIG+CM9gjHSfHHc
1ipLlO5kZT3/U5rCUIo/KcHtR1tVvQWV0fls8KHQhKuHwSzCuYYU1DtqKGoHQEj6wPztjz6GiJGC
DhD1Qy9Qzza2+Wo/FwQXQVxk32tSrslkMwphHlXtPaH7MbTSiGUTwHQtNZAPM6uw0Ic48nL7X4NO
+3JBhnI4fktgebppbGdo/bEre7xa+HEg0z6+pFCcUKLW2C47jTdV354zzQbN228r0B91zfO50cMf
4p3o9wMdnO5txRgxJJViiOvCfBO8e17ailbcsYxVwUbvTiydCMUCLsfIOYQt4AFbfNWtoGTYGBrV
BJKacwc3eWxes9IxF+vgD9aU9AqfN9rOkHDhehnZG5yeZ15yTyDDZL4bVwxP7QXKfpqgO+Mg4vgD
KOdNY0l4imeUFXtKZ8DpR7Bnh6rkLcPLrLC2f7l+A0ZaIuO475dTZ7ntxcikhdiuzcdrxHpnCoEv
DGcgv35mUbz4+jI0sR1ueyfNCsVoUzJv0zv+Jz8UuCgBbmPgP4g+NUwEa3b8lZhqEBvpaXnyuNti
HBV8EgVqiVHOLoATUmHZbSzmGSe0WmvR1mHxQRcdmoWIVQYb8IMxT+jWBFu0d4ks7mEZc3ebYM5j
2eeQ5A2FNK8sbdlcXHn3yYFjMCwBYF5OA7GUQ3qHKNIAa0ygq/G2wAb/FOmIHNM/nqNh5Kpn6Uyt
ZLCt7M4QW8tef2ve7FCZvNzwi5TeYaQ4K34r7sGDeK/xhPiRyYNSovlh9WAeHFPVgEePE3lAPOSu
PiaPJwlmMP6VkEP3IUDl6osHnzBwKFGQJZRvGQSaAlGm0mYzWAbk1T+ja90T3KMqtsjTYEQd9oyL
LujDGv8Rj6jMiXiJC7CMz6wlulZfEvtvnXRFJSl128O9nxb4m2q8pj+pPfKdf0lePDOu41c86BM/
YLJDmlQxiSP41IUAUcPutJa10Jte336R4z482gk/0wsCU0P/goY/N4APtyQ+s1TwPhlAgDkm7sZ1
ghsPtox0v3z8NqIIbP8Hvv/mOx5IReNZ+H7UEI3m9HunniplSgRO1053RJezlooQXnX77CofyQxl
Gd2W+4lZ2g27femK9VOQtNdhdev2azhYt89HaJ6aFCCWUE6VFcwADmPuSh75HeDcXnIJ7mKcgJI8
j0BZrmzriLg/FxyOO4jTMtGEL/sR4SfL+u0QOaS/o9F2nRY2wsqh7n0MSjgmrONP7m6JWq5psg8p
zdGA7dPWbq0lAzuFOouTeKC3NKy9s3QcusKymJsDsnL0Z08fznK3gPtW4AL7Cb2yPCrow7DuGo5n
8a8t11GdAAG9M1BQd66xi40k0AQ/IN9lvdEdwMSe8vi1QuwB6sVASWRsgCWR2OZ7L6+tKSv9PEAc
wIC9Gqom978svg/iOFpYDPJ1QnWoqpmOHVyjuydOzKCiSTBwoZN9pQCv+JXDSalpYknXRLanrZmZ
UFyL6+H5Gu8qk7rS+dd05dIHj4fKojzeB0exl4wiXM6vJipi9N2ik/Kg3LkSs8NhgpkJ0c81uWrk
52jJmx6mqL4SksY5KLWExkzclOKBD1/JGXBUPFAsBie8HaT81wI4OyB2QXOwgPTtyNm3N7zj/kLD
bNTaGhx02/cWREWzv0ymJjeWyXaF9u9OqMRhxY1fh7lNIWrj+VyoXdtA8lZuFpBTlLUx1/LezHD6
u8uIAedyUkPm/Bchuozm3qQxTnQsMdf+952ECzCjdIS8EBaeSxQzeB8kuikaW7wxCYiF4Vk+7+76
uhitgyP0UhA/+IuhmSox9aj/3yBBeOj+bELanARqwT9cOsLFpjdkfJsjIBCKR5svWivRte5PVXxh
x5LSENxjWaQx7mhMDqkzAFHfTwoAUl9auBnfKR+AI6GiwjvGaHUnK4e8I1zJzvd8CvkGfuaDIKSS
LSjZ+kGmHH7EPx8/MGYAUMBxIic/gaTvdbDz3Oh4Havfh8gWHR1kGXJqAjyRPbJJIeDy1zUQzB+R
5o3HLO9+lHLzgsrUcz8Iy5zFlnls0Lg99U0Z8/dwVY4kQSB9KzjXpEmS7Va/ZBpaxoNDt6KrD6KS
oj8kOLD6DAapHv2w8sL28NQ8GoEtRecZzAIh0SaoZf6Jp40EorUFrAPUqzfdulJ8UzC6ldB/LOSL
pFCx4agqvEDYj6f53cGA5QvljePGuyXdgkIlOgQW0Hp/jo79BuP9Tzw++eJUqMYNmSbAX6HIHAOK
d5RvQ+ujen/4WfFj9CsaSZjYnTxy93lDq14CDwuLYOjF+wYTrZSJ6xkwywnKpJk+r0vIJQP/0VZ/
2vgd3jSFrCrQbhRVgelA8uQlYmPbR5P2/1ISCblTmAbcqGfOwep6xWbGve2rtvpA9qrKJDPGdy71
0nDpHgK3O+QnBxxldIYILErUaAY5FLzHuZf8Ntfv7FUqlcAK6g77VPpAvZBMnrHk6JS2tCpnuSLo
QXGk6obHJpmujJFYjT1JDfgb3qU+nynroejVAhg8/8Vifb7n0WjHT7RmN/OVYBOJfYfINFZVfVoG
LND+Z8rpU0GAyFesX/8W3jsC86LOZu1QcaARui2eeM41MRpuWftitdPj9OPHFiz3S/EreB4mld27
F9noyg9G74woeTmDpDpS/Rw0Yk4r1H6qSGzSToV8ytLdXtGIV4Un/3WIzeWG6xT0ySECXtRLhitb
pdG8gy6EH831nunCG9bzFTyyxAs/5EGr4Q1AYeAOEOJP/WbsWgrWZLT3rF5QGL7pviAdbeb58gHv
1PlKWCAEt6WmLSS1GaNF6GnhjT1IHfcjfHaSvBoArGn16nLTuhGSPoJsl1YskvfU95JMVtF37ttc
ogj7ICYqL+qgWFmUikLdg96hgvClyjhxrtn3V/hXtPIUmFE+eNNSzgvmtvVXHLiRA5iLQSZvUOQK
SArQwN6bcdeOfAdxJDePECLrpPnYsH2KCnwTudxJTvaxoPyLGZYhGvp2wvm1w54fqJf4PU+Pqgfe
WRM+oyXqWdL7Ti77GXNK3xCh/lDWaaphIlN+KBwHCRTXfeLkIPeK9Gq5jarYvIlrBsfJQfoqBzEB
7ZFTwj9+MnjdHBlbx8iwbIJIs3Ct1Qw49FMF+EnBmUvg/BQkLpByaUnuAJSm+KRehyfZofMui1tL
RfdN2mFjwmecz7QkQMZ4eKyn31CnjlgLyO9oVXNWMCkGt1vWvdMLPUvkWBqgUc1VEQzB7AbQXYQq
e56eXCbsw4CDHVBaYfCnfNhDHyf26p+AIJW9xRQ7W7F6cQfB1Wdh+OHPIezY6EX5e6P8uv3RCaXy
p/PSdA/67pqN7ftKBPG2ZXjDOVgsGhK6jK8Tt50YCyR2Az8PTIb8qWyNSOKW5GW0X/dPDpVe5hwa
YaXg0EUc6BL6BQjVS8R/bp1Aqsk3fcSZMxozw1MLV37zMSIrJ+V/f6Y5/XtEfGyZBCotlpui1TIm
B1dMrgL7Ce5PCvBl5siCtHdu7c0pKAgR1Cmr22D8gXJtHx6ufBnG6yudQpt9oYue1MhgzE3FZUZc
OGAz+omahMwtpnx5BdyIQpyVePoR6nItfnWZprsTLuDK5O2/PznFRsPp7CZw2ocEBuL7KkSoHLzs
50K9Q847wnVxdA89ph6AL1a3bJ8CsLJ4GUL9ewyvYusHB/eaSMbIu9Nq1HMpNLh9iUbJOO0bTcS1
6m0MCNY5rrnpUNdJ5t6YFlsDgB2H61fLAZoPp9W77f2b9uEiwLpK/dL+8oSASNJf3/prhdWEsb7T
/XsirFL9LSxQbtgjoWPX+Sln0LCD4RMsnTMK0bgWH9xx7JXu8Ta0U26IRVNbAFSb7NDjsp063NOq
+4KX28ZCcc7SSl5T9rl6uU6mmYudN53xN8QvE3N1bcUEvv3HfCTAcZteuJqnylmb36ieIZNC8McV
qXnRhl00dR6jAY3b+i3hT13CZBuYv3IPlXQ98EG0ZXGmQfsnMADdV5s5qy7d0FjXmCxBgIydHTBE
gCR13/Q63Anp1vATcATagHKJVA7GtUXRYnlvRqJ/EtgVfM2nglBI9hJcVZVjpt3CPsQP0qsHrizo
a6iy8rqVqMjoJtSmw3v3rHm5jCwfkMSrfODeptJ4YT8Els9X8QQ4GdjIxTxYe3zirJB2wDF+UPCe
d40Ei7sC5ydH9dgmMclqzsjEcxiFp5USJqiqe/56U/TWuHAC356qvjfCcHs5dlzjN+78VkOylB9F
YzqKBhJoq46x9g1wtY2F2uue0zdLbqYeiYrJSoiozxo22Q9NB1V12Tz38GyeOjHgQ2FJpSYUYPVQ
MuVmlm5o07cLoezqrS+wQ7T80R2b0v/evo7j3mwTnUx7kmsAw933i1w9DOz92axXXUot9zauo6Bp
flXsjaBpJ0g5J+zQcSqrWUJ6XHU4f9a/xK/PyeoildgYNehooMbrBoooGF3yGDkLITdUGz/bZtho
Ngc/ZJaj5zcR13XPQyJZB98QVT3OULhKNpUaOpq0nfPWobI6rpRV8EgW4VEwVBWjEM9HxyR6/Lar
Z1pOij3RBayxFMpEay+6w7iHDqjULB7wCYtpNlILjoDRVbLbsHiZKirf4MY/CyP5N4E4sb6L0U+z
2H/+sWA3s8xmse5fL1ioVYavo/0B0hipxHgE0Fi5IOX1yKT+K08zJw8cOxgS/OU8jBpwZqdblCy+
jm0qAGFCsSs8hWAlsmuxk/GcmuZGUM8etvQ7ly6gP5V+GddbNdwb2QIsogzKuSewccKbTpfpXa4j
1xrJYmH0QRJLuwAqYh15iO1LEaWUeSRlypRftx6+gDK8JK/ZtOtSb9om9YKpTyuc0CW/58jyUl4h
29D19OHqV59zbJzJvwrQGV/+DC775n9g8aC8AcfuQ8mJoUhcwn0uDJuVh3t0humiyy3nX1g5oOQY
vEvAF47EweQhwK6m5DAlxbVWZ8ICBlHyknK9c6lwWymUiD45PfCRLSXgT5KTwS5iV+AaCHk5IaTe
l3FQyMzdRjrlSO3iKqdYonoooKvKIPrKhN0oE/9s4+i9BvSjr6Y+a/eTYfT0oR9wDQBcQuDnEzVh
uiT5fOILBZKKfeX/pmiW/Ntl3ZwS1spQ8XDN8agriXMQuyMnAR+HNM2WRZWOXKxpHEtkT+kIyfId
VUcjCUfe6WaJeGGb7WXvgMJcTFJLYXD+lMVJW9B0n+JGLYYe3BZtqy2DKYQF+CINfOpTwVCFiXiS
PWcAo5GrwVbJ0TYhlW/EDAmcEose7smgB3uV6vDX0YaDmy27DrXtNQJEaRVEqZfn659F4I4/ZnG6
3UbE9mu7d6xwFazYCyq/5w0hm28HCO9R0TzkkR7NixTo0uDFDkqryJE6HRCjHoajX4Gz24UqEO1B
tGrvHIKgzu5A1B+gT0Xp9SgaRfh6M/bsxy3lOznvcqIKNCd13g1kVeK5zURYNWChwxRUCYxU5sA7
UhRKclIdGvJJpRffwO+gGhxpR1/UO93/AFO9Jcp+cQFnSdmLuwfkzeipGjycBoFSUODilWHIBeln
eMX9vTkIGwpvg+aO+smDtEB7+P6aXY1A6s7u3pYQYKWyCa4sPwYKh4ZcR8ikUl19ep3A8aEpWWm8
U2XcC28LEB7aF//ZQR9NQUxt5HlgaDXTgDrqBAP/QjcIpUnd5K1ZFbshLC2ZFySJj5Hm8tz3YNiu
Vrbr0IGM6DcHcTAuSq5BLhoAgAglQeVStC/xSt77VEFel3360s3r4pTD/19G51/sy+SKptt/CNnl
4SrJ/ZwNl4+Lkc7B1k/o4Sa1id4Pd+f8o+ee43OnxN73YlLnB0kti6maM0vWutF/wQ5ZZybyNHVJ
7vv9uvp8eayoNsZrfBVdseYESaW/MnriwAukXusIr04Kqe00hoNnmblXsIOZ3N0JYmvfsFEZ/i3A
4alVIZNjyL3hDJJ5lw3zsfzQd2YOOh4GukjaBbu8Ivp+9drDCG6BNvbkb/CWCWWWWx2LaWiJxZn6
7BLIsIYwohZB7Xl05lguHWMhs+hqw2ft50VRgSSYvSAbUPNchBMQrUIOYCsUqDm9duk9JbUfcVc+
1pmGrfoXtEWCydR8jDdSko2SMFd7koR0sX6MCJweMXpoepdyw4ea1YwlAUIKNtyy35n39R4/r+4d
VRU9nnQJt8jkgUMVr1lHoE9sCjaCU8JMnCHjalHPB9tETI5UyG6NBkGBry9lWmEL5ZmAebBlLcpS
W+exWqFHgaFO2hRZzNkKNqbea2ULxLIc4TAJmQmD9hP2rZecFg4Y0u5sCpO4hfnnrnrA0AZTg5jN
fjlNlFPV08cPsaB475WsJdI57S3dh/U+QsOAkNYkJ9x1in1ZlCML5CjhrbDmHBMFgxmnc0Lnp36A
XOdWGg8iMdjz7PPceysUNBXko25ZdGrG+8ItkNna5eLA3lozSLYGQmahAgk5uIRCWOmjIxOEQRES
n3g7VjxDJbxYC3EpRvQxU2aCOB51etcG2oIS/ht0NkdtAhVY4gaZ9viFFMsL9hvXmBGcyafdCaxk
RHA1RnEffupalyhdhn88OsIIHjjsOZZfPTBNiTB+R3PGF4icJ2XOdy6NCxzZqJ9qa8d2ZKjF203V
ycacTiyozYIS7o4q9huDDQ0G9DJXdKPYgJvwFPz0qSnvQlfWqVznyj7DLx085IG/NOVocfmzl9Dp
2sIWNn8VZnFsesuEU/7fAuiIg3tT6dc7lua+D3yty1jEkwA3vulX7r6kN6IBCfplmw+V6Fxuq7ky
dQH2xCTgWLq9B6DRRj71WRQQ0lgH7NvTOSIgjKPOi0Y1w/koq0kpQHw1v96PN2Lrq1guLMCtwZcB
YD9qbvNbDmbbBe+LnVnAKpjyB9PET2ax8K2f3m1HEYwW6OJAvl1su0xDKc82HO+n/HkZOAMAO6a/
A595tCT9dxNcQBN52EFwNOOwqD4q60GdxMG9M2+lSurkNMFMLq/8wn+RoVVHUSpHKQyX50tW7G+l
S7wuH2Eo6VakvrN5HtYGx7BC46/3TQKencGtqGV8Os9F67l6NF8NwaaLzhZC/Ygh1TANpb8hFu+G
Vq0BbMfQD8jlfQylwguC+arry6bthiNQ3BeAxbnHp87beMGv+tLYzzEN2RCrG7ZElRYaYt76GbtU
95GvjSjUkD/Q5GZE0V7E1pWjrzlsqe6++c+nW9guKVzoGqrqgd/VFKmIQuesmF/6NoJTMBX2tjAZ
FRpU+bxYZdQMgZMTSlCeOrUX+mbpu+ueuoAYTkkTZaA6y8Qr+cEnCi0Snnw0EtaL1Q8f/ksffKQQ
HwQWcBkFWr1uiWY0/vZlejZndSIXoRlhGHu4KSO/LEwBN/3sTQ5oVbuRt0OC8B1axU4gA8SYaH4K
fGu0BeLYcXVKne7UIs5dGFJfjQANrL0e2fnJEoQzCH0hZwT1B8KlFomR8csQWVAnMVlBDFZrxUe/
v9WFYbVezbCMspoF6DYDRHiHA9/94vANJQm0iTKcBCvNaiQQXnKuqOztTzk7BonOkulJiuhm+6BG
3tNMt1rcFzQPIvKy9ySrR7/HKmUhEUghv63Z/JEnV6Ah1CIKACsCdo05FQ33dkOT4UM6CShbYFY8
5uu7TPJB0ySvieil17PGCf0b69yvYAdnqfYUf1vbuse8CpwuZgCTJhX05byq63IqlJDqBR+KApZl
SDPCLvi+7Y/qYLAfqSKLJ6NL8Qt8Khj5gSOojHWVpr/plJ18kdl757/3xtMf2ejmX9usykTmcN3j
sFUDJwUIQaQjQ+ctOUSuVUUfirR67KmRKreS6pUCYAxYzYggTsrzxgobluPmxRAQbJP9kWzd1sYS
mYaDVzp7sj5h94lR3NhYD4as73wHM97qTW5yr1iu/hwD/a+LZvYoHEi6OahSzXB4adMiKhwfJtma
AJDwJPbtZZ+3WADxZ2KLyon7H08Shx8HHk2gRvcYd9wT+m8iHWFYk5eEW5AwDMHrJ/gE4gB5DmVl
9IR/vRoq+aSI8TRJ9D6OTtuREwdQdVFz36OTsCpsu0GUwabMOC0IXuM14BySj6HOVhRN1L+R0nKb
TXYZKyG214Kj6HKmdT2epPNBzwlCltyb3QlrxxKKUovd2j4HQl8BHbAmknPMmaIdvCxz6DBn4YmL
nuFlXr6qyIO98AbLg6Bjb68OPx65ilQScIvWw2T/ZJbAbKZQFWmxjZnESkSN8B5cWn+czPQ6Smzx
tPvcDrxrnvqeYm/MiekuBy3Z7GHCdXU656DapsHGV0NL5jpcWNZTVKLvqKhqnLZ6ljM40j9W5JFW
gk2sPkDPonSj5q7wctNDS0NxRAaPpJw6E1eJNcSwaH7ZBALkRet2q9fI+hPMlNmDrMuP1ncorSdL
yUXP073EY/W/dnCCqT+cu4Hk3Nt6QNEU6mgvo3hl1pgiL/i1raC+r3T5MMQg+b2e7x0QfNO/TVlA
LAp7vt4xGhy0lJnTB1PUiHilH53p3bBR6a//Tx7g4U5a2beg0cw4vz4HOYjqo9MoDHSJLBMbV88t
hP0AzAZgql7+XNGS81TDMNU+8gkmVKH1W65o8BT/FnmMKzVX50F4ro4zE6TARY6ZBc5hMlkznKH1
ndOwKUz6uLDcmBeKwicsFxhbpe2lwusk8gRqH4ueIeOVWEqppJdoiy/aouArKj5ikotLReZli+4l
DyHTCfU2YCmrq2pK6myUs32WtRRLycmUq+GmX/MZ/KwqxV8BhcaoyigMJBmSyAIrGvWJywCvUvv9
x/sAwVLryd1lRx1aOSoan5RIrhChaRPysfRwbKT+Yily5l9V94q9ckGGzEYNzw88Ir7RogvAndlP
x1L1pmKQxm4ovyCFquGGN/ZpiHnKdQLfTlECPKpKqEAsEZErbszGeLOk9NTRmAF4euLfdFBDFtcK
Jz5/0rn4HwJSuk78mfC2maAJKhw5GPi9pD0ktPHQRDoBuGP0umA70lnwwWJVTyVs0SqWk9QL3DBB
Y2C2daB9N0zsu5YZr8sr2HIfCpRUpPNeP0r1jAZyMRX8js88WXebdw0+h+pj7nzo8j2s8Yy0UqiG
vu/8MUJSU4Bh0xkC5KOy9mtKzTzMb5XC9T8BAI0chXxUBbvryaYynOqj0JEqmNO49y6xYeWE954W
VAUATO/8eEY7bunaAM07QfKaYIN6qvB7otd4iXzMlLT7AneWQG04+7Fb00fC5ktK552Nf9n5wJTy
uSGP/dc1kg+p3N1bTMTpJJOkt5fDvWiRej7xmrUkJw4dcNm2DiP47LUqztudVyGE6IDJRcmlgQEN
Q9VVGkYF7dPCWq3QEo0VdmBcB2aQEQ+iCbQn8JuaxLz5s84GWPykvj2XMOf9K7wE9RlqPIV9RmUX
T1bXeQcEIN0yR0GbQ2uJwH46kL/07VTGoUWFF+Qsla4g4aYy/KVi9CdINJQI9LsIfzcnC5ktC1FJ
aYXcC0Rk8iMwdtqjYGDDrQoCOCL4+PVZV8CfPTR/bPNgTcQGlgNcznlJEGaJ97RsN+NLc6sS9k3Q
XvJv+jo0eS7FvIBbKRnne3+63UZNpDDxLd+rL+ob4qom9fMxqQphV79orDqSCo9W+BYX0h8AGiSa
bK00DkGkAxmAs15LlyFquU6S0M1X358NzBqnCGMPr2cW1phcJ/UBBD2WASyHS+n0QCGa2/7heSZV
/eYUT4os60B2UXf0q140gGxbRfsZtHJuEmYi96ETFEabfYgGfWlh88lCsynyyC3EUMu/UlbFjw5T
sdk7AxeDUVpgyovkV+kHIzLIRjqx9AYwuBfKt6K+NJLa4SKI++1aYOVOwszO+RspFoYwsdWIoYd8
XPZSS6KcsZ3/ZWjUD0gQXCF3ONpP0HCPV1iCIX6MD/2W7u+fSj1wRsGLEQOe4m+F7VRISr0PSqTQ
THtPnzL6cuSGOJWfZ/Pq6eweGHSpHag426pLlYkZ8QIr3Ve+6aiy6lwp04ODFRMwBaJ724P8/Hkz
NrPt4pqZ4ws00RtZaC5CO8BO+RihnJ22eDo5XlFiJ2G5gO4gpZhHaJCkrsgg5JAsxEBcxj6DcLiC
Ibi71sUwRH7Xz/+QS6i4kgU5G3QyP3034OUamCqNpl40Ps4SnGd+SFjIynzPtndGln3/qf/b8jur
WrPaQsicDeLU/5/baH2tItnlOBDy+Gb20o/GD1G/pGROu7jHAdgHu+z4iUdpYuDIi12ZgSfGF8t6
m1n6BANE8rcX6slye7ARt2fZ099d1OPr46KpNrKqEilHP+yx0/ybL4j1+bFcun2RUzf90nHfwMX4
01bNvh0mYLY883UE6w38e1o7bfJ4A7eY91bABBTjMz1R0aNiy7C6ElwGQrZBo7XexIoeWIOCFWrW
uWC/ACfaDwDmHyZJLUs3YA2X3C5mZ/4/u0X5zbcObyCYrfXvcoL8pFRXqjxchTMQLAr8pqf70s5k
pHmdfwgl3SVos3kSnqWe4rl42enr9Phi3RbZs3BolcPAUCgRdtAcnzWGyijERlO/hW6G3cZ5xP6V
9PH51UV+V7YUeXLOWI0NuBne8Y4sN0snVastYQYuGxp7IJS9MhOHY4LQ3k3ZCKC9KHW991RUuGNK
G06sOI0Dt+J1waTQSSerGkQWFBDtbBch6jnC8HL//vdJAt2C+Qrh6W8WuBO9YNOJt03dc5YUGCy9
cFmpksBL5ME0P9SGaKKAKobuG9P0eI9HhHmk4O4UpnbHf2Ro1AiDasHK2z5Om0jbxvdj1qruxLbm
rsm05vEzQDKhUMcxa2g7OAQt4THDLsd3+kv2DJqPIfQ9mPsiULKgTCiXIaDV5LGnW2dDSYMpEMp4
A5WemuTVPWr+A0XxLOjg29VDJ2Iynt2/5zqGR5tivUuvqRSlEXgAvbJmvVKQUzoAfoOnRPOV6oLU
ywWin1V1z0BQT4uULPcZdFxdLtrB2wixt/gSBZb4BBIhhAAFAtaa7/WcH62TkkP9ySKY5jqRyJa9
ZKkNx3x4/tyLk2yVtUNwTnZnTOnFzeW3/j/K9CBTiJhjKWPjonCZb7GIrat549IK7FrFlb+NAPhU
BBYO7tdG9n6S/2lc/7G1AEw+rbcDJ6dgZdDze9ElDQr/S/ixusdZivEjj9n4CTmoowfBJXDjHGXW
voWQCWQV3WQ7qLELXnndVsqWnunaCqFed5ClIN3I+U8H30Ncdgtxi1GH+aQvlcPFkurYiUht1LW0
m0YFDrHfLAr7kfQD6Qvp7mUs1gZA2z9nhx3+Odj7wtahgE2STz1FvYT8RotarbAbEoTQ4lcqcnPh
QMYElABpqRilWe5bcVONeDcbwc1pzqCVtalCA0XDrVMh0x/h5euOlrI9BhXbfJPDXoyMX8dXBvop
Rv7Fj3ahR4FjHu4zbUQB5xtk9xYyCgQcm7fdwjOxtDLxWD1UpiJPUCJy7AaIqXNjEhFkVrjKE4wt
IfJ62/Z7YAfymzGAyGViPcBllLlVzLxQ78v7L8OftIdFEtbn4pa1+TnYmAIhG1cNubGn99Uqay+A
TkxydctWo/qzVThL0bcNQ5Jx0z9pJ7QwSRfrMRffivQRVZqeu39lU/8ciBj70/gOe32szEud33Bs
oDlb/9Oerik3PFoim/9pkTYNfT0lmOebodb1lQJIRlQGgkGhnNQ+4BPrIvkTU1HtsmBYb7LiI+f5
91qjDbAaCOia9h1z0ZRdyC2qYOob+l0VbHRyvNIFrOPlEub8ElrEyskvEkrN+D9B/VwtzrERxZ/q
1MrYuMK8u8SMD6tGYmfZg1184qh4orlYlboAQyd+3Upmy1vOCmVEHiWogw6ESh8gcILMlHDg75fa
JOSg1E8ISzvUKO9FrrdHva2nlDcnPPRxP06YVaMPrslO8rtzWUz2x6xXQ/kmNEyO5mosLq3FVlOc
TPLpTIEL3CZgDNY4UjmlLYZTAxW2ndnSIGp4JbLEE+HQbn/TXQ3BSTLWd+ZDk/3dHMKJZPL8Gtl8
ZGQxq8Fx7PZh66XotRj3zVyQnh4u94/wgyMJvnKKwnp0i7aLGw+dvUSwNDqwhsYmQyk4r1aEGFj7
WW3ZAlKjPWmhcSnfWZJJD2yqtX5pr7A0+kLwSE9EUu46e3bNHOqjL3OgweyQikaoFlF3HGpsDy7Y
gxh2YNH7ezx9JOv3FUkKUD6WqwjfNxqVLqeeF2PQRSl2ZokWbDrex02cA72Pg14+gIdej+bQck0t
yU/JVWLltFbAF2wtSlte8uEqEM54ArjSjFLK9Q1LcAZrR4Z3ecPbYLQH2E4KmnhPQ4pwQ5CnRN21
+Hoauw9Rc7h0xne2f1bKKsHdFMd/ZLnWo5hXl+YoL3fZgNc3vYsCubuOoizccu5QAUeUImFb/LjN
3q/IjgXv+q04qTb5g6YPdw+7TLjh1XTIEFG53l2KSITJXVz7y1n3HA7TYn6xjXmg7KyOpfZMgKdj
m13Xdw8xNiRDthJU1Mryh6/dCuH1+/Y6Gq6caBnUO1k16sniQUf3ZpaPEmviB0zEffA8b5UavfrH
K5ITkcdyw82fIPh3jTA/e5p4MaQGcJcarGQdcs87JWIiHCLwT0tK8RKevavai6JebjFDWkaemW0f
JbVWj//gJIdC5TjTi70Pz3Opwh/jGY34SGvpH+hnGmgJz1O+LDLKjhUNb27fMoETNqowXysoRN90
BsEBjwXzAlyqOsTnVVVA7miFEs/zhEWeBGnI1CfOOYQEPWnc2WQtVQFFNWCCZAyAeYo5KY1u1lP7
VlHF7qZRY18H2BWWpHES6xLETVpAheNavG9KX29zVc3xQhswhEDCEEwtfKoXg11z5HoEAvQoqMBB
JNZW2DYjqa55r2tTmCHvVd3v4rYJLhsVGPFbBhgJ/h/Z5daZUwfwooq/Lb/I5iwyUb+Z8sj1TAqd
5RdqZCCH3KLTtj4Fm13HF8ENr6qfdTEoo7NUqQ7frNePIi6A5f7J4coiS0OSzwMxaqILzFx5blL0
fpXTbFuQBek1bNvPCTLpv2q5bOcr4awIs1djultcnhPPnUNBWqtESpl8OXMEPmBflKwLIidf5mw7
GwzhZNy+LneD+/HKCDI4Yn+UoA2KRYr/SeLQ08g03a0k/m5Vs/04208i6Wh4SMSNyLNJodSHZolh
Fo5mz21RmZQ8nVlxnR3gSqQvy672Ws2AfrxUCsAiYD48jhiQTlJ5Wz5PyLk0V13+BCX0W91Vv5wi
IrAE6GSJibIwV70P7wgyIyn0lf+c7DsDTja0kb0kCPNpudZMdlR1S0PKQHVZDhJ7qbUqMMCEtrNz
PApKcW5kfz+m2X1gDQJS/baQSIqnaHDWMfPC/6cGfYrco6yeW481gp9spNvCncke1c5JbShq/D6I
loACTdy0E4DNAX8D/qjUmnVWShdhfoo41N+HrwWyhi6rDCSwhuLsyVgAJqeiwCr8gFFpA9E3wqsV
WcsuveASyBEfy/yEQAkq6Fezcd12gxaIIc2K0mrcXQs7AiZkCfj01WJQXqvIT7W64cQpjFfzQXn2
2fc3U452yHDA09V5/cA1GNXXY7Qe3FFgwSW6BhPBnwe3nGmU2n7rNHd7glHcKZldKyNYYOfjvnBb
f792gcNpM8CS84TERjkyroeut3ORooJHp84fuJx3JGjIbhpaj494SREHh6nm//Uzd1uNTe2T2/2v
44aNnfszj3Mg4UAuRmbb6eiMv1UYgZbiCuE2ZLubOffAI4uNnDqn5jP39J9sAbwCikw7UM7yWd+G
D9jhzDFpZa/0ukiTCUiuFcXAvIKMoFA4ZelOjMkL0gng3i33IDQaNIOS+IT7AzTZqcXY2WdX5EAP
1g+FlhIXxEoYfbUExTd7zFsFvOOIrr5bbzxCBw29bvq/tYJtuzDrEILF+DdaKtzrwYuK46XaFLNh
/rh239523oXFwDKH/DlP0dbFgtuwj9Z/VryTtC5rXS+9s2qSEWDtpGbqFAAzWLLa3x+PAT9VCCWR
refx0KGgo2QqXouB7XUK56Eg07NNkcALks5w+IdEyRfS7RfCM22Aw9s3dhEPuptPewbKOMBYXTou
L+q2eFVFkSMNivAeCeB2QZuNNTGzqt+XlYVbazR2Z3X1exwJMq8ToF5fbguMAvkdFJ9P0adOz4Oe
L/OtD5qofbVc6k8KfrzL1rVmg4vyOVZ34SQpgSA18XV867N6hmTcTG7ZsmkyPfxOCneyBye0On/m
SaDKO/8IICcUCOGvRy7fSztcd9TIUfw+abQ0njrd907g1VH5OmNYXHmjOYuXRxAXzu/Vks7bgHkO
MvdLI108f0cpevapOsl+2676ooS90UyV+qDAQK+rCVdx+8CWVrRTdU6hutmmFX53orQFWcriGI+A
R/V2vakDdGN2GpiEWYfdvT4jCDUsnO7DdQjumUMonyU+ZuIQTmkLD1ygVYKrRPb5maD6FpGdLD9i
2xvij+PcDMVvndRynKjkwiPFa/T8am/eQ2vUjWpl2eeePwVQUE4rh7bP//X74sa72e7IsuIy5dcl
C0jWVTPOeLnjwPfUY3VPieO0RZUyNXvM8Mz/7oJd+f9wT+eWxFEC2DMJagbILhuy1BVuV5hZAMVs
uRLV4RYwFVCQCy77fniOqkUcgErHEiA/Wk6upagzAKPhZTdqGv+y1AHDE47/VOHwit/FqafOJj73
h04AptcPrd3sQRNn7rapHf5Qa5PWnADtjuETDh3xl/j6kE6yDTrplunpt35GzLocokLDlX81N6DJ
7RWwQntAdVwXoj0JY0xpD3n2IcMFNFdkhk1YYtLdi9/0PKYkxDcK+1Z1ohiHqEjW4iWPN5G7Hxle
4UPbkhgfi6i/Rky/+IRbsbUDzJBzdHVDoMU3kviDprXY9Ibfi5o7ONnpyZQvT1tSwpp+GCulL45t
VeU0n2c+UrQrbnKduLdL7PEUdii5jjODmGCbo9iC5JtUXZIHe57XFw7cCsNTdNEPFNiB8UrzGXGD
+q7XzAfv2m3E0mGHfmdqB6oAr8IZRS7a6+jv7Go3wjkCIBTNKDkHJ9liM3KREuvRpS+B14XjO9xr
NS2WV0at9Ba877Z3HVTNj1gCGepv2WU38gPFTWbDC4vPr7VoXOlogRnercAE3c9cmLNnwopBfIyB
IRMk2tcr5AP90sjgRjcW2uuAbAje6Pq7we4d2vnM+wv/XzAY+O5mTXRIGam1XVzPWM/LqUd5BzDS
i3n5Askn8WYqqxzQdpvlX/1grRqQUQT+jvPQP4W1OR2PhwLfSjbAqZH+MeZWuJKMP/o4VwsRANoz
CRcJ3stzcxDw08E5BR7ssoigEBIUnO9TXgVhkxJphSR9EAuCZHA6+OdqBFbiAfAp0nh5tJJe/T9t
bm/DfEfjwK/0nML+6KhhK/Ceq6rOCUAgPf+GBQ15ZJUFcAakrAnyvTFqohJVBfDgVvd8O1p3A9M8
Sfuu3PmCg6oRUxzN/muKh48GUtPofWlUu1MHuBP06huECvoElXbmxi2tgLLRyUXgkkCIZ6SsJWAJ
Zh8EuZwlX1groSSOiTKzK1y5NH1aUT43cZkUjmCImPGCAl2YsgXEb6cd5zzK+caeTImcpewlcxtW
PfVwhufXC8lpOSZFeGDKfWC/kQoSHTiXLBBMYhTIAB1AZus7N8Lv4T0QLqgVWtRoeW/orvk/+zHC
MTkWpAdHF/NvIthv6veJ+zjo4HrnngDDathrpa76XpgoKeA9LM3rc6GGEEbi9yAT9QZx/tr57ccc
a4sidWmQvPyvUnP/KBrNj6/Ur6dyW8Eiz2xr0d6UTJ30j8cDWRxTlYBsO/RijjfXJHwucRkVbL1r
v5G4IqsKdYRIpsg6cN3drkxgmhnejVdFhTq/AppGzw4kzxJvlnOBAqmL0Y1d9eae5EoZ5swVBB9h
FV0iI7BzMrboA01R9rqZk/T5uRUxbhLH1tToYDJ3uirBhHLsWvdtpw/rwhx5vITuRM+a/YOEWc9O
59ccgp+yAiPjYzX60ZnOb75RD977T3xblf9v1bWDIJNesRKQ6TUAj7fYxrcZloIoDpmdUTutWYF5
Efsm0wvW8ivrz9eYEbE5MFQNzeoVNpkDw7R5A8KYCdizFmYFxWgrSFmBJ8+b899OtsJ+MBeUE1lD
XXhG+sFLX1gazs6aC51t54JrZaAkqBfOBN1Np+H+rZJ3ejFVbhG/xBT82YO1WW+HI3r+5BwgTlSg
4VXNtgd1zwoPcY4ccCB8pRSb4QQeF8acvO2PcgR+J+28PaVLxepmo2qzJbE6vHgpn6Ey4qMPl4h9
ghZbHdCX7WkeEzopthKi9HwaZJyqPaqGvbIkY5D407T5PeUJkgXe0H0qMGN4uQPJfVXh7u/hj4ms
OI30Oz7Gq4WXaoLMuktm28hz3RQWcaXte8lq18pJdpGT2sOBZZtkjoyPmOpn1dcQKbmA/3iqFry4
kwlvKTXXVnercj9eqhsak92enSs2dXkIvATnu4a085pOfbud673qVehKhQVGbT9SNOtG5FavJhtd
u7lMC6NecyO/aE1o5NoCpRAuLSY9FcO+XiXc2OCq0IbsJTh5O59ddPOK4p9CmrycWQOs5EY4BPKi
IR92DYsq6EWZ/PcCCpoF0AYJ2HA3eYQZaHSWb9H3odpMpKHXCW1wYBV6OzlPdDARn0OOKouiQ0+O
X6UnJMNTz3F1C7+7diZA96VClFnZ7+e6ZwJVO0AMOhhAowbvajlyF4MtRCkVempjsiX/EpQFahMK
QHnkvoU89nYTa7qzDxXMmsF6+IQMKWqlr5CkchHIlA03AsQcwhVigcV2M4WcJ3x0goaiKQo6Wncx
osQwJGdA0ZgDDDGBD7EG5Kktu8kJDyd8uafosLMi2qQpqOQwlxIPd9VzOOaNtoBJQI4nkU8AZiFh
e5e+G3MqRxcqQBlZPf4wuKbICaoBohR2BsEbVDoUsC1KnKxj8nDSnRTYxPVVjaEKQcqKaMksG0lq
MgYQb8U4Bc0T08LhCmTgR3574oCJxQqVVv9rzFNSWt23fnVO5bSHgrDy0LZyzLlsX8ztsbjLoWSM
rcxnVY5SwyXbw88vNgXuB1yS5fyqVCtm0/ve04HD61qg2pvn45cT6rHjpX2wk7EKDs2Vy1xfYNJj
6ixJ8W0aJ9HAmjykBqL622Fm4R8BheAWZmwxctJkvZm3yPxBx4e9c7BjfpemNPONwLGwSI73Lvep
wgKnYhd7sTeOjg8VIBXuybmVQnQTMB0EHQDIGpLmsCJ0ddm6ulDcLuSdwqrjW38T17kOkypYv1Ze
LKJDbYpEsXPAKdlNNFE+3lJLaeHNKZCs9oG80I5dNZSUFUHh1y5mZODgsvn5SqxwswwgZhtzdXR1
QTng2sxOjc7c8aH7X046Um68uOBzPBFHSapE6r21BK9uohHL8SbrWwwZDJunCREgKdRvPbOdwe8X
p7TQMUiKoap2R1t6Tu7wOs5A/dX+VCVdf93d7rhqXs6IELO/6vebITQkVVW8zyLAWM1dA7/j8XsS
YUvTR+PEvUXPWMh7mJYdX0ffut6lrWmkc0xkkKz4VkHsAvmyWEt8wiuoXUTPvJ7AXInbjmBJ8+mN
0I7uU6AkpvvCfXAQ05sU5iB/jUnRdJNZlGj9pfrZ5O2++ZdNSqp5/iyNVfrE4qdxGv4NXCpBK719
1Sm7MLL+p1jWBRc1jUkyqKFNv0k0UhONwippgKXEtKvYTrtVH+GL/P6KokoPtd/eqSLE60iW23sk
Y+jKrr55nr3TCW4MLLAAg+nm0pvYTNj6dwWL48ZcvAcBp7FaixHA6JqBVzJji9ZOKkJSV6fC81gk
5nr7IuuhMLo+xI35BnUWMYK7DOfIZWpx6EyAv7Gjcb3ndK404bq3sA0DlEeE+NwxpuvDhkZXf/fS
+52w2w2N4wJBf9745bAWQXvy+MMuhk/ssPnrV99CA4SPlkgWaKrloSBtXvwe6/+XHOHNqaRr90OH
sQmIDrWfu7HXFfXfBAsx0sdrjPpjG93sI23actIBz0KoA88zJ6xVvcWkrgcaT1VkpgpwJSneJ0Nh
jzaYEmTinZEF/yKS1Y7J1376PJx9/jhAQyx91DoOeCK/WIG6HP7EC9emSLtqXtbHXI1NBjo6ZiSi
qTnIU97IpIQPuY6DKgvVjqikPazGBhq43FtD7QRgO5K/DCuXomZ2ie2s9ke/Rq9SEiga4WrYZjgm
fp/7J3s/Cz0YFvuqh1WhPWPpcnoMgj8pQTjEgI9E9n1/jCpiq6HC9ZMscYPlS6DqsXa4vzVJX4CS
MSsEKwW6FHijmoNZVEZ6LBfrIQ5fkfRzILTTmVXAD5sUTHt3XwyJS9IfNXZ+bpHtQFr57GWRnRe7
0PcL6gMgNqVrmxEY0F4NPnVpSk0JiWm89TUW9+LhhOUsQZ98NTIhY776V9R26Sy4efHW3fOsc8nT
ppKfeLu/soJ7yMjO+iPyQAQgV0mP64h/qx+z8dNp2tA/ai5RfgJJaT6dyapNr2VKyzPG/Dsxz0Xj
4P/MGLeN69EH3pmo6O30n6eiALrGvCK7zTlCSYUt3NytjUhpw8rngwfm5LKy64lvwsXatRpr+gdv
SBUv4g4OnEYjHZy3/4a82MoDvuxRHDR2CP7NLg5KCLPPemWPBh2VhXuRorlrO/dhmB4i6f+hIvJR
6bt6vN0LbnrdnoVzH+unqP4acjDAQgKva58yo9rSpo1+ToEkrZ6t5z8crByde+wtVN3QqMaXadAj
t/Ie7kEb2t/IH1N4fhtP1g6FyNA6KL2obxBht0242/FjZLrjP1CDXikYffmAGcP4QA7eAqy/UZdp
qY6IBMe3klXiHyJxGaOupp0KgdZwc7+CPEIZP2huWLoKQWmSaBgs2D2Xz+kKa1iAimkt5vnwnftE
qqG0ZOesZ6LSvNuvRpYqM6D+s+FqTshFGhmLClNY0JpayVV2wMSAc8HD5ZXsYmAo9l1+TiDfrKiS
Nug7Fmrl7Mmegt4FvvDtQc0Dbtb1MRj6wSJWEIp/jN+GVVaaJ8iXKfwelMHkx+GQYkMVcy8gEZei
fJ3Gmcto4SdcOpAm49uMx2PQ7Y46TMIngIfpEs1czYYbeM23ng1VP8FCOY2JuVd3R1oZxs3Jrm2B
7Wx1e2XGoj0M9gSS04I/wnvjkiiv6w4eIuV9/4Bf4BUzlcEK3F6W1tj2Cx6Gd2yIczQZ8KCpWGVU
aR9TKp9r67kw0WBEzlbJB7M8m/Vbg8YtblXkTFvGqmIp94nF7lVcR/Wif0EZ0TPPQ4roIqKudoNO
Gj8fsFM9C5birPly9WTIBP4+f4Hxok3uOFfy3jXoNUZV3NcnlLEj4JvV7qEnO691ZvvvFjAqUBc+
hK1H8P8BLDiaYEEWp92Wt9uHgCdXG5v3Dpi2cB2PGzk/cn0fUgXB7WAL0EyeXSwkjgfsx8Bh7wPn
2oaDaSrp/lBvlZb/w1NncxqRgFN7My+fOqL75FW6s8xlCuxX3QRr9GM7GLx9NPbY5MOlAxJ8GGcI
/MsTzr8Cb+21dKud+a9iwobDGV2QawXyskgZ+GgDH44okoi/11LMIejy36WQXuLl5T5GqNyfqyBK
TtvFEPRAAOW/92HYEj0B/CYdlOZaK/e0G+FsFdvwOB1vMgcVsXH73oEzsHZRfy/rW/TlCwJ+rxDz
6XwizA22OFvRhxktF8R9aUAka92dyyjtW7HmjTIW8MCU8qiLf21do+RmuERMLjNblaYgSDrWABB5
LECDYMadsT4Qp1Hkb75+pHAS9Uwq0miwUEagnotFoQ56oDmtleEI15+QqCg7HjPiDguSieaz9FeZ
H3z+BDf7mAu8gbNgWDCTJCatxf2YVat86jnVfkACSc+K7T3T+vaHyalurpreakP3v3BvG+YoOlYo
J2NDU+DCsJ0hgNS6KvOXop0pZliJlEhrH96B0TnUKIiXIu2eubEGYptT65ICYmctCJ+2ger62zJt
jnjp2Fw/Mawb/pYGsWhz4q5H2BiADD+m/a5cusYhCQdXvaGgIL7xl+NrLv/qcFJ2tWnSn1TjrFXD
kueSWH0GXM/swXwWClwffSvFoEEh552ybtho3gZnoPusTb3DN6qOAa1nLaSmV2c7zhibux679SJI
RWEdC8GqEU7esqtSDkXa2qh3CyrfPEwy3PsR3kvMS6ZO9KMuu+eDZaJk83GlUKCcYj1sUKD+L4om
C8TiQGGxdFHE702eYWoV/IneNkITX+zetsUpJTmsACi4hpgXiqltqVaGZOgOvWmNrG5h2E8ZrRne
+9t1iS1JwSkwjL+HgoLokBmVlrdypRTg9GQTWXeO3MoM282dkPX5a9OrdL0aluz8fgT0S36evoBQ
3L9Q2YPvwY/ENeaEpCMBi7ck5rNrC+J8z2JmVFSg7si/Em2fPC1DfZutcLTq4RyUOLvtlEhHJ7+7
3VrXFEbaWoZ9lDoEHss1vHQnQgXU+gTeXkRxiAO2Fgea64u5LS9yMqPC/P34Wt2JM6Mw8tWDHpM0
dHBAu77cqPpnWzG2fhYIGWS7g/CEOhWDLI0nHBvFseVdkR9EIgWWKabbVtwJKtU287JSbDlVM6qM
FY28BI+OiyjwLGuiS1avL+m+83lnt4UPmf3VUBfLtOsAIAB/RSyrk422bn+wzgJLOug+w6c6tnt+
TK93mHIiUr/c8uNcds+9dgDTYlNYlGT7gqYHcn96UpCtNPcp4F95MStV5LKp98cY5dgNf39ySEdD
ncxBgy2m6R8kivLgw4XthEn1k3YsEkR7unutbUP7sL23ZqAssiicU5J6O6mgdpwkDdQv9rEwYUy4
IbOYmpOu6tDG7yW9ZrxXNsdj8NuVE4Q7fbQebWKZj9+e5eyOs6T3TmTkGk/wbxWLdYNZMfDDFdnk
f2qOjc3X8VTMs6rCxipZjXAQmTgMTDJjoVf0aVou36Heu48p8YI6t367V1nXiw6HWBH+GUrmNUVW
aRAow/WtHKzmjtUD0G/XraLvWnh1WvMQccNc3Z8zuysnqxcC1QYVmCh53qOlVzmJrKuosT4id2Jq
L93hP0jHIUS+RLiuec2VQvo2QK6Ywkt0gyGHEptJRxtYVevsCC1c2mjZd39hVTs7n3/vz87YUdNq
fovRBd55LFNsmmizqMbfWLDhnbXqDKNmk+SF+9SA2mvnqhBYc5wShUxtXgqlU3jvucX/7PKRTU7Z
5bAOQjOxp9pxrOPeFavBi4kdxw2HlmCQWSA9NbZUj5ESXSBQaUkREoOWo3/8gFg36Z8CsZAQWXCX
l6GOaHe6n4xZDVGE3RIjx3haXV6ewAL56eNM3YRILo6abclYidf0q/z5GynO/OCXACl/vi5gqGn4
Z4ZHUQCFE82ch1EAephhE6hBIzCWWp0j+cJlM33LXgWzDvuKkvNNpCIWhlrXxAsCm/bv9UV3kPwE
j92wgLNm4RFJJL03hFtLaBSZyIzYAdgk+aGc7AKRWEFfcDsVWxmxqJEoIKNUhF6i4NAvQghthIfH
o8u6+cStYC6Sl50LqWW0MiD12egFX6Dtrf7nKcCG6zzlFCQjgGw3Bs0EQbX+jHSHa8S73Uoc78lP
hXZ7hC99PGr7RG+TvLtmtLXEX0SMfW6RzrYeh9QcSTiTr09CJLZOHwKvtov9c2H4k3iDzHsdn4AK
EVQDR+bu0QfdExn6S83CXiC1/GipIJEqiAp62qA0Lk/hk+U0y9wIWfDnaCKPYrSy2mVhryu4QyPQ
uimovqkATfvQD5nSX81G1FUUH6xXtn14QSD4ji8mFTAInfRWws6S9OSPR29UgEE1KTl1J/dxwAsN
0fwzKokhfwAqcQEPHQdI7OkALsy2Vmmwk7vkGu87iOttdpjnGr1LK3usRNFMaddB/yw7RrsButq2
J/zN7KwbxTpZ/FKsmHXlGnfxcBZi8CsAYhTzQL75a39QwKIkjPczJmcIH4iYCCXtyMVkDSQ5BYaC
4VIL6ORsfhVuW+VgGNHRJX/rSY5E8IUocIg+cSyB1V/NCj1Kw+WLMLj7Q+mGNeZk0xnDJUEjTEQR
nxQl+4yvKW7X2CiFoPSP6U6vwYRDD2WkfE6EhT/lmbmg+pF+LbWYTOAG/r9u1+jEr8i7CHnq6x4F
j4Jeces+Lt6eT4LC356Jv0a6Hl60kV6YDygV4iMtGitA7AH9vmvejzHz+bbG/HNQnqmkBCWHq/M8
sBuGJrZ4jCRveCiGKxuKN84fI0DDz0WkzCGDwXQkTuteHz8wwuILR9zAy9qTv4I7tvr1YUPaW7qQ
qtHEoff8awsfuFQcuf6y5emsV/GhVEJNzmdDM/5W/8w2B6GjqnjyIJJtbqXqPfxURMcYhdZZ29Ve
sCGlBchiBN8kUid4IdTJVwJPFps7iK+PLqzIAWjzttVAkR1N2pO95QD+pHElvKM2BhdYP77AILIf
D16cffz9Azphaq2ki6Tcwwx4PibvBROwUrahekzucrkQQc5Gd+nOu/jBYEMNbOtQSZJ4pNdQu4Yn
cft/wMv6yFpceGN82e84rPxdWx2vnl25JH3j8NBx+PQP3W9zpLEjSmsXWii+vhj01WQneFxak25T
bOqUYC4Y9oDmDo1PY3tZRHGbr4T5cZ5MNXLnHNmZVKkefBz5a8PJBXyj0Ud6WU+xJFWx5JV+ogz/
y4gjMdYtJCcy/dItA+S/R1qqOMwZyY9c1A1VylaCo15rDHzb+4DzB7gRjcE3Sb7It8ZdEqty9Xgd
pk5/gY5U0wAo1gVTmLV3nreM1uz0clMZGCHRfqEM05byynCK4qAoRroi0HvvamUvoGA5WffAnnIk
8V9M7QC6A20lXwkrNYef/OB52TXYs4rQEzo8UXHHtAikj9IX9B/QvC87fxO3AAb20mQkqK6oFvcG
X7NJLQ1NwQyyrg1FtPYqn4MnTXbQdyhXt9CGuUKZf/y0NGt0NSXP4HhFWH4DWX72Glm7alNoEMTp
fWVBsfdD0glg2LuodJKwAdqmhnF+H9w7PJJxAuh8zB04GbMLS+GGqItNWbjCY9yZqSRdxl+b/+uq
wwsWx9h3SptDBswVBddona9xKP4fxxTd2Yg84mPxIfg5w3Om79fe50SoRdH+HaN8bDjYjURaCFxy
/kUwQ/COEfyxw83VhVlw+cuwTBsjQ3GM2jc8GLidV3tbOafSoQz2fDwuKXTaBQyHsNanfxCuDuUA
z2ecGWj4tqhp6G0Y+nH6I5llmgnHVcYy/uuqFCUrMHLaMgNFf+bEEwcBr04pkmYZs8OOht8hXjYS
Jpzfbs+wQUcW5FsTNeb3coUM03jSfgiXGTmQRPgSEkThm2L+mKNEKMelIqNLMiHm32qdQTrnjPMF
iYVy+vwIxfxjMLi5jbRju9I1vNBFsGbTAOx6UiHkiyK+C2DbVyJnD/Olo+piT4f31ahOJ4YXLzIk
6DS8IB/uaY4588ekAGR9arDWZwDR7aAVksAOc/yDGWgjoQBDyQESYnuJNizsho7Q2rl2pq2mKIeK
wu82MDN4rxxGoGrPy9RDqQJycgY/jqGVvRGHEGpBDL9268Ra9Cwfp8zoTalDXPI5i2RgKyIjUXct
DWOF4cIUiLIV15C1HYyEiqBvE6oEJy5qcV6X1HX41UBwo5j9h2VAnp+DwZDPj+DVbHu8NwuSuwX6
FdqigtGoHQl0vete6JGmgDaqmg+caOXo/j4dlYqDHNtosvIx73D2QBKMOz9pHF8guoTNcgseZJBW
p9qRrnOXjdISFbW47VmSfGlX0iee7wZ8OhL9ihvQq7Xf+zczSOTJ/YWHgnOqoS+Eu4mkUO661eHF
trgkBDJFsyLmu7MVZZtG/B2y6UK2wRwpvTTEyPhbbjl9FBNQJZl7vT/NCCey5YwQO5dE1rcHHKRO
QSIbc57H9HSiXdzUJWlwYNghgAW7Q37a+c4Ol/UBy3z3xxnHkiTaWQ/pIc2PZXoxsaWOMFcRz0gJ
eHCUuyFhhREDXuKfwp5oeuy8l8yiydB8ZxXQD/0gRCDnyzgeBNgwAaP/0b/TNGfrh4CgFZ86dM7O
blcbsVlEB0ssRWHrUsYszwB1+Z7oGadbVsczGXyUbrgf3wElK3Gqraiv7dRBmeFCVAgfJzSYZbpm
OAHUjtI0LZJEbF8Hc0l+7Y9DqtiI3j+TyhaA24tbjtIzTVeRxGku26ey10+pX88U5xMKhMoWhIvc
x7G43gEujsA0Anpl0Oa89Jy+/aHrAYjEV7qXdC5iwcbyvYDhP3ZpRPaYJMjlqoKB6TXHMWlmfolj
jxI/KsdNZa+k4qX856j5YDqePnNs+OHLqV7Vc56AcM8W3fNmasQ2m2CSs32x8TBsWG7UWuQSFU8J
/5a3Uubc9+/KFzrZQggT9GADaE25LG3/eQ/2Zfa+JqWB2VpmpuEou1DdkVeWXV8Q5k4InXMbHCaY
Yhq8unxU3DtMdjZVWa5u5qmQVgxh6lF6qUclZK5ksQMP5TOHE6A8GZQAitPs0uSIYaaaDj+IMkmE
50c5K8Ag8mC81uokwayi4mCW/K+jtXfDRWd3o/b6+kLeFDneJVwmdhFs7drJMZCAbrYq6cXR3bt1
tXjNlY4kiIh4xTSmGtbzZzshwTFULhS9lwjGzRnXmt2TeX7LhmA7j1QXhL7tRWiWJQIPVbYrhb92
+KbkC68Vs4Vf/vRti+SUo6ROAdKePHBWXeZbyfjSt30ZW0udQ6LidKUbzM7UOn5T05uooIdxico9
amB3ye5cidggF+BZOEQjJrIevRVlR176Ize7/1UhvUE+FwOSX104fdR14IvRaqzm3km3kpz/i+Zs
xdQV1Cmsr/aUM6D1rrjvXNOXjbQ9DOFwkkrfstVMjZwR4A5JyunJYcEgTRj0lmS9aPKyIgp1Q/rL
8DpUxiMUdzPiIoM5Kjf5Kx25jY4tKsXQbJREvKCdWRmp5ZkYteF3dO5sjcsGyRfwCCrQbhddYQl9
qI4oMB2cdcxn9gIOW5ezSdaC+0Zf209YYgBWPP+6NHk1XlYw7triMXfXIq66wg/q581Z6PqYu26g
cZqzqgJIbLCxqzPLHEwnSaIZ90ICMy1Wb93iTIfcvXfKdfqbAlqqohEdCnmufhRHJOMcP2POoXXd
oO0YOa1zfpZTrbymqSwz+fWNrvIplEMireFSC1ww1YH2Id+u8NxC4aQOeCkv8ygi8O7W18PAxxPX
pU2f66UPDgsBmVpi23NFbspT4TIukFwo2mx//eXufLk+TBPHVgWOXwhs7s8VV3JDDH8ASpeW2gC0
wAcoSZWJFVjrU3KBu0eQV7DYAdDtr1DQqaEVIexNvlhLFPYdmEsJRjHIMeLxiHWJHDxh5mNKCTog
Mg9ADHrTz/psk3sZos+0Y+hN/bgV3bas1x1JJdjNSl8OWmAudr+zqlWl0S6CILqIxfXxnHHvbLs2
zOnXDIuMjcO6LJLf+M8fP9xpJfMOXb1sYoJQiWIVPAhEkl9TnSbmNRvGEbsJ8yPPPd+9UIymJy+C
ug3HpVupnnds9AR18LPqRK1dpZQcTZ3RUoZpdfg6BbahpYDjC7KXHZyXGVM0M5eZuddX2C4UvenQ
J8oSKdxZXEEeJx5LOed7QVP+WiuXmY6eS2ddQQAk669zErTCbOq7nzpk0b/IImGIRp/O4gAUlpvz
WPSvtKubKm1A4OR+oUk0nttKBCvbK+guZdeP71VoTAMHN5l/TqTBVHtku9IsJVLJpkimr6Cn71zc
KaTb9E5B3GVYravCgEMrG0FzW6OjPGifinNvkD08aSFtWLfkTMxO6WmhIYAHqeSku9e1wjTfBAB4
7UtpYGq3oBHRwNMrh7cSNmkE6Xz2Rg7MIVHs1WkB4JNLi4DqKE0YlBQGQ41Puh3I7/g6k1t/VpIT
Nj/woeuiN5Tp+FKGk0EVGLLYg5H5anQpWK7Vvbp+ut1qg4nMW7ZbCExEQEbTuAhhgQ6DmO6BkJ5p
pdGPTT9obvLZ2P98yv/8cs7sZsED3zxDw8OLC5KA2MgCjX6ijzl5qX1i3vrCDx3Gd4sfA7ActtIo
KeAGJV1+qyihKA3OEAax3jejcT2UP3rhQGtpy78sQ9PZMvjqQ0BBeUbusZ8cH55sherIHqLvfScD
+Hbuk2C/SU3mqW0Abe8yVus8/G3M8zwdc5UDwuNtKinDr+eglrgfS1ZtHT6JABfDp5qDbyweiDV8
AmX5fT4xuWOFycKoykABXg2sch3ZLLKzMgIUcRrcfSnzWAxDfD1LogsNZ993gzE3AM/M1Rik+bnP
hh8Ubfl+Nq0jAHR95RtrSfPNmd804LKbVP7TT72hrouSalXW6Y2yeutQ3I6ror5nIhg2HEEcEN60
7jLpYlA463y+MbCLFuu96JzSg9huR6gCkCihC2BGq/txNEeICWewhBAH/kxJFPJ2QDqRYxiueSr7
OSBBeHv6ImZ4FR1a6lAoSIQyzlTOP4CAlU8EWltLFNkWiE0svQ1JIDxB5XO56MFWkkhaLyPIWLj+
ZV21NTODA53KFJ4OUVmdexiGHqX6HBumc6riCjPfLNWtRhY6+OUE9I29y1spXh6Mj3ifsMWTWp59
NVDxAkTAup/Yj3RExQbECgKTf55OC5Oh9Xwb5ER8/8Ne2W5o3z/gjLW0cc7WXWaF8OvHm7yZktlc
6Yh5sMMsrOj66Y7WAV+btddXG22Stb8EeYZdWdYd3S8jbNmxR1j1JNN56Vxl7Wm2TRCFb+U7qxCe
PW4TgHz5MJ5kEjGKQFgyU9FqZG4ZEVB1Hn78em3+Xmtu/wWDv68QwNHxeMmK+0xZtxKG8QO6PqaI
Dc9lbaCTslRp8WYDJbJW4ve/V3Aa5J/mQpdsp1o5mAvZaGm6SFstiuIQhfPR1bs7NryFNq5tIOIu
L7MqoyBMruMaR+ZGzX0iUyEV+P72fn9tPDGk/moiN+M3bjRrAu27IkjwvQvOecNEEa2wAadWbaST
ISmgg0JJWGme5QMNKJvO+/tdYi6UN3OhphibZZNhAdgdflUb02mJP2SUlb+J4oAtdMUBhqvPR36I
4N5l+i/9JooVTQmrgeugSHsjrUCLRIRmy3opqFyiPpYP5DkHlJjF4UgkysYWr05CLFYZVVhYcJaD
Wd8zVOKF0E4MYFL4dWjt0wlD6XNJZXXCIlwp7T+okLLDGFuQjI2c21DgdL/bkeD1oUFO7PaLr8L9
88k8H2BwkBhpmcV8QVIOpx681+5WVoHlgvOBdJG7qnfpAtJeG+kAnLekMLtZhi8Zk5Hiq81ru6x2
ZoLw9R2JoGlBo6v1giWFcl2mbfheSpdvLfqhwK7Uayx7LIdiYF+lHtcsyxQIWQPyBdCPAm2JAMcK
tfv7K6dA9K6lqblkmZQaSVC08Ppw6Ou0ptueKwHbHrHB2dpuJo74+dk6MSKzxBC193g5+Fb4iBRU
aroxE3bviX7SdnOqLZPpVETf7KRSL0ZKTEbVZ6RmrLXjWntFFBfUr32xd4xOe0uzp9QN/4SUJt3r
oOENHhxRtED8hTCL8RL53N0K2E7sHnK7cPtUXV90ImBCHRHItc8BCnb0iGWqpDeU7GR8KQJG5dL6
4P911CAiBa62HdgdPSyxUH7OruIPCd9phtfZF3Sr/dOFXqigm1pIJvDG/sJhcGaYvtcozDpfPDjR
Wo3EXySequ16pfPNoKuYBqC1KQ9lQ22HJ4GUi01RLdiZuQgHlVSVwlzmV6zSQbJWOb2U7sUmzArY
cMZxYXipiZL/ifroWT7dcFWxVVA/vNREobz9E3F0q7LISLJrM+j557+LvmVCJhLEaynomnFeziTo
A2hc92gaFL97H6b4FcJbl7N+Os6RTOYVw9ABmFGTVC8EWdXuH/nXANylZg1O8u1eoWRqMk0qaeA6
Gh99zK9BZmYyVxNZZAThKYz2IErZoAIX3e1W2wJ4sBIEbAudUqZ3yCvc/k503mW0OYToPlJ9hB8H
KIR6rdFustu/ZK389TdcgdtTQpvoFFoJ9Bzr4/RnOLwgm2vNyXu0GKLvHlB80Eye+10b2MbTsmpa
yTg9QUF+C/emO6lj6Bf5Bmh0jXy/PSD1qw0Bt+btrDggZAaP8FwSB6Fwllx/xZ0E6jbOQE8P/JqJ
nE7FcbrG2VaTgQEOHIjmW1NjTpYELVzCIT7nI36M5w5qk0RGgJAXiJSrYAibDPT5OIQLyZY+tfdf
8Z1fA8o6O4QvDSa2eHIennUQNE0U5Q/LmK+71uZybjuO3yv42404Elsh54HuHcKphJpxB4ul2bJb
y3AjMC4aly/PlnZ2X+MkVwzj7uwYPCcVVAEWOc3DtSyG9ARp5eRv61R24RkHyikjoSnwJIzmUHyM
Rc839CHWpSakY+l1sNBgP+K0RSVnJNaQc8qPj+stZ5TTHndsWPzQkBLvywunldIXiBrlwkCYkVYf
HLvce6bVxR242BCAI+mYny9GCj7Ey92uUxeT5rmWCSlWZfqOg2yu8js2n1yZqYw2n5B4fka+SpG2
MgmZ5A5+ZKj55GpDi96LGQNL3V2hz4jmnGHyi1m75pLdDiaHakCUhXfmNG7S5ZU0caA4Zu5WLFZ9
VmjdUy2dKhrUsT+UeMzi93iI0poykUAWQa6hTFn37rluIGnKk1LxxDeSPUpqnsWOjnA77yB2j2Xn
6WVBiWPOcGm2lPfgv5jB3ttiwxMmyiJBWldbPx3eHhbyOpN3/8uoGBeB7nNp8PM9UynQa/NEztVU
mfS03HQ0cheyYLt1YXoxuhHbXLdf7rHXEhSKOzqqVXWi64gC1dWEF2ERj4TTjP3sLRcphI/RFmP0
E/RwiwN0hroLYuMmHTRVqbtES0ZTs+TNQFVTyCKldMLVPgoUB7ec44SfsTXkxWoHjU/AUQbbg2Xp
FoH3crEC9D7qtFExkP5sH9Eo2IFx7GzvTEzUVouRxrnOFYCGgqxIHTjHzd0kPpaQALCGF6VFeNpE
v3LOZBhhQzel8Eu2L6ZvSUaIydeb24ebOAZi01MhrF7jaVksUA0lIvII5lPDwv7zg/G3zzhmOk6V
LF+J4ffq7kFq8hK76aeu3Up8yVkyuXqYfTK4bpXBoan41t0tFklp22faXgD7L1XjU3CjM8DS1o8a
66A/HIrp+Y5YrsxZkbewqhD4Sse3DFDU6fNPVVEMT5H5HvIS1WldDuGL8JjGJ8W3uvg6CaB3Gn0E
akSvTO3zdrWx+50eFXghutqXSr4Ovq9nhG0njQYi5tkWjNqe2VM6PfjNT6N1Y7oJjDkh6b9zE27k
X9K2B7LQ5dd50fbVKkrXd3NfkGM69ka7lvu0Mh7ltyKUNQaaNbOxIQ/GRdAIfBIc8hVAf/k4lVZC
qNIbNCGC0yEoRMd0tT0wOUieDcxl2GYNey4CsQHtRqtBDjW+X6sMVVIzND73T7vi2ItwOBjcB+jt
wvsXQbT64MbSpKGc43ZlVq9eAjfGKYvF9ABrC/UmSOaeIi9NGXOFAvBvnB7tcwxfhYsb9G7KlGmq
8WVtlwd8yZzrzVSSkPFADqcBySXp0bKyEQt1lPJcyHBX+4TAlgJ7AXha+0dw3RgzpnUKYeex32J9
nZ7Up3bb0rUemx8gRM1620oao5uxClassnyYaDLJ0fK+TDaIsg7c0VEWQNKbp0RrTBLXnKC7fkNq
ZQMFKxCXtGcMLsK8D9P7e7bwaeqhWn/ZHk47uvW6Ln2APHAKfhx3GmBcxjsGigoPxF1bOv0682pK
AI862plQN0Z3Ox6INBwf7ZMEo1LwvSQALpE72yNvaax+40vaw3DFFdUXCIkHTeyxazKKcTnK/RtN
nB1XDPZyeEvPL2AClPUBPywDvas6U7o70Gt9bIPiHqfquY3HNp9NGYbC1RBu5yag/SVNvSIJS+X0
gpcJ6UzS8cg38pmriIg+zW4gBGU3/aVpu4R4aas8KItjhtBSxAb2DOUHMELiY6GbN4EBfpJycvQU
rBpWiY+kWnQwnLE0DtIG86AGkIGmQ4P2tBxlhlp5pmCZoYX5WLS5FSZAnXM0d+blbClwRX0nJVp+
dA2gDi5lj4feGmjGrlMQas6Mxo7ud6LuxMupJ9VWOwAjvLwnbzGmSzX0/K7XaQ6d1ZacWDV7o5yl
k1OqVQSJFsyuS7PA8H7qxEO8WumNC46yHosffz3aN3lORZCDhaYcgEPY0BjW/NKBL0lcPk0HsPCI
QkbRYWs/DlGsIo2xFH0gIl/6U33Fp8+daDlvj3Apq1GvE2TE7xWxv2ZC4RmZ6hDP/meUqxq/BLhx
/wD4J8RAgIdO1pJxfvllXXYJTlMeIhEmEkAD2tO86agqlZd5Q7QLfFgUG4tDqHSix5LUx+YZQiND
bkmSHH22DT9SHv3caGrn8pTqnNu/tXSlPsCmGgxjCUsvDegMC7yRgqIMwu4Fs+FlOLdGtHHwpXLT
oBB8587qqynq1FvcdOKqFCVEbCj4CRov6wTX3d57J9y+DtCiEPFSa4rm48f069RBPbqncoMx/kTq
FZivnJn1g75M0RODbp1BMQWECe6GvWqc36RLmSwdLrYUZROkqcdiz/mFqNvjxqfXXrSvdPQDyWrm
ow21044GGpQ0aSPdvlcnCywN+j/3Xv8oiwBeZdvY0HzMNM+Q+tLBgJk/cPXeK6lZ6iHgBLXi3b2j
R7IqFQBE3h8OUW8xi3laqfIMNTLc+Wb46MruG0hA2yRnjR6s6g355Aw0FnfKT6pfhin2WgBFQiXH
gGNAORiV2+YcA1uXLMIx+CSifcFY5rhYuaD8nrvRiQ9RN80w/YXxXgJGQneilT88EkPkel+Mbqh6
tmC9oU/QAa1r6IZJFjBr3swlj9ojOB6wZpWdqObrE4rH5z9Pg/HGZAnumXuxd/e38N0vszqIVPuM
guDw+bMPVPOkV/5tSPI55lSQYNOGQ6BKmV5f/6t6eIMqmwblsFFHTjZLkIiIQK6QigjT5LeLSOTx
nTXboIDpVspc40pC7bx9T7O2343KzfyIqbvixWl5wh6Q4O3NC2sC98HFy0OkUbcUFI38L8+DbnIT
cDU5sJpV15JH8Mq4zjfj+M18sw6RB5qsLz9qP9O23r25t15FEz4kVNCkuHdVkfJS1o3XZM3TpnIg
AyKxDmHENrbwvvJTkLpbs+BO+eFSX1ZesMzplk46fLkbcWIr4PpYuITAf3cCO1fy2zecqcNIhmaw
gmdyxif5sEpKokmR8Fl+bO+Yy91R3Dp0rZtUxbzt76gnABrMHqex58M7rKNqejqOdb7KYitPoc9t
qT2A6HRa0W/Jl3Z1YElj74Ek+cuyNtnek6FGofUHVpj1nTC+fw4z9B11q8Wxmm8llx9bP1ixfWGY
MflF9SbkNymrRQBp3J/JElPEx19nSmnjXJZ8YxtCj12sWAjWK7mepRWHzrhSvRZJ1filkPapp+nK
bb6UohYdkw3Hapr2dbqxwHYlaacoDeoavm/rgRoUeyu8AfGr20xVWaqHHGZXSMlcBb+oJadHM/Gu
o0K1z09S6d89ud0cNWkkuNNdQYgs4CpV5tTgBI4G/455BtCh7aU/hjWd2mRDnpZeRoB+1+ihf3Tk
asoWsCW6mBOhqfcm9OUsUMW7FhZiTHBCZ5o+nt9Qvpuo0TpIzIdX/bWD9rnDOxm/EmM9DBaQLUuE
90exab+YoAcTCjj5AM3otwiJibfkV5GW9JujSDY7X3A8vvo2U9bK29E7y0rUBvADPcU8Yi0IbAGR
G7py6pDM8atnsthJXbIi8gQ3iZlrRKa1dcMep+nBzpAi8Yb6gJq7WwOjgoeWKNviHt/VmeVuSfG+
ydq/cPeH8DGkIhOOzUZTKLYGWgadiPctgLsWn0ii70CMqQrjjpNhm2rree/H9iIV8uWAi6I6NhMP
3mgoS5APiZA8G1ViMiN2DqcP/vXaGH9+LbYRs+DZGBytOwyhocGQhhd1NFrc+tOVHzyJ56s7gXx9
XQIBY4mXspChV4TxQY7Er+b54SX/HiQfDKSaRh2zlR8v4OxVNJZMh7HjSC3Me35gs4oD+FZl6MNX
DfZD+ILo+F/txDK0lQ/W3QtKAAj6td8ICPV5EJbe9M24LW/6IIdU9xyTlvd2AqOM70gnO6J/pX4D
vzs0kOmL3GB/ACYyD/quNzvEeA785CgHzUvlSkM8pYww2ELeiNzaCgQ6NyqgP2OMBTe/3HjwfiGl
eGYExWc17XZ2ge8QYwKzAN4OWCs0VGnJ/3QyLGBT6k/hVuFZsUoHKeENaIGY9j0RSwAddCYO3wdq
VDGprhl1RX4Bvpjuh30yBWmQhSKR94sCcbnThikj5OczEFysGCCz9GCOI+cnyLCNoM5otbFb+kma
vHA8NiI2GEtB2bEqfiPaw1/lz0dbNbv1gbU19EMTQvPjFqOTilZoAPWIKvctTgzPew9BZDlAwdqM
Zv2iYbLq9ImM6z8x0HfZcUganbp7C0vLvhQG3YMRFF0VUX4Xc0HOAtaPZM5YtFg035Bv9DgAL02c
LV7fOeqJjtCfgIWJHTLksce3uhj2zSS02EtamQKkFH5bcYZ+61EfvkpUW2HiB/MsPY77wiE4AdXL
XxOvCRbjglzvZNbJXGHmoruZJ3NbHSyoTt10PGSEuz0ApNmTcZ/bDyRyMRL9woDsadtIJxMJfqd0
SQFROryOViNRjb/ehKbpM2+8Lo9shFDZ+IPqqUbUHsMPkwdS8AbsONcgt24mZ4bqSwyT8CC9nhBg
YBlBdGiW0UUET+GZvDbxX+JQR+TJQts3SyvrF/j98Ylrv48AxbCRaKHSE8XWteeehABvwfzRD5Aq
tQ7yg3a9Q5+b0TZWNRLnObVjOVlh6GvF6qej84QQH15Hln6aFb47pW+TAsENrSx4hAok3kybCIvn
LiNfwM/0A8BBjXzLzVfRzab9aaKDOBkTURAHPTE+FLcWLa1zsIr1nf5xGSg+mJ8Q/bRYIZkCvzCT
ZLEfJmOmIOWQ0wYxhbsDhUpnyhC2MGe/1XgnY2Gd7yaY6YtJyYr/zn0tsyIzHLNaLY2pJZcPHRuS
neQ0QhYoAqU8xD6k5/zEJyhpHAIZfcFV+NR2cyS3FKKG6oPUuDUkbT8UpxY83cVnm9+v+a9hwvoD
Bk1E4P0BJ4qs/Ao2Za1GTITEhaeKqHdBOheQVqZ5LSwu69n8vIlSF6KcwZCyCy8S4iYGg0+NtHJA
MapV+VoTHtGz8v7gkjLfLhpb3IlSxswRoiWEaI+QkQMBg8J/upLakIPuHr6bzLdHnnzS9Ko4X6vR
mnmZWCeCtqa/mM0xjIsG9qR+d1q6D9MK1F2BEqwmTupAMzTuSytMmCs2E6YzkXfr/rGoVGgR6HUU
3VdgAOvt2iPfSI+SH9JJLElIpGf9L79g3DnOyHvi1daWTzQMRniboPUHYJ3/MDWHbCbBG9vdychV
/8MLewPNdVmy0xExfDoveNflT6gTMCEBF7lRhBA0vyoRJQrXQO+yGzYs04YPSAf/VQMcxIaVo31A
dT8Mj1SMu/T2XMoN4zTtsBGmXdYoCPjx+BIXQ+ZwiQOSHwXheaP865NZSXHk5PcgrFONODyvQTAI
n1zZFICq2O0AvpFXmhOZxZUNyumejSFwerrWBn0UCYau7mneA6QjciC3uu1uac34m5XS/rqKVrh9
gU9AqHDouew7qC9qYn4oswf4S6eGG3SKY+9MVs0req+TIxbMg5oh9WsgHhLPsg3FDf2VZPOrv/Jr
LxApNYDo9Rlc19E4KMDjPHal9faRuS+ymWz2A0oKuwkCP2GoPeqpGNpg89jyNjH2Ps4OjgcfWeQP
gDRo+1pf6H+M07yrAP/HLa3syJQgvoMNYSWBKKdRsXgNhXLj3O7VDRQIefQe/4d/Qpwrq/sh0kM7
QDB+2xbG8VVGJA6ld/fInHObMAFUdgrGPa/0StE7z9CLhoUHHdt0WrRJkGNn4NRIEMDAxK51cFSl
aUlWiCO2ItUGTcbGIvyV2dV/FSUNsQqYY46bVEo7ThmD2IOjz4l+IRU7D/hpqziVzfRkXJ708yN4
Cn+8f+qiNVQkHmJLUKymQOxSJave2rRpN+rFKRAL5YFjmmFt8Cb2oQmxw8TKHmnmOWKT+ef5Hkl2
B2CKf3VZpzF54W5AEUSHdNRsJKhFFQFZnmxArOaY69/PNGIZcfnQ0bHykyW9Oh2Xy4SVEt7C00SV
d2ifmZwcfPa5nx2/9pCAJZ4fHUDpaPg8pG/DJrVz7FGJNm/xrMVuROSsRtNMk6JUdtTXbqUG52M1
ZKtX6rgss9qoZXx2wqZVGtIJaOIKiaGZljeHk9Mycg7AB27JvQLAmQRVVz9yfblTRMigh2x2wpjx
Te4Kag3gpFIPTnGqUJDnSAT3xo9ex/01xiQrCLnrzSF7Jl0KbRLyQmtC7Mjq9tbP+bMF8Wn4FJ/h
LXmOmKR+mm/KHb/hk/UW8bbLSY7FgiAytqFc57OSurmAjp5t8ZVAzoAFXgLIZka7Z0dfrKp6mz9X
h3bMxv4wzEzG/p9CL6YqTMYC9lpd6YpGmBsBQqHKFZDlCEnevRsbIZ9/i6RrARJY3bHpkDQHB8jz
iix1qz0hq3ofY5JUQBLnLsiHNfurMt1DgIS4VNssfWmbZ4yyITNdEKnqnmWlcGHQ/zK7KtQmRJy4
PMXxQx716RG/UdmvXLTrmMPttyqENt9F+NX3bW2fXkCmzJ5n6GnU3sV7LVxOwf+EAPZ1Fwxv2mjo
YVAy3bxOi29+2S9i6eXB2o+nFEc2xPcZZtw3+LwrfJ6STE9n6sej+09TI/bSdqCvEdMSPE4KEYNB
je+bmlQcGvG8nAZHtSKpldWoZ3b+Y/ql2eFZ5jhktclMp3eXn1YoI33jqJe0uA3QSnxwbBRkJJn3
I49TYvUi3UvhCc6squ63Mf9mWK6QryEoXXnJbrmXsQ9tirHhzZRZclYR/e55k8yw0Xgcg7SqBRjY
dDkxaqiKTo9irMLdERWxirs7GP0rhjbb2Phl23mRHROtv4xrceEG+4CWlPLg3CmgjKOFSyFZ11mr
atakorzkaJsLATsRHDiNGZKDb8aDqySKztmlG+r2QnS0hxvV7s6Vtiu1dPGBuJoHUFq4VukmdpmQ
2iP0NNomijifVr1Sh2nFMEOeP0f1O07s+e7rE+89ckImvOxD4tK2QB/CZc4ZQsExcsU8AAu7ltOT
AYrsR56Cf+fwjTCAr/eQPwFX/MoN+zsJ5XMpzGH3agCSQMUW9ZEyptWJRUjYCF0XZna9KLvSrhnV
Gv/6yJ4t3MyoFpnU+abDpXdZ0s8D/54kD6iye7xvIK81je15vbVj3SdPZCwxjCMkvPgio8k2HyBr
tyHTlSIjIoagD3qoK4nSSks2wn5jw+ZBVhkpdw296uLRU8ry83lTIiBwuDZfsCZ8dDDAjwR73gdU
UxiHszZvii9NTpDQxOwbbZeHwWSDi3RRDHqenWWSrxifSEkKZWPfjN+o3YAA0GDel+3koL0qNZHx
zuBLPUnTUQ942GlyfUz9NwxTI4hS0kesczG1/0WFFHIIU4Udlb2G9f+4jkgyORjELCK8EO9oOW9O
0YBHgL4eqztUVy+sx3K9/prsJb2V5/vvkQaPIhaGZ8FOveuASvnla2df7qL3NNV+REMLjvkrSn6n
fv3c4XOdJo+6yMT+6cvJde2HWu1y+nWyjSPi5lwm6xAi2S/rgKLK3TTVkUQxjbdFwoR/veow5583
O8RzzOwh7Vc52j4JSf7qotPc+X58mrKdc6sHEOV4TTvYU3FQaBBRr7rx9Lax+pOgoY1AvSB4rjWb
M4SqVidmV8ErV97KcTWOFPinidUPp3wVhupUMarfjJLeKEjNytGfMKg0FF2iCgNVzQibBoGDjCqU
YN0wiYZIXOqOzIwCZ90hqRRHxndVtP9QD4khhPUvxXY+g+PeFswVxIaHOGB0Rb0qu4vcgff2m0E9
0mDNIruc1XZiNxOJzpWNhbiLXZSpl37j7YSDDYP/ab75JyyD5bjtbjLzCteceLDSOf1iigT5tiBZ
4EXIWEf13o4kmNk/dtESjkGxXmS/4WC5gk51G4Rod5/DjDn9m0yM0lkgB6yNn8RRpMf+YRyv2Fj7
spJWDc/BqGFL/WYVAEBDTkn8dMt0geIvD4ls/j8FttnGaGN/Oy7lgrjh+d3aa2mshTc6Z4/2tGlt
H4viKQPU7Xbqls+qZvr51Vrbyc+sgWaTneomQPXdNR1acrbSgqn1UUz7Di17btPsdzSsvTSZc1Qa
TiOLWKP8N00LunolrlTGGCNzuyQqLZPQbIdC85XKBtuZfAwaKt7oS32ncaPn6sOlQdFJpBPpVHSs
LYwxd6F7IEm/O5M1px8iOLMCuXqdpAJ4qQ4k/sD06SaMWlPfAkayNcArxkR12dWHzY261F0D5pbT
I3MlhyEVJa+8kjMoQsgRLxOqtIU/84On/IaWkirpER5g1tpfOex2Lt27UL6gXigRD0e6vqlx3HwG
nuLE+9XtziJSU2OcZb6KWRQ4aaLNfu6l/B412n1ZrGgkT16N+aoU84sGsqt6lNLDjJtlaMKh1XtE
QMpG4pk47xtLvZ98Ooms8AfJNkJqwnm0JbxljPFePrHw7yg6Z0Gz+defOyWJXl4eGPwnaSwlu2o/
lJtovXCMS5//fxB2sCo/7b/MoSPyrB5blyz9yo8eVySDQhqfJ4lacfjIsH9gcIIFJrcm+2l+JwjC
8240X0Ic9NTfgXpgQZ4rdt4JZ4rUkN9FtHxQf2IMetsHNExpaMo7BjTu1MW9Vhayfrte85xMeeBZ
/lT3AjymVTB5diI22TFOTKJysj1jFiSCK4+2MPjBCUEby1BbyHs2tNeZRcAjfhDsCdrSsNXSAA46
z/87gr68uHosrJa8OYG2h8RRRu7oD8obe7fUNCkXlJ0S6xCzXgh/P84RJ5e8b77ijM40zdFfYc85
Jg/1DMc0sSbGtYv02JUoYyqY1Ni8TsqgEiZcOxT0V1c8Zds0rEMDIqv5H+2ernj57bZ62LOUxScp
zWi20O6ReIY7UAFj0X+EIKuQO7xqJ+hXiIiq23ZCP/xP0+yCLE4yxgqoi/6WNHLInNSJrDaOXjbr
Uat+ZYIB/TN/lSC727rRg6dvnx+9V6y9AcBF5fL8HVZ538iCQcfBuL0i1jiFO5YwFyhjm3hNjAL9
QQ5EMO5kRCFd28DZZQMXn9g082PZvf8lvHUF7GTRm7A9941wF9n5DHRUAMK+d4JFCZKY2Jq/wN7e
Yf1bFovdMvtT21EdWIrCvLU14E0xiYYwvLLqD5vKDnuMhkwbFUpb6Nw6JmPUDbofGBtU/EtWQPUc
jKSBBSQy1HfIqT6DiXmPW1OSdwUE1bPTl273up6pW+v1O4KPGvPxW6FB5aNUqAOLnhdvQRCxDNLX
xSR/piz/fo2yI21E9RoyUiQ9VAOeP9EDUwTd3pSk+l04nZG83z2WShvCPHMSpHAa2yqxL7LHSCUZ
dfm9OWcBtyJ2xM/6wtBI8OBSn+S1R9o8uHkuwdYGfNKz3BUEVnIbgoLNXM6JfLhOzpO4UoMQXs7n
hGPfxn02AWmRr4zp8zNJlg4fONMICse7m+WUldLUSZ/ZCRqFodaE1Q0XGJMV1iup5M3VWCWe9Lar
AgCX0kxytjibKaokThtPWRxomczWykhX9zrfrxwCgDnSFybh2BerFzRmo9bYGKJFKq4Ky6NtWoDF
xVmP8MaOPPXH27JKILv+Ar+MCX13CGjgm42nCIZR+85Kd5Zgvv1DtmArdEiGCDOcfugAPEvZgxIB
MjWDY4JbosJUmiW4SwtwC8D/apnPpVyVXVk6TiAKhM1HYTBf5UiBquO+JXkbR7CxgDeRmYI3gy+h
MDX5V2fg7IqwdObsTmTsygx3cTsGcBOK1WYdITdgw8jL5Ja44YCL2W1r8eLIsWLidvJsWW5PzSy9
IoNePZNI02JOQ2gBwMQQ8glQjxmyTIGmAgu8mFg+X9IzxjsuXqdXAiqcQkKtQTbIA34X9QzEOdvr
uqL7IJ2y4AcCXMkY5Vva0xC++cnUslaggSk2baRO8cHHBEwtlKxrIDlY9CSbaQUjhgyDRTtNrwX0
tj9yJopIPwO9jKBjq1036JMR8Fa7dE4yI6Mzc56PMsZsqxuHvQMbYrzAA41xW5F9QQMkeojQC0ZA
UHLnKcKkj8rkCGIu2ysL1K90QZNZrpzUfyMbCMQFSt6dzUkT/pXSEOieDxLg9TFXJyxsHF+5UCrI
VZ3HcX9upf4l7hL+qtBFmEdbDKWGhxjotu7fT69Kp0UKZglDu30TH/rRAxy9pjc928kMDv1ygw8m
1SecUKwJIH+ufuKNOovroRIxM4gu0/dXeYJKHjDEUDUpOCrtiqx+fSKmweXVA/XXxa2ZoWUAtJ+2
HwsFup6rSnIX2K0pk4OKoaJxQFtqZDyZzh9cpO9PV8/DI0kAlEz/DpfYs2WubZYyEacpSl0rJWws
RN0PGj2lsOGc3BEhz94lqBwLFO3ONPqgq3cBwhMKRL/QDh/mm58BgRcMv/v8hXP0NuDwwD5BuzG+
YOS5l3VgKjL0jx0vwxoKrxA0uvPI31FX8MlSTjDsmLsKlzp0qfsJN5gnH62WIRR1WS7lMI1a+5Ga
QGHFYzcTCQ5T1B+CMAgOXpGZ/opgwJj3bE5SnW5Qjb6qhYiAEGhow+9sbAoGdMk8AuapxKW7Wq2l
jJGMlErO2HsEz9i5PIR+P/R241yojFdusCYaVdx/xWcT4mCm/Ez211vQCK1bPCqECEy2CJ8/1hg2
m6Y9OLhB02G2oRm/d2gOU4yjhrR0sdEleGsw8zwHvvqgPbO9X+q5VfkU/wFt5HSo6LesS78HT/d9
mYSW6Bg7dtwxURA76C5cRUMly3TmlbgUqSx+uO9LQMPOsG7WQbFI5XAeGiPHbutJr9boCHb8lbCk
2WFIELQwZw7lwOURt5seuR35P023W4lNqblTVWz2tWDWSes1qS3+pEE2KNTUjJ/wcS9zzuRQgfKn
13QxcWiFGv8IV6TcCT/rPM0nt7niEh7HpOxSgOw35DgSkF0PW5lQh/OXa3K7PRmRZjhg2zZwK/MT
Bf162x/9fNL79g8AS0wDGdbzRHWg4ECeA2ifEoxzKWzARRzArWJJ/YD3Zf///e8i5bpossGasjPq
9axZP8xsnTVELrdGSH9eBrU/hzW6qZUZcamH8AzSOwy/dqS/IwX3xsPv1ve50OiUl/mGWnSJySjq
OruiDtTSKV1/orEiw7JhgtDSUsBVKA1KOVoCngD3O6hJHUUErJqDlV0eXhz7BazqS9CkNzBGp/q7
SOdlL6V8zMrcKfeif+xHcXEJH+R/qJmH94v316iuXm9Sd+eVwRBfLUDID14LTVXaMPnX9TJzjjPb
Tgvgz3eZjwolc/VleIvveMxXmIFKEiwJh5J4QvooWTAuDGO9LZt1jlvLwn91NA3bqWlu5+EMWsg9
XY15MsPK6vU4p+yOi05v0ERDsANbmT0MHptyLR8jwTWOQfnnWYdIQP+e6MActKp2cTnidYkGSD+S
QoFrBIt7Vpx2vkfY+uK9NniqIYhueoE7mfn1V8jODdgJU7qnfKOTVoSYvnRssz3XH9oUlEt8Ud3A
s1UzCETCe/mqCxkNrjNFor//mICmeZCtMtqvH9MsLQlxeoTHYQLsMO0CtLdZzqAvtevbM7TM3DVh
z03kAHIrqkbEMWx2/4lzBn1R0wvDFPDJKs6+tEg7FN2YuBXewv6Fypl2d9kbKrImwBlYChZdTIuw
3Syr+oUL5v8edBRqq91qTalaXdjflEeOuQ+7IejH/HU1WuVLEL+Lqkdp16AGvcee04pBJRwv+WND
Lyc33UIzPDyrflleKIKD1yOfX8fvgGMQOd5vsAmivf56RgzGy6usqoEuYENsI7Hdmze55LfSHFYn
IZbrtNl+e6QkKBOIjgxrej8sgMumSrqRR/Quibji4ShbWxIQw+adCVdMfU1Z8+aZFbRrnrFZ8JY0
TVnUY+NHxFNM40yV2AL52En1CJ7VsIFhlh+kUTq6B5Xpt6iJEMe6obCvwYeATvW9vMcHWkhqf0cs
34LyYmeGoKZqrscyVPq6ylBpLrjnLBKCYokNXFLNV5AX47SZPFCCYyI+4+WEebkAfGAEwHSovLhw
S3VWjX/J/kw78FR4z0fVjYpxnzlBr45E1Y/ZD5x+UxZtU/Gymn16cUcQGByRHRoyXboeDnAg7zwg
Z1OJrJVdGPjbMrwhhXZY/xqD7w1uAiLeGfG8LaNhhdhNU8cEFeqQxzTfvv+IYRPaevEty9jbgssc
deyOk1OeazzuhmkO42YmUxRu8KEkrWBDdOYhxWQsg2Tb0FYFhnKrgt6MBeS3T9UwQtiXpV21Qtk0
ZKg4EqgsBAnPXKt/RNSi/1fNhhvg1rBjgL3PN9KUU5XE9e9MGXX2UNupizo5zf/SC19ZC2z475qc
YhGxGB62vSjn+U3ds0YHSDe/AuTaKzYncDNSBkQQ+eciMGaJa+HeTKiKC7C4GVVgAchgw9Y+blJ1
czTkHXvVlEttRgNpxDYe5LDy+W48nHouT+FxcV7/UlDHQ18DkWpU1wR4ONjPDd5qkP5GfGwYwh6e
ry3UgP89MTrLRYvctJDhI/wJm5BHEISvwiXRNLhr9xy5cEF69qgd6e7EHilbLECNXQiAEiJe4fAQ
UssqHdhYUiA/tBLXt5KcwqzLh1MGXsPeaE7FTZUDY9VNVMDBuaF37AMGEEUPmVITAp9Sz3GdxdIq
Ygym4oHcmrdxNm7A7Hsz5ngkNLRgUmQxu8XDfBlefpA8NhFwfjTDa2RQt13QvjDXAtgiSW+kjCJd
DDQyLADe8vdcfoA685J0WIE9RAW9TbLQLdDvV5g2VxktdAtt+Z8T9bTEyUt1bn5wOibSMbzbyPcs
WFmKt+CaGOcfc7mzNu4XmXcC0kxECHtK5LrBZEK8zTklySATMlK/NyMWguqCqWCpxYux4R7NE+xj
S6B0E5Lj4NEF6QmBY7N/PFuMPJqmUlobubDVa6jVmXtsVWwOJqLQY7V1CzxJ+i9qpujpcsKTOTs6
PtmyHCZ013mDyjLD3lyNaIidRYtifIvu93sOHLJAqdULBzf9o9E5RZGBR5uG5Uyz/3cdN1hZE+GK
V3Aa8mn0XYCOpn9ZhpNdNn6vOVNavD7dBIcl3zyDEMlkwEaqgnlzPLiBPeqTXGd4IwUjoUouDB4A
k9LCooBmBGpZz4qN8v98yfV4U+HN7JwK5Am8CLYzmw1nMTZuOMZy6XKSlgoMitaYP7IUaQvLwxC1
uePHXFUH4WJKiUr+6wzkeGQfvuboWXf6eMsIVQT0Y6SsRbC7qT0HSlrdtqRZXiFV8jvVhxcyZ8D/
jIHQYD4zLeiBAO3QLLjPrRbb9KOsAetx7q8W44JiR/0VuZi8DeWNxdhQ+x3MMpbJvrZJFDFycUGa
l38RWnbC/ndSvNlXyLu4BRunD+6AbN0K0tbQ3RidA1Uvl9mQn+y9P6u/MLu+oAVsENisvJn8M0O4
kI/z38z0K0ojt9XN4SF/haHk5RusazxVIxsJCu+AgKOJfmyHISaUAo61ZOZXgURaaAJ8fxSTtM30
WNKtuPHSMSAeeAy9BeDAcwVQeGRdunTtV5woqHgqZo+pKZK+JGBQRxYv9BSg6J5QY9RZXJT7nJcr
sPpleUMDiZrz6g6JTSY8t83yMdyixgP+YLLWFaPTkcpIxNXq9bTOl5gyNK/Kvge7nUyZKjlc7w9c
QTKOgaHtp6Db3eRBZvP4sMr9vXQTMIv8mTIIfuH8GU0IFNlmKiHxSdZ2eR2PB7T7EPxABvJRinJ/
RAi0Wv/kBSlXCK7a/cVrFA9B/qEKjH3UjkYNEjJVNcvneDTnmXBMuuLHsjhFtysL6RzSFdftWq46
VmUAo5bqb7Vdvs5+6DFlkqYkks2yUdyrTgT0Z9BE2aAJwuxcc0f4BtvWzjZ+3zlCpVOa3wb5/5qm
eF4C9rS5Z6/7J04feKcv9WYi/fRO5EUzrwySOMxoRxo2CrydB8nADuTEJLG/aS0klGRCfeNBEOCY
NAMG0TNGwe2qOSVtFU8oisdDV0+4Znd6ywCYY/7OOOVXnAAAmD5OKvHZH7iOGOb/bZlEkpQ924Po
jrUTUbUt1n1aD/tqFGg1tHzl/eH8l0r8phbcRC2rAZRDGLxXVEXHLdNllGIGTgrf12GClbxRFjOl
ZI20D3/i6Wc5OfRBD9AsyfIYy6XxD04IBA5TZUQIvpEhz+pcu2X4qPPBAegOv/6NKWeyZgynwgJB
xMBq66GhE2Fp0Q3BV/87xpvuN6sPJjAIHI3Vjqff0XFDWBlXji7RRxUGZ0w5qQqb67RugmpTFAF1
wlnT9bqBKMkIxtkMq0tK5Hew0/nRLXdFbsxeebhnkx3EJ9uVjFBwaCtfDyUenqs4ZMndsaZLhEFg
VGR22/K3JL0iSnS2lXfNMOXne//iFcc5ELGCFZThw1qW9G+WcyygLtAI/2bYcuE8YJz9mWnxDtdi
pLy8pblSPYKANtstet6fPKYurh7Zd2qDl510IkArtfjdR7f5i45VH8qi483bCciYWiJd6S39sRfx
40XEi50kcmnbWkXXGsRoWJdM3JaFSk7jFUXVUu9oRv0NDhsDSSOKUyrxaJlKXscSOUGMBTXArAzW
SOdZg0gkwDyLR9ocgCdv5qXk+Lqfe8DMghgN9Y2fe6+F1OuzKiqsjnrfYOQIBJ2CzlerGvTonnKH
ImpH7+364APodYKTwU8SuT8KBlYStkz5SaDiMXGo34vfQCvhfQKe+IwfvSc5Sfb+h5mnSNc3OX0A
fNauWiKXR6n9L0LOXbKuyznsy13f48uiblD+G4T6QgoxebGu/pRpMZJTG4TYAFHfsuwqWZ5M2oZC
ud7VmhM+nxK/JRTwakiQracBDoI+Suu8qQDej2hceuf6au3MwpyDN3Y6Tumxyv23GJD3lOZ0jidw
leKxtkj0S3z1At3WeBlAyHapzFxW8km9xZmwG00MQubZpihCBYvG7UZyIyLGd4A+e/Vy0wL6LVvl
c3KtXQzIGzxW7lL8s8rXuDgiVsgIPArc7Amk4e/0sKrikMw2e9oD/+nzzeZ10sto7wWQfBSL4Mhg
oPHjUG9lbFQVfa/CeJJhLlGaDNuUFe9L/RMPZSgNog9avSrzGUWrdGGTk7C6TBUbG3A6uwbdxtKv
NkVbzsKusg+8DuNXUJN/ITqNzDVH5NI78e/IGOp6htrEQlHMl9kO85CBHC6i3gn4SDNHdderIu8d
1CMagwgEUvdpcUwNqlZ2qsqAVeOnRL16cci/qIvt0JxPP9Eu0qZc4Vtc0dAYRvDu7h4XQaf1ydRk
I7TkSskQaK+WqSyqwgdBcq+gfIkQBPITkABF3fUbtfbpAtq1/YCfhOxc2TRIJ07Ewn7npCN+wRtn
9a3qjN4ljVTLz9X50rO1QMQYlbyrzZIYOQZXk+jH4Pm1/9CQxbAmLY2WSPngA7XSWgWBhpZ/kmgE
RzITVX0MXy4mjzkS2MxzFi3+xdgq5fdBhmBfi3KRO5LY3MrsC0Bu78jO2vJFYsZrDtRSPz0+td5R
thDMqMXUmvR91VClNGbCovCiBuTZfLjbKFXpWNSwCeSKVW+UwH4+s2lSwvxoBDk4BARjULKK+4wa
+NcPMKpD3pzwLETwg0naTjkC6nlO9U2bpJmguAMEfW3XkAHhV13hhpnIUmjPA+qNDSsEz0cVhEIC
h1DwhV51Gdp/7AV9huYUVJMVCE1C7RVK2q6aunTwwpEKJ79OFB3Llii2Yws/pmL+Pt3OdRMIFA5/
fBHSSVZv/jdUDOYEX/GccrPts7Yg0w7zkCSvE3Aq1T5ZxeC230LFQtObxJqozJaR5TswQDdiKr2Z
8RDOdCiwDwXYg3vXq2N14Gf2xxZJSEvf2/fdVYEVIaFU12Cpa+Ojp0CUM6VBdaDLCyxKotqB+enK
KHxhb8KEE8Io2sAZc6g/1MD1fkCjy7sLOHx3qzG5a8UoJhkV1cFVApsJa/pMFSsfwRCQiGyYQD27
jEc8BRQ1jsoUnyLfHLig4BBFpXf9wm+POJJy2giKimMCEu8TaC+65bLi7IoeXyJRBufLooSynUxf
SKLbRZHNgIffqKV2eTinC6QMT74lynqvfVmVW/TM6sAX54Lfrd3BZQVw3gl5aleOYcTsEuZ/IXPd
Rx+R6wGclZB9AqFIW2ZuDczbaw7AUMRwwDqL7/K8nTaYf51xrEJCDDkCVa5Pco0K2jIz4+3VY6yb
G+SdNWQh3rxtMoXXV1ZswTbtfV+pfzpMVDx5bSZTUCNxZuHW4zdA6fbuInnfmHBbLLdkcBmznFoL
NefWPwixkg1ACcCFlV6OKdo3HH87GLxb6y8IdcUcTkyNL+Hi2z9/lcfAl0UHv384Gk4CMM1iB2wN
MPCsk6CCnlTKx0c8wH9eeXL2QN+ZZ40y0sAQyOwTsHUrxSdJ+xvnEihvCg1bZLAuFfibelUHTzBe
03g2NZuL4q1cEyHUT+XFEjm7OlX8qomyrA5QScP5Ca6vrQhj6Xn/3Oe/iT9t+vi26RTtZ0eqj8a1
JWxcu6AENI5noYjS5mAPWQZOrcTGtUS68+zVGW3vJuJhWX2IGXXC1lFjDC3iLAYtTQ5Tji4P3UlR
4O25kDtyXNf+vWYTVj7KztEIETRyY0SMeD+4KJNh5Fw3l/rhR0ficNu8/ulX6kHFq3Y1q3FV+Kdr
8vYEfkKP9ZdH9U1sRpfpMCWwEX7jcOWQNypGGsCgLIVRG74emN0QsJKLMtYPM64m5XxJ2tcRQiXM
o7H5G/jBysFq+1zy/+x2fOs/9hphk0jI7f/AzGQvFlEG1ByUQQvxJYs9HUhmidjm+Ue67sJQs16O
SXe12m8b8gYEhyeusyBcO7HW3m/feqs6lZ+h/UcZDxAolMr6+X5SkLepTeAWMHO4zqqNgN6RPL27
C/0XNW5NTp04H7y+qr14T/oE1x/pMUd6j4pVpU6dGLHigDN8mMwFv6sZ576jD8RxE02G/XlrOsBo
BKMK5T2utG3Vy8gDAKxV24IAtLo+ax4foCIKkQVPytpi0wnacJXygZhLJNLs612fdG7wydFrEdU8
EYHvVuWTdeeq/FzbqdleSRct4Rpq8RE0McwMzdztOS7ybP37vUzwT2ptOu85PMDZdwM+Z3pX/ijF
u4N55HRURC65qHGlq3biBgaOoG9iO2czovaAMAhJzdlDsah3vYp70VKvaieGPOIwn1AcjcSl+R10
kxN2OGhyWnHdUPENbMk8VlHvxs9SDh8oZbQoBzpI3wtq501VtQSjw/cfWqyfTOuFhppQd0oRCs2b
lEo1gmXf3HvNArxtthWTqXdlyvldcUSHZGwEcWO0xQMjdJHQfXodUvOJTBRv+MuhsSGfYnqWkniP
Ml6Ej+frMvd9rhtQOuHxvowMloSudFil9YS7rMxTu93WJLTkgF3+CbLUnlfjkL2HRjFCuBQxWrV5
ZxMQOM7G/A9IiIUnz+H6KxDUt43gpGUgDqbirQ3zhlj0RpM0ue1/RCuIo0t+p/Gn6f4pO2uj10+z
dulY7EmLQgZ5EK7FiCQTVqrOBkqUIV6mvI4txWS3zaBSoksYhwYFes64wkdAWymvYb6k/4BERjrk
ojo7vg43KZQmHYK46bFmwvd4yKsqtPlzhCmBX2ps4sq0tjdinDXE77oXsXBJK04Veqs1Z3bm9yK6
ATs7a8qPXtorRoES/eD5guJIaXVh/YBgbYEd05K+EkEXu551oVNS4TUiToep6pKfdevRwUv8BiV2
HE301ST/LU9jACfzhuI3ER2MPj74mZGTXv6xCrXKxf3SZ0qsDClzv8keC6TFNP2HTUSHhFvS4uWr
Zfk4n3OEeIhVrbuT2RHdyH9pLhsCuxsssOb0FUIcI2XFI0RsXA/HPOtkWz47WK9Lm/MLurSuJVgE
2ex9nnxyrV30ELLNoJQaP1aSXUtBgQ0xlRyxvoBPMyJWC8MNpsjabszS8ZtIzvEgP/fbFcns/j0M
44OhJOAq7CByVMLA7+r5feRb0ydRFXrVJUqMYuXFrqHk+m8f5SKTsvfzjhnso9quVNGMNBnp5BFa
ZqrebEDf1iJG8Y9DMn+dP+6AnApUy3+rVOkBQa4Cl+KkLOkF4iVTBeHRFWrKOIf1pE5PcUKTgJQO
KduleeMqtHV40HkTbWn/nXuMevM2/7vC8o0nd8YfT6NJynNMHAxDr1ZWmda7TyE4YuR2g9JQ7lv8
vlX31uwwoOaYQujIjYgxxWjRNEk1G19jJlV5/JSzK3Gvgmo2PbhNe5/EB4wQ+zjDyonlZ4YrnmUV
MxoDDpKZDCqvS82kWKtDHjxgR2l6kWNhzU/17+9zOiIr6XKLthQJ73Jt343FAxEh6LF12oKE6xrL
Rwb+tof4MJ0TD/M13B9dabFLRHychH1EfxVtPhpPka74AXAaIm5XjL0+WP/4Gfz/EahdQl5b4Uyf
L7OZudgcg7XCDHslaTfR6dx7WvQxosga3JBJM2gdyx+KK37VzA0wDrYShVrQDrs9KHNJHRAhwo4I
aRlCjMvlkMlmSwKIXU8Uo4h/W0KbKV+GyvZGsnur/aB6gKEW5CrwumEL8i/By5vk5P/6vKkXoP8P
cRqR0iUybP/hHoLVVORlvRitzcsfCtk356q7DKVKfsmovP7sKvi8wS/vc6h6Ws3+lIZQWSN4A/yA
RW3u+HSD8qQpyWMivN0IGV4G8sqghMa8gcEtbw9zRI0C0U0x6SPz1pfrQj4s0jBPLJ7TxGUOWp5i
ukFFEQSt1te3t3i/w0Tdr2O7bovrI6wbKdFhP1zLBsZ2DAaoUdlIkAWZz50rhnrskH+XeziK2iIa
VexnS/HMK6LNOvHqZNH+Cx74Z8Nz23i2Sd/nQrjNO+fMbbrNUpOYGlLQ1/RUtQ/9rXY4DF0si6Re
hVzwHaVsaedytl3PHMZq1Zj4bn0feQsth8CakJRL+bg+5CyayApPin6qg6F6OIxTmGbAF52dAD6O
orFa7gVK3aLLNi74swV6vsZGoJ27Hna1hlROmGH0k1Fv3GkYaE5xysuV30fwfcK26lYfIzrpUR7o
49DcF9ddkDVY0kNYYkW6pZ8yKdkQfy4uQK0aMXyCVCOr5XIUAM2DGoZgJ1MW9yYP6/cREOy8X6HU
rvlSwLD2HJC3hC97qMqdtFNzgSCqV+nGvwvhTt8xkmhjjNWEL8Bzdfn32wG+YZz9tRlN0T9pBESo
wrkPkNkiCXcUwIn6i6cOu0xXvLDAloufzu63+lhGCJFcAz56nvNaL8WBUZoHGtJp+VTivNtm+YNl
fjJEwVxrN6o9AuSrxyUVZh6hqwIf95/71IgS0R2GSHuI1AQIVZ/M+i6hno1qfgn5oz2qfk4Rucdh
Ars0wAYaA3CniEzHXeXIjA2bybWicNvk1kDY4V6g6Txhc76PtCizUzRusqVE6D4iXCryHG8OnfNh
tfTgNH8lkTZRgXNNTjbT7Enh/Nno130kQmSPYRSyKwlsiyoRe7p6qLwtag++3ovOaeimbQ5c12YK
l7wXBN9fjlntral6LNLH5IVEQZcSqFgh74hMilk0+8lHg9Aa39r3LEq6mLLb7LXpwizf5FA9Y41/
HCm4CFBtZP+VIAtf1iXu2ARM3AGpVVi5fn5J1F1l6xB5wyJeYXBamtBu7iIpxNUqVB3isWrrMvYl
hf6ARd6aqpJNAUaDMJlEhAKAbx22JxZykBujAmREjUB7NUXtlBnOm5T6sl7mA8/ytpVafTFfYf/c
kxaNdbIfbwXu9s1FjR1O4PgrQ8JLYhCJDmR8iPJthTowookZET3c26+i2jVhXpcPahmvMBiXnR8G
zg37nK/xy0TXzqlUA3osXEwYV7+5b87IpmM+nugOAZqqYlq7IT2zRaBAEslFBbPYJE9DTORhp72s
NDQ2QTM403zlreZyFXjmQv3GFi3YKsC+9nXgfLeZrXEeMNG6l3BEij+V0wqX/0RqBLGyJO1hH6Tz
fwBCgSfu1d4C2Xi2C9Aqgjxxnq6dQSNs/bc9skJIhK+Oh6OrBjYItlcAUE0AZgvNekfKFNfRh+mu
fudZWdkXwVKSum4PZzPa0G9FkgyjXvekAMo5yIiIIyQG6RMGF+9+9eu6LfNzxckEBWDrUEQW5xHj
H4WmMHEqp0Zlbfn1qGvaqqgiBp8U+SX9eISMP69qujhgCKNGSh4gWYXwBO1bmHFSZAmNpDb4u39e
Af0C4y3gdrz+IgabzipUSvfJd71ETvEnsDGkxoI/krBj5sP5kjQ932xouoHKnj0DPZwFHz50Ch5h
3/+7uO+ou+ZgoYCzgtZ0lkY2THzylxVpmpWFgNBgI77bgRc9ybgHh+UY4W8QxeiqAc6vvqTBMk5X
Q8sPaiyLSls7z4uZh2zAZqCQudk6bx5P3NT11i3eFH8G2WkY3h5KcqHsK8s68FnXIJpOnlNd2gzy
IhTQrNXvZTqvQihnHVTeUhZ7Wgz6M+Cm2+TkzOS45Y6ArWl9eJIVqFeu0Jtx6L2U8EIQg3AQtmNp
QfE6T7o8dIP++I+wdUvL7+GCHQd+g8D0NpLSQOExIQvKzMZdgNA3OLfg+n3ycmG/6JSipavq7Los
oBoh9fk05kNASKjTqxw7vMFdFi3HzHDeO42mIiRrXAKL+wqXwurcR/698tEbdjNdyixZCcLOJZwW
f2h1Y5C5BpDUKeVvh5HsCIQYjrTeWhDdgpiXf7kiH0FQ1DaQ405pt87IiAsRi/W0pd8IVHa5xmX4
NzGDVV1yLj3kQOGnRnhwWdFou6r4e9Tb0uuwA8p8HRz2qo/8nhbxReoeoekD2dGpyeF1nQWlUXOm
Pw1JlpYkPD2P3wBxjI8pngQ5Mvf2tv4o/YpOKd/zAaKfmW5XE2+9ltpbNcO2I5DeT4+8Lf0JJaTB
WzM6SjktzdqlBcOTpS0w6I1maYKq5N4lnUR41F/Jmv5blE1M/cjg+i//iv8mZ9mTPXR/pbYfnHHo
oiWJGYhdr3DZ4G1ogoQa/otvVLySPv5Be1OJ3DNdICDW4nQUfQTRIwIfVEUrRiewiMl8TbnI1JPP
CQs5XPYNf0Ps61lmGSedOQFiqYgWrG1kmbjwkvaE++KgQusaR8wYDCQ+jIzjs0Q5arDJph6yzrWT
Ov0vZr3kzHqCCaFd/SDrzHhG7YHcFU9ysoEcxW8Fdg0cLGtKkMzdZZUEYyYT8cxAsfPWK9E7rq1x
XFyzDQXg+MjIBZ9BjJWm72rOnT2E51RQN4+RuiaMs7jVOFzK1Wk4ZMjGOVCJLCo2G/OGcNlfzynT
l4RBqcjwwm4/CU+1xo2caK/BnNfLugMUKTvJUPr7O0NoTKNq96oIw4lsKbLsm+Fzakd+vBuypYRK
RgF1lOeXm+wD9EmFSMiFLI1zs8BbJtQ6y/8RF2WpCZl3EWYsqvNjZNzYTVbE5kU50J6KeYTesCEl
k9GIlkKp2IB03aBgWSsKuPTwWp4Q+X6H9iAU8O8lis8xbzQnYkiyBpfPxI6L2x0PSTQJLqTl4T1m
BxQOtlK5Z8gC3Q1QV3Ea1P80V0je4dKk76f3DNO5kF43sAjqiAzXHi5heOPyl2CSanfQjcph7UBC
eFlVEf7ryeCQJPczb4H40gUrYKIRbm3zUdXOSH0KLJjipYo4Qzk2sOcf2RMwaSIeBidkQ/lx8trh
6reiPpwTggNtjz+NuQKDFCz6u8j12VPm/mGMom+aSJgir75V7JJ+8QYrCA/aIZKTVuub8fDZLI/D
PMP3f3B+/cAAF9SEhxmyQqFQY10EBzNGuD7qmfH/vsk8qbS2b4Hvz46hZjryUhUEm70hDnZ4X80z
hAYpnCSYNsgJXFXlH+nje7JezO2xu9GGuLDuac+kgJNbfujp5X3ptvxt+m2FJsW2sqnFhiZtjEuA
3sUNhVYkTXuLOyyyWfA6dNV/exvTBCTK3EqtalFgUqwLP4aG8IKAHsvgQ7Fjz3PPnnExq/Z1uX9F
mSn20gaqzcYP0q4C/Kmc+ZPKYhN7vRfu9dYi6jtuNaLNaQk0/cm99fcSSelCyRCILc2FgOvOZXro
1cCeQKYRPkredQwSgnJagofOa85F8uRBxwbtTdH8atMa4wc8LXPDU84L8DxBV5gBQ0UOJsCIOvxv
QUGwcGpET7RayOZ0HHkjL413AZS69119w7IOMZX9q8yqZjDozYrfnbm665KOdGdXKyyWZcAE6uvN
weCAF1k+TJ9EnBGWizp23YMSWgJ+1lJ7Pq1lCMQUO4xt49SwHTSPLwg+sFvux4dsHUsI0kLjAdcF
ExVnJMQV3SLlslGIqmZvg/BCkqx/It4eGwK2OaoT8vwhm97vRvSP6V7Eg2hOoHQJrhx+/e8hgwuX
5nwt6Hu2VzMvKYtFIQHK/M/nyc0Ob3KezUdda/nHHyJeC9GlA1BcKsWgvWK6fk0EASaXjsD/hSvO
/gv8t8TefuxepS95VWBJbhs33dIGJcnCLhaYD5P/rFrT7VVGMZXJTrt829NF0SqlSRpR7yVT3vJa
B6ekcuLg76X1Ywh5D9BzikKJao4dG9q1HWEpkkP8gaimXQPH1C3SZYJooMMuE+uAoQu/jeMEZmX5
gz6w5koXzuAdGUgqbqvH8jPJ1EplhnxfPBvoTE4EIjBEd6rN3PajSDOLWJijBtg7/juHHNa5aDU+
fvtGWu/dXymqioJD8pRs2lqt4xC6kCcA2qif37vaS4976rabKuJqdtgWoal5Vxd4ojokBw2ZFZN9
Gr4TDyr0N/ic+vAyGk0R/G5maI6rhASopqctErDCa2jeXzrP9Dg8JtuVW1o9v6nOiLuy6+nWHOIy
1c5KpNg6w8AGyioc+XXYOdqrXF3E2NpwHcIKhOg9WEEl4tqn2lAcGy8Xnqd9uzfBoA2ZphbkWYkf
ZjKfI/CqQF83vBjXk3o48O3bOK1lCXEx7/0cml2J40LASrexxb5o0vwlvKy9uAu+8yb/mUG5skZt
ge3OuynxG6mmO6bD07QUV9sKdxRVmEA6Stk5aXk1zBNAOeo4Qk3jHe288v0YGpW3N2IYCfCUcMn5
8UDyOIBkiKOoWmd9yT1dUH/2uCotvLVVwjRWSnr6RHJBwEy4cKKWbufoEfYFrmRvB3IxPMOScsnL
WTKF14YGH2zK+Uv6wMIou+h+Zj08n19+eO1UZcnaB7jlPF4qHUJValfSsZSHyTe/CPYzVTFhqIK2
qOu92wy7vGPsavoKoxzSnKXBUbTMiuqEt4SYapmnKoVNj0N4gO7rgAuUbWBAGDWKY+IBfUhUOGC3
RylTetNMWLq2j36lrwYU+rPY0v330U3aMQQMzlAveQJYem9G7fZPnfCgP6KM3d3SX8sdXLcmhT4O
4sAF1owj4hnNpKL4wM4Mxd8GKI1nbVzA/QbYbb5sWLgZjfu7s7pAN+Dx6Yrpr4qErS8cJfqt62q6
Wc0TNkhowGak/siwmnpAbWUMP3hgagm0NibxdIAxpJPguU+zep3pSZK7za4hBX21PbeJXE7FbHap
Ln0xhg/f6R/zIQQvVldOXy82qEEVkL5rH5Et6+7WiGsNF3JOCl88IQjX7bFs54aDvu7zKUISHHdZ
S7AcDdVdbUZwTZiPPWrtf2/yBbnjSFhsIYcJXaZFeamRhxkcGqqQRCOd7f9bhOZuDX/UrMafKyfP
VwsKx9msT1kXTgDcs16gFCE7KZPJM60qviWSP/fhagqqKKGZeZep6CXl71g5aGNFh0d15ImG3SRQ
jh4/jh1nU4EQElTcf2atGfpVKkx9sMPXZoekL9uY9oJv83NWBjmvifdya75sJJoRnonjUczDyBhY
tc/7xVydMQA6e/Q29HIEF1n4Et5ittsEPQPckDcalS51aE/hAmUNsWt8u9RN9cq7FEBix65yIwTs
ri+oxAgyfepOs7IB3Xi+qkxDv3Rkw5LP1IA7ns0RR6iV3xdp8dFu1oTVzEaaMcEmXsHumNaJAKY/
hXeIRWUtEmjxHxBnp6SPpLfq7to5qa9znBZmpZZVn1uo1yPWbGavF4MVUJlm1hppjbpLG/Qyj2ng
TbBNKWkdjY+0NXYekg58o94CFZ3jbeqH3iJYh6/+Eq57Kz32hLF+sroMd3wn0zmfoRfOSfTBmSlR
8eWn1uKmi4MAA1BAdkhR2nwXQETNZUWNa4AAv/cLPDjsK0tGXrZ5v318/r7ysk7Sz7oG8mkzJfjr
STiP5RyqqelrS/76uK4vBFsJgTuy+rM/P4mywp/p5ENfGxSyei56S8M7ktqgG8X69agWuA3qqIkS
Rqtgh3PTJJ7MhVgczd4ONhjR67tYPswVxAcQb96gu1MNCgOWZrFiH1K/OoK00bcSeNUgOj4W8Ylk
PovWiWT6QQwWRXVq2K9vRXh8sbxvDDspZxdZN21qmosTfvzAJnoCh5wn3YyxBd7PQ7NzsOJTv49+
3t9JYUcoQb1wqPpCSYkQEK5q28yglPqKSahJ/qH5SXdUqXXR8PQMNytMo0F8fcBxZucRjd8UeSs6
aV5O3sjNPOjHG7SanyUw7Wvk+f8sFVOKSCSFRpHw8ecfR1wnvDtEYksVr3P1zysMtG2lS8TklyVa
lYN0a9IWFVZj95I4EzhIOHLClOGIgJe/2urn6eEOg0Q3NS7ODQyjXTZrOfX3dzHkXaMiiIxslFUK
qiq9GG+eCu3oQuD8pa1k4qkD/KWX6RjLynJwbP9nytQz5HTk2sGpsu+Jk0zIa+G6T/0VWdugNdL7
AI54MT02z8oDrkCNSbFjCi8kz6fs6qsBV8Lq6Go+9WyKsNi6J5t16HTwOuHY/edNRjkyhDMs1Hen
poWXx975sIgkQQloONBDWI/WRxDHmt+qy/unDsnrtTswfrTNCjjQZ1hLPMnaFWfttWVsow4TMnO3
31gf5W5XW5DJm0nuaEMTujvJ03/IRLPYM0gTh9yi0UVu76i1IoH/m/3I7SgPAblooHNfalq7RByU
kGtS683ogEUrdJxo4TaGtGf6hmbbz3k50SNVNIJx9TqUW2vOKnAHXA8Q063nVOKn1Wg1jUJ30qvn
1S/cAn36s1BN55vsvZRbZn5RI9+ibd0HOGkEZcpHIscwe1DfUG6wdufsq5U9fQgiHF++/hnSnl6G
ffXqhCsxTpJM8QLixX6GqYB6WXojakZAeD7CPu2mQ9IKbWREx9SWBiOt4dezMIV3FvUZIZIe84HP
DhOb11rhVEEq7t64vZO4GOnVxTmv4j6uLkVn8gtytDGp5bnhpUgRkWHm/2U5ftZn8Wc5evphpQfu
e+6E2aLemusOBJM8Lld24vclnk0iHjqDtW8+MdWPrd/StEgou6zpXtESHN+BBRXeZW/PC6ViAJII
SbOycuUy6DTGmgbKRlIeaz9RWhqh/KGVTe/aZSXwj0CzXYb3wjMGj7VB7uAi/M0Qzm5q7MQIyfJX
F+w0Cz2NzDZE+e9eaZGCQSLYJhpzikU9EfqlMSUfmoJPC4+8yirVSQGvmQFfBd7+zF132c+DwaIt
K0QzyLYgpdt5DT2Cbgftt2Up7QGVm0iNrIGI97vL55X32XjT8M5cqxXkIHLn4Af3lu0AS2RiTcJ9
N35OdRgHZ0y2M8lUFW8R4FEBxU3tKt9ldxVkTAHGsVG1qteBFIC3w1q45gzyB1W42q7q8AQnmOUI
525wjscNq+2IOYFoZ9h8OQXJMNewOMjDI9qlzRCbHywa+Ov/BgIDIFkuhBAZltbyzm2R6xMRZp9R
gsbO5g8ByPml4bMYnMb2/v8kFuMtUxB8Ip2IAPbv1xPYeKHFmB685QffgO454hFynF18qeaEAgwu
bt7KuezqKXUo0OO7Bq5JfY6FeEEq0G7AJs0zW79nlW7rYpcxE3sbL8j7uBC8fMmrS+ZMbzBGuH82
CLxaquEcQ7QBgGk84xlvnlbshCD/oGL6IfrV5jImkhJams9oWDkJU5ieOx6/Weszdn8Gwi3SoMel
dlDsCFCxkfJzrwa9DJd2gxzDCZ1d3wdz3aF9DSJmS318e/9LF33W6VG5aEh4RrPR7dthvtztMM0S
3sF+dYLrqVT2lSHFObK2JHdeiAAY5HHldmvRn7/986rzhxcd7gZ8oX+28c7Bc6wKKf5SQVPmSCjC
Ef+3Q4x0mzrmVvKCPLXGjGEvU6pGJKc8oeGlM3RYB8RGqMdE/Ufjrro3Jw4NFIhUU35U80Z4txlB
pSYTgiLsUatNNPUlCGzyiDlHsWlyeUlDRP0/jvtXMZhQNMzRPADetpk5qHPJwcANGg+d6mBYgI4n
d7EpiFQ0WdL1PoFgRAkU87N7UT6J4q1eFxPPW7K2jBge65M3en9C9TBxq3aNrFohzj4Q7xiGCh+3
l0wfqkcAbzCLPLT2Lv0gmWL4u9OO1RrwJopdGgDz8eT+79CLWy82J7p6j2SQohTmYJ8XMQSmQc9j
meoK3qKuhftIxsJb21K4rdfIe8PKdk02HYMB9e7ufzC09njjddf3Jz+SPn84WCws8/4SJ7+W+aA4
IU3hMnlHgcOUzL5Vg8BVqCHXy/FL9qtDwFx0NZdWmOWSd5wwLuonLKCHacevK5NzFeGIbmtYyorj
+zMyCBxe/saZTxTUAoljYHngZ7xh6/Km72my8ACbcY7EbosUVBiXtEEEk3MUJDLm+0ttY68CWqsG
q99X+c0H4CLHYdUaMxCo4ll/rcc1bzARNMpYtaPYvEKY7xm7eTa0omoycEpxz9tJqd0KfxIWXydy
XHAo841knX1O8FrEs6a5evqiDYnzQEnShRmVeKEsKc79ox2n0ENrRG2egAyfowIJNeca/OmAx8lZ
0pmCSYQ6OyH8BlbZq6v10NyL1zmW94ZEQbHLeqBhKOTTtp1Q6mz33SCU3ikoOVgAAUPREiE0kIY4
WkusGbjIYl5128vcE6SpTQiAvC1v641o3sAITbcKqargJqFTSDsAhPxeh1MmF4B39nBvHuB3ak+u
A1esxiLbLqNlsaVt+2NOGOEWXIYFeCnGEuRyZ43elU80MSqCKlKqOuD6bb5r+XQma88L36fjE53G
aJdTXmjAhgGnBDrEbAMbhlDz+ubp3yMrPE8te0fZXurpAFg5wXEFgZTswDP4K34E5sfFNDi73jBX
A3BfG2i/DKRQlkZ/QG527JWSlItWiWF7vtAkgbK940gfEyHUo7ymhCESWBflV6eQDn6z2Hv2Lxz+
3K/FpGOAU7HfKDZ6f/YqmGQNuB76ubdq3pW5+ajOguvxAtjnFkP8sTPsJPzgv5uRwxRXhYDD5bMI
feFby2ZDRxjNsb9gY+l33catvEDXOrIZJ9J0aC5YF1yNogKg3Iv4hBOT/SG0zCBxCMIh4aOVU2J+
7By0UnKqD9qBRDluUO4ah6T87I6o7p2NW7AJP+I4cTmOyPNkSI/S7MoZs+IkF9h4VzTgD0qmh+47
phNblSSUQcvNr2Ww+6Yh9ujVejasP+lHeya8IfI6rgk4Vl5Q6CPLlskjcwLqSBBcbgyTFJ7ASy7r
U/HqUWBIl7YQUbl+Wfz4os60/x8dxaA4s8b41Psde1z7t49aQxJfN7iOXul4BHzGyB/9nE2K/GRA
+EEMnqE/sjkytLK6nl1cMDllxqmUTXo3JN1a00/jikcc3L3EIxdekiNddtKtE282HxtrR+2d5Okx
1169x2k3JJLgxpHbmiHro2STrssvZxbxo7t6EZTd+CAYGidSJaqNhp/vgN9vtdzNIGVB5Fenh+WM
2rNGSM5C2HJ1Ray+xbPmpyK8whI5zbptTqm8l+iRPv6/RJslqKLF1XxLnjmhtIEOLCqG2WjJyl6T
nBhDQrpw3T0fASRoMT38RsRymeo4WXSNb2iK6Yg8AB57x38f5kjLf/WGw1NsQ9Y/1NTFw/F6oPrd
zy9x+yWFYtH3E7bMq0PBKhA3vw1VJMlGNQ83ApR9ti3SPSF4cbckVspovAScIsUcii3Tr1RYUDyp
zkz7H5SYhQG24wZCJunOnovk8nMzrL5xTbuDNWy63ZdFOV/rz8YkY9AkgBiA+wcW1RwiquG4bXKl
zGo6XtyjR8sFQkAnUbpPl1jmesnxkaiObvsvNaSJC4kfAyZYaCnwNDWzRUBjf+4Hktym5lbQBO0d
Cc7cZZiIEzeam7kvYSVD5CHklJgKx0JY+zEI4pBmRyOrtMGBJwJGY1qcbESjr/VDfTN0P0UEF7F/
mz8qLmXi9bdt/0nH+UnDXN2gLgEguTuzturJw73i6ahzazwZ9TBtkxm8T6PLLBm9CYnmkiwsy14g
n+vjVJdxznWgPWdn8GdHhP6Dgvz3FDUiFxcH3IQ3XM21TifRkKVD+mGQTwKydkOFC0Te8GOzeqwZ
a9Op9WmNuoIFIkgQ4seaklR7o3N6MZUkX4B5QzWK1R0XPQRPR/6CgRuFDySKiOfpBJamyQ2Gmioh
jToi0Jp+vqBD/Z8sMRqMabQUMwBWTtVdhkaqrbg4veMA/0rE7PZzP9kjjAylmzPg8pi+hyJuQHxw
Bfu2C5MlNQNWtLBPL1kzLpw4vUbAxQq0kXLLDCqc1glJBQ15fnudVCvCciFmWOxIrm9X6rvo9H2k
d6M+ttk9Df7OT/fIiNNCsOQkl3S3nFbLY4eg4zh6Oph4GFnlIGvjVEosC0S2d0yEAQrWoVQznKrl
dcxY/j8fexxsiMFYlvALBCfzEMvIuNfM3SRp0OrxBHjiKrtafvJIqlYjaJRm9h867ji7CK9hcxdj
OLytX7Qu85fnc+Xwbwq4A/V5o9Jizl81us1Cx5YH83x1ROi///SbQHt5LuhGzDqJUqFykI0ZAmKR
O/wLh0uxaiw16Fy6ye/rNuRk0BGxy62Tx4kTHM+eUxNHHopfFYC3nXcGkZ7efCRBMsrbBf+tn7kY
y1lDtfD2j2D3Hgjh5/1IyGKK76TvZ87nxXX4TsDaBKj3zYE2WdLNiTRyrdXT3ES232FreR0VRUna
T6E9jJWEirOFqV4uZf2gKQA7jWHOukt7NzK+wKPYBx6CimmL57N+czPiE2EuZIHoDaRmbQo0+lak
0JKKNzCP4rWWd17WrJ6IMhBIGfBSov2zEXb0CJG5SgNwWOPKzhGhTpqZS8GAir3RpNzkAXxOAS6A
cvq5/dyyt8aKnrcH00qUPPI+Jf36ImKX3cPQYLaAbjENsukwRC7C48peFxxOJNiSlEEyUg0av4XE
96LAFFXAxTuH89ME1QhwuRDfgwwoJiePHujJsCVKmubO6Og5hJE3RQwOHzM1gHbBPbqICLsFW89R
UVtKU+vinv5x0s4s8U+ITh05ajdOftfHFzmgtintPyr8Zlt9XADP2Qn9NAYnprde6yNdnd4v465c
JPTR9nycbwpQjlEa5raa2KpBK+wJwn/bv2+ByzzhsWooKi+Bt1GrBriIe5LgkzehcdfCyXw0M7ve
mbaJIiJvpmRw5ipA/zO+ng0dmIgaAF7nhMP4UEQceJeAq0b8y7iwEZGH8x+GD3uEK4kY5im2JvmM
p4EPZeT6UUW9JA2gL3+IKTb/HbNP0It07y87LuP6hIhyE92WdLSvE6n7ewYCt9bSda2Oo+5JdnPU
iPGeAvbzB68A0uo6JgOqKUoR/7khKp7k1tJQKePxTS6EGMhIzWYFz541RhYOlubx+BT7FgiIyMYw
2bVkQgTUgxWynmvJrrF78e/xGSC+TlWZIHqCehMAzuvNcKGZjLB0kGtQqqnriQIV9EuAFab9MPAY
TOjhbq2ukxanMqOo3IZdpQWEklB+Mu/eyPB+ua5N6I3PUz3wU/jNot3solaBWGENpHphMd50Vyl6
g5lQhuEFi19ZtLTa4ecWJdqfT5PGcZwkIr7Fh4FV12yn3SGRlm4b9LM/yBk8VeJ3UKorCKK3yjLt
C8K3WKsu9ntx0zTSDjtFoVJ4dMF7ESHckxMyFrQp37VCBEwWpPObR5BjnKkJ4Vm9UR8Xk9nZf/W6
RiYlkBM2kc99YouORdJkCcToiJtuBmgRc2ovAEuvyOyhM8NTpgyvV14R+B3Ydta1iA/eYPqwwJfM
n8hjHRywfrNJ0WtQuSE6y/2zo/u0Au/I0JEJbHjLRMnGfD1p9ThZKlg4Iotlwqx8eWTBny2L7OC9
g/c459AV4ZOhhSTvZui4z1/gEPuvjEfHkey9S0yjnlPf7WTxKTXFdoJvSTTshFysJrSQYWjnrv2K
yWPzUAa2K74XD7WbfaubEVVXoQcDu54ypyKmWw/ErhnnkpiYYT2PzxqrvGaLy0+fVkt2F4i5GNLi
gT0nJru5GK8qjsuAYbE3fv1HJcMtwF5ePyMkzPtBVtDdAGmWJVlmM+ttEp11WhlyTNunKQIsl4So
Pb27YcLVhTM7k11hmBR9XfJt6Ylx0+qhdGrFxBLqPaSd6OEaVjUzzKhh1IlzdyTV/bk8CNPgDJ1K
sKdKI6g6lsr3febxEpmFAmeaahkqOS363gUypTh4w3KzUNBLnYh34Vilavq2chK2IY7u2vl2QTNq
avd8OgHhZzu3fHtc+jTFqUpobmF0WqA+Rj461b2tBigLiK6fQ/xKBdHIzM528eOcU0SkQa60GgTM
nAix+aefkchLtmewWfsDm+G4gHG/yVWl7egjvi8/m945vbdr1wSh3JJff+08KFcrDNTbFlhWzlJd
AlENirZ4JzDMwFpkZediIsSNIiZWuAbeqcJTriVToBjGFKFkOcUkL4O7z8pMP7dDpY+Gg/A+OnTB
soAewXgI7e+oJbNDhpH82SQ2iWErnRFLnTnCDuDvVWj7v6Yxe+utUQPlRMCjJE4of19VlNUc7JwE
X+OTDqcr52At3J8+kPKhmm/kyr8Y0RJrjN1i4WhLVRcbe8TAvZvlPZQAbVTBcduuSZ5UY4N6v83z
JKU4EezpKYwf05cqzpBTaZ6l6TXQo1QdtFS/yFrfdHtD756rXr26bcSzdwlnu13tTPrU5I4XJd32
FB6zdnV/Q3vYNTy6w355Wa0zWbMc6CQgqLj6AdiQ3WlWqBjjsM5XKUDKrRDTAtwlDaEbLrPhtmTu
Ipp3R7hzONEzcgJdTwIAhlxNVCNhi+m4Pt0YdpGDmdsnXZdXVlYRnh7zN2pONFfKrShVP1vAHru1
2vVZXk238alftV3nuxXhZPqLqHxNUy0jUzGegv8zFzvnOO2qmOSsSjwKICsWbRxurz2WJVq8Ch2i
TuOXeTeTn3TUR30Oty8MSy9E8AFPSYRanBPqBNqo6npNu2gLEM2bG1qG7ku/jWTxOXwwlUbo4wHg
R2LNtkLv61NwZigVcVs0MOkqKfCBh41SmLh8UltU6oiiyaWfzv3GDWRTRbrnaHbmsp6Js8tuQ1SQ
I+Na9yU43bfmE3lZ5pP0QVU64UGzamOOFxzWPNboEFAXdzVw4YTnso1xmYcz8rqBmcEEEojfU8MU
jEgTE74HAF0RxxAnUb1iuX2lhTgs3duJSjmNVBflYC8t+eChFRETKIELhfF8cP2ZJCchiiMH1lEx
FdZEmaz9UhVWUcwmExOAR/KfrKXvzFwVnahlNBxS9dRilTxAQeDGLPCrl/I/8TIe4B62A8ANdIWl
8UHJ/iBaFARaQ2XD4o804jdBosIYZQt9GDnHT9c0Ga4dkOXr7+6jZJ/ritI3l+f3Vzoq1hlVuCXc
3zXGahKy2iDN1naI6Mqn7SxSTCptl7e837SwttWnPRDDYnvCdfxz5MsFLNmkYJjvldp2ZawdfEd2
fmx25cwl/H1mk8wPirCcZMlMdtYdEFhAL2OVLZwJ0iK9IX47/tcmmwCPi4IdhKPDA0sUSVNVy6mX
mdRB6df2/TlsgLevlEkzguradgyG6c+lua8HUiSYjYUVIHoyoIc4beRJx1w74Zdbnt96EOCQuLaa
QahbLTPskqtlzsTy8do2rMO/Pwn5P4L5V+o7NX7CBxQu8/RKq1VKI5kAyuTpK80hqP8aA69vkG+W
p2sHKDI55EZZkLV8TKZzQnbQXKmFvqA0kGgPBl1zsynq2SjQ4uIuE41jdcgwe0b3NfTkkZSZeP8c
JpcCPwjw7wQhpUNEKM0bxe6ow9BM8HGWcTcYEOS+xw0IRLaDpwuIONaolKvNhfkp1ZbqME+wWBTg
buiW9zql2UmD30dku2cIGoCupssyfT8bSfnQxZiDrDU3WSiSNZpBMLOqw3Kw0AOm0S+dnshXm4iK
TU4BzI0XYq6WjIoijfsZGtH3TsN77fbJB80LwVi9X9yn3DaC7jgkFptks4QSyNRnk7U1tCoAjc5u
9aOVWpQ6Dq6+YwDFo5BMRrnC0HeJ2kNIcdgjNGOCyMe5OIO9sWzWc4Qtw16m5VuWyshTrAbSiYz0
q7OEDQVi23vvJtiqm4RPNDIGArAoGEzfq01026Z6IKZPWp+QeFY5q7CaOr1pRhcTYQREtCwdy8PG
PBfZteo/A3NVHEKqs4rtoXns2oD/0T1dB2N7CcT4GhQjm4aShBNwntdOAcF+A2Cm6y2IZ/9hBm6T
iUx2KUSNX9LkE9WiXuEOkhZeI2Oo8A4vQeZ9Q2G8QvtKfPGCzA2q1XIVZcdjYVJ2DWB1kcy5PwsG
pnBRwtrAmQ/Amaq3pxrlY4UWV2GcbNuM5PZb2qPcwKbAdunCQhBROadnnf3OMMVmhgUQNFEXdS1q
QzPXpoOKz8m8/mr+M0iVxAiXCLE5FPCyX7Grp/iIir4R+dGQ+PlCYGL6PlaN9tJ1UGQuiEPgz/Pd
mf9nbHldFR8mpUtaJw1bgX9Tz1FgkUCmvIs1SNjU3l73qQDJWrDROYN2bs9Sxu8Z+I3FihgJknPw
3VXFPzKEHs1kPvukY9onYNy1ChEG6xizGVw2kz0dfrqYL9NIWO9FRkrTlCpUjBdZQuXLTfhkyp5m
AiWvVAUueUgZVTNRR27WLx7uSznhsBuss6OuK3rw1BPPBGpm0iYYbE45iF5u3kzljbEfZABneJ6O
Cfyn7z9VcW/B4pGUOAbq3kO020Ly/edT7KXvWVi1NWf/Mygqmofvll1n7Uuqxfev5f+RuHkOXL5d
neqEt9E2a1SL5BYmrBmuzmKE7xb83CPrYJzY6of/F8g9J4eh7yjJerQpTuV27XumSMsPhtJLKX+g
arHbwXBret3YRBT4Mf9WZdufRk8UabdwjEqqF0E55nWLYoWab/S+i6xQWwdKaD1XEq2LVVGHOBmm
ow6kikhYySkB2bt/sIZL+dXtzSvF4KqFTjQNlPUKKm35Dy5JUxUfQsmLga6tCJUWgRCtvWabEb+d
eX4AOnA34gl9eOr734wJY3wU/Q2cc9aIhKmRufiuW4nuDvfnp9Vll9pgR1xNnwRtgskg+yHmHKAi
VGTfWCYEcdijCY4ltjG2LiajpsWaJIDyB/udNvPYJrTOIOYhzPFYv+5oRef7mZKSHYauDPt/gxls
bk1IIx3NpvvdwLxlvVYfrSpzcFeZ2kRzW7l8fioTcg0x63LWa/FWdw9Z+blBtFphjkK/1k9hcDuU
YdjbPaVhTsw0mk9vBRVAnHRoYsuK8ygYC4Nx9jv4ffrLeKcKJJuwLutYGD1wB3UDW3PqNvNNjaOF
pHHuuz0WHvmDt+3Ai8Qqb3PpbEstlcn71XzWLnlEsCqkkb1mLBEmsL4a0TsNaz8QqjCtvfPkiU4G
Tmd6kDEa/7d4v4RHmSxWXKn/zpU634LNd6sEAVKkM9KfXIVAq3Wnu3TcDdyLMXDuOabQ/UNp2nVs
Ok+pMo1fZMXx5kmiJM6Q67RX6PeQDg5Ae+pKKbj/W46ZQUoSj7G4bWSt1nd3/ro4VPjDs3mN8nKh
05WV4i2PsdQASFzL3vBzEcsF9JYuY9J8NV5ucNQjmJ7Gw8GJBpp68vEFj1q6fmzf8+P6xkgvBYQS
wgUcrkUMi8ZCUJ+bmdMq0Lcwm0AADWqXRlilN/saNI1fiIRpfyr0U/JRy5ZK259qvcrAR3WaqMSz
qT9QKJb+kdc7ypVExcU2aSA3yUNk5ZFXLWnctRgme6GAR+IZnoFMhHMO4bsGymghjg54qljy0Qos
t24SX/WRZL76C3gpWLAtib5wyDZuFMuoc+cgNWiy8ebXXaZ/EvxQyIFXfs6pQPzpLtSAfo5y8J/4
624fSs/9CD9H/lvl2u5/4dhv+JYJjvPgdDH7xqFfNCeXRFzEdgVGVYBydRmJzJWT2XLKkz9US71o
CiORbiQR/yrews3TO89Vg19nEkhZtgbfwDoD3KAABqITWmEDU3QJN0H7J+HfaJ0Y2dmTDTb0opq8
JEe7J/+CFcqSwqE8AOYVpfsM+itBycRCwka9SJi2JqB6ZNndAznXtGX2ImfWCOJ/6frVki4yxi4K
Xovq8YhufrkRGbIivlw6GFxXimMPykD2trumdEx7OqCH1vK/M5bVgJNl3d+9o3jBbqF7jQ5YjVvz
GE68yzyuVvgLiAYEde05u5fHLgxEajyBX/JvEQXO1BzrYnZ/KdIqZpb6TUFn7ZL0tSX/npXDkhcj
jQjwTFSuaBs11qilvHkpPg1R9nUkPxdSxUP8eqWADxdHIbm931Ukh9u+StPcpij6x1GLp2PNdM48
q/cnq5Oru+/ijASFAhi55WvHZ9lMT+Wl3rgYmKhkwIJbZ7oTg6vzfAQFnQccFYNhf0TZeaxXbAWJ
yuSwpKfmQurQfzQJFA24dtkqfZMdjYR4dZ8qv97woKaswSNYJmAe/PUyJNmEzh6gDcaAp397Y+hc
tm63adNGBEnnHHZjaMmDSTklkDgGmJjrBQ6pNTOjc8ChedILAU501cRGjxWWFKN+7esWmnGJ1mhd
CvCnNCKcusNUE/K09dflzOYDEDN0JzI6DUJjoLMEhv1ILzYeqctVUkaZOvVB0oJkc5GQlOYHlzlD
G0vHcqzP+UfwLX5i8OdQK1E9KmQJYCQCY0ZK2cpkfSb078DlmKna2mDGZggcnTcw7N2S4qCjjNnB
IMQTNxqAGYHNbDChiDK2GyoJZ+SdjCyvob5A5OPt0LGHYO6Bi6XLe0GyTRgWcWPD349EaHRFv2ar
TC13boLbcMbARyBHSajr/wkUSXEU2V0EQhV+y2nIuzkbVnNHGq/RimNz7KDeG5OPft38xhzYxjQJ
SZ9+0XGEr9w4WpiHrC1ih8oCQBSgLtLkUYWMHlz+TSLIEHRwEOnYpRe16vnkazhJ+xmAfiaj3psz
2GMYOfvRS7Yb0ujk6l1fCpdvYkvjDhV0ZwM9Sidx4u5sR5WTZJW6xu+wz8+ULjj8fSdNPqM3LW4m
5Nv9Uz1sx63An8eMQ+2vvr65kiYLC3EkTFiDTF16wnUBHwJZLofCSm33atzLLcxIOiW+r5NG1ta3
9W/IOkDXGLX/TgSVIoNplzfikSrYt4gumLLTeuRSSvlGeTZciRteJFvM4n9VtEQnyL0+kZhqGDNv
fnnOSNvgSWQsWM4EZxwrQnf9pJehq0T5T8qvI528D9kPhvxzsouHj1kRdUFM9NT3O6d/GddB29t6
zR0n2BN4cPhwzisuQFHbgDRaberHm5eMUJodigqSTLKVCuYqcVZhV9jG0efno9Zq9mVyxm0XfMd9
ViWyfDiySjWAH/WN42kJPah+4qWXYT33h5cP3JgUPijH1md11x3NmZ92XqeXsl1prkj2ggJoJOPe
LiDonJOhxaFszLqkpQXMozGYeCBpXq1pC+fOkMsl4rTW9J1kgpWRD0JFEqLEpNvRRgufclG3awy9
mIyXRALMNBStCoHbj3JKRKIm8bwnsexkt51ZjoN4ucAeOICglU4tQT8tydHkPFPwo07H0jO5zzJV
buorsuL6hpwF4ZHMaThqOYwqRKw5UaEYXA93tHFqUS5z62+xZBvUWjKsF9QYuNo/MDZdShEtlt0d
h7oP/F4kTfGuhlYNJiJ5WlYURsHphnlQkm2rgmLNCJbpGI41F2Hbj1ETnXR5NF0ZP987Bn+h7AuQ
D7LgHPi1IBh3ZCLKGSCMZG7FuiUTCQkRRZA/I7cUI52988iUcdqL1Siy243f8rm3/E5uiHkqirMd
43ekD1AS/tyYI2ck7X/cDILoduV2SjHUx0X7vg2YkkrMT/HS0JRcKykmahroSnak9EIhQaMf1Y/4
IjcipAxXgrINV+x0bE8kZpmkPk0QiN8LH6qIRFJrndSYpeBYcm73LdgLvYt2dNPbz7FUPCO9guun
ggsJClqZ3B9B8y673rzdKVgxNsNndF1Qxwd1ubB7bC6BV+g8mct4utNvntTyuLtbmQZAVc9N6DtS
Ccs/pBD1aWuTEjmFh+D0JxziPteA2SEiIFoofPZnIlQQ9vOBkUYOwVpLyPOnLF8ctVma+VJ3dxHc
yNLQepTEcE8lx+d0wXa0PXDh1rLLKO/BQRtaUa7bYvx8vdDrLvcY+6eDtzHZ9twajm61Q5acxsK4
DMVv0XlvPf4k76bB+Gk5znsJDgZ8aJFZNMYHfs9VqjQvPG5t4rgrpIfB9d7+RTZ55oBMlPZEPuMR
P3GxP4n8EfPUAxKnG8l+8HRMRyWqCeZKZBe0670aLayl9r62SsEsYWiAro0JSgbaeFG/NEN6b7hW
NZ8pA2lzSszSzI6cY5wBb5PxBjyDRD9ig+8wGgOSoVuQ0yxJVdfk+/XCWhGYvwlQ/8YlT3CuKKNt
3Zz91NvBXSFiMcDNxhA4q+FVq26i/wvH0oW+8D26sLUv9Np1qVn6TX/ZW2CCmgTDRv7xKH7ik0bK
Y8UFNdElXCsNMSGM3/FMmgBISkURWeG6p7jG6pWxh5eYk+jTZUctwzHEbDxAM7AdQ0WtPhmhhxYf
GnZqJudYBbcdJhPsa3Ff3t1M5QoEKb8kApRRp2EEr/2c/7f4LxvYHf+w8zVjMCztvLx2uKYn3TG3
0oSdqS+ZdbTZ5++OILC5nE0rTg56fQ2QD/6LqzNcg9XXzz+WnK3RhQ2T1ERLbvGuiSBRjqpHIjsJ
JuojNJiqkJCSnibT4jBNHRhrvBmJJ+hfPqrgqQ3fFZ8jjmxyX/rHwHvNbsc5Xu/eZxadwBeR6Eyc
ruRb8eB8AEy5DglYYdtOKTnJA2NjLlmxx2nNkGoG4LiEQuTPNXKCfk6eDzDn6djN1HmWtY3mU/St
mE2qtDN6LBq8ExoiLjqj9NTWctrd6ALOoHVU3qLj0icbdWnzNyVbvUn0PQMyQJpk9iffF/qFT1x/
/b85XQmVVa7SZgg8recrjCESLfTVEJxxH8tARF7z4uXSX143qIaIqdDZuwg7zhDxxzy6dMCDL6dB
6qzne+GQ7etQY0qhy3H0BtAaR+epohpfu3nhXZqjUGJ3BmH6dSc3DfbiA7vBMuSLJtPPDc98j3Eg
UQzJtnTUPh3i899Ti4y3DYusIjK9KDOZpM+H6RGrSqPrZP4txXntRXLI/Bf1f1iQHBiteYm8V7kK
NxHE/175DBb6z5zBdoyReOCkMJX05PAwnYsldh5+Ou26vsRLS/UakEZrolD4BtEqaid5kxW6d0Nh
1tPNnIY/uhqdsVMWCAV5J8jZUFPYRdkw7qzYRdct06WbOrBQ3bSAw0DnpqFcfzg4nDYiMxIQUpXQ
QqkxZoaAVF8wP4mdV1pqA9zvrpOYFBfqHkOCrLfuHDsvZUKQOqf8R9jmDiF3SLgcu8neSqBISOJn
u8GXNC/AYihaP/m5Ta+g9MvLyyzBcMmdGk0KnET/6p5hmNnEuN7oVMJRfNJVid9d4vv6SzmmsYYi
p2abl9pJMLVtQJLqQN6Fzlj6GWboIPlx+MLpBjw+Xjmx67loQnqY35dtSOhOgT21na6qz3LFCzPP
4Ff9HKV6E6fqsyl1y8Z3EkGpbPN4YVW/omjqHY4vx1Vrz3tKTvrLNfjydEFkDc62JxJ0oSRbWYgE
rHGX2EU+0hi9K1pcU1MF9KHcH0mhGqPluGQZYBQvo+Kx03p2o8/WYPd8oFvcvHwijGz84UsIsbgD
uRN8pTOObkAJyyZrWAELqCt86wd45GIjq2GemHAh2R/JIntL7UvBIHxUQHxbZKvgvw30K82pkgFb
8muANvhZaou3bAWxPw44CEsMST4ejswV5FfKcXKQeqVECYk1K9vmXpNJOGOlJGbccobb7ThG8XHr
9pacEJmKZX4avkqgzIAC5korccFktdTaplyhUM1zQgbC+P6jMHEy+joUC54+J9nhLeo9l7O8ZJ5w
xisOGGgziNdo8+cZqnKZcPSb6OyJ+pl9BHY888ngLabTpObjoybuDcmkZqMg8WDkaEtb9x9VpC4i
pb8KgaA+l3Rkb0Hl/wG9QwS+zBo+bI/83g4Sq/PNkmRwq5e54uF3jS0jNnqhSLk/Tpuwf+fmnvIR
RAZGvGqQFVGvA2yoXb/f6LDaeR0vxTNzdlHPZ83ynikggadSIgjZBlv8voULDvfuPyDh+zPiGmUm
/7cTcp0CmCww+pEvR4jte1S1X0a/Yd7a7nSMRyxR7pmipk0fzh6/Vr0GlJA4CVvGM8/92znjc6qS
+C3roycm1IkvBMt9WcQOexLePZG0gCDMvKblup0bH7KcAPDhfQxNyWb0zfLWdknr8J9jUrdzp/W0
FzmFw3D0WmYT0vhr+pW/Yh76vDbQWMvNiwtJnWNFCxWw4scMkgrQ/KmGeiR97hz2Z+L3udEOh443
6M8f+HUG/r+5zzw81544llvAYFXNtMAT6LEz3lQ3apXz0NnWcXrT3jjxv7rRU1kqiB19zFr7qKoT
7wwpg6jvFPt07f/8B9+QVUQIT34xAYiulxepfu5zjaerzhSIPsDc2Y0g8jJiPWOwkRkQas32GJOv
LIGkxZlSCcYc6boEyKJGUTxkMX1qq0iqpfSM+29mWwLeSijCuHJEVoB15eb0GV2InF70dkAYj/Ht
TrCMjSA5D5EGO1GLVQ5KHqldNwAyBX4ljvfAVNyvysBZE4q14uyKzTKb5tw3AZW/ZPeoT9DkRstt
Hg/ORlDebNKCYM9pG6yoCO7zkOOBjWyoLKHIGwf3cOhenJc/HVI3dUaOpeUfhKsG3ItktYnBHY4K
gXpNxf3DPuCfWxSBsZ6eD37V9SkbUijQd7cg63ZL0K9GfOQgIR+aQYcPssB8YeZOzw8iQzzqro9F
Ic5mCJGDURMXgZMeiordgwJ+m1+Q7T+fRfegYJUqwXXULBqATuJwLm9NjSKK1cFq1eYe+FFicSuy
vx80oY9NXqIxMP4siQqpPkKIWqAzOfMYm9PS777jCdgLqKwvZUcl4a74EE3EMAZzXcqYbRehkEK1
LwWTL3akLyHGDzL2gs8quhAQvnnhR+YBObOR3aXdXdT5JNUNrDiKh1M1K4b/iIaNPc3QfpyTmKkD
A02glZffiwLO8Yp9tVdPjGGAyt3Clq7hxs3rRW43x84rW5LB5Y8sJvA8tPmQ5NarmPgwm9Mu0n2a
wlyTRlp1UC/ZX6e3hyA4w2Hq/7UXANR0azId9Q0GPy5CSa9ImThdGOwalbQyFZzX8bld9baCLluY
rS4vORlTXRwDe5mRUJg+FKtfSUIzGAJojXOu9v4KuQida1RV0Cu38OC9JFl8/SMQeE5p+khMNSea
T8tqmcSMiLhssT/lkHgTVVbKAH5MBN0SrILR81IeWLFv/PC8DLy2V9QEuxL9RCLcSI9jbTMLAngM
sa/9nbDkWS0K+57oEpT5v3MbokM9aTEfL+U5+olcrxYTKdM/r46fPKlb8KRaPeH3z/YI2aM0teFL
yge7VJoDeojPBeQ32eOquSgveKpqvOYLVAI7l13Enfk33o8go/bsKQoN3jaW5/OAO0xDs8hUk21E
BA8iXzOOfE4Jnt07Gl1UxnxUrCPlz/p+ozpR49aQoedrl6TqB5E44ITzAlDS0I79e0CT385PECbz
ADLA5DpLM7idURGwtVYm31nEQGXYmvt+3fyge25gFTCIQ4KGCT74+E4z+JKdyPmQEpON2Y5otVxx
1gQl4cmUD7TZuHQ7vAstz9XtAn7LdYR72xdi1dMptWh68WpStoft13ypQ58Vb7jU3ItjqgX6xuf8
SCG+Rgnz97Ri/S3AbqPDFFAgvWqwucZiNOPCaz5etsMPQhCg6ILSH0wbn9yxY6R+KHI3NZAiCtti
Nq0BPQ0doreSE/1iBibvVZO7lHYuRssHAzoL0eO0V0hgkVtsORkoUraAHRr+cIUoBMUQ2lvVkqn8
n+I8yxG4zDdUwJDFBoUIOsAN11l1fjlnpK+oFdztnC13r+Z8E00un9tPg35wq3QfjzabtzpVdLaG
KcYr0eVVnAlPtc8OtZsXGWKUdZV1JTeN1u0KU3wTMa25DYoU3vV/YiZz7X9s3ELkYe8uqUnZhFdI
V4jt+HptD6/Us8kHriApqQQ7BNi7687yvQdFOEQ/OEvKLVP26MKYGQnhmdKhi2KAIs8e24Wcv/q5
DYSX5A1TZUi5ZTK+QIotIYkcn35nGSlSOh0+X11I4NFPHlBUbdOensA3qPzk7rkh+Xzb4caQcx+o
3GnKFdbT5yPxA4IMNO5+qyW9jopl9jAserqe0KOU3mgMpl6PODN7Sty5DcbLrc0bg7g7H1chVD1j
pJfGNTbTwyMWS0w3D/Y8sl3UjdaAoYkaKeR9mlcFrPZeIdRp6U3LMiFh+ERyx+F83+U1SlzSCYqi
b74IQVTgqOyyZGFBZPBpeEgMoAVYwhcQrNMviRl58uipPgSkqYJTYEqgiQaIdIO8YzvEMBy69DYb
PUwWZJ3lb7s31JZcmt1Q06SiyXOMoK8h0iTS/naUHOGmcOEoNtMyToM+mU3T/R5sDDNzs6KyQZ3y
z4bLGCldZsAXHi65jDcbrUgomAQhh/lnaxY+tIQyCkI+ziVTD1lpv9zzMWjvdH2fYGmlGIVrlkuG
24+XzhguaBiJXeHHgumLdYD9KKJk/Yl29UcppcFeg1FaZ/aQAYNjHuxkfkS0ERqcki9nPfh5fFej
SjPgDksUi5dShFYlbBk7Phg2pe3sPs0WzEnimmeMa51lXWDRvrSBVVeQbd4Ko89gLFua6dEvbRG3
vL+Px4OneRVk5m4W9NgJ8XyN+qhXv9VkptMCzxMy/zKiReoSmTOYWbwUxQ7QHGk4y8kDvkuK2fht
AFGej7IgX24xRqw2UhUOlf6LXBgI2B8MZCdNyZ6asT4YyglqP2Xab+k9glFpqcvvXoLG+9B3jC8G
7fO7QVs1nbZG4RgJCf2EG0/+/wxomM78qlt18d4HNc10s6R7qRRyhqdFR2OooCQiP9Zh9eghbM2e
w8SI8zMD1cyjEu1alGobiNlBk2+5eI1LkoRr3x3XnzhoIkBFDpHQDmrUi+vLYs9m7xavQhZ/oCPL
BDKSA9f+hHkvhNBL95Ex8/jgl23UzzXRaz67zKVrzrrRYAYjg2JpqlNAI7gwNGSn6MjpwDY1AFvV
e/kfwlUZnToW5YAu38uYuGpIeyC7wJT1LTuAfaHHgv0oq0077CIE6XYx9k3KFWurUmKVzOZixVCD
l+yHGrhpLdH0d4dxpEGREngS5CQLN2Scmh06UiQqBkQDPOwCBkqSkx0kyzAWXESX0yf3LBTuER58
9PNBiCncK9HzrlT6cYYPU6FyCVrzHkuXiIq+mTquDF0YXrYhsqA1B/ZXmFf2Nt6kRq/4CsLq4VKl
/Uqoicaio3/50g4ol2X/WC3fLoUdg/pTkcv1evyFjE3HNIfztnJznxIhRTd8JKiNxLms1GAuQXkb
RbWsdVZfKqFliF87K1W1jkvUmxj8Yy9NZKwU0J72UKelXSjlKhyPQr0TZ/GLDSbo04HdL0Q4sYVN
HMJ42hy98iiHW2jLxAvXC0uSHZTGU4cdbak7y3p0wV124IHv407ETNlAxET6w25I73p1c7XJmXta
VYPWhJ1fWTkAu/TrMnSnAU2RdnjjOudsmxdei1dOxlG5cbKFD9PBTI6+rpkh1/BEE7cdJyqE2tLD
2PtoJZB5wd8KxL+emBVCXIxJDHl+kS1GUGGzYWlospXhmWq1TF1k1Kkx/L4wvbXR7eo7g08cNiNQ
yrtnxGxMIR3RA8nyjRHFFotpgJhg46YJnkrA6Y3UJem2BCJ5TOU6F3c/M3uGUEnIbbxheWINVt3K
S9Neu9lnPgv39kiJQCaEjgczP3AudOaWoOcEdSGOwTAOtAGUutHxte10JIzOr7+OqNA+nT7ATmHy
HvQ5nNuxdTlGzTOuD7gjtTM4ze2nG+SG2r/E3IwadrHzrIMq0MOnbWhu+q4IYHeOTTG8vIYZTEH7
LHMNywUiy8ZvcPR2WHbsZfFygfZPoWWVqHZY6dtd1fAvHrT+iJXnVoXB/sVS1neEXvHJVD8OslTp
HYr3y2fmXDjr17DndL50McvYJWlxyqLdFBuH+0eRJ0DKYeGGQnrl/1kGhImFNiYFoKxiA4LFjdkO
mxJHSEoN3A5GV6p5THRHkBD04lzwLfOmIIT+N3ORS9ZsYBHx1XtqLC+5FceA0dIC1g7Nk36TToVm
5nG77Wf3KnXwwAQWB/jj6OCHk7rTbUxtKuty1IIwqKdmeZTzDHhafsC6FBglKIGXxO8UT5OvKQid
jzRJ194676Ghx98aHmnT6JjCHJ8cHhspVlj96WcrYSmOP+HepivY/iNxs9N54FM74aNZ/zjc81bw
xzP0P2i2azPm0NlLhdBy3AHF5taF88dR504Qkqoj5dlUm8ykbNPUTX1afIl7mOoE0+3J4zCLgRy/
MmWW1VZL240A0IrLdMHl45xy/A2ohurQSotxSvhZWezVJ7ZKwIijOb3a1g8EYnvPilxgPxlxCH9B
L7E7QRb/hLbqZVcE2Fuu1HAhDprCnSAs1/G/ivGZuRgNNmrMDGqIEOtxYQcky7OUY+irEmEMgD1G
4MrhMY/VY5DRMnJZAVA+V08w4xHpceyat9e5VvbhSRE+wCJKZBsL4ZiL42IroD6h/ES6K/prW3gP
nLxDfl63nwhoBjyvLmlJD4hks6eWb+ZGN6wcoduHMDlewiiPjLCZkVkGe+qWuj/MRuV6nx37J6nY
1vpgDed2zoZPF/WrNjWn+nNJbm+JZII6sC45WDM1P1JGq/jjvdaFzzvDbQqrDAl0VBHmYGyxVwCV
Opjabba77Q22aITAdjADx8CLlRVYX8yJI92m8bq9A78OGHii//+UVuk598IfApqlHDcz3lOmpkOw
GQSO5Q4rLGN0cB+1jvJfsjfz+U2UX3DKow5yfvy49xW0e+qMkkQiZvq+1W7G0afvhptQduHFm8G9
HMiwh20xzwgas1avaGevfMqOTz3n1W+A6qXldlPrUCFb8hvATRmLzl0QB73buxzGkpHSYwLL6JJt
G0ndxe6JwGu0nDOrYZtDB0DXNSQL7/2mqJ0/RKJrFSo4LrOm9twJl3dRwt0gV47rDxhOWjUQg+lD
ljYkjj4znfRhHhAOeDib/0Be/aFsjWiWfff9KDFOsMINGJp79GffyW07lkwhKz6F4zW4ZjM1prtL
s6mQNNxZ4z0GqV5ebSegIqo9dLXNicAf+9nAcYGbxD9NeDfPirLRwbttgT+1OPkoWArkhxV83xKE
+bi6u0yoaAwARWe4GIkEe7Nadpqla+TUJGPfJf5Xwkb3j7sMRPe++gN0y0Kk142Azt1IrK0nypW8
hbNwNKGnqTu1/VfdHVCxoz0uBYhP96I5o3HHJ7nJYnaTVvz8WYd6O5j/NktST9oBXNNQO6C+MqBU
CBi5Kzpg7AtwbjZbG74MvQ5n1rItu8g5juRzM+nqnXB2gd1Hw9irmvsDnwmCto+EqJQ+SXQHN4GD
zxUKFtXFRhnjfeOfmbaUtUn+PEInB9Gct7SJfMaYj2SciGLp1gAErVsa4vr/COgaNBxiTkVM80mb
YEB7Px+mSIqKhMSTCFvMd2Y7S/okYIgiAj4ndO+YbK+xqMs7KpzM1XPYD+o/xr7oIjfq4k6P97YV
9lfuqgtP0JCT8juQpvFL98EXtxrspSLqk7BQ7v+ABa2Ovx0+3HMWth1Oj+cID3tyDQS26BYhZNn+
7bXW5AFCGYcG41jse2fFFF611glOx+720aoEI4xnZeEJXPHN0e8gWiPUj2DX63jSVbD9LC5s+OdD
YnunqzJJbIk2oFAUliVPmyONrrGRJLMgokvOCcsVagwwTqdhBD2TP8iAnpgyYjwPuC+4F4f1Fnrs
UuUcoAwQ+kJ3vEWIOiJKXirsMpDA+NmJUKTWm4/KvEkhsPL5OTwtTFLZNK73VWgNlude865RyG1l
LSp4PYwJcEBGBVWMHxlbAbAuH6dzH5xecc4JKGQ+fp+/GvMXce55FHj4N+UXnPo7Qv7g+BzMJsfU
eNtu7Yi+LAG7rxgx4EGx2CCXdhSmJqHMb0TF8XUczFnC5L/y3upJMwe49s52rb4TQtpGUSFhIEe8
dhj3ZI6ac4mko3WYNcCFFdUAko7Ck58hVOfahxXedmB1IfC6BstjFHR7AWRMRLRDANxGYHvAs0HR
4CQEy45BBZRc6ldYJOnV5UI12EM1HcwiMt5YmBaeUbJ5hey0huooIP0IUGmiy7DDKxlBm/XVP5t+
D261zQCJ56aT/LqVEK1GP+FFrfb8arnqPYTE4vCVmwxxfZAcZ6VL4eqB0JBPan0Lf3KtIWTFZXt9
vRsmimTPBZBrzWKd29L3y48U3a4sxmGNNwvq+sSzh5kmrI5wd1FuofUuMt/XkqHSSH5fNWhsWjBB
P9RewDO9eFsQJV+8x/g0WI3KDcnTuwHGAGC3pzLF5IZlLfW5sJRDU1Ty52jnBUDpjzqyhw5Ta7qg
JQARUnbMW/gyoIAIEvXk+Qjfed3A8og2anfx2BqJqMMWlY8XT0M1p3IF3elyTLrEIByji1KUhR3J
GMR9C3o/MzqBQecJYmxiu+L+5HG634HhuTR6BHa0KNceOZI0dl5ns6rqb6tNIQbOOwA4EMOGD3tz
219Q1pZshpZP2oobipNJNtoRBRKq6jWJ3tQil8BlkkJKGBxAT16ZDJTdKw1lBMkCkuylLgv+54YR
YnNh5KoZJvJvHXq1FwdiQAIpGZn4wy3eBOez2tD3/bbcocxoHdHwITBkRrOvOdm/Zjc3PqkvLYJ5
4OBYCAodPnhnmV/SR+Nudl7AwYTbxCzwRAf2pxu9RlZl3ShS+SNB3e37dS11005T90BfYFc5yBpq
E1ehL2+JPaN9qWeNCQ+KpL7VhY8/Rsng6yizdPTF/LmOHPEQm6mIjo5oDqg9FoYU6YhCVXbTmgO2
MqpC3rO99wysQmHfNpw1VDIbq+lj9JP6tV8vRAxpUN41WqVtN2HzkbJvoL4Z140DDuFDl3VOo7bB
dBu+ftCcxwKujuOc+unfuf+qV1nNUK9FF0lXpiAnPCDqWGUANHQ5UqtrGD0clfyN4ldtnIhqk3Cm
exqWIdbyUry0+esJK1w+7GTfygwyVRnvq4bI3AOA132S2PeiLPfzdnr4PThN6209axJBNE/XOt80
GjqqaY8aHAm+21MsBZHwpjdW8aaVRZk54xJTSVBvzuaT7Cf5EIDFEANwJApgHc1JS4bNdYop8wmZ
T/jpHOv8dB8gZsu4ffc6UrkYZK1z5RnvvOvxyosLxy8Cfqxu+rBg+YB24iwR7J8/8+oLcUXh5O5x
25/EPUTzYgo+2RolUOF/i86JVHFEGptEtGJCsmRafqmlLSymIcEzj0PdoTExWoK2SOlOgZET5DSt
/3BHe3piyESGK+wZuaPKJvZ/YyGsYrATpcqRkjgY7y+oXuj26WFKk+fGewrVp20s0E1wWtd8n4dN
6qPb4OFWPkE8G07Mz28AR8Rz0SBuesdpXzHUF96t62ZE/jcXKwErmvbglUfH6cOj6LKii4xz/E16
xDSKz6VrP0/p43yiNWU8RyrSm75yBg/WNAVMyb4LEcTvzlDhRfEg1yP4EKhiqugvxnRFP68TN4Jq
f257pa08XmjkhVD3PTQANGyj9QvgqX/4DBeE/iLUOgEZNAmx+2mMSIh3kTZmI9O1aR5uq7Bj04bn
TUEqGaftxBypcKcxoqBw1YHErcSotb2cp3Hmn1dFwjX8UupJSKTdVKqfUTP3xyRKGr1tiBcD+Qcc
2fbneBm/C4A6i9eiYuTQbL/YlI2xnrsiRFuJOydeHfXsmDrJ0SGLTmqfI1k9qJ3o9CYf6UlCsbY7
Ms2wZ+MFFzcLnQo/mAqlZvib6LWh3Z11TyllvUAn21k4/cgoc27EU+1KtCMLAiPmT3PamoRxgetT
2Z7OKoo2CV5Bsg72zGevirxm005wBPAPiFG6dEX+rq6D5z88rrJlOTbclrICMiExhQ5ypLqecv8x
GcajKgUyNnkIuQ95za5EXZyvLTKVXaCprUeN/Xw70C1qow7urvChkG5tdWCWGwvpn3C7ID3HbgG/
t7Ke3Whbf76eU/ilITHTa9mA/AhPTFLhgt0WXXFG1VjNp8JHsGHUkPe5Z71XO7BzdTkVJ1QRPm6C
L+pg256eQcrlRXhcJX3RVC4qO7VEc+iE4EBGasHr2N7hb/eCvbB/fHbw1L6hWsj/qS94gfmDphlf
LjS5prcEBPSTGFVkFoQvg8Qwlt/qGEYuYaUf9ceqNRhH0Npd3O3AARTR9/Mk7R0/5agQPsXM5Yme
TfDLotI4j1klK3MazWGeh0vPyNcloh6aQIqW0mHuE4vWM0apFCDpqMV9wdt3AmyUmCPG0PE+tkdT
z95LZ5LPnul3++eIdcGHmq5+8cl1IOl8w5hc+OZnb2K03jgBYwiAkQrU1FrWiFV6KXKhGgpbZajb
LguDVfQjLZ4D7C42FkrLyj99OzdkUcOseLkZhEgE//C3xPsh470QJxnl667glfGCZoKLC2Ng2GQi
R3a1W8V4X2uP+yrG1PZjZX1NHhEmpLEVfWX/G4mbDqcXR1PS+XVmFQT7dn5UWp/u7ONEyHRWH6EI
EsKtNees7ccnZziARiyhvM228RJehbn2hygeKgoWv7AmB9nk3rx05z4MniY2RYWT4OfOrq2AHRiJ
djvV+reT1wNuH8t7Sg2p+0qpsqdjMZP9Chzen+KNfhiWpPvVuIvZgsinZ2WeQuuCda/X89YDB9fo
+A3U6IgvsDWL3UeIzW2nA7dAaju/Wwd36pylKVmSMGX/AOK1HhkxXTXH+S5xCGxWwLTqzXX1dUxO
uhscmE8DJkiwbGPwJXF+kg2eD64xahwjaUaWedyDoIgk0kH/F3B06o+7uReO8QlZxMe99LgxYvtp
iUpXPBXfzKAQyLvCrsEhi/X8B4SWLx01kHuNKwdXoQp2KmEHww3YIvP1lrSIJrGrU+nI0iYFO9/t
7xX5YsKAAmd2D5UK3oledxejlaVn1b7Ce0tei2igy7Axal+YHsvkwCYAu8nzypaiJItU4PrGi62c
J9J6nOODYeunWGyTKBcs4LcIZRKiB8xZ/9Qcj0NDadG4lGrcsz5/BEm/VSDzPSsNLRX8fbkyQ+eL
G1qwwaGrmCRnvo90kTbPpEXJwO2BNf6GgSg6wKPlJKEJJ7CS21E9Wrt344XSn9BP9bmmh5wevnS0
hBXvpelqbi95i234CY1o0AXs3ZekDdeboywquM4QhGIPbwbCnRsHGauxHMgjFUMtqz11HF4XDvao
iTT3sYaHtfweCXFFocqsRyZAYSRnO8uvDiMQNLcbDE0DIAR0tjwkgFWf/fn8HY52YF61FzsBTg0r
PdyUhsCH+GeffImKNfdUH9+Eb6DLd3bqQNS9UdC1VF4df9eMe8s/rsCdAhxSfF3wLlAtNoIyP9A8
ssffzUEUYpEB2INVzCEfCRN83VRMJKbGEeedfkICJkWCP76AIA2vf4s0zy46SEUDktEMmw1XB17D
wmIudRlkfO+JuW98rrlJu6Pgnx/EV9YZqCF3FJCdrrVhVVYQ5NG00S8ZBy9gIA2to9j0KQPVqu+X
uavfo0LfJFveXXkjkNaSEHdI3ApyXkBKwwktlvbi+ObidnX0bRcSCg6s7+KY07tWnjSKkq/S6bEZ
pqvV2yvbvoMUN2HW6kYMrHaFmBwXZng/sETXzRoV2aJSSlk7xebCx3CNSSrcMnbNTaj1au12s26O
4Fy4D/hzUFcbqwWFAPDU8QDIRN3qLBVmhsf4vivhQMhPkdm2j4lack02jB8tp8Wd8aPRY8vuWgG9
WLHj/ra2CrmsveUUJ1rFROJ+xhfcMiWSKeySWNqHb4HnX7ba4ISUv5dCvSqILpOedp6KhK7RJGWj
DoTc1ym1RdPpWGAJZn4HrE6hnbgDlV0EHLGlH6l3Z2/S9jzSz+FulHyz2PHUQQhwK99g6PbbHMBH
NFBK6MP2FQOdFRE1fYVCzJMwgXNhGknEa4PUe+zysFyxfOhU/bxKqXsg7kQPa1KQxoiiZd7UW9GO
KNIEM0YjYwYzw1PV1I2YdFBlY4jjVjztBrVnC0W1kzdNWbeiEmj6pnT+feeUhBjRG79FtsaPYtUg
p31ODdd08cSYeXh+x/iE6FNKdDST463BKVJve/53i9qo6TMMAJ/4ZaXaGzp1x4krer8VECpkjHZb
jrzQyT84iSada/Pe6nwmJmQ6gneSFqyRXSm6BL3enSo2sKA98plQhqw6dCWGH0S1UjYv2KJDGckU
lQ1Fv0ZlWYYSnvpYg6yDKNBgDCdQTD/jjVeAft6pVPa/PbzdAQN7nxb9zOeUT5LRiKVnKQRv39fb
b/oEo7AN5YVoerAe27UgSkhkaNxt1WW9CFvXCWCJ5Iw6p/Vq+CUxJcWRBXp+5kkZVyoXJH0gzhis
7F68Oh+u0LSunlXhT/zoqJ/82PV9KidrQTFIEbqk3t4IygqIi17u/PZ6d0ekXwoq1qMjYix8xee+
aZfO9xb0lOCb1JyGKq73o8w3+uC6vTzEXjLHyEkNc9vvczE77iTDq53zcGOMWn7rYxADvXxNOG93
5es8lWmXTFfsr7Inl9z+wNpdvm6EgWjFuesXfXRMKlrNhg++3RD4aZvBUdOg+OXPFUOOoiDIZgdu
3k13Ru2V+sS8s1zGVqZkt27/f9sFxn/85hgSChf4kSKXJz62GqfupWLdc/PrnxjQSKxWip05m6H6
C3TpnbTmrqgyF/hGCSueREZWDqxXQJVokpP3I2S0rn3rX26sU0nuvUuIa9vwPXo7JT7NeCzYotJF
KzTbndB/4CdFseDGoH9YQ3heTydTIhlKbyYReYGPqYNwVOFj/3RfNreB+AZs4Cz+U4atgdh6PlfT
dNfkxQjdUGl5MrFOZjKz9MEhLTB1J1bAGPZXYhnWBbACmQibZwD+GeNsZTmfNLoT5OFudB19/agt
yTNHCTKx6H1jDaCQSwNfSF9ve6R16M+wh6kK2RIpbMHH2kU3jVUZ+wm2xoXXSXBRMV+ii57w/kMv
MV06pNKRJe8IcHnAmJpUlWL5ugW9rqP+d7kCeLNvE5X5Ye/HQ3FB36TzGSuSu2aVDdrwLhEtxuFB
6SFLoWF/DkSuU+LkALGW1vP1ew3Kdvy3InwTc9CXSEtBg5z+kgj0olxkGgPIbIGFY6Hm+nQ63vF7
3p88gJ7ysjSzTJSxWsmnUDQNOEtBuDGRgqjDpxXThGH5zcGb1Jxs3mii01JYxG0b6JR012osh89s
txFdNxmB85AO6w36/QWcCnFcBp0cRjMNbfqWmQGqLIOQtEXSBczUn3hWZJ4AR747ZTn4RDsaRZ7s
bF2kG8tjszNxsITLNTaVqtbP5kLbAxpAFO4U5V1w5E6IT2+xofkzFwlka921OxrjCv4DF7N8avIc
7Zq3esFK+mBH+5PUIquOqB82qtAafsHd2rkWE2I690Px5xauko3zB/ePTbd1w5U/a7fvKP6j/kkt
khg9YLPawDJR2NcDKYtDQuJ/QUtZkEurYoGTEAMXiYGj9j7UeyDEgiOIOce46EjAx7FYZfS7POFZ
8aA1wiVEMFp8/LeDoOcmhn4aq1mhcihQYZCiWSa+LnDTnoBHDBrOjur29GBpuIQYwezfSvRR5B+b
rvbc0y/V5r90gb53qenYVQM3VgW5zV26PyDEiKLbqO6B6kx9PLmpcZ+cT+jFx4FzhzeTyBxc5j3S
WLlCywAhSseeNuAWLgzW+2lx74FKmcZrSe7IgkMpLbX/YeJ2RmPvhgjseNolXOAad+tRDOCONxzY
u3UrNhijzSC5CiZtbWufwiXF9OHxICwHJp9rxSXK8RlJDl+qk7wNd1YJG4BMT0bAEx48hpOO9Sk4
Bof1WnpLYJ09Nn8pVeJpZb32EIJFd2GJFQVpFbRsNZgb65xB08TqX1x3QnWiPWsACWZGTi3GhKZ9
i6xDmxKqwI8LYhUAbyhMBe6zhmWaKCdtHRGEuXWXFgXaI2TVPLdmcg1Uc1Mq6436ZzIEtOzMeYtp
9t/3F0qIbm7aMvSFx5AFCv0Iqezwx6xIBEIv+jPNlFdgsiEKaGSFEUYmQ82J2hrFmlmL7eHyoIcO
FJroltFSSc2InXt0aXqHvIbcY5hqt0xhJZF7hMFZK24sYyXxSo1OCr8C2F1XotLXEFBELkK6i9tD
8qsJ2UpSigOMjIIJPWMqyRarTxk7Ydecp2AjhpDHKzX8mdajqTmfdO10F8g/z1faPRH4OC3i3JzK
j/TfqS2/E3a+1YJeZcWXyB8QF6hGGxLTv9BlQcRlFBHDs55pZn6pATGYsPfLsx7NQ7y+IiCgWETU
dAHlhljwUAloRcRKDvcNVC1Vq3D32YwV9G3DMFaw7+atwMZFPeDANA9iWKemSvSAOLYt2H4DnvfJ
Mr0OSZ2WWrDTO+XsaTNJ1p+89wkSoVNmTnPxdxPr2a3KMUF/6akUexVFP8sf9j9v9D59NMXLHtcY
dsk1q7jJJmloOBq52xdq84E+VibprubTVE6km3VfU7TmQ2Hv/kbzz0rqt9yUDdrbPTKzu2jqDf+l
U36TMtnAPgv0Fj34aCcvBvHXC3JGlBauokFIGlfkmm8Od4oyxSQ8ISFH0DN4CtNEbnV7e7U2o32y
7HyW7YGLPDepQknxyxUUZN1CdWQ/WmALvaOKtJWE1mI+XN3TTA7mswF/8BUBq7dkNW7SzHFHjxoh
ikyBqe5ZHQIVP41uv8/st0aTucsTdJ9WNvzQ82uUsXLX96/zxWapbkpqiXFG3ouN4lfiUvrZYPdJ
VlVAuHJSx3+wnVtVcG6kSufXIv2iOpy1x8orkdXOW+eIY+brJUSnFzyYBVJE3oUQJ3vmaEdjeGXS
aN/ODdgcc1PsjiXEFHf6EY3UPZ+OCDdu0mmyPZq3dfCP/g7FTNpJ1foHVxaRZDtWSNRXNxqAj1PF
Os2XS7f/1DgclYc2hNkucudLmIvriQsnJffxGeObvlQB92s/1iT2njRJKJWy4T9ChxeZM7PGMvDc
na2cxYuwYe3g7FCWspPhuU5kBt6La8x5NKDpnxbXfbYUZqcvRfoIoeHXk5mxuTWBqjnCngnA9Omr
s1t5tIIlL3X8sCSNEQ7S9Qi40dchkxkuuP08tESdZ+5jM7jOiv8PSBRS3hA5Q7Dxv9D1Fp0QXtAo
wOyiXg9pSe44bS8HgkSiSQKWJQoRJ21rr2d0zMt7YSB3xwqS/AKPWdwRzUidSUchaSEXTKleCiQR
i/gGMeUtZtT9hjSAJfzSJrBqFHZNNSNvOPzaG0iutXrliMlgOQgtQJXB35an/ld14OMlrDJ43LPP
7dcfb3Agijkk+pDjiB80eZiKjYYP0UaOZFHBUOVP3NBek8vj8JGHP9rP8O6eSHTnW+/sq6KNiArh
v5ihL+cVRQX5+qqsxicxaj8zFvBl8bu/DDeLuaIc1jcFiGAvXwkpxbVfLJtvjIYibiKQSwhyOO/9
8bUUXyPPWQaa0W97FO0XFWoarRY3VH81naBmbqel4gaFUi5Tsc1I0vahqoo4DB7vx1qh2oAWsZsa
ASSZipkJOaGxYod0MSJI7UdHd/ZoG6UxfcpHiEbWPRUIqj+/7dHN01yCjCU/ffkjfL90r+tcTFTm
fpAaWIfgxeshzEbiBnP+NnwyrxbSnk/Syt+Q5uTtLaTTttBaBw57PjTRn5feXKw4VLNS05eS0tIJ
sRi7KZYvmCOswhe0kq5JOu6B40+H1JHCdif1i5InW7m/YOURDHTb93PVv1EiNvgV+nA0ypEBUZDL
EMq3ejm3zVMuYBg5pVkF7iFAkdvAGFAtYr4010UqWICtNLDuQEg2/xiL4k4z4ogoFRutVn5/RhJ+
gKqQrdcmnhN++x9IvziH2Hebe1g8mglbYC17LYBlENxy8DeFhDl3Zs4xKXH5mYUo6OYicGlEwEHj
Ww6hhz6Zc2YzmuBeolYay5MdcPrnyv4O/Zu0ytdDkNm3Zo2CIeNMtFIejrWWbvrbgSSONO/00dCP
cvslkE2DK/gJeuMT9B5ISNqL93MV7+WGqZgAT2MDnlZldCRwY4uXu8JelQapUvlkIcbZDnpWrks3
Li0bGrZCsYL7HstI5czuenG0qSpKwO75rAuK7Wo8k23wkD32vjq4VkpWkOjxCDl5eXuxc5FF0Jnk
FI8Ja3vbQjl7SPmIA8bVG86eV8O/s1bZFDpijQYTTLrFzdkImB25ljaSYkvsajiqWjaztC50bAsZ
27bYQPuFkdzx3cSqeign9l7Pt4GeWntBNdRgKkAqzNZbvq+/IkjkkOxRSqsWmrol8KSWA4mG7I1j
3s5Zv4TJPs2iUXCMkUOfYRq+NHGaw/H929e8GSraPTcxgmIglGXjnT31pSDSzgVC5j/fHL83cpPl
56RQY7J4t+gXLikBVP12JZqWZt5EoTIqD2SPKRclaqTJOm+Wx7K+Wo4DBQf2KIL08rM+fgt9NCxQ
RKiBU5eAVvO00YjaqlPz34VNcFYjCWH6uF/uYRhILus5/N1yGSRVz7+/+0H0ivRZ2WOEAZftd3sM
//yLsbLBggQAgcoTMKcTwnSGZAYMf8skMdWW2Tm/ve5Ac/86IOOGLhTIlhXD4FmwLRVn4f/z7rpY
0o0dcW+/CRF+K0kemBehgfrj3Mq8rVn4CcHyACGp9FsXha0tzZXMAUDPkkje5uYxaNjpUsDxz5Bk
kuD+TXEz0g4Syhcq0jRfeWXkO0mv89Tfq7Fa1iksySVYHlaAdB528HkMCbOteRDtyAPUta00dZjH
LbvTVNR38giWK3gKgn36BWyRhvVr5p/D+YGK229pk23syE1bArTmGcy8O3DKA9qbsloDEYEuTnvp
aNBSO7/JqvAOzrJAaVD0uo596u6okNg6yzBFatl5owZGZQjDlklHGbs2SjtTCqx1O0hJLzzULdbD
a9t5mzUWeJqFWfrbSdCGfxW69Dw7kSk7OfiCqcxKwC9fnEm5mtsMN/eFwWB3OiMWWMiUj461X6Kl
VzTPsMzdsmofgze3jpKwwIkuMHjIytF2FxK7wO/1zGi5kZ4JjWaydGD+R0NQunDN+1JKUdriDa0r
CA4vZfOv6R/5ZKvkJx2FLnGYrKuE6yFKMfMgCguZsJpUH3GZ0BdJPAcni2jqhLBRTpxY+rn0xKh1
GaSy+68HtiVnDjgPKEIYjEfh23MctfvfOFOBO7WzyMFY8DMq+0NTkyTAqe8uM1uq5RRXGG7swwsi
z72bOBw5OLbAoYU0074SMCPdAPGTskaa9kTW8SMekiB/ytn135E3/IY+vmR37svMQY/+ce6sQvEI
4KlT2daET1RsuvlXuyPd3pzQIib3MK8cPZoklS9KwiOLAPxcUxevYt+0RpGe+L+k8dqi2CIDDmcW
prrVjuoMvI43ZTDCVq9r9zXEE04Q4R+01+zu/4ZFTj4t7+YHsv9CxRlrmkSXO6aghnQrGbEk+4Xd
7ES6/cjRpQzRvl9bflaVskgxHA5K0HdIevv6NFXIYKnE5g+S8C470BBcLpC650dCP3FOmYTfhSka
8G12RBmgzweNBTPxGKT8hjEhSC/LKhEXtMJRJcKemgd5YzHNApTgJ1SsZNy8CHaxRJg7EdeEJvpn
3KwJ+5+3Bi5MBTCUKXezt3nF+WOwWgiijGMujO0PpKAgK3N3mP6nlecXpPg07USdC/tTfieqmXC1
fG6Li0eiOCcpm3SiripxRs+pQOog4eziUkLNlD/uXmaqSbOyKEBYSn175QkMN+tAVTzFUYioCpCK
deleV4DbI0DyAImTA5B+zFFJDcmUaOF9NQcBB0OrWekZsh5qRIN8vYrIZM7vdEuosiBkv6Udbbbu
Y4YxO7ywwTpo8U6ndOAD0zs4Yfo1jMPBTIIw7aYS8P2ntWygY+WdagMChobLcz10HoyKEs97frgG
aqNWkN4Bn9kI06UOmC6LMvvJHXkxVZFvAqBQytnpN5UFZBjoQsCux+YYmY1/rnOPXly4xVuIxg4t
e6KkzPeQQUNfBG605S7gKFsZ8KTC9hYegnkUWd73bZ3CN7jiOnLrweocbV52zQzXNeFQt//QyiYI
rqvJGlH+pPixVn8Apa0Y3ovkAwOoMsjvA2WiIOq4O4//PxSdSY+kU5/lb1NIshK4bqImdGLkO0fg
8NjOWd7sl0itoSdAVPz9K7zA7IiikEbpjBxIadmSl77NNeE9gvQRowit+tRvSlBbzt4aE4AYiLK2
rAXXsRfnoh1aYtpgoihrQJ4m6ITaXTADw6VI4qBLhezQKHxG+Epw0GGcAMRnIMpV5Q00tIt9W46o
Rc2BesPVFQl1GZA2kCg/O7K929ycQEs1zA6ddkanZedsUQKQcNunOYjaMA+pvuSjl4z9VNsOd2jl
8vX2zxVqYCq3o3JJU2qM2BHRAI/XsSIXofxE5HJt7g8panmLeK7f9fTon/Mhjcvr7HDUk5ErR+wb
fyCDZvzV6QP16ueqRDW2aDFzFh2H6QFkQc7E9lw4jsSSIxvpe0U4//4Q+nd1k4RPnI2IDp3H43c/
R4Ub/PUIgDEqm8NnNSHB1ZYATaxlsRmefL+ZPsz3ZFDBiIq3XY3Btr0gfERuEPp1C23q0eo+R4su
rCj4lR6+4bKCNhHYOH6P3XJ9XQN+vE4wgMvYM2YDdJErJdvRHpJj3jGjKODon+WucOWqH65COEii
QABIbsaPCvuvk6GMxjM+vSu/+qvjS+fN0uKvezqo66nJHXE/hSPYXPJ8nKYaRAjZYOhFBEG0rIwI
luz9Io2iNXyS9xBHuKwA9q13ermWykubqusCh/AP6EDTr/cb0gC1vao0fKqRgRd5QaTeDTXJlziH
a/Y3P72a7Pfc7nHeC5u704XKYGKtxvRh60KbE50dCTcSCosM1+XUU1l6vYonOLp4gvSwv30H0Uxw
Dp22sMnGDsHU/yK4jX1VNiUct44Sx/Mwemv0C8KCy6nePM+8wK8dR+lAsv5NTHfE4+NOX9JbzCnx
JP+HgQ4+ikGrEXlngvzAOR4/yfaSQuozcr8pIqXWJr0PMDmzriQL9N8FvgM4r3UMBA9TiXxTwAET
uq18g84GxZdU8003SsdWmREZ5r97mci5zVJNeYAJlWwymdCYNJX3wy1MQH1s82FR6yACo7p9qJuf
a7H7RLnkXdGFZvCTdp5cN+qc9pkSDEEaOIPRgLxcCn0FU5p14MUbBOB09AwMHk0q6NsHAZRJOLyA
L4ulLSvLPQbYTOSjaRwM0AunaLYpQXD64PUzGDL8+LE2hjymVDrNVzWDdsARZlqTGR3hZAirItFV
C/n69bakL4V0X+MRvsdXGErScdnovk5xvSaiqLBQK+70TJqWxtIsoyxJRYMKwTicgASsYpsGIkrs
chtviwNw0CNHK11oetC3GC32y4fi/NIrH19b/bi9rVqD5IwhzZR1FYDhh38BkiKQMc40Y4CQaCpc
eAU9dettT95UeQe3Fq1gj3t7GvCJGbOdOZmzzXxIu91aX1TdobsfM6hGk545XyHKGP+LR7uCdxUl
cZTy1Lywt49y1pM1YlsKyyzfZSLSpxjeS4xI1QkSk0WKJDDspFBhYyhJSXGVhs/s+zm/S7RGyCBt
Xb9SXnlKJrXEFxoHhHV8fEj/cC80xydZ1u64vKoNvXVzp9XAcMuJXkoB8GWCDufKtV93TeAQL/fS
CQJ+20Yvmiff0CSMmaIaKNrTXVQk6KkxET57OlkMLlCSGmHEBueNsNxWKPBgM/8/ZYeHkb/1N6Ba
eXlNQJ5OdIiNNUHuCPz7e5u0qOagfsj7JhuVwnt5nYT0VjQvpa5AaHRNLO1WPCHGUoI3f0R0RL4j
QGMOM9HTnPZo1sL0hYbjimHHJoClCEHrPBpZjqHyxrW2/9stCYvT6yuOip8xVaz88IGpbKU4DoWa
LPqpkk170Oopt4kQQQS6YGWuByLxo+XwVBMPHUL2gWNqFEx6/UDZ1sB8FkVksB3c8whdW1kQL1WQ
PiQMeiJN9nlWOT2KvPwzC2JPyEreq6zGvUPaF7/a+rD9BYceWo/tmh5fQ4X4mZmcogRU92WVth9G
cAbaE1kTzACe5Zg55gDPZFwQh84nYuxNt1rR/C6R1BrlPbg2Q6m94+wWjFYLE/VqbliXOlvwyu6T
wh46C6k7VYfD9dLAP4Ik2N5bfX6j5zp8/uYR0Qh1QGneCOAiGJcH6MvAUbjNnQ8oNvjBRl5W62n1
RD8UIYDVlqwR6AASPqy8fpR/aTxXIRisyf+COPZ3+f0+WQ0hi9kRhR+yspvDSB6k15HlN4HcfGac
6/Mu+vv0iZPIiDMg+yzPP5OP7tGY4PD69ocEiGIrZegq4RNoAi9mXL2Tm32OctpiDzM+KG1TufpV
0VNXi5zCfnvGkhgQsPpmB01WD7ZVc3/6MuOLU1aBiBnI7Q9FTOZkX7TssTHRYMDgpZw3ZTa1qA3s
SzYZEscMH0XpPnohLMuZhXaxxkfWCWakDeNuD0FoQS0VrroEw+cDvBxuJS4iOyws9A2Cx9d1MHa8
letHamiIMFew/uW9M1oQAc2SmAvFR9U1id5gOxfxEmyo/SRgfHZ3pV2uPKh+0uLppMnSWxs15utJ
CopXaEH0syAkNIX/ryhbYiWq0ZJonDYc4xx8FpoC5bB/Fw++LCg1Aj0ha6UAi/aLpGYHSiW7U4E7
4+QrLUL0u8nLnX0lvfGbDeFtR0tnEK9aN0QXzl1eYEARa8FyKFaMfNBcKF0L25sg9SyaGCduZ3R9
A/xhz4dQMw0k7v0Ti+3dXsJQu+j/OGtKbcgsN3qf4tqXDosAlXf87G1q9EygefhCP1FepQR7LL9o
V9cEbvTOqVetQ5NdaONjNaVif1rFn3s6Qr7mc50EG3atljZ5QgjXYnqmAgc2qKI0PCtaLrb/+M7W
aGAI4spgtWoYoEXVS9pgvaWO1f4IdhJEyYgCEH/o1+e7N2U8k1HwNAavrN6YP8X2/1vc2q6Fz/O9
qS1ZY6eGl7+wQOTRKbtAQMdWlALMbYCJAPDQWlZ1XGpcIbJGPoYwfCsT07i7XDichjEHAqc9ql0q
2IU7iAHMiav+PjspD8YHQPCckS99hI0m8bP7qHMnRDIh/1ZHYq46DqICv4eAvdiD+0+5XLnFq1+a
JkGaRfF2uVEfPeBK0UNUa5g/TIWv+D96Q+t1sKurlWMGUKfd0R8Jx52Zgj8AczehLQYzzC3oQFII
dQ62OdRPrZv52aKXp8F/kk1hRkbUreL9pJYZ0zdGeiVumlr0GPh5n8rOi2w6wiu03VAYuuFy3q1E
20waE4XpHrH1dOsjU4nrxmQ5/UVXBw5a3v1tj/AZjLmnuQA/b0SVbFMPB9nre7lMdIJSnh7h9iKv
5xpnFDypfTZo31iFrzL2JP7wk7bhdf7L65bLWCjmqA3fWmrMSgJICL7+JjazdgPbeUh3GhTZAjKj
pLFpGtrHWEQe+UbHeY6UT616sOJvD8a4ZVfcrk4p/0wIzbngF/TkK4uu9xSe/3P8sBO6cMq8TxNU
G5MwHBjCJBMEwN6qlNYFlqO8Xo4W1aZen8YulaTgXpAZGRPkOFNw/Bcv9Z9BF3ahY3jci8CHwI40
OgkglvapTKAMD2X/fSReJWYubgz71L6PTHzFtoA9JfzpMqJt+kYX806UvhRqDItXGcLPLHpkse97
x2FzhUP+n+f0rMTWmwFkcJYyfrf2c1hdV7y2ROp865iV/cXQojcD+Ha7/c7apJwmuKflRtGhbmpR
xwhYgv3PgVwBixIil4sg6M/xUH62il6njNO3rd9/NVoRVUv/Q93WFktbSL/P16O1VnU0aISzLjr2
6/GUsH80WOVEMWuUd0n0IGdpQ1NPCR0fG0NUKX3Dq0Ldwzi5Vx1QdCUVsM6LWFKEIMAITVW9kK4a
TgFFY8yTe0fz8XpXr1h4xqBwulXvqArLTCiWSssW969O/Zmv/oaA9IOsdzCf+2DM+TRwLNx0QJYS
rU1zHdiE6BSovk+XZfc5bF55i4K1HcIjGXzaMDmoDEMUjJK0zr3PmXqFjYRhJWaA3u2IFuvsHbg3
c5xlUEJgJZ5tsgk7SdZqUnTr2wuwLwU6bgS4WtQTACEjhCeXezxDUjLntDmjLKk2j0OlOTN5FMlQ
odqSRTfir1ksUV+vqYV0WAKJMzf539P4WOAZODggK2NQKN2pUuD1LaHwykAL50ehgmqUQx0WZ1YC
XKwXgmPv7JWU5az7Nd8noXoqdTuh2nvedbMimimHw043jdgX3QrkexmLLgWRdhrKpuokv0yuLhmm
D3Y9xC44UDKEBDZxNplLjnXv/txzdpFqK9vkEWjChXZ5PSrcqaxmpegk27MdbJJp6mfxMoZ3FXbH
uzNh9/hEx2XHfZf3J6dSaXodZMobJh3svk5vYRrz+HcB3T8fEbafjOOxharOTVhaWX9V0eugkwmV
uHYdZbwsdbRgge7SGF1j1d4PJdSncJh+W5PPIJN/jyJPwfKKF12/jY/KPlUQ8P5v6700RWCYkcFo
DkI1JWCQWFWZbgt5OzhnVz/mukYHa7pgu0jGcWi3GdvEv2EUkXsYX6b1IMt63huF/f1A8gINZPvV
c/urb9KKShMv4vCk9MyuNUmpsvKtbUK9CfulF+LFSTcsob7gtEdnbHfjQ8PC48j66PMNG8Eyuy3H
oqc9mZBtk15q1SuwBSM/TLFM5YzSnWA+7woPIPwNFEgekmcB8v2wh/BAqouY+3I4fyGX7ADaHIwk
myUAlURnKWyA4hPIlMlFUoRatheIYiyy7zR6GB2yd2XG+n+Ckf8FzUszzdx6eY0cXTOXP8kNVXxe
fGWZZHOe3zYbMVoz9V0sZeQ0G6w0tbz9aw5j6p9a5TJnRyqOkGmptg8KXmkVPJ7gJBPQf5TPMdoh
7SmUz2FC87r12+C5Otlk/3527nFF/SKIGtm0g7WJX/0Ngm9SEkNgRDY+qTFJfSRQaQ52L3MuL5xC
Gjq86p1P5ZMHQhHT64zIyCXJDDI1Hu345aPtzTf3ltO7c0OwW5PxFI+4KSFJRVyo2t3FoJVPGP7V
VrFzaHKki78nbvfBKphxrkvRqwCeGiA8SByySXQ4zG/rGkqAPCYdM1zlp7PRLBxAeU5TNENIirk7
JNVGHqysyWsXT3HIANwmBFkDMGwRGmoQ4jkuLIfkO3xnRlVxIEeEGuC2onKK7FttVUPo2kJCkhqc
w+sFbesZYBMVwMvi1/Ja62dbNXQsorCSYj/isAhWarftXjzzrWTguUha42BGVef6xTF+lg0srBZA
DVhEASykY/4Wx4p33jstLS5YjXjR5/QiNPy+gVrlfIkRlU3Cbo8+2FO/dW5PVpxYQyoTwC+tjae5
VfwVKNDH8Js4MVrb1cCIHrzG0fotAMaaw7n4MSrUWxoQaCb0G6PXCMDbGmJCvpBYrBPrGC8aU6EG
y+3nIemOCAXE4uTlFBhkw9+TfUdSjSTZBuTpnBTJDCNVqSL/1p57tArMYBc0vtJe3GaOwctVz70Q
ZWuPQpSUVeLL2caGiTxFr7npfHM26ot4fAHz+HIm2g2o9u3iCBMwAyKRHFeOk46asH6T/DrEYrYX
OJMh6mFs79Yh4OCNtyO4Lw0be3/xNj0PuIaJA3e231H+W194TCzyCA0/2v0qN4qmuJIxrG/bLIxh
QjsnZaC1FO09KfyXwridmDaqDB2Bkya114HyVo7YixCXGY3dnlI/VZc1i/l/5xymRVYRYt2hEnta
Oov5cN+GIvaHH7J9RjekLQ0c7UVI7H1DmAnmos7T7AUGLOc7XVY4diu4DuEw1lkXpu0mwzGZZWB4
MhVwehyrBCCtlTC+MpFNSHxg7UIfm9DQc4HKc9nTqEZKOvxJnap+1DWFrFfAuSHagbI8E8fa+4YT
J4xK9MWAK+nXzO5ygwuWsRV6s7/Xnqd1WlvxMf0DLBo4FnQW/w0xGbzsuBIqkg1rDD/u3IxepqJL
QMx2hwhv4mEG12AMyiOme2SHMuJfYA91k2V4P0aMOjC5R58rsYGJdnSkQF0uPk/Ic/j7Jlv4KzgT
GM//IpKZ+Ozc+yi55MJfJB5vo4YoSt4otjBTgBwNhADy6B83aviJdsdxiilDrP8LXmRxocx6xDcY
7Cllxye+ogLYkgMan/XiQp6ItvoeibXZzHicvdAbD06TKSE76nbaIgN6BfpJnbDYFV+HvLvEl4DB
8I7eqswwRmjntVAt+bXFTi91qBSoV7r3mCMnWKQ+nedFD1ZNS9e3fTpU8Sj+xqVPNBpryvSDM/0w
yyPmv6SfzY/HOn0Zxi/R64uum+0mXk/5rW8eSFLt5Vkh0PFRFinzPn8sNSUQgYrmoFWv/p7bCvg/
GBG8g9+sjMlIzPvOHQwFX3YV9VHVSzkBfbiWHE29qwIToaUmN3SNaSG/24QVdG4Pe4YngQkeyFFa
I/MIjGqHKiWQHbTuLjNDZtzWgydhX83RY4t5hzHRg0mdh6t+rQsptYg3UqYlUg3HDw8Qs0fWKN0U
EEtDQJ695oaydhTDmWdZ2KKFUwsv16+Q4l2+MEreL2IuyhuA47ML411D1T1OMxwFFMs5uQGfF6DV
drUkXqagejGF9E4cjnKzE9Qa8exECQXECFXMEsEL7pIQDVuGqpUuKYKdzg9lFp/wodZWXS+Xhcs6
pmfeiYYx/NALWOeymROZdCj9T/hPk7vRGNiaBjBe1mGUFXlrVoszfVCw/j2ZJ20R2G4m6QsULR1t
HRQ/bYC0WMVWVmiI8htkemnNZ9QeQmf2whhpt38lrfihw6zGyxO+0u8u0FIn5OpXoDwSO+ExaYmj
X9EG8oSzsv0D1i7vxKSo9l9XmccpaXZudD4oxyROw8wuxa68IQVNXL57L6MFNC1o83majBrYRgKW
uxjuS+R0IqLrxRbloLYnMWqFByyKbqAJCTF+DLRxujAxQHDdQ4RiHsYs7ylm6G7nDuuLXckvadKH
zDPQIW//z0xmd+pbHclqSK46XwG4EXK27ANjJqq9auGglV8gtr0B9+TdS43Cx79pqMSQQNVi8FgD
4ekpDC65Cf7EGO51yxq+n0ALbzZqZqAl5Q3eH0ar0/5wRS1QJqFkKxvNv8Zo8gbvM+hzHUJQRqYA
qENnL2ohoQRzB91oAMAyrzJEDxO8o9Rsqc88xKguBIr7SpaUz4QBbH0MlY9HL7NhrqKv+WIcFotz
XjkSqwwg2Jks3ZdLBIvv5AS1KfLZ3j5sO+DOgkQVEAdySO1TwC7KfdmR0PLNNeqq2buTxTD525g3
RXvg1e+vRfWp4/Z82YTzh9bdSFimYkk5FXcrGGAGnNUzNWno+fQEsBbkEqz7+r0DMAUKSN2LA6ks
ub/BrPNB3oKRMuS4Q55mZ7CKWDm/04vBXCBUw0KMun2sLEct/pqOmBGAFcdvltNd9A7he+UyRaC0
AQ9Nru0Wtt5VTmYprL3RM/cpAQPkHhrm2bXDPkDPmXweywi0SAQcgDeA6HAA9iG5jrQsP7mFup6s
GyGsiiIYZiG+exIkUlPWOjo1e08C7OBeYxrLYhICShdaVnes773aW+BtG234nQWpf1OAQqGXywhP
2EJpk4VJO25Hs4Ywh6rJ7xmgFfTKYLKFNUSsb1JWyVOO+6hE1xYsoqCUGd7YYcf7Y7cUI4mXMN0i
1cgx/UwxOlIC40yFFid1pOG9nPaShawt7aR9uVJ/pCPOfJVedh+IXCS5e241crv3OrWp6zX4QgFq
COOBXxxeDB/bzkjI4RLr6qegoZMrK79KBXJnVIIKXHFUKVi5I4RHO0bqXnZS3r71Oz7h0EHcCFBP
y29h0XiCaC5FnWZl02kWsLKaV1qwwM0cBd4s+rqURVp9g5XAypQhVz4jNkEb2Dnw7KAIFYg8uhVU
Tk4YkOQghTBOxlEJ8ST2Vw5a/kjTUS/+4viLpasxqtVrm+SoD6eN0Ol6QfOow6nvJQKRWeVzWZGU
eLuU9mDJJTEKGycd/i0Jte1n770l9BJPB/+guchrehuUHkBL7E2ENIwSGVh8ze4/++LU9KUKbzEk
dSjP7nPhxeMFjN4vB9NV4y/5oH9j3yUlAug4mKitrCWgsmSbRZaTZncRWWapEOkqGojfobQLsaad
+YQtQtp1/BgOjf5WMZbmBfPFdyd9t3F0LAIrr+xRiM7WEzD03RQDd8qyNGYZ2m+XFYchdUHcrxPw
mh0ze1V/d0VVBm1ONIDPo2Lknfw3RCVg2B5QXNV05gae07WzY9aetAIwsCp0QRvCY1xjIP5HsY2x
Oe8qh/Tda3y4OpBMvMTPvSxCyYHxdaW0uavZv1OCXM7oFkNzjcEPerErv8dGwtSZrL91YUk4wuZf
Cb2KxAlkJqIiLD9QIfexhWtHT4yWVGKUBj0616U6b9njNQVFXexRWZ1Is+bHgVh08fnmYl7XyGKd
uXoitF8jRAfRbd8oc1pTJN/2G3uIOT7cwZhYEc7KDyJV4VGIfD55O9SZEo7ZmTtDN7um41umNf1V
vMVq/y9a4afkcgkwilDtneYjtmn7s737bjBOXWkOFwJ6rVkRaPOa9Uu7urn8nr5wAOtQYLWzBo3g
f4+lic9lNZavBPWyYIX62EUzr2aFyR705Xj8JsMAxFeRYduqUashk1fPf1J3mLqgHovBGU6pe5U2
TC03ZMZSpdE/QI9xG75q+75XpXDPVKV1aDfsJfkY6B1AIUNxF2gMcuSYmRk1QPt1jpgu9JronA1g
hkxeogjOV4DH0nBhcEQgZYo+oEmBL+us4iFhgiQB44ME46J95Kc1KpnrRpklGIv2v8n5L99nyQAq
SDIIDxKb2I5+s+T9uKfy0NesfkfZu3v6bzsq+TR1wpZ0pTtaSV4hYCGNK7oaPps62GTrrIrgx7x8
g4Qvynuj2V94999O0VxSGeyOC1N/QUk0lg1o+Ecuu3+6+xTrL5xC8C1o1MO7/RAhSnKDmqGviTod
QyUctpUi3gfdN+6Z6MUBlM7Xb7NIgH5eRumPBPp7wr5oh8JeUDjqNY1QxPy4O/EoL5aaPqCxyvl5
h0UitZQs+vm/bSUAVti1NKECjv0ViSyvVvEQ3stWLlbl3mT4xqsaCHAAG25wNTi4e+pBPiVhD3ja
LjqAC4ve9YtELj2sTm37J3165RPginHb7UKMx79zBdF6hhw/STLHy1+CSH24GtNLnr9fZnKFobfw
tsSejJ7GCL1ezaF+h85HJu01WRdCWP6nY4wxs9Xm1K+B+GyNAUJunz06ufIAF25HGQfO8lhLQUSd
inAtuBMvh9Aj7kQkY5jHadFCieUfN9oKr79rqarhCLGFbXpS6TnjFKnNIT0vY/DA1/SRlsVuv9OM
Aact4Ao1Ygw4sW0sNuVQCt0HEHDKy+cKb/HnoxWqx/ptoIGfO4NkFHMxBav3QofeLlGr/7bUKT6G
5NiYkXpCU+ASamzWTTCBK+HxFG6uIvM3a3vT3e6uM3h6LGhfKblI/aKip7/RmRuO3ykML7WjSbni
NLlNtlob69WolUFBmMRDDIdEGHGS1Xe353UD6z9iG/slT7P54b/4gqZ0FME8T/R0VAtPUpcd1T6g
jCQqECIGPDVtgU4b8jnHtv48FgXC+KABaC513kM5m64847A76lsjGylVhVNLnFANJcLG80RvKZXX
f1/a1GmkbBSknX35skATsvsvA5U9aRLLdVybaWTbYzzSlkD7tJeQcXITA6U/Ny5Z0X/sek3uIXDK
m4JWf0Di9pK9/h4LrzKVUwO58/PnOQkOq9PuWO9HJ3xG38Yft9S7Q6twZglEfIGRMBHrPbiDIMv9
2jAHpmJUtXnuF66JfW3Cw4261I2nIIQUW0KnX7cew1PY9fRnNpAhEamITyYBZyVVMTq6sXHJ1WuO
qYBgxcDCGdEWykkN9yvxv9VCZbIbkd++g7bZiEfjViokpfajOnt89v4iSsEsic5OQsRJqrhwbPNZ
1TMBviw72DuMQg1+Kao2UszX2guNCG8DkRdpAkQ+ky4SRUnn9hU1VVRlCYeaXSlCNLB4cnwBJT71
HkIU0XUFIvIaOLmAc7kXHiUTwjnXHCBw4cp4FfH0X2fAPXarQRwjjcjJ8u3jYMl0tmur8C/Bvoy3
aw2kyLOFglB6zMnIIXco1KFPONpjsMw1wN0vS0F3wdtbxwux1r99FZDvHyFMF6bHPFgm9RWJj29X
Z/1pow3GzvwQcodpd8Pjj85lTrqOnn0ZDt0grejoTBpZws+ExVHebSUlfmpTgwyn5UJEs4F2JYCG
1tYGo+pSl3+xxOSb1x8+XXm7lMLpadRBWI4HzXtmWuUYoH+JW4E/6bDYHzUSEOH0/32SsNHck0Ey
9sBpeK5Gk/4DGTYGCV2TUqPdVD9gAQfuOHHlcdS5oAQax+GpMS+xJ5BcfayrsAIdCk36FuNr2phS
I2sMUBkSx60qpiYAnqDe/ki7oHkUpubundOGVWkCddTTkU8xEcsEFgh1FHPeAWaXCtqUGfszti6D
XwaP+WXgbln/slOes0eqyqflJi4ESz6FLkg1HWZIcBmYiRS9I2ePhyxBhN5rUFkcA1TokgforIjd
oiB0Bl6CmZRsw3wg7IO11TyFfnLhJh31fJmLPgfpJ4o4FD+mxP16AYixqp/WCqgfKIxrKHO7P8Mw
QBO8ylEWmLGp4M3COWnBSTlsoDveWCvYj5hSIq9rKm/QA7N4TI/T6wsRy7q4uuPsZCu/awiaLbaa
AIthERixB+18xt5449572k9DWIhH1bg2T/hp7KZe+qyuKcEZQ5lDcb3EMqG346XVgx92KS0K8WrT
4mVPpBFKahWPVWHVJWAExzdGuQpgDwQZyIF6Jw7bEAKWYDvYOGX32yUUQiRFwiMryI/rWq9bdSSd
szCJ1g6/0Ht7DBWTI+w7XuGtOvmKQEj2BQ9m8FM3CCbAUXC+hlSfnAVc7BBYxOwOUeu2jXCMr+RN
l68cyXL7PR+4KmVOPKVTueSdwER7wj1GbwVILFOP44JKBGi4m+dp/4ECheNIKMW+NvetW0FtEIDM
UlfhjiuT7wKYdee7BK716stFAdzOacViwb6VwU+zJbY5cULSM1DFpr6dLfstac2rOyXtK1VA1yFy
tq3Nu3aSNlYRmc5KNq/OBMnZgh5EfL0Ekueir5XDVlxw++a2Vv1sS2S23TNJY4/yEpKoCACg49tB
h/Ly83amUXXv8WL9HObuse7dFnGde8R0hFrPVVD1SmHahR6FuiPRkMIZuQdTHZZYIsd71+WbDVDG
Y4C0REdDUdTNvBZhruuxt5FyxSi33OP7k9cai/+msRKvAcVx6/qmCUoPjnX2qlh6kwh15Xi/OJpt
aGnyM/rcJfCP5UX9leLfXkfansAXODpYvZRAh5BEE62sqp+b6ov/zhjw+7BLs3tuoJdqIoPkzu+t
QqtppY9rWB2zEGEDpixMvIkw5tZ4ak9b/akuLigtttk43mo+1Qs8q0aRJnf0jA09hQZNZmH+RlLp
YgrQNTEBCGtRwUwkicPD80UYB2TjFBa8J1rV9HCPuCRvRb1FThedclNThm0788ZUi8anyQBd489L
RBVfIImZU2+78OgoJbh8vawWA/p4lsBaGDqfVJQMmqSBfk4Nb4jf1YZCN7UT6HCSA75v1NjEqi3S
pLW70Ytj2gwy4R4/hhk+HglE3AznWr4JZmzTS4mS5xtZfPkpek4B2eHXpUf492CmgC49bLCR1dEM
+9pWB0kyB9hS/VRKkdLeF0l0/qSn2Nx0yJ6yhDIVDGOdL/ItBdB6tt7SWhRG2pm/hjHzC4nXPGIs
81zMgywD/tOrHpQQEO9RKpeBPSO+hVhIemtedmL8HXpQQy6bYIgi5vStHgJm1lupVCGlBlgcrDO7
uk0oT0VxPuMlZsvl3fGm1yvoSXECp0sfRvZIovwo/djWFsVsTtyW4vGfpalNCNx67rXsDbYC1VxQ
vFU9g94v2qhC9fA22t6NyEtFT8TfHCumVshJNJKOd7jpA5tXz8dM4rxGt176w9c4uudN/PuC8L6T
9eYv7Llpq2Pj4yHu5Cve1hSTpxeCtip9cc4hpgK13CS2cTVZfyeYOZ2W4sndPuHn8FFsWk4Exc9y
o4oF+NmIBf1p5DVfurhqgNyS60rUg6m+IWLUyk1Jl7s+/NsjIhTTETFV1gS4lDmW/dic+52d20Dg
H7xGNnGZE/JWNkVJMukN7De1wtgiGLBtpuiOj8OA9RDasLaFI1LuXU4gogVu1dHoymf8duo725GB
yfldJSR3T0pafveOfQZf7GnAKKy4tPdAbsFBNOXLASwrynQdYi0ofUsOW5aFBLgP+n1klHFObWo1
/nF5Wxji3tldz0+649ExRBREtGRhK7E9Tr7zgW6N435xVemOqX9hw2Wp/r4yLntgHk3UbennqVve
tNPqFMlT1HIo+5wnZfRqMXBMyYodNuSI0hpJ7l1araW42PI7832xNCT2dGXSnj5ui188JkBjGrHo
NORGs5AprE22auo3zvdE+TkQL1335OtDl6IUoc8uBWT1SvsCe5rwhi1wWYyj3QXXnNyfjJP4y4I3
xLtenW8vNYFI8c/35vuR77HhTBJdUvBn1h5rH7kUQMVkqQhL5beo/y6lhF945jtphQqObXEfKYcM
xWhTJqe5YjF80lXBzvw61nu9/h11s87yfQ1KlqNMAAaSUzy/0NKe8dbHjdhymhez+LyqpYm9R5SD
8OfEIrD5nb5UDzgM+yA2X2ej1B2/FDniXasZlpP3ZbIWF7PcdNzPyT494gKdOpHNliUf1paByoqI
pr04y6KawMWwI7TtAY0ozsa/fiFaUYsbIPzuzCpGb0aEX7Z2sM+gMH5vMGnTxaUBhwXElt810g58
RoIrlL96GOqmhihogY+CJ0TH/EPTtdNTOugWTJAXn7xuzNcL8vH7vzOAJNWkOi/8iA7oZ+OGgzRT
Cn+KALsVW3uvNi3CXwNoUCdfyDB+IN0hAfmDz7t9hi9sLJftAfUldAJ/WBYsJZfU5MHflf1FDWZi
ePIpklzYNq/CI8EowDLHzO8gpahvLvmv87OieG6FVk1UHnPMSx9Wvzg5p5JmlLMgjpIoAJfB/A0q
r0BDPRfa8NpKlp97k39uGJmEKp1CeZCE5B1x7wC7A4S98ZRkM9jq2UWtzjntZxkT2mv8kXkFbE9U
jsCJxivx9SlWaVEL6lTYgZ/HIXXgvv01sZgWdZ8lt2+0x5x0eXNAWtWKvTszQwF8nt16OKS5wEOv
WEQlclKT3K9Z2HAqzkJSUelUNbyAm/p5vHXVSdNeZh0G9CQTdFMiEGrYc2ornl7xZ5TRJAIPwtcD
dGXVCg5X8USUQKbd4z0tlp9OnK4I+0zMnqk/2n7EkS/LE36PcaObk5EBhKECvKscksGXCqYeEssN
RXE3J5+VrQ9L6dsTuBslS7ZElSR1GNwgTmITTZwmsgIMQmjRoAQsiXSicqPGoItnjzMliiDaMenM
xEhte2TCGkGn+jIxPH+Ydaf7SWFtGlUQlaS3t/g65uUFGMq5GV5IA1soNal2lEks8V0ZR6kW3IYH
Mcs5rkeyNInoKlerNO/3Fd2PJMPEVkcau3cYTZBixWyT2soG/kU3gfeA1oY29nAB5ZD93g0pkOnq
xfPBEyMJHk6TE8hxmDjTpe9DabdIt31jTE6kvOQHHw54yAAMB1HTCXgcQVi9J/EigZ8orUcXbMbS
avCYQaRwJp+/yzwtlPWgtO/RqL+uQbjZ2P1m9MGFV76cE7la56MrPsOklYqS0TdklNL05WYRItz6
9qcJcMuKBb97jGajlIUF8RGPwdBFIAnd1C4fDaIvLnwy6LKkrClsaPOit2jQSOR0TN/kA8w73eAw
Z1PghhglT1SSCR6j+JH5uPjRdnG52V8yH6Usju5peMNxoghsYQq+gkBShKbiFE83zwiOwRdDGlOU
hoMZd64f8BWSKBuGYpOjyd0llAzRooYXdfn19h/1wCaIzCgoWZpMQkTtGc2sNs0ihM6rruAmNSXI
Q6mR8tH1ja4viyDK4kD0umuGp0tFOa3qEAjzme/npjMrzi5w0qqXtry6pPksTOrm+Eld708sBgqo
t6j/Df9q8JxCx2gOmt6Y16Nnu0RgcvJyBZU7eCSVQuzEKCXNhQIl85XNGp1Cp1FsGReVHp4wi9+I
kI1DggxfJ9JgIzsrSczSff/XhoIX62ZPT1uRqelRt3BJv3rKu0rfOfHOamnfJDXshjvlAf73/qO5
syskynANHkd3C/w/VcTh6623UJzJDMXGfWOVMLwQQ+ZoQfEQb/rUlVch5kL9IFjbjpjL5FB+b8dK
NQPSeIdnQpUt2m6ivvmkzTHt9lmIrZ327RqUPtTOVVqESTZ2YNyAju9MS5+6MrR0VQMK5oLNgwTH
74Cg2NHxoTlLYAEjAJOgbO3hi/kPTBC967H7yNL9o7JbSs8uNf3Od9blcSYUKzRg/F2wfwuRKNhk
38gOvsDsatgSLr2t93lywVnRKX0vnSARlBZhBPbLNvl6y79JjuYilomilWQw5ZXHdzLLhMIdU20G
DUiyylUtijV4lXEzO2jjKT6cQUbPMvoO5luVnzIIgdUWRJkNMTs9etMAtgRav3Gl8Td9xAAcRGSx
owbRhdFoYQ4jWAHRl7zmYPsMh3BYA2bsCFT2lV4JoFzwMtFVgrauHShwXIOzmoC/kBsTnTRDN3xW
IyU/B94a3mfQhxbivjcm4WaLtba+57ZjOOmmRnRz4n6P2o4/gha7lIs2sBVZ7cuANGTz10HV1D4c
F6sE6WGXzvLRmX6jsP7SlSSR/O30fCUh0JPRsDHLgiK3cT6o9bCpHDgjQv6TDv5btuGFjm+GMz17
5JVP8UTstR5/ewAdwqueLNOAJQCGarQVnT0iQM4g8CKy/60gVIKjF1VKqKBRr0/xWNBjxC+NaqYm
mcVnuve9PPkxU2Bbg9lfbIODivwNIvQEXOK8IG/V2Bcsjy1NA15+d/r9r7Tfm2E3FNT9M0ZJ3e6S
k/vIi03wYNuJNwbRO0o8KqKxa4sJ4Tml8GLz0A7fUiayaScv0wCR7lpmarrptYcetESKUTGRCfe5
zLszEWGy2Eniln2mUMU2eONCi6oWDYTqbJkMXHR5wYeU+37si4jUVcHspsNwUSqf8MYGMu4y3V1K
vCdRPjWEjQPq3Y52f/TBIobXAKjuCOU9kIa1rF8ajwd4RA29Aqj9ko/O8OAx47neIq8S7sRshZTb
fL2YBTjqSvh/tETdNxa5VDS0ShiNbhRQF/TGbWVTox72QHXC01VfsfLef0C7jaUqXth1FsOE+PWx
VwbnzNmIJjsLPJ2eympFSJkRK3zFq4M1sPI07nwjBh02/2RJhxNNC4GSZV47xj1oU6JCfcdn/26F
PF7WccuEkbf4m4tZTxFK5qER1oi4XgG6gdTTGGdzrr7G0qPcZoe97HXvjK9OPzTr3AS/qGXxxfhd
Q21aNNVMydx9AjxLWNDeRg4IQkcqaW2tVnPG7TkndI4RRDktLCSHE+qtl0eMZ+t9NkeO6vKOijvh
/401MuaXWnv9Xm18hu3pKCjFLN7a5+lBvJuZFo/+V4mjv5Jqe4pyveCvoTgz09GVOyOiwYMQDUT7
4uemZtzjvvWGybbtQIQTVPN6pKsy0l6mg2ZfBTaXxZHBu1O5OqGwIPZ9IQEbJ5gAS49aFTPyBsER
KMXZ317PG/4G92GJwCuYuOXO69qhdMl1cO9UBY931Z2GnvRVQr7JLb+XTMSt8z4dNyjcOkB1PL2x
PyJWU53DW6UPuQc/8ElHsVvEWWitbu1hwXrTOQa4NpTKVde2QG+EpyzMJSrUWZMGsPAPh6LWAm5H
DVIZRo/BsWoKGuTa6ldcnsnRw56IOjfvFk2+l7z3Y9fNriBhcUKDaZdrbfecLy1JmGzn3++ZMu8H
KbsdwTxSoSWIh1bV850tk+IrdW5p8PiO6ii843WzFPTON7DoVD/TI5bGdWW/8oSFJ6Sy9WUAaw2X
HVd/XzB8RnLTee0cJvuSYU67taO0COaayuABoN+GMSXaFPGxH7DS2tSTipaXK1G6+EyrMrh6o/LV
S/JDcsaKVrV6TELdu5+Hf9tpP+pV9YbUt/CBsX6T/ZoZCxYrUR9PRFyOs7+hvirK4T09Gp58ZvbD
u/j/vK55JPg2YIrmCdCNUnz5AXd6zT3Mc3IvpurVI6Z2gDJ0sxXAStWflDdXvnN3PV5ESRc8rdI6
XyUr8Yp4pEyi7O1ao2xpoOdjugtGbDMpdl4I/4z64yft/PF5+8M+Hu4IvVikk7y3Kcr+hkJIxMWg
PBFVLq8AjDI2Kgw3wNX6j/m9fCDbcFsEN/1Qb/02FwOBfsKCjbRkpEpxMvTYxk864w6gHgfKLkV8
1uf5rfzBwxCSvm9I5vfV5wTacBaUDx1BsrcuSmbjGlxcnupLYy2j3Xv/yVzIOePdPe/fJ7NKs5Sh
4DfTm6jS7AHjs2uLgRRSPx0pVwBj8rJiYpUpT7hPvaDOATuA+hAvJq6iWDFQHOrecCdKelTkZJrm
G87+J0OdlUzrswgMEdRS7guSMWSO07yB6BnZWorcSBn83ASXsTZUCB1ogbDOuVKs+4+XPz8ALrL+
XUYvHBXAE5KTMrAqTHheQS6ze5B1uGiBCMMG3Eb+IAJbQuWPRlM8fi7N0V8O+xtJeMw8h4gzlIJr
nKDSeNvuZnSiaUoe+V6GxYMYKN+rX7LILDnNKT2RebmxnxFhy3e+NynFhPFpdY5JXyrY9fW6l5sH
xOtc+9QlcPH6gAJ25QtqpwVk60wgSWw19PZIyntLJsbJcfBJmiP0COto5QotEAjw6qwPos9/cnKx
1McqozkUd+O4tMPlPvqZx7lbBA5oQuLuDuN/w4yVAvEntQRMAmZbEktjY5GBGy3726QJF51EW+af
uWqDLwR0dO0Wi+cazNlJI9j/wxzUllCH6198545HTvW/ZBiJ+WGHiTNCOLMlGZ4YvweIoeixiNuY
AEZxWfjl3y5UBMAgzfuxtDHDhZJoTdZnVFSZUV1nNLdeRFtqeXYtCJElXr/1juzeJ21ADFGM4e31
71WR70olaNar9IdHtdq47CmaGmh/Djjg/iaZ9u5y4a/jHU1SSnqCfCuPpZLulLim6fPUsUSxJTKR
IoHOZbspZAQQOYI0xXrEgWHq68P2Zr1DysbfWGbo6CxiEA6Zw3ZBgit001ykH43+y7RpCnHSkPPn
5NwPnm9ZF3i4soKlTMBIcCAi+u5y2w2qgtMoise/w9aSnGJmtcx5ATREUD0STpERoaSM/bGIAho3
aU7w7RKaR9FaFTfo1iUN4V/HNia5NI9aLWoRhAjqnOr2yCX8gU1U+0VRTjhWnX2Y5veh9CspuzP/
UOQzTARPcHXrsuUgOt9OOX17z34MMwtZHZ8u6omGkMPCscRyQDX69Zfrn9Q9DEu1p9q38PiQR+hr
TE/OvyT41FEipCk4R6ksxZU90nIpoSuAWILNGHW+FhpJTivH6jnP9gKv1P8S6BbvxLsAAh6y7qMB
pkX0zhMAHnM33WgAxxmvKWtBGRcPfknlBRDX3T+XTnMRN9omNgsoiZVjsgQLFsifSQ696kLONQW2
anGUsz7WjBiudsQR0WdhZMBlzy6lVVpgm7Gu+NnF3Qztp3mH7NJKRQlwpSMZWpvHJqwwfcR53EUl
eW0+sTT1EGX8hO/mQQ9h+J7OhW8msmCf/ZjwjVXcoPMGevS2sl2R9KQl/0JzvJHeC4ccTbURGB1j
hSMhQvXh5u1I/zFrezlpX6/6+i87pvUnLMx/NB8huOu57LKl8s54Ni94jX0V1C8MnRGlutnC/uTd
rZ9IWLWOhnTrvQNiFS1Zxb0VM7tiGF23wnTyVLM64ziNPE7Pd/ZCvbhmBG27P3uaO6y0vBF6jQYv
tLX/tFNNcbbewj/nB3oRgTx1U/brjhOYQkH+RuDZ9yCHplO1zufGkoewIR60MQnvLAIphMWcZR2e
9EDmQT8eLfDA2S7W1VPlwE1uKn+7m8KQaEpGz1zu3nDqMfXSGnNcIYbCi94PjxEecZspXzIpTwOQ
37ZbaCK64AIPvlulv9v1KA2jWV3EWcPNEsnO7AEEdSqA2l6IyyKVQCrPyCEQL1VFKVghb56UQ/y0
Icbib0Dtydk6alWQ2R5vba7hurZ57U23HpYgLvj/Xd468IFZCnHWZe447Uo2YXFNdpl0DFsp9RAC
rqTivA+TS0YIbgqNSmwzlcAtS6wMcq68AUCvKPe5LnjmwaPE5tB46KTE3BM/WrcK1ufSe7ETWe64
ZnytdS3Pn0Y24Aximp7BFsmj+uEC8wznjdwFClu1GwUtMPYrD6x/xUowuhOTq3D+IF6wnSHd4Bkf
MjHr46PMb+OtP85BWr7I3lX7YUFF1enTarIoASWKIE9pX8L5oE/efpe6Wgd+P5IPl5bafKacS9UL
3LutWJ4yN5eomqJhE69hVWH3RYIbx2VO8k9/j69c2XfmCzXgeii9+lCUxUXDg9dfWpK0NRxioX/S
ezoh716tA3omCI4xGOSpouMECOIEbesObzH0PqHovIT6KC6b/8O/wndmlbZxtDPaHM3nwPjX6qum
xSSmcxGHWpuvceyEoR7+Lwi9I7PGZYO3UWy5ZaRhEAev+0U6xNvCiwuPx121dOtsKOCNNdGlw7lJ
YTRtUauNSv/B0tSmTlloMgK0rSR6pho/377LGBAVTgil3EUE4mrboo6ZtE9ZArlJ8d7rQOvZ7QPC
b3b6Pgs49g4HLSz8RA/G3frAeuF4x4U9khA9Bxp/LymhnWKDJVdi2KNjE7sKketFYSIMa3xatlKn
6QtnB25gatJ+vpSs7PsvAysLPZsEOXsD9HKVPUQ8IWAtWiDmhLxt/0w7Z7D1F1qvEZGurTSKb3+E
8oWkDrN9mE6T/s0uwM4X7MxSkmiYm3x/Pk/8nU3uMBD49DCv57Ed0+uyPEK7h39onAZopsRns+zF
0ctbuhPZR4bp78o6oZR4cCfnH+KXJ2KaEnoI/cqICQ8aG2Op1He5kIEGvx+u/IDtChZheolH2u7v
1/s2izUFH8/9XrHrb0HId9o43EuL/a3z1WJ3GexNrZvZjok6+mYJLjU8kr+S68dQE/stn0qD42Io
ST+3xqI2baCWNWkd/FQuQnOA1AR1HEVWxe0W47abCnYcT4Iv061rOFAXtg83Wn3JPiLAA1AWwyXf
nV2ls9D6IrtT6HuNWe4W3DatPRKfe+f6f+v7MpSyGdlDSVAlyHkCKL/5qvALPAAF0OLXY+7qnmzb
eh1ToU+cXy2+kk5EbbVXWKoeeMeS/Ve7WgOKIrFAro1ss49qwgo2ltWtlMgu56pZfUrtcjzRmYG4
rwg275prGWouJpWL2meFzVyBEZe8Ll50bECMXcv1kp2NVPyPPN2ledq2denkz0WYmf8iVgKT+VHq
ryyfnyrlIi4lR6hy9Cnb0d7GGjA6U5YwgVrS1zGuspWm43ruBicPkmHtJhIoSGfpGowad8xWxIYX
xhhVXOkwCOCsMMn4zQ4cbVSPIjgABfBFG81up2SZE7jvcSBeyUZeJJfpArQ21uFibm+KpIVYY/e7
DfUlfZmU2lNLj31TURiXYyAl/mppnebN66NiHLql+eU3bhoavzfaHk/ehiqFNZAz9tcdo8FTqFrP
XaKddTIjcGrfjkemeY1TLl8vtM4XNB/uLaAYpTm8oPBMOWzfc8UDtP7dInow2FjW4rEvQarOHACp
IgZjRZPYnjeDwhH5AoPA15hdpL6RaPefabOjkzLprahdWgIMXO67KtUkNhAXnzGa7W/vsA/Qyaa2
vtPrKUrY4xspMXE2NJv4Pr/FXOWt6WfojxMbodNs7qdFcr0MYlnm/MLgD7DIO+gSrf+03/mevDcb
fkBlJJqgbQ/oi4zegYwGlpPZnQFBtZSKHAar6jw8AhLm7l0MqjwVNtMhOLNbycqDreG/VUy9TGZ+
HGPBNuh1oQuvZFd/T10hQGFyc1mkHU0ToBkQPHcH49BmUsVUHqcHfBRhRdoivvTIXeJRsOWmzxqN
/5ry3Px6KEOXHQnhDdtsoPPlVLSVXPek0nTKI/tzxIu1htoUh8rwEgni+nV+/ZNkHgcuPiLnowM5
c30/iuJA1+kGGSQL12JA+DYspE4BV78LoxrTL5Tk5wbxjQVSmRdkPGKiPH9A59KBfhwsMkNXQSJb
PsWvksX7kgekgaAuVJlMZqxX3+jrtQSDCSIkSIkTxuH3o8E6wBHjpyjwU+TI7ip8JMNdJET+PKaZ
6FKithjRMxnPwwOXNnDr1jf8bvzlkuG+zDLe2CV6ulTnYx7K1EmEFuRPH+dlD9zC7KaCaIgcNJeE
ADVAyGBBITrY0qR7xcgOrDo6h1ikz7lRhP9x95JBIn9zDSBhwLMb9X9D8zn0DCWqVrtCUjxMwvcI
0QtS0jycdauCRxdS11c2pEap5Ve/sEwlgy/18E+32sHOC32nlDhRvuL4aoYIDN0Cemx3s7KdlNCs
aqML/2eCtRZvd6KV7jRh5Mz5Fdxe2Zcpfs2QAIpkOz9oSQiytC0bpGgMGJPrlvqJ1bpp5rP5UHQt
8g2Etw5ftqNNHsduMW7jGOIa6P0AOkv5dvQeEYTdfNWpH3sL5PiZtA1AzB7YyAwFxema3Z92IJww
GZTYe7lKT0wEVzr1Fs9o5ESDL2zIVA8mu+oWRBRjXRzCUlMB+vdeksWoX1LQQkc6BsgiGN1tUMRm
EUBJDMW4JYC+/ny0vQaIz1IS5g4BIiaLaix2fhszFuUWo87bo6ABmQiCLpv/+2qsrzAJGC8PlIeT
w3rOpaIL26xT3XXOnZkw+1pwNRECpQ5Pe2l0uEqMjl3Bt4D4yAlbVw1fAsqK8dXoFUA1FHC18T9V
F3sq2NqJ1wUklr0ut7rHxlN+rEG4UgRoy0bPERgJ+/QKZwpmw3qt55ZN/JA21ydmZDGfKPHz0ffi
1LyFbrL4ln+2mK36zNyXNprqy6EF05WQV84Qszjl93NbC8urhfXk/lPbyS8aLmhwQs7xVm+ufXhd
AxMRsOXwUsD/vyZ+XVd8DTzjeDblt37lGprGv4XFdO+7s0HHrSe2upmcs5R4F6PjmGDrLcc3I+KI
Gc3xHSbR/MOOjfbQ2zivdGES2TtZ3iOjyli60CiAHLASNsK4nsNtU9mT8fki/Y+SFxlMW4o9NXmL
Eq9H8qILC4VZPb13UvyA55T1x5xxs85prFMwsZVy2ynidLzaVm0E1h/ecy75knkueVwgIPnN4HrW
bAExf3zD7qdMrd2U5tWkwbwk7VSvRnBRg5QY6GdkB4ZGi+UvfL13BxnH2MRizQ2Ck+/Ph9RDBE8p
v89kBbW1VPOB+HP1Wfki9eXs+Aum3i2b+65ameHT3idAcP5fova5aDAcToTla1bqFZHqjTE9Zo4H
9OHSoNwgHaKufCU5BGVsxZjp+TxW5GJq518lKKlALu76gjaGdndb+EYMjBcuTkcHeXHG5Mxf4gAJ
jiYwZxkKUHTZWE/PQWVLIXC/X3A8iFOTIWwT9WT6NhVJbvrsRGCz5GkF7LfX+sK5Nl3mm4K0h280
YctDY6S1J6wXr7lnUMq5U8DL6hw3vVUMFG7iVNtmir5JDSPwr27gH0jb+nXE5Bv6JYwNAfgTfWqM
88r7aNlmyfbWacc2ssSYJynUlLm5PcW2zGAu19pHL8oFrD6pmDVQyxsjtK4J3LOFNcKf6ROYua5P
ErAJDHnMAhqWauW4JiMjzeOSo/SYT5XCNADSkkAXvehWkZSq9Y8Oxjv94fRaJ5ah0Nye/J8GFT7b
QW4b7T3eN1VmMAYtYk9vnMni9u2kQDafQhHKTsOcA++SRBFrm/P1k8HXO+Q/Te2pHTWF0ev41yxd
buJEiW3cmQ6uvF40b8OJexVljtUF3rmYiiur5RML0Flwh8aHhNgLRAksyklgGlERQ03qeJ/zYgIT
NMUN9lFaQWB4It4iTcj/xV18kLW04EZ2n/gWRmHKnrGmINSMpoFMZUrNqIPysE/Wyd7H8HYxXPUU
SI32k7QwrIx4O4GLuJKezUVgqLcpW+ZnmBEogCuDRM25kMVVUcz2/DB3R/GOvqwOgsPlptYI9Llj
21Tn9cRVQGc5d9sbFztZa0elpOp1g0zq822SAG68dK2rw+xAv7DCN/5jtRkgYd0fdntsCyLoKkTg
Gy3ICryvMCGlsnId9KtjiRIDvIyt+XBNxcd3abo/SK9ju2pTNV9sISpKQM0ZJBrAIgN2FQELMCRf
x7Nya+E+NRiytGESdq4ULEsbjNC7y1qd/RMokjcNCFRQELCRvhbmtBuLSOtrNoOI3XBbOVkoPclX
Zq34FLZzv9a/RUafccq684RfRQ8Wumgd+JflJ1coGd3ya7D6g/6j6bVxGyWqgavNpRJ648nj+8kg
GKc+VbAVWWyHBA8zh0qW3IduEQrfBeRnKf3uCof9U7yUHi/DCp+zQvJeNi/zkCRfU+V6bURmIdFK
GF7bZJaZkJCfpeDx1n93evIRdhopIbnwCxLiZVFaRsDqH9hfrZ4vw7WH7cjyz0XJ3SxWrBUi4O+V
ZN+5c2dY/BUwYTxuAvEFhKdCgNCTNgXxU9VlK14lucfQb8E4sNetXTcngWdkASw9r4JLGmEYpElJ
jY2MsimCLehac7Y/x/Uzp98/nkTnESsIif0dN5c+ICKSQSbvwApuXlQ3+xp664dMj16OmVIBZ0Ra
CcY+zahDAurDWN7sMdg7uBcsL5TkQrp3vksFiTjoy+oznD7u7b/9WNfvkaYDDlbAZyQezY8rUYhE
0Bp7p/8eJ2H7jlBQiBS7nPssi0tiHN1yAU9TlatyJkjksthepHQPtkk7W0CvXFJCd2kI0ehwJHwp
zGqrndukmWS4gxPSwU2ZSOZ00s8cvhWiqtc/KkPo9hhyT3BPQvqotSZdcX8/NonnLk/CKmWAhccr
OuKqlM0B5ImLtutKqcabkWZHXQhEAX/rm0oSW8RW3m83j+JqngOOJZMtKnc7BqgBUt4r/o9/CUvT
kPKIX4HJeuJ00vmGxd40y9BBZUWMzEyJW7+LZPNXP0E97ngS1d502WyNQ5fDFCzjvzNiDGcSQ1UI
LEqFuGhF0d1W6VZOJhckyPR7gczyWvw5m6FsHZEkgmAqmfjfZzmDoCU6NPW9IkYQecMpXxYQXkNG
urmxn3IsVdP3eoZEJw0Q7JnkaNAORflW+6zQPL8NF9hpy56zNv07RaSvu5B0UKanJmmOYsc6sxxR
8isLtuZf90WSAxTIhMALCcyiPeemen4Fr12oNLqoznPHLXthe80shMmIRnTVLBBq0DhF2tb/0IAE
yfJl+8B0Qgo7Gh2CMNTkJm5DCzkhJsSH+6zF0GB3uPrKA5r88rRXpTcrY2cyM5qldU78PDbb+gL3
5jE8ldG/t0YsRsj3PPcKF2tAvQt755txzJoZPnl8E0j5EZ+pG8lVPKozCKI++EwMOVJV3IL390Ic
/p4g+m7K5VdbEfBY1ZgSNmwrTi1jYs0k8ktYjQy/EIksOz3liULRsyf9KwENpcvyP7FcbTgbLcNH
M2GtU3hjOk7YUaJeCJ9USmUyvSpoIavZyJ3aCOhV9M9NighmYqY265vjHKcOC+zXwdndEURitf/C
ntwhmFXu1aJ6yx5Y1T6NlZrZwSMA1Luz4mFexIGHu5q3odgfwEOYN2nBLseNh/vrfiuGHuadl9PK
n5cY+OkKTXwU2J3j0mVlrL6/5rwFAWHH18gu59QIETP1qd5Jj2NP7s6piSYvKmHwNs4qF7nmOuEA
rlmLKAicO2cuavjY0F8NseEBykpFDnyqDRr1CBKsls91UlYsh71COsKz0kdTgYgS72Lf9iwg9+1t
tgQWX1VpYHPjYZFWwwjWRS1FjH3sUQGG8xMnfxyFa/JUzLK5ZyAlrvR1h8h7QZ8/QLR/r4DNUsv9
YIIQBb7bDZVWtI8abIjF+GGsskIsDF/3fOHaLkPVJL24K3a5G+FTwTSJcLG7cnsViZUUoKxHlvlr
e25TYT4JaXfcsKIavxyB/D8Ac5q79xuWZf9hS+u3KJjTNvooItkHdXSO+4O5+Yt80WKTC+vnoHth
vh4q+S/lEAmQKOP7cq+vIZh8YL2xmO8ozLVyAV1+PErE6+bLTk7EA5iBw/3Rv1O5i5Wbhj54Yvq2
fdr7vCTuYV5GHTFBrMQYdeQlQ6RgUr1yBJJwE4ilU4lhN9DoXg7iZ4CCqm0i8UUOx46jwG2Epjkr
o5+E1vQnGiASxVheM616etQtbvoXT4iwMuL1bMam5o4LFwwtNQke909tPujHNLX/xSXO2lD5oKXO
QKbDmpVZncNo6Jqy+3l8XwHaJVvYE1lZQjaxHoGCYlpSIF2BSuECh2PQbnQyLl3v06cfluHM6rxH
3a5vuCRUbjtCb3HjfuNCNErlIGtdQrsqOwIIB8g8Usvn8QRo8UDCT4Y0t9+gVPK62GvvyU+eiacL
clrICP81UgEEe9GMdesB9f/tWwlId1/95xLBAd328HukS++vGWCiJFw7hk7tn6RNCpC7/N+Yb+S2
BpwVbKpZXEgfTBXSM/OVKrjhfHNEod/aqvWTw6uSeQzDPZEbqWGfXou/t7a6ijiQZBYi8u+if3cB
ox1vDPEad6+QdnbNISPCBzNpivYF9yR8cQxAjAmfx9yu/8CkDeSNfXc0oJwW3HyEXzS++cXx9mGm
OkLASyDadpTBf1ivz+7aROFqUCsqbLw1ZRf01u2MT27WfYaiZws/bAiPYu3bgUGENtQJmSBW+/YX
iVXyPFESWPoykBxXk8aKAsX8YofRMGKufO1O8sm12OvB76gTcvsvdNohstp1lIlu2M8mGSfYgrp3
xzF++IT8TQaExS5kqmLNBE6bgFVcRTfSojU0zN+h0JBW+uXKmS29yOYOjAEMTTE94tLgVQ4HQYVU
ahQ7qHgSkr+NYiDzETC6B1nj0/WbgMvB6VddJydO6UFIzlvlqT+ljneuWkML8Xw+totf902QLQyH
8/Fya692KeOgMQIS9+TxxK26Tu45Yq/S8zlozLDVKBK126OvsZVbvyAHvUBWb+HvqT3sejBS9fR9
v3McmQsGoEraKQVmObffqQlD+gAYT5ZGBAV7Iw/ykpGecATqPpWKwNEucOpk41W3qinP/69x7E9N
zxMr1zPDV3cGFBx9EgJxaU8kQL6U2rAu1bKC4F6NT/8eGvipwYtOwWSDxRyvQJWBritxMQOd7g/x
WBf9TUFwHH0sSGqKBhwRR5POhwirk54QTlYnELqePflVRunazNobvhqvn8a1q12hoEoJsJegsIsD
JEAxTXJ/1lWjBeiUm4L52DfFtj0ASLUgOUjJHFosJBc+KapXU0j5v4MWEf3ZrimCukdt2MEJBn2z
vLwWTh5pWpDkkA8q15FNsuVPNDZ6ooDBaUXZj5bNPU7TIVFkzTj7ueZVGSDuesg6GiZ2ILUba72G
d5dZCm67fxqVNZYwf+yZ8tZCGiFv64RgNvOXNNwaI/lFiCvgwPFE2lcctcN0VAX83+57IzcF/zOg
vTsB8BWyStU4tOWVoLf/AZFYYnN1G7ASQohmJt4Dc4gb1WRQHVJDfYlALQydpA+w5aWBpjsmYyrM
FFuLtclNNQhgyuC1pDqnmb1Vos0iANrWwfRwdYZY7V9ocNdWpCIcA3Jex8B52Jmc7rf8h6SUwppq
YCsKO43dtKYNMqiNZWUEYIexiQoAFphWEukm41AX78aUU2xu6ur++y789DmuHVXm32qseVMFhopt
SUdSrv1aouYZRJRmgoULvbvhHMSsSJLZGFlAIsWGgf3FLl21o0OAqRwAXa24JB3C6oiK8imLSBiG
NiP2GCWWr9q0GQxWP5oneI7H108YKhfgMmTzEfxAem/iO2Y/hMP1bvExBVO6UGiqzZvOtS3UZNjg
mzUXbyQD7g9uUYfw+XI3CU7eaunKD/rBhNdft0g6+v/F18KRix2xmtF+CwjY8moGlZhUL6y8Rqq6
IzFCFYiE4KYoQal7dhCpOvDh3+UpDA6PzPYxsTw+N3XWUEI12WdWUlE8PvzR8QScNdHaIihUJ/jh
xOcmCk9wPAS1UAhuzxpSr5eqklFbBmVFGcrK/tL5fR0Chz6r0OHNW8Aajy+q+cPX9QJn+YjrOl5U
Wok3UvtjQNvwKXU2OL6zVYoiT5PbVF6nHGLzQWU9GoIguPoLef78Rf4Rovf3fVUzgqSooTt2DjOd
FhEcC87ULrjCt9+UIVIrm1fRaCIwaOr+5d6SeLbvaxZTrMx2qqikXiR4TkNSLYfJADg/hzKBmrUp
BwVAr5RRmxzgimjWLKS8cLnsFMy2PJOYnqgn0HuV3sOLLKJYYwpnBUjGMz2ITP6ey9yZlT2Bl3Zs
hY4uvUlh5Y0ZwzPqepKhZ0j2fG9tK5sSNv1MQHkxwSs9txq/ph2tK+vhBrU7bNgk09wdLeJj/428
w1eI8RY2pQVR6LBEEGn3Ug0W9z2Vn4V5brkF6r0lpIZ875JuNYCWTkKH9GAdaGCnPzWpDOx0A7xl
/oQ6c7bzsYUrU2wRdehzk1MTcNBnJl7bqzoizIB7DJ1tqez7XSslqTJ/HTDwhZHmc8FBlgqix1e4
QVmOPXMA+TfFILW6zQu0iznOvRoLVQ5IUTK/Sgl9USkARb/9UBr/FHMsK0Y/y8t0ZsBCWQox/TOL
REVG0+699CfSmCYetHa+6742vB4LT5NVIrrOZcn5zpHCGUJCYckhwGrBCXC5XHHAz06Ehb8yt+Cd
35pmPiYNsMY+tTpwJ4CYA+C86njAZtniKoKKrY8zg/wYURRHG1bzzTvVwJ0kNLJvB9+JFFsqbSxo
9SxjvwKDUUkUkc6waaxN22ePQXufniIPdmNX4iRTpZKlBOBVQSxS7uaK6GTPDWqCWSKOGAcyqHXJ
F8OXDnrjkg07EwSA/uuGnLrAsCDhL0KRTBcOjtqzYLMYHAD1Cj/P30w96gpz4LOVZ5kvNFrDJr5a
9eP5TyZsp2EfHt010pzoudsF37J874AKsxwUsbyLUDoX901Ku3srThHoLj1PHKJSfie6G8uprBxe
GVtK+ZR11NyzKP8prPK7y5UwurIxdjtZxbxrsrPKVB12BKjlVZ9O2+xZFv9jlLoimXifSnbAo9R2
zyCBh1/r+9ZMe0FqjHSateX3xvFN+5P7vQ72tWBfdIb6+A6aZLOsNCvMxeuPf+zcB/Lx4bUkNCXx
8c5zdG2cFfSMaIkrqFzAAP0pLqVSdiLPDPzqPJNneBeEFwtgaPIn53l1WsLNYQfgSb+EYzvYDEo8
gh+jbP/5X3JiJoMEPF/Utx2gdGU6rYGmU6VoOub1T+5x7EK+/9X7xFKwQuwgsSpBClalAj7ipVMi
cOJ7SDhUEbON4HYPn9RFi25qtTRaI1x71DGMY+TjKGSgVnbDXWoJFnBepRQuwuIeYYC4S505230a
8Z2tp/Qoua/m7qVumtXOQ4L6CHWOAAEikqzhU2jzIb5OPdYf6RIIhSDUWU/wDdAjx7pq/4srosNv
aOUDimeJD43ZDQKCYwXwkiIESPGS0IBIGCk4iiUEbQPI7BxyXfYiTkkdWxNaAJ/I2OrN1e+1xMT3
R4EEu7HFGB+LpQbaaUOIlszghHtRrBxNnaZZUqoHVN94acLcQfxzMjKbsSrU609eVG+Jo62kB8ad
5hU93baNiEb39klbGQSP1cKWLyaocs9JFq9OyjrmxiRu1LVfT+lIUFfeqRJLDf+CaWzkATIkAoO2
M5WmNHPJL9NJThEc0W8mCAXr3lh16DsktKCUbTkQFnVsAfdhcydqK6C/pkuUhARdlrmy43GK7WGN
Dr+AGwlWkXzsWitVz1UGQJ2S98F/v9ZU9iW7fFuozNOoHiA7M/oXGukaD8OqzeX7tkh+Gvrw3Xi+
+sxsahqkBeq8uiBxHI+gfv5Qq8cwfEyzl1tuiTaGhuCS3wCcuWGzZuugVIDNnI5VVObAqGjG0Xxu
5y1rRtT7NnXlx9jNjBhi0mkL0VK5TGZrpq9Mh9LF7iHar3u5AiENKLqQVzqW3ki3mELXvIpU7pdf
eJBNl0R/GJmfiXC/HdhV+SQcr3lBBqDVuP5qbUJm4oVNtWvvfKdL93Yv9tuSzRc6jDiwqxbE2olB
zaAvt/NurvxetUHDPUwPrYn+mFAIhXgzRWV9Y77K2QZv2xBdNMfnPLUjhx/Lj0L85zGEDFY2HcPU
tCoLz91e7aFVMbVgZeP+wCbbLmbEfoKauf8xXhcnNBLqqvMF8BUFTDZSr3/GlXKXP7ypRS7NI29I
vXmZVRMxnlWysn1mXSrfKju3mlA5m7ydD30FlUJdT5cPup+2wWVRyLd4A8aVHcmvDy+TSEkScxFK
cYbWGDyn3NgKuk3o+gCdllUXq5gBRnUunjKkD49aZEq+WerA6Upi30xrSSwtf4SrEkUoPzL+9bMu
/nAzqhTfOBQVlYpYgTpA3O2i06G/1lQw+xCZPKgI8LlQ10TrqdWSPRmWOB29XBfHmarCAjtIXvmE
m8Wcvt9rboO4SAqeGNuHgEGa5+NrsQC3DGg2rF78dluUNxf+Ir/dBoXv6ZCqElhL+anl7Qhznu/C
mMJ+sbedPB8OHDR9Cj5vJ1EJUIpIgnbQQPVQgMNf2zn4ATCH7+asfwwJ3O9PEglqfhI/bJ7rtQ4J
sRGOgzGAlNINWZ3wIzdz9gHofbMGl1TG8py9zGcxLzl73HB3mTKJYRndo64rOk6efS4ycm5n4Rsk
MNxDTq/Ur1IR9zW0BmKuylzXoSOopSFt9dMYSuvmcw6JeS4JPbtFAiphixBoo7cluf03+HgAcMIY
v9+paFBB5t00KwmC4H4jBfb0+SnMm7yczhlirFsQT6sW/EpL7sFXFiCeYVEv1VxEFzfwdjiMNtfS
26Blqm0kKBDMr/atdXlqXvgflUz/akvGniouvVlRi/A5omF2+KYp7Ei7tYiHKlc3soAG8nEpzlf1
5oLSIL3aJp85ZbNSedqES21cKrhOycS8/bNHAPNKMJQxIXmDM4vMpJQv9FcCQYT3PuMc2KjPWeqg
1LOT+GTViQoPJbSJw8n5ia+5Hm4qK/twP0bOquCekt5XIcFDoE7/2/cCP9MQFYZNLYby8xcP9lPz
Y0ICbW2Ist8SGWDzgocDqVPAGd4wX1EA2C4mob8Ckga/WPtkit9QqC+jxDzxelBOu2mO/wfAZ++h
HQ2YJ+EzJvdyf2vP7aHMqA7xkt7PtTqtGZKgZ4FWExNck6iHfD0IO8qcBrxMeU8WRLVDPvU8clWI
8tNrI9cQ9EuKzzVReDOdT7KM7+fEi7Q339Usb8mX0X9JuAUA3RkFffVa8uDg4+WcjY7W4j8lhAie
tPsXg/abZ0mZKLRh138jLpgVB/RWbND8wvtCoJN3Lft9K2mGi4mDU245s1fs7dFEKxbC2FoHqbXg
/amL0cjWP2RKzZ64pbqYVqiEIqhSECJa4LU3pskF1p+ML9eU/Ir6OSrauRrl8B0lPYx2x6h+AiAQ
xHEgJksgTySfqMBfHAcsWVvBBVWeP2Lqwd1eNm/2cD6vnstOSzN8uU9juJKyQQSJCpGAgcxtyCDm
HZFZO5N2qEL9zr4FR8uJA5z3JJJG9pOGqbAoeL51wN6GokhvQHZoae2LuZpCtuMPF0bGkhS1uD13
pPPyZdltw7i1epoCqNakNR7qCRsD7k3jtOPPiibT1qGDU6Ce5v/rED5W2mS6a+tiidl+DWAE1jDq
zes6YN2jfCpe++WVvjAz9Fxi6oazT1JybAZWBltM4prhuk2lr+isBDvdykBQAi7mPbYbh7ZYTGrR
gSl2/53ScEA4KiERGF0dimVubueqydE/wdn+iRTnOIyC9k9go4ImU9voIPm13BjuQpXdSODXTjcS
btPNWte+EO0q44M0F/asB49NMTnO6+t8Z7fOHke9myqO+20DPTSb3RFVYhndGQ2b+M6IUPdIm/mX
UHQ+t6XzYI4A2jYauHGgbPf48UyoBVed6irdsEhQt35830iAo9lOblUEsk3usy/b/BmMWGuJv3Wj
4Oftc6pY6NaNTzKkpy3Z4uHxqtPwveaU2vq/oy7GHBxBaHTKhtrMeJ7NxpVSCFeW7FDc/6fyP1SW
Jg8V+2fjuDLtuX1gy/qB0BJSFjplhbYeu4DB5gpL2jDxVb1ALCtfxMXOJlozvS3HRJNv9Yr21HTQ
QUpwRJ9aREuvKAjLwFmy6gGr3kkSohZHcydj9mdJzvM+6nd7/F/+1/byWwevJJXRHLII4pawaIV8
H2Cca1OgbKpv+4q5OzxTK3KutqvsaPx4CS+CgCsCYTT1DAssq6B268vD8sgPerf6scUaKxjwi9bq
rMcDus0lF5AXBW8OVvDA3O0IWPlfj11IffgDWapkL/gwYQdwGJGHfGDufccEkcZK8kt1mSyJduip
8eLvniLNVmeruVf24jSTMau3qtxvPuYGDzHFo3eEwN/CXMhDW0SmhY5T98HnhX2K6hFO2aBKJUjC
asXu5TAOH02mSm2okhaoL1DWCsga1yVOpmEnQkJWfzTWxUP6rOGjLr856296FIKTqobRM8i1+4K7
pMdvahKql0wLOBRGluJJppfpM/Z7gVsBQsqDDvGlcohDV8s+o3Y9tGJcmlUxHTALTNMbRPMgI4uf
NuE8r+Nl6fCCj7wFtXlqQu919Av47IkgzUmC5ZmX4I5UVppwSvX9PLjA2z9ePBq6lnRdia1PHuqo
o86wDR/dOpwR3FRiuH2ArouTSazTg5cRKiBDKSdX0SKs1T3F1fl3zK0ObnNpys01F8p132BbdVXF
U6YPg33pO5Gw+Eck16gi6pM5G6YHhaDAEbSHQm3KhdX2K1dWkKCZZB9y/xyT9ddqtWq3PP62mDcB
izGE1leOG/pNg+e5+R8i9z7m5JyfuLGEC6NrvQcxSuYa5znBf+m6WJKLemBL1TtxvFsUBJxMJOFs
abGAHEXGyu85yLn2VHbp7jBz2Ru6hvJdmEIlEWKdIzcm/zp5XlDE5nOgS6/EGOS+q1vz9NJxObbb
R16INu25uIS39RU8Kqk/C6VNwN8DCHq6LWS1+mf3RLTh9wOuI8eN48Ck6bxsrDSDGJBPE+A59wGz
TGAEYbwtg+GCrYSdLzmIR8t54Q6YzctrFBR9iCFWOziA2qR1SWE09jXbEtUqhJ/XfUW8Nz/TatuD
MPWPRe1vyeRbxH4xxIB50sHPT9D04sLvp9AQ2LIqZLWSVcqqSGgN7AEflbrsItmoCipJhFHLSDd/
vGbLLZsc5XqVAuaFWf9xw2Vng2ikH9Rhxwzu672fePoviE8pGKoTUZkmSu0R93vCftF3aVq/3ovo
Px8QNCm0tNFxoLx0E0WhWurDxFgD5ZHQvyJuafRRG4OvhZQG7vnC0+C8GAAD9GwJR7uIfZlke5ES
UzX9MmjqX45ZbZpp31HknMjtCntoBUO5eyUadLZeMFHCN9SGDMR+lumAqZ50Dd9+2VDdVp60tZd4
DffDlCBrohoNziJZbHJ4+79b35uQUaOsRweNitz6Z0qA94LebhW+E/dCe5nDPyI3Bliv93w87+VV
gW5hL9rp1cb8kWwOgzkojufxqdnFDZt4OvGbLJl+NliGO8x31JjimEXa8t/BjzyiHijuO0zGwC81
VflDq7vLlM7ZDIvb3lNYacv7tk0S1oOSIOn7og+72oYQbcpRpsG/NpmNNXuc2PtkyBeJughhGi1r
X0UnRB1wnZktIz3yaMfEjhLZeIFVGEIz0i+m6uAegkvDttQzJG7YaOVEPpK7I7UoIaIDUVmjw7+D
4gcm0LP8s9I2+tyDctn+lcUWx4dsoMdTaZ6vg/Tr7AUAoX7Xs2StIgzTAmP0O+bttNeoCxr8D10m
JWUPEIMt/dZF5v84RsGJWKlLiFXL4aBXg7kGiGUrqj1OX2d5jNQ65FdBbGH4x4hQQIJvKShZVZ0l
mNMTziC51Fjq4p0+M9OQ/gcHmbcr/lgfLljwEfbTd9L8W77Z9Ph8tHH9N8rMHL48AAoXXnJSIXwY
hH35mbBFArSTm571YxzFVtxxiyWFaDGVorL2HUsdn3IWWImf67fTgeaVL6w0mAbdLNoCbmynNvCD
c8bcbVloIWioSR4B8jcuJF4arMISiA+35fJwO64uAQ8AWuOtaz22xgWA8CVAkBzRfz2j7AmJHIO2
AfPO5ah4bagb4qwuP+96tNiCCsdyqnztuFjZtGgP+aRK7VnyJG14xu2R8bquxWc0b2dJgTeuNJGm
B+WuM5o1RSSJ+NwC6zs7Kv6ONsT03vnt6urL3XkXF0b7j1oXurB2idqzk/nw+CC/7uOTNoCxBQ89
JcxiurRjstyPFRgmHBS3igpeMz9ZWsvu6ehRtZ6TUPtnJYmoBm8AuGUTxC9t9R9sttHvknR5lCfz
QC8CK3CHSnhNgQxLS5G8quutdlH9DmTdQ/8647RcoMB5NAaB7PQo5HElovluMLZfbsV1ixlyIo3P
vLm3NtZ6Tl2N8WziuZ07rWuJQxDDlQlypMb1PiNCFbeEcbF7UX47v9Jbh0/UBUoSSsCSPjJvqTCU
ra4E/EObG5okih16hlrc56cAE52nFQDxpCmVVcBlhXWf5NN26hAgBIYRtS/HOJ7eGFoJH5TArrYM
Q+riDgOToqnynbtwQ97TAIqZGFtOekZXFeyJ7ecTJgrkUMLqPwp+cnOAl+saLh1Ao2CsOxQDlw1g
CWh9BUL1cThpORuR4mJtz0HTuGGl5Rs5noTS91Tu34L/fPxg2A7tKm/TdF4ej+xQjx8uwaRhiMSp
Dtj/4ocEJU9IRKkLr23iAXjr+xjHJrdHc5IjHafgZRL2wAmSBg9B/hVSlLrKYy4nNGVz+5kY8Mnw
Q0t2UivVSsOHR5k+ITSESeTarIwprLedMnAAnJtezwkptFkKC7lR5eFXs9d50BS7NdrbdNXyuPue
SiOxGqjogAO2ryAU9SSjmDizpV9x3yPTsoId/M7nw79SndlXCE0sZOdMoB4aIX2XkB/4c6fqACwq
LQJZv/S7i1wiCxEGUuMtyZW14sIXgZboJ/cBRZdvIDD6F7M459Exja0Ay80i5sNZuJQpwsdicjo7
NoHC2EbA+/F2lbXJvZMuo8o2/yDVtuP4JO64Zy9wDrHw+5KoQR+63pSXN7e/3NoORkChPj1h7L7Z
HfLlSC5rm/FYkXnQWiYc8WfByoEvHnTmmbdTeTi2iUCn5+65WcVca/ijVA3oqy6lUCeNbAMX0h+x
L2SWJMa/4fgRDsCwKqH95zEbdF7QZGgQvULxBdgj2ddhMQpU0H6zqK16bfkKJSUylrf/R2ues85E
DgyBLZAdTZcVmVuLglaF574ObCM5KmyHO7b91ObGJ4IF3ndLWaaFMuvBLWMTJStbz0Mxyp07KS6S
krMx0v1d9shZEGrcffx1Hz8eMNRIUXDKIgGBhLsuqP/glfpIdQbp32h1xrV37yfz/2fuWK9r9CUr
sFTuMwmIuxTVWfVwUmu2a8HNwoSrW9f319VEinKvGPddndWFtRU5gJhtH0G8e9Aj4flglfKZfKKo
L72SwxVgZT5NyPKsnHNYfcoVWxKqqHdj+mW2OrjFaX0zcfP6iXk6WwXUcULq4eW9nNTCNoQCCYPR
Lsopxc/fwyMes6ryIJRDXf5BLdOn4Wb3xkWw7YScyp8/Et01YehNvvtje3RVl3wJXpQtOoKgpH1u
In16G6/3gAri9Y8wlw8c8aUO2gPtSQQ8M4R6AIN8pGco++bSDUx0fXY/oIP8CwT189erPljwR/et
yZTRJ7fAXDzmGlt4DR04N5E/5Ak22yrZqOMKXp11gE0vl20vuMVia2ZPAIcfCsbJqtGTHz4Zq18d
Yz8b7ugaJAxKq7en5ZukbKXJaxakdzV7UUgZzHYN3EDOmCJ9s/KHHEiLi2kWToFQJqs+Ti+0DABB
wZnBGC5/unGcDAe7IV6HlRpQ7c/XP/4yOgonyciFWp39Irad57XKB1d58dTYDqlKuiZ8LqcPWHXM
KXZcakQKYpQqpnV1BTmyIlLfKAsdnozFr9tR2vZuu+bRLUk+Ro6xObylWu4O6GlhY25jttoprBsd
pOnbyhj94lTVonIM/kEBASJyAbxIYKWb5UjlO22pBpD2fURWNY43iQkZmZSrJNZCZewJFzpwlMZq
jcUfKP/Kyw9pkwpwiOdRQWdp43iBcOEheKqzd7AuskywFCiKzhpyPHWJVkFTvm+Uq17YLDVHoynK
sHUmwy7X00NxRsDs/BwAGMlUaF0ziCys1guRefe8Ry00yS1mGsRO6S7LK4qJFagUAU+bo2Xm/iv4
x6ehz0i/CQIXgI85Rz/JZfmeOYqUqSGswylUwowXkcVgznKEgLN58hpUqwkCarsveAxs+o9WTUJf
Xqb2v+36ibuY/xWCyS6MqUzMGKJBDD44WQjPC9wFpP2AejadGMnsugr0IrN1NSVwILU46/JBC+UR
fKHH7LFT0wo9pHf5fRnwdZXV7AG5eaEwAkS06PSyUvffJ/kSkTm3zyAKJAcYNvigfVgfBfN09hIZ
kTeXN9fntdJ2m+aYf2uyCFsmdqDvuP5wZ3xtd/asdf4hTlvO7bNxbK/vZIjDl18nt0batPnFThOP
K2cwmamIN4U8Ob03SMnVBZZ9Ag1bOoMeBQ7DB68ILZL37qGNxig/Qa8iXMzwAloTJSoOCbaw03Rb
lQWDwg8VdsEIx3wSxW3oWiCBYG0DCl+w/GDRkf5aKOOjD4lK640UGqK+DGb+r3SqdGzyAq9JeKWF
i1aNzHH/FWs4o1YSOwYni7PjKvdl04Fh1FTpgpX25FX+JSO8/QjNQ2zH7uV2UxmRb2mKvVPwvfzr
DKA1JuuT1P+cPJgJrHy8Ed0+xSJzZCDE1BDVHUAmuYU+W/hpBFROq+bozCDlj2uzAfzH4O0IFy9c
PhGQjswauUBCiqzyCPyBvBePj+cRuXTg/u0ut1l0Px51/Cnf0M2Cr7hXU4qUekIRcZLixHm9atSP
KBddn389drcN6tDmJzsipo9X8RgVOCEsndGREFQkiUGjKyrCz4hhSrn6Kz0PsK6lReMHKCKwiMOn
09IjqBmno84CAYqKD8k9J0lf2dxk6u/Za9Etrtpp0xk7cUuSVYchcl0PevPCvLjTuoVm7+lEqcx9
ANRA7TV2frdrJB5zFBhMLk8QVUipIKVEexCCt/oYXbc6pcJq2HzOc8/hZdhUjIyyCdPJ0bunJ6tW
MbBflldbDI4J0tWQSinrH0uxkwENZOHM3N+ysDYepuz5UmHiQ7hzI3xXnOTzBvOhD8PZnITpwpRD
HUekt7s+YTffaLnu1At9syLJ8tw9Z6+OJ8ewUEsJGVhaxLJ9HuJlx2wYS7AyDAl0D6VwCrcRj1Mz
e0ZR+oZaWtiDfWxq7ZJGSDbT3nczIPgd4WFvaUInmI1H39fFKl/HprQGRyu27AJEvcbTtCxqaCAS
QzJ1C7kohWxaJoiidUgn2s7syb6vNDTv9aupq8mvsvFSzPPWmCYal+OEASSM2+JI7xarnZfTO9Nw
gNKlz9xYd68xxODkVvtgHt0K5XjTPgB/ZofaJlPSlwMekzOLAv8bhpkErWskRTVFDkPs9/1Dkm/C
twRm/iAd7CpMIjdsFgm6FCvbErRDuwqkJPW0w8GJvMyr4wiDVUhZLUAG69LT9M5RyW/ERNNSGT/N
X8dyZV1DRHgkYoDWhoqTjYb3O8yafRP1WJJIixf+6Yjvr0LUv8O8XvnGRcMTlFkk4r2g8yt4JmAS
HX8VVJakpIO3i9cGoTC0YDV3LfsiTkJGMVT9BnczlXYhvQW2YrbR3OmBDfNPaTFc3zBTr/R6zhbd
rRkEJtwPf8EN5N2ViNzOTrrM/eDroPmfyndsVIZ+xGaV4cXLfnYR38U4kgeHagwz62L1t2r0H8mI
/0eoXLmkKkHeEGHKL4ngM5AE8GdNok4DL/9b17Pck1WS/t8UWB5GEVYvsmOU1Acg2h2r/q8xKZnV
F6WsqkLe5Jz0GBb4kZyxXQQMHBAHI2GuYu4C3jTzWWLpCASeWfJBPLFOgZ7tKyaDO78ciTFO0TO1
JDP6+A4DjG5jngXDLptL3s43HAcde5tT64ehVetKjPPTCYs2rSVwC5OPm63kBdOGZ0O9JhKpYtqj
SedHIJdPvaxwUU5MGewgLTZx8EZx+euaI2KpR2Q8x51IEvMp2HCz8knhwWiCuN18bLpwM4Y0htv4
PPjAMfpqF6c1UgWA93NAtAOlJBIuQ03bZ5GU0kn2BegbJ29xTX9jELLN6kk28fRdHU+TY3gg0sRC
UDP6NBIpxD6v3needGx6Xe1q2gpAdyi4K+MevhR9eCbVO4ZnOVAbvk1aDPGP8/uok6U5Z7UuKBUP
+AIZDj67VlTMbI4+mWEoo69uLWcLOBH/dPCIEPH4Si9USO098oLK4UgOV8cqkt/VYjWWCrReK07U
ciJjbc8KrVToqrfcA8ag15lMCZWECdUPax4tfpK3D2RXqGdCnuk8cBeDrdSy+h36t1Orngn/Jch4
wsvIuaubfYizglC9yxY3jRfnnRIp+NhPi/12EvqlGN/+K2gHATxMKSMSAAwbnEOeC/WxEt1VDI+q
4EkA/dbFhpH73woNfJPvvoEvb3NanyuBa5LYy9JbIF5sRPOKh+VjDhdbTn03MFLKDDn3AQYUzT3m
9cAPYDCMJm3MEvbWmDqy5dcuLbNP7rehaFMb8VyZ5pKiNWOE1P8MV71x+myHAnGP0l20oxjZrjD7
cFpBUNuyTL3VzZTGDVb10t5boXeaja4AiNJs0QzSrkiMp5vahWqmz8+GBtjh2jB0W3PZjWSrYInh
wNddnIDIzvdDQPdwnAvKUjSxX8EsJ+i+3v4mj19EUpSDyRZv5FxrOkZQ+fHVnqs7stqm46qdLuzc
1xm5L6B/06ZP2WzqG/44JuFJ20qSTNvVN1EZ2VlT8zZzUFzyliLmFTxN3rPcnfMLn4XHI74RHUst
CESwmlCqwLL+t7QM4ZlQRtDp9Wqtw9grFDvB/iaGxAfo4hStC/vMVe7bHjHVAQ8oXCw8z6eG/kmo
449dGK5dYEBTzXBi24L2+hZd4brcKaFmUY4p16T5NDhZSaVVb20jkFAaqCQNq/ojTktMrl+2YKAs
imVyZeHBVSEKDuKXxhzRzrOR42NbIEAxXvWvUAF1YxPwETWl/UalGAqaUb5b4YL4dcTdBmtIq1lF
RbKrvyt4OIZvlxgNfFoDmwel1Mxx2885EYUkEol1cCciTzJgLByJtfEERy5FP6+SDi2GtNMg1KII
gAgGoyLzV/KuWVT9veOG07KHp8+GR6Iep13OSQEZFIXhV8em7fCwUI7pNPi0qxZgWv/jeXlAeAY+
MTq0jmmnZe9SIjqartAW1V6NStArpUTiMCsCmoqCzhO3FHjQVNAh4/v//tsBfZha0D3Pj5wRSqtr
hMyCMdYOOqU4H5S8OoRxKLwNr9auxcGuT/DLx0boyCtNjfOJ0tTEYtXLN2STE7Cu9wI0pwfWphiw
MTBY+R1YC4hOAXW5W3VrAu4f7Zkn8FqT0teJvt2kTXwhsFijfipb/Fhx6g8smPXcKORgPLWRgm5t
x8l04VOEJHxE8rtR/q9qGumwWTdXuy/+N0ongYCQkEJ2TT5QBjZ8T7YoWjEjb965EVjDkZ8qbY74
KqhOaUPFOWqNKt/vVX+fI95sy03iG4FebFU3zCcH8xbJWoBGjCJkgskN3HeKrrmgBTlji/i7JhT7
kcJwpkQXNe2bLqxZiix7LBfnwSSExuMPVLNVrdRua47HIZB7hryLOaFAslUs+jdD3Fq2R7rW4ieD
VtOFLtCb4/fw0uQxu4urgdP6NodWJivE9v4xKEKeD/f2Ux79MwzQ3RBa+B1Tq1BsGw2e0OSpN0Gk
3nN3of20FsZsEc1TmcNsCmxQ/Fg9K8h1PLpbYpUEZwvzC2D611J+Qpr3rgJtcP3Lr5LW+kfL0WDU
IT7yTDZ0oPOBWq5urcd4eom/LR7nSiCnvIc4ojX7ZeOvWFUmhiTKJN1/uAhPxdJ2SJzBvmKu/5Uc
EW7V9UVOR6G9CJd5m6TNWwIFyT3Ytq4n1rDf14rv75a6TrFlG7Oq8R08hAibnRzrDq1FrAoSD/1I
YUxHQAuMP8tIpOdwNORF2qQF4X4Vr9BpISRSBYbDqxmlyHvI7u38SBjCpIHesRbudCEAbDLsQRnl
SppNgmHKVlv5u+M+XoRs0VjHl2KJQKxkBwTwgImGz3oKMjBGUe2bzJ5ogIXFpPU6aDOo8yFSytmL
Yyz0hL8syxKjaFOxwmkuZjMYoU0qnLDD2gAoA+BR5o7MLJOiLb1WpVDUK/kbiQa/2hyoY/eUIAPc
xm2xbGCGxiTTT/PAQkmQGkKmrVYEcTFL5K5PMWDBixPKISlphQe4WLMvB0PxWJ9cckApqy6q07wt
YT3QFpAA4ddVFJBnFYif35Rrnso1dDJtv19JRkFnL0t0IlLKygabpLVfqkkvcrCzQbtPWx7gyMft
G2yVvgfqmpiTDBcnhzSmIIkqlAeICujetMeJQrlGPTvCksLh3xs/jDwdr3srNgxC8QeVRZdmmEy7
L3hjwcxXGdRT9h303xkDU/CG9lY4MkDobKZC5S0fDbjPymRrhtGCFY+ITFMw5MM2pzjUenfn061W
LNP6rNSPF31b5fYBRA3rtq/uPwYjx4YLBeLPyhxcaAB/JY2HfYFF5Dwjb4S715AXH8isrZIA+U99
wHJuFDcwM7C+x+n5/niJ5KWR0gyQLUmxXdtXi1J0+KmSpgsjjsT4SOPAa0M0PCzuf/jS5QIyGEOG
b+qWTsc73Wx1up1fYElC/ea8LylinvFfu8rE58RGiK+ceQCMg50lOmeqSRVOymgQZvOkZw3zKa0U
ygM0yDfWMy9MWRCObvIB38IPZ/dvmhbwf+3gXvZI1iF9S6amDREWz8gEJcO9i5JFkAuMW3BuNWJk
i6Vk9Dyqy3DAzc16RLP6XAj66k01kkmXOzyGN/pqdfbHh8iNtCAN4nZQr+NCPS7jinjrBor2/a9I
dutaSPclAjY5h24swFCeh8PuRph9t+OEDWl4wm20uvAbiAYgW3KV3U4vPizcWivXh7oqqrhq5aEP
s0DNiEwmSaMDUp2d0xaZSvIStTtAu6An4cPJuETLCxPoI45+U628k+tVY9liAMz8cOtMv152WohD
z1QRYie+j3WYAlFiEQKY5Ju0J+rX/AXqpitm161T3g6VtP1qzOjP5RWwajn5rnrCPCxuyTCcU33f
KT9smR0VscxFN9rPVJwoKBZiMPHBQBoF6Y7nJ32ZYoFF6/R8hJ0s59eyI9vMk+6XEHqabRv6mGQW
XaHFFMpQzaU3ZRTderncjno3dF8ibYL0hy0zskT6D0sjoPJYtiQBG3nvm+OohIMhNZIfQuAM+Kbd
vNbhDBtsisr7WAX/uuz4XAjXynI+0DMDosne5rjdsBb8h17tTbYdW0NhW+EK9G8ASJdEPFqdwcCU
cHupuQv9zbz1qsWLvEXXIlZ8Lk7/rTxGBzwT7Y9qWPIF//MTro8xHauS+UmF1ECvhuho7HqSSLcQ
oqiqXlSprw/oZgrMjfpJNQOJ2R57DF5kk8RfmFvW7YGq9Is1erTnWkXQYN9X3g8BLsFXRSiQJGmA
nSrNL9GheoevQ2etjPfkU8teSEFmj0xLKZe3eC60Hso7QDeBDzjqVDrK/NLOyMZGi8ODY2UiXzHj
Y55kbGb7ObYvzxJ2p2VNy2SeoG4ki5n38r5YsfVgz8Ypet2eTFvP9fLdS56w8+ZWcs7wHHrwDPOy
Bhrycl9U4GGBNS1zuLOJpbVUzkLwMbbv3i+OrET+Dal2S1THfkstZroE/JiRzCrSP2s/1BZfN/z9
Xta2C5H0GEmOskkV6m4E14QoYo3dkOx2/5/Q3ZON1RvP/Xc+QyoJBhMlNR4ri3JtUNg49gS7Xp0d
zZmq5s++DGxlaXhMSoolumtYOH5+1YT3GNtdbv9dFKmwxaSoJQx/u1HBg3WH0s+JRx2ULslFLNl0
DKbX6iDTqCm99qxcZgY+XXX83gB5icPof7r1mv2ckLfJwNNnwvzilYEn2lY4rsMiwcpaFaTPjieS
+mMZDlE2+IwVGEmIDmrn651zuyOkk80eoW9F2kQ0/kF9jEn+0nvAr3we2w+m+2CObw1XGbYJPkDA
v/wwqNJlQ15w+SElecXSeoujuTgFPE+cjNAufzlG65XbLeNuoP1HbG32v75Wovtj8Scr0ENLsPlD
PgSYbtgvKK0IWRax95dt/MyGljubQotdCR20T1p5IrLY3JViABBmusNxDHebgzZ1hgTv56CDIIMv
KKM/UdqMaqvttx55OL3RvAeYyQSlC90rHHV5SVtPwZEBZ1laV02bdJiPys8ICfa6JmGatLzyzIQc
7G7eOP5q54XLdhrqOxso18/VJYuaJBAm/RKbOa3BGGCPyg3p/Ng8gWPP+HnVUo8cp9xfm1wr4Djl
KaCS4dU1Cocgw7Poj1pIqNzSMYqt570qVCP2uRD61j3EgbNikw+wLJfoYxwalCld7ykaL2ywd/pu
uXMXpsPz7OcVkDJIM2yKeO6/Qpgs/4jO5MJ9jq9xSsA2GhofhvVjc+R6o1OqhitKl0J2kkI/x+M3
8dtWDeF5kjxSNijn68R5G8jhjuMCrjVN/DeOCtCJZYUeZuXGL0WTtMnd2Zo9kvXkwpDFUQQL8M6x
aEPFJsKTUsD7A+VZiKfgeINVGrr4ea8r/Nforg+kv4vYBoP83JA93+qcrAsrkqf37IupmhpFKv0p
bHJM0o/0T4NvkoAB5D/xzzHKKlatJPnQVz1BrdE7Kkhd8MQRnZSLzWKS5C9WQqglsHNl7OQBvEpp
icYLzICmDqe+RFqr8fNYUKTl9XkWROEY7dQUNDADStLpnViPtuzFA/3Ezxry2AqieHy1nNQNcyVg
Hd9eeM6a4xvYm6n9q8UqZ/HaPt5669zpuN2mpUZ2ci80A9i1dWwQzyZ/J7u4MmEdMnp5dNf4HJpr
XzcTFjMqxZqXZdi+yVdiIEhgS+JJvlb7vvZBoKpH71191kLjjwzLUv4Q3wbuf/BUiSwt14pPzb0/
ij1d9xarrQ1rxxOJYS57nWIE1y8xdPus9aZKFHTPmSMe5e0VRcX4JyfEn4jynvKxIGI6WChByQM3
VNw7JBjqNvoJb/ap6532WZkQ5i9CSJbbTruqSYCcm9j9b7H/w0pvMiurRVhD2cLyNDit8iYK2wyu
wuIZjBjU1RZyoiF0EM/6OtEgCGlKUrgZVVZn6Wdgp9Lyt1Ofr5AEtLiIuFYHdErCYfYenOSpSMdw
maRALHD09GOwvZS0x0OVu3glNqNfwpyUaYLYNQgLtZZwQAkUnQ75/d9joBdIzhzwO3XNBDoyJ5Yd
T432X1FqwqDQmy8D3X5VLwVW1321E3KBWiks5Cy+VPAobtH64nSM0IQDRe7Gtc2VUFKDBQIdNdPJ
46ot4kzGp+B1oQKUxZlpoMh/CmB6YLx087j1t6mghhPj+r7BTqHwLW6MyPQWmGajZS5f7mT6GGLn
8WBt1s6tKju71ZlWhfvN1vWmH7nOc5LI2yllh6LTBz/rIIWDSZB9Dh0dmyZFJoFLfuavc0pD0IHO
A4oOPT9YjHbKvK3H+thM93qTdMW8DK9eiEF9CjUZ0EiIlZR9U3k5g/hatpXk5GfDvk7j66UXkiiK
k8uvKSAe3nqv+NoZBTeBlxmeDMw+LDDp+MrR+X6LbFuQCJqAMjdT/8Cl+ZAqddrOJcq3CaQ0CRaD
HrPPSLq+KSJllruLfm83qqkQyHWz9arPpauOoEAjlLZ8AKQr1j3X0xoExb/Xa6r8zJGGvOAFuHaq
hx7i8lYphKY4Nhl3sl0FIYqG8BlVluKdW65Qhx6X92hCKmMrRSQgPH0AyAB+GgwFZVT4kNwJrxfQ
FcfdWT9tjGrWbnPhp876KTUSYeLwpKxiGig/ssbIVDuM28gcmyw+fvO3kvGPoNhOMYK2G1ig9ZOM
3JY4OkIOFerQ3bT/AxpcIAvY6p3UFV7LSWgznLmoMg6LtbT1Pl4QawNZd5PYd5xmVn1NCrXpKsdE
SkT1t+RpS5j46C5TGwqsP4ZFr9AVRrwlm7RtCfVESs1+CCJw6wenZ4g/AbN/uYEb3Hf7scqMVE5i
v9fzC4QBX4eExI/H5v3oWqedUFXobJRVrsnY+gt5zzpFxZV8XHb3OLgBshm7Nrx1dx3tT1xs9LUv
IIfCVUyya87OTQzhadKrwYoBFXwBbcX6ifOzpWyBfAdXpwoJG2Jfwb4qyTTqI0NaC/geS41tcZej
OLvM1So70+driZWhiPwAhglvGrA6MoLfORZSHQSQCbRXEB0LXVrk1/kS1d2GE/t6GvbrN2jNIsRH
jqp6HmGfm3y0XlCyIEYCgp6/w7eGhMdBu6jJjqZD5LPfxZiqWNQLPwPQv0eAU6XvhaSaBG51ySGn
I7+8/kJit8ISoFP2Xf6GkED4ZOTRXdFCjmyEaqq2GL81IE7OqM+lDN9lz53M1YveqcHBITlD/5IU
s9FObb084R9NQu9r5wMP79rQi0lBKjxjZlCyTi2iMcEe1B+xGUXCi/t+uLaiTOpDOxOrMN+Rlol1
UEI6gWfVEMq6PEtkQF5IlK11rwbSESfcPrcxRj2nbSy1g1/ElOZsLHgycTE4chBfJGF6tYADk1K7
pr1fcKPoBX4zzEIWNrqVpeaMwl+DOrvc+gmorH/YUbTlkUlY/BMh1gCcPv47Xd7TxzUdd3QqrEBo
zUL7amlrN7y89MXCLwBqZLB8m31rrbuLSLRcYovYNr7zbMlA1MhUizlPEzSV4/Xb7O5TaEkjLDBi
MeGJ9koWrpVl/x+JpAtV5b2dI+iKtXGWdHalaCqAt68ko/yGuCv7kkXXr+dJFT2bDtFW3skAGQbY
EBSx/eftzCBmzX4efcLdmfpi4So7QgVpGnmlm9fCCdXMp6GRJEAwxX6rGDtxK/xpJOwwW8lATenx
LbRtfZfSyMsMtisIJH1NZNAf3GKei5oh6042liqpHt6DSkhVwMXepsMyi+ADYqjgAg+A6beD8tBH
ZNyzLXlNsr6mrrJ67krGMeqDUuYDXUXZUTxvHhCyCdf8LG29KPn/UNoESJRrZeYXeducoIPR2kcG
+SDqOdU59F8h8lOyu5WpG25zy9mNxnnq9KrEKzuOU5RfTO0kJZ0SxX/y7qNuiX09GBQvCgFJrIYC
lqsqiMJXwvz8AEVFpQhzOyb+WtnOflVR6F/qoYF2SfnEYP8CzY9CrTkNG7of7zWkqDj4Kfe4u6Ir
R3JJHnm4AucylJFcfTAmJ83TkRlU8LABnG8l2/f216PTIgDiNYzwQ4LpMeXrVbfWCFLciJOW7+0Z
f8Qpu7S2AspSremWXuErAa6g2/u1z2bMV2SmUdqY8OsFjhGfur1+rZqJd74Nc74uMKGIF/QJscmA
Faoso4aocpOgSUHueJMXyQTItLpfXGzOAOE4Bbhiok+Uy+XJSRlAgTqIMgSyN/rExpfKMWnZvL7T
/pknhywVuFUpWe0XnpxVVGViV2rziouvYfwS8mhICorUZIfLNWiVtYeEj8BzFslGM7/p1aTbVTFP
rTzFYgMW9FZ6FD4gKFDMmBGRNi0y6WxUqPmDTIBxq7dFQWeYKoKBAEwBihh4CjoWD64zM5+nlMig
wo27viqchIRBPQMquC2nMI4FzJuq6K4duytvPCZ4U9ITaVyyw/m+CHksDCv2WQmv6f3jd5M4r3se
qLcBcaQB5F/VdYFbXaK9j+PvzZSD0e6prrSgzqrDOGXxGTBljzh5dCVpe5XHr84iFcSC+ZGf+AMM
SzgXrORnWC1fyIyHADP7uA/w+QUmcXNC+iM43q7J8W4gis0R2Df8yOVJcg7vvXay1w0JBpYZyOvK
zkGH4OeB3DyjA5C0Dftl7mSxnsDOtJ9yvZ974sIsCoaRlTfSkCuvN/LYavo799mk5w/rSPjZYRRA
JlSVAHIA0dlq5yU56x/xib489pwJHnI/2mws1XayR2NzrsxyXI2VS22aP4V+tM2OtnLOGolE0H5/
iJ0PoOuyYVO7SUNHAXTfm/MxvCgLKNfNMalReZ0kQ4qY6d9vIdNiLp1TCFcs5Y6uK+M2htxUuksi
67lsdkpAZYoikuhiOXUrMyq0zlV5KXeygsnAmIPXeJfucaQ3DTWKlOacxXB5Z58Zo+s4sYEKSw45
jI2jg7dvZQa387Zv7VjldHZb6gHhkJX7Vf/SyoRH/jlMpEGY5q+3DCDWZcCSZ+rYw8ohfc6jmBZ/
6n56Qo3pXNGlgykZjSmDjW98J5nYrPWQq9EtsiVdEQm6eJpf0y5vTt9a5ZYAgbYlO05tN+EznN97
B06tfZhA0k3KoHqUXr9DX8fWKtVtmMGJhRznZ35b/DlfEyyuqTZykfE7J+QSrs6BztjWtR68WOtR
KpZ1RKG1jrG0QpQyj1zCLwg0Hb5fN4wofVZUoXfGYXBQODqV2FkN9LX/vG3WMc+siW88WyM1uh0W
m8/wnNaV7ur6mbIw1SEwo2xjoicCrcMl6Y2VwMJxujbQ+9cdJ8UMQGEuq9NHPIXcvKtb4wb6OryY
ZonPrsMqenjJ3pSXq8AQtxO/TX9d9W7IAC+IAigKpNXWQiKwDcW9PsIYrL7bnoHfxsyWF9om22Xz
uC99NWAacXHITxTBEGl4Di2Zt2DKJ8MZi1lD4BkxOOTH2fPFQ4KQ2b5OW6gGePuD4vvK9gTFQ+1/
Um7jHa0SKuB8GjC8IzYef33CVebf9TohsaOAx2j5W+Yi2C4N+1VvuT7lrZUJe1AWxevNX37QxyuX
9t7qYMYiFx6lICoa9LAk+DCoqKOKp1Xxuu4/PVTA//1gZ4OrNeK2JNkRzhChYnCPYjozLX/opMbC
6+HDY8PHwFTJ8S7zDNYcufCl6zvWMOD2zPUKO/bQoFsDd3XfI1Qg2co+XS9Nvz1dfRGRMWEz/4x0
XSSYHNIlHmzzgusIM16Wz7W7Wk5xj50ToGytxOH5AOcZwx+qnp3EiYj3A1DTur4LJ/d+llZt2Sv7
zwjMwFXGKxO4c2xmTKNa6UXfEChQb8/2SK9vWdYOD2P7CyNKtlfsIrRck1XRIQD3WviVuxu/qdFf
wYyyvvaFO5KkSIRLzrt7JmjsO2xR1XKhN6hAogOcKFdjL0EM8+WbWCdFn0Z5S3I/dZ7vrJI3l9T3
jbm5/8sr3LJOqzAETlHJvoFWxVbIk1PBXhJr9+j7wIMYwg1bXAH9/kl6MLoa1caP1E4btOHcrPiE
Cqble8zUE3kZeo5A2LB8e5XH4AujmRqhrWJ0bBNImKN05ErSAVRQXBrNUbteBwFeEBAn7VN447y3
0Uebqbb2rNOvl1Dt5sbc568CCtWes0MpcrSo1kJhBQviHZKskaAVgdWw2JjBA9ySdmRNYc8t2ttH
ElJBYdxBE6TPjDvLQxn68/L4esvy1prHbDzOPnDTu8tjvd5lTqGYDC+LPwFu9hutLbLXSlLiL/mE
N38FqBQp8NJ/U5EXxy6pvQbiCWT6Z9rqu4xo70z/TE6InsQTQPllcrTNq+hnKSmyY8G/Bht0sG6L
DDj+OdNwNTYhLdNv4yBl4hD249380y76VCqHIlyyP4bjUCfIGFmV2R1ef7SjWdFMPfWCpUKM0dTR
qJVB329C4gRqPyzHL7WSkmQe2SxJos5WVS9EZ5Om4cn78cXemZPSunttb5Ytmf3+YjnGRF/pQcQ6
HlLfvl3WhG3gK13Y3RwLslxAKcEeN2zx/lcJtFtTdRCR5+A4I9sYOgyzaST5LhKWSEOzMu9zxUWh
hyPpJkh4wZSK1qc9yxxBttxuIaxiGbV41npIk3XRDLnzFpk8zOagzYNikCw5lvjnRTA8jjD7eGry
meAas4JsJl/Z3HXqIEdbN/yDny8xORJtJ0+Dn7Hk+CtjvdDdJBP0TS2XVNZjZubEgSJVnPa5XOqz
nUBtHwrEIFpazkNy093kJSj7BrG2c4Ger9XzCJJPAD2isfE8Y+QplrBQYlBb50/bJASI5EaLqRXI
+fVpAgj+Ozwhm1+oE3ONhzp6h0rlsfvMsixFJuVbXVtADe+U99v5fVEVK0XS0NN88pv9dWpB0xRu
20qFGJXOigqM3gOFU9CcYIVuGPUDwMHmJpr0kH6RGuXkfAoSsE1XQgjnVIGEkAMBVeIgX0flloQw
dRAGGoQhHwt4NV2TyySzIUZ8rfhjBcL3a3jp8r5HpY7et68cLYeP0TpqhFpf/TpwQ6rlhrKA3JLu
zv2V7H2XRbSmt6VKFwGfDJnFSLTDHzyIvbZiSWEt1YvXIu9N7OiF0bAu/kBT8w/rWEZ7wIb7icib
azcd902CZ4g4BpknRL4si5a8q4/Xyxr2QiYOQKLfww/B/Rhn4nPbD8EqiIJS+xJLrziQ8Olep314
jVumdb3yFL+p9CnuNo0STeeGuEKTqIJAooyfPvBGiiQfo9ju7qDaZyZXZwducw9GOgiUke3OSJ+l
MY4tnKLx4h3nsAAWAGvLw/LCz0D0dA139PxWkKl5+HX0W4HFJomCiEeIcCD1nWh+qQlwZhBgifUt
gcNLuYl703Npo6hIoKcgIVlu1uSsO9h2eHI+egimowZ0YlLqiDxaxFvGncMNEBm/tKC5em1z5X36
ja6nFQvFFnM7ZddTJSVOA81VT/Hbks2RrukVLlBUm4ogOL3YXuA6DJzdj48swJV+choBGQaqVnG7
cljn75DgDHqYabjz6ZljIKo+UC79VS+XWFLTE9Mok5Q6TpDC5wHxrxN9UCL1WI/1Bwgm3Vk6UlWH
gdaKWjBni4USdiFcYvWVtm/hJNMcwrTiyODlN1HX4HnWCrp6ou/I9PMCjEKg0Xsig6goMKH8ilxv
fYmk6X0nQreozMhVAGZY8wJxEsllUobgit3HF8++jO3P9/0ZDdruCaLFKych/GccgpWKER6tuHYh
cXW6Ol+V/Y63m63P3PEpu4wxoCnxGpwBQqMQ2U4sBwYJokX3UHzY+Ndb6ZjPM9j0zbKaD4gGPX3Q
B6gSHZLz/2yMcqwEal6Jrx71cD6PBHf9z1fj2+KTUUQxs5JJDBJYeRaOkBwNxLe4drKITobywUGD
fUE8KP0iP6EMmPMn9doP8RtHsrxdtw7TEjvJSy+p5Q3/UrDV19PzdgQkX70w+jl5wkgs+NEHt5fu
nuL3HedXmnbREOLULC+/LR0BOqDghL4R2AD9HlN6iWsckDUl7v2ar0tD316mS54TtqOiwl6GRGPH
aMZGnTRRQjknu7LOCODxkvpIycn45ozLF2HYhktlV3/0sRy3u59bJd9Sy+IM41QnQqH2uZro7kRO
kNGpvA8aC9TjDiHIfYrnPXKx10hmpz6ZBUkL/xWQCDGamIfmhrNzV6HiUSQZy1cPp6QYfoo+c8eS
efVLLL6uUrNOWBXSaEMaI+dmXzyVKHzSMBaEnY27Y5UOB/PgLjgte7N4cwMMvkgt2MK5X9XbPZhz
Kz/vNvJIl3izwfl2FuJH94MYeORncs5DEPwwE790fBhOwWw8JU90SkuB8Jk6Gj7hj16NDptOFVZH
yZjRI7E8HSoDxIi6/Pp3YaapCpd3qb1sO/N7GxB7Oj2+rspkmSdEO3zYw9EAhTvMlcqyytcfBJie
1r58dIMojsnWTo2zPuVeu9V+b+ezwEVlUIfe30JSiI66IGFFcqYOmKCvDfBFPz9CXrZzbt/2bGY0
yZI4iY9KzRrMtd+6T4YoBc53P26efEeEZLdZrhPv2Dmv3C4ISyS3qSWn9k1KRLaC8FjHQZ/+KI1P
47lt0W4p3d/g1Qki8RppxIyP3zqv0emBFEM2dV3rMbjGdldyTjGH4+BVXzg3EtwelFYa3mJDOJ+b
xldDfNUmxdZHVzeT18FvEMLMmct3tQ1cXcbYCdGqF121MWLacyZdFgOeCm3i80TXV1l2MC0tPLeL
ySTDMRSOKfygxlIbKv8c7BPD5xXZyeBeX+JmW2oXmrbyRjvOR7MKIKU8eFCfckWhRa9wWFixcwZ/
EHyEZC7SBlYf0nIaNmfjTUk2++GcKQGw8gLuRTzDosvmITV6IOFOCm8NJQB1ijX5BloxmRvM3Trw
jeOZCL4ewE9sdM/W4wLPeKOc9t1Dp6/Lmmma1B5GtdeT3dczb5IGD4J6JYBREPbLstTNNklrXg4T
a/tXdfehDLYXQEINGuMSpWP3If6942b7PqJ+H6+quYpcptYKMghsUNmEbLNHL+VT1HhG6dPv5jOT
TdKogg/Q23wiK8qJxdnDprxvI+r9KLTOXy/F56DsTT7z7g2YOnnBa7+c0jsyRVktA50bQJiadwy7
4fJiykUCldi7BNnkTj6Haj5CKyvofvdoZYf7Bz4+T637HxxFCRmPmGCsRB0jwLEmwwQc2KfgalJG
o27hBMaZyky3bn66HQSbz5rpdWmkegiDON4Yy7gwEiONcnDWOEEGb6F0mqqGkev3TAXHBK69bqc+
9ajEbcQVMYYhl019Ey00jR0wrNVd9qsW8NJUKD83Q1kj/NiBuJ2WkppEz4V+8Tv89exaxNnP8Z6t
bTp05AhS0ATIGTueDhPXUM1Sx7QwqY5kiRcgfsFTfQMP0LlVP4EeKmEJhXnxReOOCZcWy62lbl2g
JJXl0WCon2rQB4qIkRl/5rfdaAHSH2ZhLRFpmCEhaGw7yyM77xksbkWVQbMzydnI5EFzzqf2ZcCb
J4kh4GPgxI4gf10sQeKcZ7rhu5t91vLZfQQmzSWm0DOJhQW+gmAqPiddRfZP75Bwv20JOcey6VCd
bOJF1tfbONiD2PUCqrAVgJfV/jMN/mCfg+3F2ELjhuwt1jdlRcx/IcQsvvhzb8w0KDtfGcKZZwA1
Jf5yqTky1JPvhNNoaVGKVbMRpwR4PN+V2vMNKOfKLIx6CLDrcfc4Fdg1riWosQp0tSG6P6C33VFi
5zH03QnTYy0uNG8owB00CrFuwJt0spECxjS8GyMZdMYTISVOzF0swzVvVEPUpS9oC78GQ+nRzBZL
cUboVq0TpgWJH0Zg8n0hEeiiYVyUWzwWuXC+euCL4gYdJ33si88ZX6DUKUf22LgGZbjkroooj1yf
oUlNtFnJo67hZYbr7twzJfBFyOd+Q4s7XqUEhVGSkYqyQ6E51f8lbXiz1xtkjj4Z9rmR4xp0bbYL
zma1TCmh6WAOD0wNFoAjY5idsSymrwW/yBshENWo3oxxwAGxvGpkdTz4nHlUEmQc73YV/zlSf5ot
OI0LilTLcR4MT3s7gwDeGhlZh8Bznt+f7nLsN3uoEnLuAMgK1bHm4WliBnEYOfzaWzWh87BWXaHh
0K/9/PSL3W+w0yuSmm1H/ZWyA6VJ0sYNyHV4n59qWjHBXQ4YVkYk8bpq1tR5fxml0j365SkRfgkf
0jsaIbJAttkdZJ/y5PSMG3tKk/ATVeiRg/17kc76rECf3dVcJ05HabtFsjcppt75FPXsf5HfkHGM
AKsosqPtEa3PZ1+84H+5BHS9q/bI8h5ADNSRoFYml2J5nLvUem2bG0RKpOkwGPznckZI5lvv3+PE
6GjIRJT47+dGRFZ7Jf1MjoYxPSflcDXLcHVXAwHF4owuS24VeFU+PyMfMXc5HE01eVtyGuR7ld1C
Pstkz611LDe5GFyRIGFkNG9Dbk7Of6oyPTHB49QuN1jl4wNd+srTNlsRxUC4tiABKWu1+tvezS+q
i9XyUSjHb06yz34TbUTncbWYUSxWOkQhpEz9G2R6blW141I5CQeibAy+ghJq80ceI/9VDDEvstnI
KHmFuDMzLEXTZ0Hq4XRspcmhRGDC6c1ZVOJPval2rnaUsRnk3cCmG7w6clIIQtND1HBUSBEWr2IK
P1sy1xcpsHWvLp8ZvoiPE5OIqselOWNy1ZQFe9Yh05wrEDGAKGXJt+M/Nbi7SLJekIf6VGn50YeE
GUBHDBoPCJdbL3G2Cq0TWIG5QcIfTo6FzOKZbsNtLgejPDen76zkl6f6zl0rMAaGewivYXPMSfRM
zZHOvdqQXjE4F6NY/l0x5WroLvj+Q452k4ptAzADwJ6ln+ztFGB6AhZT9qzkoSPvx3awz6XGJril
CX+JFkW/kFR58waXBjS29J0AVgWJFa5A28OeEvoijlrL7wx9gGOLTwTeWnpYOD2vb6OS1gKwS4Sz
LObdIUU6Jd/3YZonnexa/XFx66VUR+hz1aPZy/xOND6Oj5iA5/Ie865gVKdsy6gDN2AETH/WeQBG
aIDjGItVGuOOhoB0X6QP7hNgWA3YpNoWhie05iF+BDtIzXfTvSH5k8lj0pevfk3Q83eskdJS8Ulu
Y8+ytYTY1t+s2d1M8tbn8/b6idNXdswBExBx7EwjwQ8Twlz5Gav/Tww2E19vc5dbFu11iCDtLt35
PZqN6aVlgTjEwjLrHOw6Z82GRrYJcT6poWml24isGV2jR2a8EO1CC7L+YZkYihPNDv6kB+bgB6pH
oRIJLHfQpEjSqBpuaHJpKGSX0WTwOOE1//0TerC/dS+UXuIRHlUfTtBsQhkJQDabVHZWN2zu/OZ9
6Kjk1jRXB3zPnYM5g45gDu0iXPS+RduXpxbjKTCvTr7zFpbJzBUINSc0RZYYhKoqzjN32fj0VIsB
qHC6CsTuaKwafDo+ZKzvxCMiRhvl28Aj0zmMBqNifMhv5jS0eetsZd1zB4tVlYMBpsUEOoHK2w37
HAUrlFxHyJSXzAwdDbpxFrB/rCqfANV9nSSnRuHF6faVruIaHqcN4sxgfgrucFy7v8ZyKJOi7qeS
qlYm8JpSNoNDJIfKvjNEV0OCiUaMHFf9ofiJrqnLiqBCzw1Tc1QCk0+5hSfrAlhl18LIJkBh/+/V
uc/mKcgjXKzVWYVDhIg0+XarFQ1eh0hdXFuj3wR7qkkT/zUYONEgc7nA6x3+LPH3T0LZpQzEQ9FI
noxdOSp4RYVcNtLuE0XdWGLXcZArKdllL0mF27cvI4VqS+wgVLlasSdWNrP8a4HNOvLc1H4UEjUg
5Rg1lrgMg+EehBGiNL6ZjrekqcnIIeHqs73bPrdKkMUqY/21nAChdlB2eAh5LngOguYfCL07NbDR
74Vy4BSv350NfNm94LO+VbOi8nuO0yatwmSBYzw6/wlsRWGzPwMMF+cDi5LS3Aztj8WFab5h5srs
lc+KAtYg7TsgSIlFqPMl+VQ27RxIYrieQI4kgxxYARLHqxG2fwJaxAPgsw/YfA8DNCE90xDNUDF9
T8ase+NnGq/MpzW3NYZiwYgNWqhj6vu8Cl6+/6ArR0oSDrte5mOASt2kS1wNTUolXLaBribFTR/f
6yDq5RfoAayWEAutSlpV01U4USKSVPd4hGETnanJODSmDihDb+lctZWPyb7ULXGfCgDNMqINHUjx
wBanACipZYM2DxSCf1ZYWC/Ueqc3otjmblJlMdYPLlhma+VUSQ/uXL+oRUtQt8si/lMNMcnB5fqW
JGkBXiM2lCNLswjUHmaoYh2VZ6/FoQQ78J4e1BLjalqfmQdpTe4gviFwtB/ifhsojRWy7CGwb5FJ
o1z5GZkf4Avtyaye1sFlL18Cs1FHI4Rp4i0Q6AqrkUpYKNqEd/EcY8QsDChbgtNmIgqF+Pk54j+i
J5fhsYV9t88/TC1ZngYE6HhL/Gd/uBtiyPvtLC8MqKcdMhUMjkH/oIhD41Fo8aE9r9K+HLmS6fG5
/mMl9KpbXsqis7Sx5C+kK/Knw/LnE58ll+Wt3Cs7yeAIzUs+DB0mjCM9czrGOuIRkYi/zJTPqXuO
I2zKShlo1XTSJVcCMLo+70iZDQS1y4miPiXNjo1LkMgdbNSb4FPWNx7iikpWtLM5vxkrqiwIao8F
jMjEVxXpEP0RmfLKj8navZPoZOZnKcm7MGOFHDyOfK4opUWUk6COIMYG6/ji2KYg6G8x21Grx8mA
eKICEZSCqwEAXXI6S4m3Jp58J+6XAd/cTOkPVx8gBbjK/SkEJzg9ktrG39LjA2Dw3OZlYuVKZzUx
8qVGRtFkOYfzpy7v0Nxrmc32WqEaW632ibJCvMSsTMuNZZmeFVhMS6bsu9xiXsW7/XdPmGksixJd
hXXLaYEkzmBo72liBil8v2ii4bu9yAbZCeuM1gZghUkRXkaox5fMurOxDMrjorl6t2YUsQmmdbHE
X4CWZVx9ux9jCsWZW7sb6E3/Flth80Omb32q93QZZ457/ei+KQd/okccbVTiMasyUNmUgDbxYxxA
kW1Vp5KlOS3ixH+/Eft3M3BuetYYz6s55V9xRIU+AizLSxbw/HfHdQszetHV8/d8WhMsvYNmeBQM
5liJJ8thpJNzqrrLHJ8GbOteSjNsOH7mUQPOD84hqtuf1etROPqBGyBoQ7JACLdeuE+GwxJw1/yX
1sE8JsafMJmNo88uoWuxaShPow4fyh64tQ1bvAgfQZNNmNXQBmGj5Bm/ftTuvXUXcIscCOkzPT6s
wQmImXn6i2c487Mpk9wjfQHb6RWOEfga+h6q1ENUsjhcnTfUqK8GCIsMxQkLoYH+QIb8aC6IHPef
wvOgO5INvJiwXQj5bZPm2ebqzPEXYTYlNiIdDUGapHqndDwmmsF+xTXL0Ejg8T1dP0hQqyNevvlZ
d9erEX7yFFQED67rDrY6HMM9Us6Axwd/kHpPjvT+ZJbBq9K5kPog/dWX98xWgWE2VnMrr+nDQTxj
4nPvhiziMbRem9IvNQ2vhzmzS7NkUaieTDGBtuE81cw12E0ROTMwFaxxoy6skAlUhEs0VMd5bPhg
oNFk2+EwlqXel8hIiHN91/A0K1jpjyUJanvYpDh/K292NVTnq7Zca9k+xPQ5o7r0RQnehFyquzeD
F36JOavxaxlDyG/hVIJlc8IQDFb9tnNpcskGH/rb2kTeHywt/AGwhDIIkAF22WSkiYRPiPLoftI/
ktY9AK6eA7Ztd+TFNHcx7JgcDSz+vZTy0gtIwdGuS3FOjDNHfq84Vnm2TzBGBSZzVCkYowh9NcER
ZJROSwvqZ7hkB0q1PRxw5kDpaV2U6w07OkChZG3B/OVkJ3MTycw4j9g1zsu7jrLyWXbjQl0BRgCy
YvZoumbBCoVtgnIygiGle7AmMr9/H5k5TXECRIvf9ocddrhZkYCtC09r0P2D6asnAfeM2HS0Stim
/myho4itMlMw8712lCPzO7WD1sxHGhy9+o6dBFnLNcfImhZko/Sezuyp3axYO+S8/SkDmMaxhYZa
M6BhqglMQ36Kzg1j1k5UxXsbNq9eWHag6Y0yFFQl7Wz5An4Wipunshgtta3SW3D/PQvav5E8L2em
AnqWbFGAQLQPbnQN4zqJxl/2wbCN2RYBuYtiH8Xo6RlF4RXsoNQ4Ggd6dzJjXuQAVlANv96wcrW4
Ts8aKDRUjuq6p0FZTw/iD3KNnisERDgOh/Yw3DGP4Q9PpqVERi0c5U0M2H34wKDXwr8CpnD5f8dA
1g2Yg52RAnVVlNb+vEggjmvjlbFcx0rZcfeXqUhW50ZldPCu1koHJvHtck4nl8RgVMAWV0uMZkK4
aiD406Um/f/UQWrrsmibIe2cZAzGOHCGADbgAnFkLukH/460p4USh1K87mRa2xE3UYeEb4kO56Dn
cOp0QFm+gBzV2MeKU2IpWr5ecGHsRc7TVcNeZ7/BSYmK2SI3Ml4A7OWTPt8zB/syfTxTU98Faior
6/1X6gOs0Eh20PIo7q7qiHr9WRBGK5HAyz/Y2CzPYMcZgaGHqwtiKAfDxt1J7liJJj2Vs7R3bvO5
NZDvrb+C2TMQojgKSg1FA3ZlssxY4vlALNYvzF0UJXUDDVbQsRMUK8nJIFKM5GnlYQCwy5jvSnZY
PN4VaTwqA3vvUDlF5R3YwH4GegebBgTSVlHj8MNUuavhwe/ZwROnjWFs52OtGhVtmSzpNF9VqDWE
6EatFJzz5+tmTJiO6d5ap0G7ZPzRD3IJkZfWkRL2SiSaSJyi/0uJt0P5oCzJwk9JZiVIOL0MBoMt
oPuaqIrJnApLI0HEynGdTGuDQnBfNrXAd6syo/CynyEuGAwUhFsaZYV+AAvW9AcSMVyGCOJXu/yu
ayyVfpyO3f8fv/R40n/7BJRfLkjQz8OoJeXktdBWozFmCaMzg4Go3PHwrfJEEF4ZS+JJ14DwvsuH
x3AoLS4DfPhaBCBaa7pu3d7EVE4xQRA+WWl0u74j5STNeNt8Trd5mVxPF2e+pjxSvLa5fxr40hoC
mEa6NBwZONVyD/n34SAG9CzWzBEQhQKS2rgzNAlIIUJOsKjErQySlZea0Cqo7w6eNWSCfqrT9+Hc
4CYAk1hBx+95KPQ3cLwR9MlvXXz1rQa3JYh2CjOR2311/dSzFcXzaXraqYv+5Fn4JuBNsPv5b1lR
kOQJ6OWORKrCCgLVjGu8bEEuPL+UPVJD9HMNcH/3kfKPIqYXxN/SIOskpu5h3OsyiF2Y4P0r8g+g
VESyb0BTTOZnGcsfbKpIRCvr871zHsZPaa9WCbyUg5pEMDn5wcxSq+yqDL9zB8jMoM7z2YVjC2fa
ec0z9SPP8enisJweIXmPumSqbfSe1ec0dqF0ciiPobYZy7Se9lls1yuf1Y7NPNSIz6kx4CkURUaQ
h8ZmCtXndmTCakdC/Ea3n8W/3oMcM3TZ5/cDwGzvEofhRVD5I4aeMfoq7J81jyzU2A7KzRyaWL8y
8i8USGa+KAywxyNdxZiDCIEv27+vCUBLwWim5gca4XlYE1zH9Z3vo23EfBTAee+etaPVMmvzt1MW
C8xv7kVx0HDOO7gjPbcYLVQIbPLClNkL922/LXr1q7qektcTxBAuYQ4vUCtZ45J3nbM2AVGJY6iZ
ehzvE3upK3vP5Cn1lbty1ORNOndaHexg+NM8ce9xpvYqbak/i9NAHGvDCKa7MFnpskPEqWDrokx8
OI6rc31ERfaB+aCjDWgbQwzwMLRUDAW7rBcLalQn1jDvoK+7nvoKEXPH0911m1pzWjJLmkkxRMw3
wlvTLlTkpJhiP5zpTcUk5akZDJanuJovdHkapYR1ffJbZO4Uqq6hweG73HfD0xAUGdi/vseFMz+V
uIkcwiUvGJaESt2H1eeF/FmZCrW8oXsbFV1oVRv53C0/mWSuuVwwsT3xncgX1oyEeTpR5s56SiXT
kixSQ7l0rOTcjYG9+eul4Q2kIbh1JNJ3RgbMk1osWRZPbbREdBot2rUjXfnrsjtGKKH98g94y9qz
zNz6YUjRtzATAs+ebRqQnIIxKqSgvZuYgfi1nhc2ISK0FftJ67rwGs1sZJf08Wv0lVBjs3kyesyr
q0do3xTCOnpUNijGBuSHGD1nNbLfaiKCyA/lvnsllYoSuuN68Ih8lKIRiTz5F1glhcVYsJQ4V2f8
b3mhvwLksSkPPHCXf3M6xz7eo631Fc9OO+3oQomuCiWt7P313/uLock0BehQZjOzNU+vbxza5Uga
KHzMTa50SJuIJvRRKoKOR3eLu1XhLKtbGglxtD271R1suG8y6NX4d5MOWT375wAWF6Nfa3qRWfDH
bf1HgorZger9bB75qD5/1FMn3tQoMmOJx6RbrPEN9bFGFL/Z5yb7aGAgj4dH+ZmgVb+8H9HxD+9H
3NsIl1DuGaPp9DXIyOWgXoiXUlz9rr5TrTjrXe17fa7RcGSebyl/gNxVMrHYkEatg4mcPkHCGvu5
61pQvD2TfJxEEYXkcnQAy9bSGslWL8AbBnh5ILQIeeQIEMQNCFXIin47hdkBQc/LMeh56NvxWQq8
Rc9VG0JuB2mlnO9Q1E063/TCiqOSQzM7909cXMvGKz4FpzAnGcaxzOIrK1uN0jgm5ot4fw+pZgjI
cGmqKgxco2BVcyB1Vhv9MklblUt+QAF9SQ13kUcT/phOOU8UbM0Fw4H8l3lZ2opOnOKSZa6GcDKl
YJrCCpiLGuLf3RWG5vUWTiO2B4hZ3otJPqTjEdF4h0s5egoq2vH/WYOR+Rge+vhGKN4mneb5jtAJ
XPQE41qO/0Y5mNvyrHjZNvI9B+7Jrfak8fT2CBkKyuAKdZBFhVU9vVpJDRngwn4fQyvvF1K3XJCY
RgWNTpV9lQK4pCDvVBUP41JR2XiBjIHaduNbyLVrqUVJIWI3xjZGovcbnQZapZiNh0xLpkyJiBL/
MnUIR5kZ2dUU7C/y06iLdqXdFQ097l/gnv+9KapmTjrQ9kAhJNJgCo9eRsd8F2GlPJiq+aa7CJsN
Sd3TUWKAeETGHUGHBkM97ZbDdHdZ1bXWQxC2RS/GJwFoGe/SQuG6CvEyaWXUEwBl6B2fDqNKbHkw
AA3lt5bv9jl83WeB48weoVtktdHEpzhuwt4PNwQQUi20Mo/IDgr+WmME/79B217ek3nI4/MMG/e2
OaSxXv4jyyD28S4dYCw482p/TiGCI/BnFDWXYtfaVtxmdMoXQ76NTIbiiHaynyhM5YHbmc8mtjkj
JeqIUPPkmY/ILcOhacxnxIWPV37UlkoSTfzw6eSgZtKZl8Zvm2MBsJyPu+ovantfF/blzkAzdTiC
KFVDO0ljsHYJlHy+50rqjtyqMoHcE/ndnlqrN6ePmZoaXtk2dnF8YKwGihKA425/BELMHk8CeQd3
7fIAm9DGfj9mX6dMwTRx292ZrmvOhz5a58pzmYkxcBtpwYk6mnNWKnwJwsPxe6r2D9pW4KLmU19N
PYyS2hww+Y2BTlkyJCXpb/a/2hriKoqmC9ohF0AdiqH4M+B3QIfKSwKK44eAeEXoRHxU4Yx7MRnr
6NYi2ZSaGmde3IX5+KRBQCxvVsGQauGCjtUfeSQyEal401S/0QP7Rs1L7VIR8R2K4dy3r1rWQAYG
O9vwL4qDbp8mhQ8EWEij+7LI4fm5OGRqJxY4gqkwC1cs2cmAgG7Q5Lr1OS4/ahR2/Xtif5Nb2SXR
l9IjpZr8XE4ixAzbyeoyKQbBQsIvlADb7J7Dn8tPNN/ck6GF1S+lC012ekquJOd+Mt2kpPlmMFhZ
KeSxYQIOsSo4vQj/i6U8dk0bhLe3eWkpKRycaK4HW/edinfGJvkw7SsRns7eBlQHL5m6kgU9AW2N
oVJIOQ0e9xMqoKB9Wg4YrFSo5suQ+0ukbqKMqJV+9Zp7oXkxkLOqnL6iH0i8X5+hMNFZ3sCwPjpQ
mJDQmUjQ5xF4geg6H8s6HY9p/YIiFc1LtRGBv+ZHszm3nGyCe8U6jySyH/adhaXRVTqXS4/lu7dr
04HCmHlKBGlcJC2RwsrGvVtc9qtBQTackZixDm6Ei+lw8/vYUdOPOW3vamL+eIkzj+ogvBr0Sade
iopt9N+EEKUpyyEdg2n2bXgq34seHKghnV28WVAXltRdowMmWEUSM4T2QzpCXNYb9cZHSemaMm6Z
Mp+5ybhJlBWyN8Is1T8AW0UpYHC3Z+NlXxYCfR8FJ4ra9uVpx71TzIJ0yR9d6UVPJjfobR3DSQCZ
K+xhSnpzeaab9Nrzl4tKvuZFYML+i0r772CpaaQSRYaTCQPEjSzcmotYP0UeWarif/l8YInDbqG+
5RfLFgZty5i3kxk/tJOFlaHKUGXB+akFi3nUC94vAp5YJvzERTVVed9VTMPXi6Wwkqj6PwvTiRal
qW/mFAwCabK7sCIsh+MGLnikVkoMxjzE1DGLKKU+Ov8IuW8WQB/FbNYCucVHkiMGYII0KmqO3IWu
FFt2NS2kUrjWRud7wbo9cjnV6laCB7fYX/sThRsHzYvDPdk7hdgBw5cHv2JUbJjFQqjgLHv5pRPk
kTdeP1+RZxjvLXLf13zMX+ZY71275xxfgLONjN/C0FbxxsMVotyCefMW+RpbG4JGAKA/0dWgyoOL
xW9V01g3C2bl2teRTgS3yAOqPZ9w/ydFt/Rbp5D31TXTItsWNMz/5qDnWkbdTRf5F2tmJTUX1/zQ
8JeEpZmiIDyTqGikHXHE6xWQhKmb1BwFhhQmMiqNnv1ISCXxzY2ctb9fSkmI8fRXYVScVH+rXfz3
cFxLpvP1ptfKS6IfLbZikA3HNNTDQDwagVcySu3g1Jp2SghWZtbTqBz6jl1bU0nRX9OlJ/Q3P/iZ
9vhBqCwtkIe5s5b7/Zp6HhpmEK82m66wTftWLn8pzWaw1v/zuGZnuoNYw7VhHHyLyebWp8IQb8gK
aGvewgL6i17lCPQRtRR8od2DQxHou3dLvbioVhRYdOk9+dipmTPdQHZ4MKdFg9LAbki/vKoU1yQ7
fKOWDXd0/2XSeEilUHlNDFWBZrzb1e1WkijVPnOmw6CZmJ5CjuiU1XfIKfdCyc3EmDgs+wmEimrJ
dLHrSD09Ut1e5VRY4OrJSDi5VMkQE772noEgSuCYn/SAvoVRA45FXcJo4lZJYAv3MyaGXvMpZHwG
yIqWfME2EQ5lnyvzj0gUsoODXiuXekb7dWCw8hmYNWrUYGwBr3TsitW8fCfBjaEgrx1XXChMokVv
gtO1/I0u6qYf7zEB74Bot+L9FQvjnqljz2EpcwzZo6pOJFOJzERVBbzNSczVuCbKOJlAcS/IT7Et
jCxz7M/mB3ZJ9KcOPtNdRinkmonqp2Zgc0MPbsSa6A70x+5UvD0O/PgRMH6xGyRzwQYunx2DRu3I
uSSE/iQUn1F+5Mdyz5QRQO5TIE+aDZqaUQd54OoMQY26s5rWqRrM5SWOTJzHKUZdB1f1iWj7A6Z2
d3HcBSi+kC9zJ9oVSkUyh5pRYzZd2zMIkxRnNiGwmw1edZyVvIpiEmSnEAIqUpU81+IkD6xSLQhZ
oBiLzPGgeofZlWoszyWMBS5ss0GEt9vH3v7u5DKAmpTZf95HKXdSvSg9Nl3Pt2zqTolDOBFHXfsT
WM3TUFE3+tMfz+vap3LOyDOgI5U6T3xEbanMxGLCdYj8M+R2VfMLuAaKBqpYIkEs7CtDWAmhNR21
gokatkZ+QIIZyshL7B0d0XR6ffRfX5D2ZLwLzO07Zb0XGAXSVCcqzyhQYCrsj8JLNEO+wMIdtAZG
LcPXWfyEjzYV6guyyJsGMIFOSZmfQqk1nMYpja/KyOyUk1VItoUXd5ylli1V9fwMKaaoib5U/E8Q
B6rBEgs5B79ul/nN7VRN0YUgjVSd6WLZVs1lxaMg5zrrudLCHJU0k9gMfDLxmYIQxrJ/v5N/vSdD
FnCGxb24qPpT0GLvJhfnkyRwZwOuSFwqFZ1TiIQTxm+vREKgzJz/AoyCPybbdLuGSM7nIq3ub7HH
D3JALWuUDEAJKs4LYgO0gLuwM2PELNsJ666UOFrAL/OUSxAtdO4nZK4IUc+xLcfpUzohADZCY49J
O7inohFYt96zhb8jstRQmg/OJITA6f2ld60YV/VNz1Fk0BM0s6IJkomCjNsoQ11IuHMEA11TXu0h
zd9eXGylwuSMLtWoougJV4sMxDN3zMd4YEIEJduh687C+Miq4M01dKncRGawy3/spNdze+MUCFbw
/iv9zHHvs7J4Uwhqt2gk1IZ6zLYe6JTw7S7mRELz1gSnuTkai7d0kFWaQCtYZDWHjxUoSdPT/Xgz
khgBVthcj1AFl2lq/Q/oH5RtK4m9K+XCBmyqAOHvpiurO84aNwtBYcQWkkbrhiKbyt7F03QVxvdl
6FZBlOZ4yglNFif63wsy0CTK2sT3mTYdJ5RvNmDkcNJIrNkYXnRvfoG6d5K8GlfSYfMdmlUGWNff
DIM2YXf0/J+1TgtyF7SDXkpcoO6osYMIqgT8UQsfIM5f7ibHyssijiYh19S8BzOarAIJXFkpnHUV
jDQVr514sa/oabx7APGQOH58UzJn5H+xXm2yMdPw8QQySDn3VpJDmV+eRSQl0xI1fL5TJpToyBO3
rK3tUdtakp/lYeYY9ntWTl3mhedhvHxeFCPoEi9GRvhuOfwlzPXXm8Y6lbrwBxXmuByo3+Ggl1hZ
G5rQkLoMjOWhJPV/mkwFQjVN3AdJqC1xVx0V2HFcHRkPOaI32W69SX/nglGcNXMhSUUkrRnJEAdy
OaL0XlbqGEl/xKvbaTdPs1rWOljcS3wWmd8reCsIMQd6bV9xOHSzBfrX8d6kSudqXzbUQVcVKZKQ
A7ih0L78vjZ88RDQORL8Y1FooZ7M2HZ7ai5+EUEhLhNq3epjYC9TW1JTij8S4zfS5EUdsXkYAgdQ
hjp5dwW35IZq1iPJvhw05zUEiPOGmOII0g4cCxrdbL7l/Py5EoDV5lAl3MZFxg4B9Vhe6ZHHhiHM
wkV2RxNQXg+I4W/wx/diAFfNS4W42QJH1Jw+mLF+7e6x9dffOYtIgOADqf/0yN6BMFtIYTPHaBIP
rFLYVuFRlolImi4B2sLD2ZIETjiIf1d/TG1ZQX+p1R/sFqwoX3GnRpUUcaWs1X0yBUnCXa/wVVTU
kXx/skzcisMP2TjCHOQtc0eBTu1wOXT1G9MU6n+FinkfnbDeAevv6vbOU+V/qjTkBpbwXhIVOULG
DFlN/RYa3mzCBO4jJP9t3u0twf5I1EyvXhtsKx9AgqHeJvY3nzLV0ulxJFJf56iAhCr5KkeK2uBA
bwGjijE4QjQ8DbwiilTX75tqutv/cT7GV2pOkN2W16dmtzh77gX238LHRvSBrImJQXZnfNNz3Vl+
HUNNtr7fgPyQdsv9wN2wsEjjxOrH31f8lNTWLxIqitvfY0gDBQcGTcDuwzIf2+edGlo6rwm6LebP
OzmR5MdWlk74V3BWr0EpXOQ/7/AqXB6lzCh5AcbWcyKLIPYQGdHeU6cqC9Wcq+nP85xM4Hej2TsB
mjU4w3RRawRaKJhOveFqniRuLmvu2enxhom6NK0KqaJN7asbMN7PJFOySvBI7D8T1id8wPgjp/yP
49BmzAQ6A3ZFofixAeReDF1av0/+g/XlqhFNylMUUi+qFqTtXdGUjoVD92SQiBdVnjPcDScCLwx1
fg5teG3/cMAT174ZA5hgAut8frALRpbXVE9AKnG/TBlvxUTcjeZK9onDHMC4RF5l36m9rPRH3Xo7
i1F8NhBamUHC2EUqfmdrxYgwZ9McInil6jKhdLwqnFjZF9LgQQKoOiC63N7eLbqkh/est9hz3j8x
y/bIqpUe77uVV0eT/RsTfc8TXSlNUawZ6hGoUxUjNbAOi6/acRpXwFuyeN4VumnGVLIXqBuUn979
2ltj3C4wDYz0NvAkmKezIdXyotO8l0g54tfpUNqzjShGCcrLEmXtpfsAiakNxYdiA11Ix57xHf8/
/Y+2TgEG3A34Odq4DFMOXZr0lDtTXfSHPzx28QbLCWcXyhN0dVQW1S9FVyD7Fyyws/Ik+qh7qzkI
kLl2Dq8cn60wx8ZyBvVxlXom3qzUxSK2Yq6Orw39Q3MF7wXC2sZ72ZEdkuHdFpT6uGVc3ndxjYK8
T/Ayh9BEDktlKz7z2tUpDPrr1TKlCIVDEXAd45J6hxf8mgJ24XLKcNiP8Qj0irwF/e2y2dTtZfxD
F1b8zMqr5p/i8xLYTQXhnbRJoRdipWqpbEjHxCSuIZFWB25Cc+oW4yZEhMAkgwxbCZRG2OfL6XhS
UxOQkBVYZwHjhYvZ8NmU+UrKCgbjs1pg83aUPQyfvf+72FbcycNP2p4viElL/hKiaYXRHOcXTSFo
w4SvMXbkOUz2UBfcwCOaPgQt322zgQusoO/O9Ato/mxxEfskB/UXUq8W9X1A8mz7/mcXR02WnHjW
rmjouTq37hdVzi06ICoUci4afcNvMA+JG7nmMbVYF+lKxqa5cx0BIUi5godTE8KMLOyBWsHFGBN9
WO8fYdxmBSPC2vLS4MU88DRPIViywe4eRRKqJndb79ebqUwfj0FGdAynz/+moRmD3nBe5CYoxrIg
Cl6PW28tF2Aa8aP/pM5HJBVm57AcKV9Yozeu6qkqqYfjbeBfOgmNI6bCXsxkN6xXboc8cFUTVaNM
VNUnqNheRhZnr3aVr/NhB8PxIP4FTLnXKf1dtruAqOwF7GPK2U39ZJV9VMzwEmL4Kk+Ge7O7NXdn
lW4fIUXjaPhkHrqp8H1bv82pHQq3SeFmb+g5cBvOM0Lv1c325hzmZn0RlMv1kWxx0UecVR1XlLZ+
3JG/yajLf8UZ8rz+JrmRKC3kP0bU3IzAp8zvV7Cr1XtIjzJfUYKntI+LIAknyDpUpDFuvkoSKtN6
mTNKDehg3dec7QOVxPgMIoOHFHoL/3AUU1Qnf5eIvn+riC/JAkOlEevxqSNgmZNXbkk6z0BDvEq1
+njS0B5fmN+LTSVytvYZgyaBkW6PT9wuDBhxt9fxP/eArWbF8ccQZGgq2X6Y0wome1uytnwpu6EC
8hQuhDsgpKtzTq2sxVBM1SQxQEO8NbZ96yNZAA6G25rA+B+bmYSFgrEnDeZW1wJykp5Xl3mOLDUi
zfl2BhIuh1uZxLohcLjg/KABF1a8qtcUx6duqbDOxPt6PwEfSwra/0xzld9C3jojATQytptqJWqD
urUF3nnVy44O5820xg6+v1MmII+12xhMASoZHKEQ7TGn/sW7eaTvLs+b1InudTnYfw4LHAqPaZCS
obP7mRDKurWUVKXvCuaDK0sd4kn82IFEy11GZKYdxo4RpBtgHAf7v3zpjcoqZyCr/7qxJlmOUjFW
qoDtltzB5wn4U78Ph6bXuOp2Ji12yf1Kaa8AQXb4Gl+mt/EZFIm2kKBZECaHzHS8BkQ6ppVGOLRB
JZ0ZaJ0B8jM0crg4/H75UC5SANKz0o9TzqBv/8jMJ/zwOTs3E5WSpZuiD43JExmfMfM1EWMy+1xA
YZbd1DxN8PECldlaKe/ofsuxLjayaDGQ3Ti5Y8nfGAbwUh/EiVwRMZ3RFUSs/qx22ON51S+ZVqME
O9SZw68vwHLCog8TvMVWV42HdJeYCFY6Bk/RVeKcQLFa10S6zi+DcAfPZPFrO4ktuvjdYr4URTMv
pOqSsjPvhHCrXvygYNvzb5RWysnbspWN8HvQ2WFrCDwLumDFhb1uFAiIZLmQuX4SQzRSDHiq7MKX
KC3AGAzLU6NnFPqWRWrzEeZRt8E+LeoAmmmSiBTYpBrGp8IAZ0eWBqa9m7tobiYlV3Vx88VHNtSf
y493yYaFW6k8bpyqL7Aa96BMY9jnLsycAYFU6waBtNOFSCrQeCzvA2/BG8g0zlkAKzrDfDTqIHEq
BKyUavQbMBSiJ1YAFOV0V7+WXSYuW9v79iREBQ3NOigrS8JTGigYgmTgrkyjIXlQ95uCbbmcZP+V
rgbxkTkkYuiBuWnNGanTXfcx7XCsCwgVOGmGJRc7g/Yv8M3z5y5P3cOY/etG/cqAEZdYC2DWeggn
Xu+h5LJcO1+fDwyH4AZrcoXQYhTtFUNWG0zeMKSGOmwADgvLjWQeWWL921pQW0ubeLzkXIkuYn80
aMg1ta3T+fkedOuvNyGjTLTHHF+eXsItU2mqq0fBTSRydd5vl0yLj2Nmlbx9Qt+8H/BODG0MKxWq
K6yjPCorkogjXhFMZl86/1u1OC2VEA4J46KM5eHrftomDXHVCctBsVR8k6gZKpY3Ns/oomtdtakj
m+IgA/9ZBPq//LKDQ8hBZlYEDCA0YlhCCpXxjPENsrk0OroTQqqFpoIupaLMYXbPiJx2JShHA9mT
3wka+rRSJ+cPTDzEH5U9us4J4IQu+qtlMO9khYCVHG6ZncEhNjYBOvAKfK0uO6r1/M4pHr+sPvJA
Oa1Y7DwlEZZ713UIjKP8Epti4b/O4LTmLEw18QpoQ+dzpXKhMPaMHF0UgfJKn2yUqd9DOih8XQou
Cw+RW5uiHjVE3SPtm7mi31NYiWGwuDi86QOpYjSy32fSF/6uVDIi+fr8Kr+3wfW6mCzuxlSXu13b
VRzvGg0467WhoVCSYuwbwhWGdYaFrIrBmuE/W9UumYZHcKwQOX7OXqpzY7aoZCmXB7nSkWtOErg+
BIN+7H/5fATz4uNykz4q9YCpp8qR67uEPTcjDCdCtDUPilCrwAaLdqP6p9iI+AfE6DmcgvT80W1a
nJPmyjj8LCVLyb7tf4cbOYeeLr++hNz13OQFO60QyexFwNLY48yjuL7s1E0j9o44rGzrR+00UPG8
97IwqdMLN3OTb5dp1OX3YgL8kqEfED9bmRt2hD8+g69bFNVzcl1cn9sg/WQrwchgdaoFepHsFolq
yDHtZVoOxarKtWk7OBo1M6qGjPqlhqu4z2QDAZfOR8irL/pqRG30+c3Ts9adbq/7g1Gw15zW6A3u
hUa2f6x9WClHu6eIrCos5HtkEYsC9rGBQxhagbimyTE165s6wejS2TeCjGeahstgR9iyrm5w/AGT
IJGSNJIDtq+d1mukofPGm45ZMJjAFloPF/EpdYGwkG/cjaQh+C2JSmWg3YHXE2OEsrwgjRheRGFA
LAFSJ1WwQ9zqx5X/sCvM3/WjCjzPWl4ftgvz0y77raB0JpjsJ2t66/JWNm7CZ/h0ODnME8v2yY4B
cXSzI111fI5pwE3BbqgqhgWauznWB0w3xAZAYP6g8emZF6HEPfWlZ8jwjpgXQn1GUMT4W9BTr16w
qMw9q//q206zP0fH9u9KNqofR8MQ88sIchM2isn/s9AI5A0wenga2JBkNBXFY5xGu8ZGWKX/2JKs
LbmgiepF3hJCnCap9pGqFoOBP7kOxQPQ69OxKbKQZH77hJBgWuioVfTYeys4sB0MvJJzVpZrx1kx
YXIaVgQENiDm5ufH1Hm8m358nPMxGSSWEW1Dp8BukcWWwCvwehsH5EqABZPyidnRKSq3QrSiJmyh
T8OL0knT4ZpsnAguAVinlr1hwHyYEzsyA368f00hlYDZ6xy2dlM5MuJFIJzCeSyDFveuFJo1UJIx
EK1OqH/fIpBJ1NGZDA58oyAroU1i7ZW9KLzO6BcLgp/mrOIZEw7p3L0Eq+ulz/dsAQLlWtbACZH2
J6o//HDyBRy8lAFKcz4xc5hxfLG/6GWEIOarRSWIM2LbhC/hw5gr2Pr6+2TeVcdGxQ2jLQ10A9hH
hunm9U2oC+rZXjHewld34LuW3X1SyJ6kpRT3VQBz9VDM44oXQV2HSUWYym0C3WM/qnzhVMfQ1nV5
5NMvHf/3otBznIw3B/wysj5ZMFqQPDk0d+esKs4449ryzG3nLk5nE8L7ftO/Q6sP1SwMH8jbnwyA
ggznUNqOH5vFj8hWrMjq8jtIl9vTcyH/o80hVzC0i1Ast0spOKgoMQNIufqHVfJABufV7ACWlnKi
7rEegzB9dpsus30XpcmJt8xfv+XHxsQjH/EZosI1zvHaLZ4ix7NC/ySfbiy6LIBvJMmYZxdJCMxB
ZHtYZJO133wwSEzD7G20sBTgnXDkmfoETiX8rsfL2LHeeZ0PTG4NET8hrE5cZxcwe8cI+rilxDo/
ovfhwTgpP5zXBB3AHeLNpVvIblkMM/5S1q8lX56rlvqWPh3+P+hVtweXioX9eylyCDUGRYfdJM1r
vRHTlD8K8AcymdksK5FupU3XqdOKqanIDn5XE+ga2quTPLyqXAAsFKQJOIORYMz9JNBvS7fEd9xt
l+NDX9fqvslKAAQMq1CGdaIO+doGQj96VeGqhtOAdBXCJBiGhoPl8k39wgHjY28sYVfFpdP0WzPG
Arzhvzm7UN6tL4DoVIM1iX1SCBuaqb9pccY3jZpVdwiLWBYSd+9ACFf2j5RjdnvNM/WN/ZVtMDTw
DCJe8WIAjcsB6CHKRtSkEYG78MWV3YOPDpl/AHSBZuYA6gIxDggJy3z1uD3A7fmCGxoLnXYDsxUP
7Yc2p1qKowY4SoI7xalRlbpTQFN03vvyJvssmTCvrba4twsPF+u5JqS8VR1fjW8VZXK/9YvV/LcJ
oBB0FYQ2zdIROHrIMCik/yLKJq0X55RAxSFQ2XBuxyvbStHQCR+krO6otLdUlgCwn+RSrqCaX0C2
cVXee3WSZYJnaQbbpjtO6q+uKgOADsXi0FWAr0ZjBBHhZi6zhN/aKsJLQjpthcgOQ7V7BQ3Ilfk6
3NCD70sm1tFWjMUgFTMWJ9uZoF8EQh74fraC5rt1q7eVRt1tbp2e1u/MDBN/xqFr39bbk05AgdDG
hoBRk/YzenGojEF8M/2btsC2URoplWPwU/FKhUdaruJudaTHwuKl2YPnV5wbp6Hl0yXjI2NTYOVu
yPdkZO6f9uxNF+LgsCtPY9sBYOQlcxkgliPrW3JWYQtgY1ZrvP+wP5yDhNVf3616JuNPuafmFj71
zoIFw5Dc2siubHMNComTCh5clAdQDmdIMkq83ivc1k32I+diRw4NmorP/dax0qIETIFwCyAXWmzD
+3QscxVybB/U1mIzD8RwNWIEco6kP/OjWPm3LfTsnR0r5Rqq1+9MJZ8TIGIGq522QQ+6nW69HhBn
JrQKGTjOAmdGM6hkBVrqZZFo1mfI5QpwasvjKisP6VOrqYVAa/rP9q1v17/91zc7gPWhkL+usCZf
iwbNbg591c8cFZDtb9bHjtWFeic7gCm1imRjYtqo9d9vl+aLzuqmf35Eh24vINe2aPgC/OAQnZ23
FhkqpWquOHC7JJVCzkoBBvUn1qmCHoECQ9DNyR3758cFkdWOUmP/iKggsEknNMnlksTZ7m34FoOP
4LWs3fxDJa5kGls14r+fRSj4+NHUHobDG/+upzAkrOG/g4UazQrkL9HKzxCTlhG710cH5JNowCpF
5vfNs0996sUZdukdgif+cjzeMVDW+1UZuAg15lkg6jYroC3b0fvkhfJ7GW2wvFOFNuv6IK0jX7Wt
bnShYluY+sp0844rMPUVdTBbCEy45ZvwgxHaDwg6ysivbaGuVh+KhG60RfBnl1j9YzELDdWgk5+G
zXbGRmnCh/4NDnMX/8wrDHCwKkGWXKXsK2/L9cvT8M2PGniw0l8E//HIYQEVBiXgN66na13bYrS9
QPGeUgX4IeVnezNiRP2xQaYsIvxftue4vjURTvrnif+EI3A3Zziffzmk92W/aB93+ltPVQLizLmW
dyqch2ly6hqeqQjVct4N0fRLjQKsmyVtZwUU3s0Q27vPDlpyzzzkBBxtzZ04i4CKsDNDnTHWfASe
aDh7HONna5s0PbXsFHI+yGVU863n+U8drLzrBn0dSpDurxH/VNPJiYsA8tmHJGI9sygtGdqU8Weh
2XscNZoi3OxYLhMX305RbPPzRLpATzWIrzH/kq9bM8rL5cOlg/AyV8AKfwdpMhJ7avzTl+IFAjbk
aJK8AftjFEjIzgqkJKFvW5IZvN91uRz1PNyu8l8NV633ck0pTlbX0FuJ1wys3m5Nkpe+4Md+CHqH
pjfDODeiJ3FzrLd7hNrgOG4YLyVbKFhL1YW2amOobf54ZOH/Y8KTM/rOKgnUwOW2c2eCq5+Y/PmC
/M26jY5YaS+tzn008cQLjMpe4GKiu0mlwRpQohWty4KjalxQw7fcKIiqNblSGuANK3kvUoaL5459
pcOD8f+bLt/DlcnmJV3YN88fgLo6O2mwY5UPlY2VnNd5nAkeFWIibFWjWXtg8Zn3yn7EIYrABrY1
K3bX2hn7sNGnryePQecr1ugAFepqndHbH7QMOB1G8C5AB9lC3RKYNf+AuvhMlIylAlPCwqG2RMYZ
4ROvd/3oDY0e3cTnk1yMZv8jbngJaXqsC1tsyplciMvdnXjxgZvGIL/cnxk9sPyka5PW00xpPm5P
eD8FXwVHEXxPvqIjVw9CO/Uk8tvLi9nHJkg90e402YG7Ckdwrl0gBzqIL4y2ZVMUuwuECH6zPm4D
NhgJPYVw+UQUQuEeF4Rmi32kXY53gZEc5PnMe8ycMZjQG7nCoClMReJoyUkUbSrP3iASfxskFuTQ
wJB8Ibk66nbSWpLmQczwZ5g01OjpSiiX1vrco7kkKQGjA8bpyYWEKrUy4F58MOA4K8/x0TPU1CQs
7jGmEkj+zLCA+nAj0wQjNHLnvvP1HTzNF1ZHmb0QUtOezltcgnLJ4eZG/LpmbLg2TTNHmaxUGqjm
0y4pmQETwdwEjGFJ1f56bN7MVbWoodB73h6pf5irZA4VSLVUQIwwFvZ9u/0vjhrNnvZPA2XcVpvY
3wxcXgzc428kHUKuxb1AYam6tCTxI4VHouPhIfk6OpBAnJN7ReNWpkLysyEJjWYKO6+Z0n3/8vzc
FHtcd+pA479XvXkbAW3vECqW3XLv9wwCh9/B78QczP0TN9AeHImWoRRoAwGGnh94KQ8uy/cnTOa+
RPGc+zinDTEn0mOq3U4MCITCjpwR/bD7j4N/47wfXYTIXAKY41bRot4TAwulSJnLRRD93sRNFzuN
uOeHSg17mjYjM3ISF7GQJZrcD9VUa7Bfks231HCS5wtIjP5gYuMglbHp8Y502fjnRN9/TukdJzUR
Rp7EoMvrKnZrJGOqtDJQRkg8Kshe/yjtYKJH43rK/kdwf2zW0O8iVlCyhTEOJRiIsIO10lxPBOW3
ZVdILAU2U3zf0FPE5ji4SYBlWMDUc1cWhiHCMEw4YLamvIn81F0u3No8C409r4J5aMrcUU2E4/pb
MwxexrYWozamGcX9+iU5GbFlItM67qzZUS8AOH093V8Ya4oKcWzEQ/ZuixLVUl5i/qoPQ6V2Oo10
rFasILIJgN5xuSU/whjV+K3EQtvGwockARA9y8jxmA7npUtEgTqXBI20plILPDJbbbVFvfeu6/Sr
FGxrENoq+FaxkSl45McAQr5uJ25GOJs3fEOnvuUuL3wAVWE5rZZ15noD2RsP+oUeuRltHOpM4Jec
2bvYR3Hie8iV9bakpZK0UX1wq7u58T3uUvXEyC7iIZDJF8N81HgkkxuzL+VfmMB7Gy5ThXrIfNY6
0IwWg4l29XsjV/hcze8Z9bkfV2x4oqzTHyoCzDDLhiXzPcSwqKM5Qwnjr3RK15PTTxz5vw00tpbe
96GPQTK99lqWENHWShRFkKLx+PdSPXh1yIzJxdEtJCf0LxXqAe3fyD9DySOXlvSi0Ggn0TtSh0Zd
pje1gL3B4aSom/l6NSahVx6W83cobSo6ZJV1fus33qrntVioOGt/rHEDWDJKJdCG8WPOXU069bqq
xXbHrnRdUUl8KemXWOrNXBDRLvUdkf3QH1Hi3K1PRYcIJNf+MaeinvgK6cnHwA7CpDWg7+RDpzaT
57MV2S4K9hqMmvWe/rn+rw058h5BD1KV6nsW6jfzgRWwFWg3zzHzb6w4n0C0EQUejInBLDppSXCt
+JD8KQ8QX3KV4hF9V4lxllcfE7pC+bxxUFGhjj1MSQdxx+ETgDSh1+Gec23GcvgX1Nx4m2VpJacV
lRWBEwYTn1QqmFkrM5lT4cmr3BHlWvzNgPdNVcFJYAntY/rBPhgLGjZqq8TNjCkfWGGsKXJYEwBq
Di1z8bm8hJgfxp38uzW3YamxmmgEBNMeA6RnOX0UvpTE6m3iPRVBhYuxx0KBVJEpiUAZpy8eSuEy
70Id/hhaSqFeOemG2Vd19lJS6b69xG4ZvQfXmEqISFoYMM740xsfFgah5jQk7+/VDsc5Iy0kzZvO
C/LcKP7sI+fcS9+aPWDGgpqbQdThM7Yz5rkQc6VYLTDfwW7LEiK3WC7w9hla/clTNZiyVzVuSWJI
EgeA65irQ1plgoB8hEkjZz9U47KWDcfHkpy6Pwxlmxvq9dsZxFL6cwuR6uUM+KB7LmGvZoStI3sv
BZ8JEKuG6JhVt1/Fl6zea+kxf2lUsq3rWImI4DrKha/SJz/3OGkJKtHc32rEPH7PrqwpqZieIxhd
Vm4IkSyeB3g0ahXCdzqh7xw3duQJoohUpwx0+NJbZuRSfzhWyBVVr6zk8X/1AvAMlcTQ/A53x6lv
LeePO0M2jNLIcMkKKbd0e0gujbGDDicnyX98GipIm4g+W3CPc1DzPtAeiZixBhN5IQwYkNefXwmN
+BLA9fdMESBDwen6e3EmzawPbB21J37UmscVvS6LS1fSHAu9cTRuxLh6BtR9K809765Ae4v/QmpN
nD4ENGtbTbX6q3VwRZv3xBZNSEEaLEQVPXfCihDmn801rxm3UlT7IDup9oSMiVkf2efgNQi9pFc/
JKERIZ6YmiLuDfoajn3nABu5bbXAqqj4b2Ffqn13d7zp+/rggPOBkoZ24/xNKAMBecvw5tLoc0+D
jeqcTU+QCmhVcwpy24F7RjHMILp6V70JIlcIOXgYqkH1Ou1BbGtCyDVvg+R6wkOH93mHO1x/5C9v
NR+deHw1FgKsGyZoWVSrcyWIQ6738+D8Yy6k/2YJaVcNBzo5emMJQgS437MXdV73/o6X5z5mS9kk
tvAqMFzb0z6v5gJEBcU5OQl+zP/O2WyJt1L4lNaJ9HOyVeg+D7YNSXsgq7UJ7HOHY0D0RUme//I7
BhFgdOY4koFFGrF66wgHpnxnn9BqlqmAQfMS+Q1Le5FovuBh3bY5YssV/Slci1rOQHcn5fDIYk8J
QNnAGvLyag0gZXuyLGRmZyFnBKQduN5tmpNu3QoCSDGwOc1XaB3IqyITqUh6BdFM3FT0IF7hIk+o
CvWFoTYl4bmcH4PN4bifXhyHmH/JsFYpbR/uPZhIgjJchuWvd1mj758Au3qD+YSu4085oxfQzXyC
9ioWe9g81782BkGy6ffG4mhSCsXms2nL8/1VmoT2j/ExzfK6nPoC8Sgmp+vtss/Snw0b0LNQ68Un
znAjpuPJ+V2YJr+TaLwxn8PiPAHVD+gHfsjY5/zzcH08EAe6VjH6lUMgLMq4Uv+IImbq0NwIbzvW
Ek8QCMqDykoZwmRp0OvVZazv1tFh+7qZDx68lfUZiP5X26dvG3oBa1h4BV15Iw45WJM0Mzd1qbKY
8jPgNL6gSl6pwB71UYQPK5Xu0A/jOcY+yRV1O+KCHJAQSUlLE17I8WrYYB4vvjcyLUlU98DyIthT
KNItZMravA7Iiw9LtNyBA/TbIviGLWtNb4vuttL5ISc39F2t5OfkLN4EjF+BwxJ474vMQcZJ1WuD
NNG8M6g8vv+P0NlB/qjTbx1h/+s7torEGBqbSJBgzmRid/ekKgoeDg0UUHEz7jldUKJLG5GPKQg9
scB4UEbYSRhgDsvnLjW//kCvO4sCBckwctK7Z7DGXdwT5Q4C/WpijittCCKrvDA7XCWsxDSjjSE0
+XtwMKub+ZBDvDofdKdzxNviDxO5NKWQxoAppJY+0H4ZJ9BGNGPf843jQyD4B3eB321FFaWcJ+ua
Izq2Q2liS1I4Ysf9np2Bjm3vRICGf0WCuN9YKU+nI/CBqWPb+orAeK8qZ8SnQ4jZmwsciQmRMH1+
bwtL44pqUGyJbFRjwIBxqwRV5E+aQs3hbq3yNO20WAULESOvoveL4kQX96zu6eIgLjQLvUR297sf
eE+7HPPbXvv1dY+0aFsivmtwDtiN9AH8lTozeURl0Qm5tsR+0AHaDe/BgRUVv+CoTmwRWZdPzeBd
Uq030JCXZvrs2io/xYn+wZlXoOIx6RmMAdKgln/F8+/LbL0dg2e6gK8U0CYySsrkdDUJD6GUMkAw
bXvR3FKB/JO4UCaT0CLTaQCotzCEUHWq2rEHGvRA8Ka+oB5kcqtBjrLekMXKkBk0+eUbyOwuu7ER
ZbL14/uSfKeqWlL5aM3ltQMXXIVAfKj6vRk4mkKA5rYf+gxFH83LYAQCmS0AJ1K6+g+HZgILnEO5
iJcSi4WV6k8rc9OokrgJaYqS2Tx57YX2LmClurtyi49AYfeh8Y4EU3qhc/Io3SVB1MPe38XOo7fW
pzmgJl/DfLVv9tZAFJy2KUfD6wLSKc+DVjxVEccMnnVP5/oNXZVGKe0zSc9QjsNgz1Cyv1qaKep/
GTr532+d3FEFG0HdKT2dS+SacJna4icfTSGsG4UNHwx/I8r3ee9OykMg4rexyW0iHJab/nEjXUwA
TBaVPsFv1c5Eddkj64992pdzi4KFUOkVYzy1gjw6KcAMC3mjaOhuzlBCAOEVBApCZ/0n0YOg71RR
bccMPAvWFHgQ9ZirRueTHiP6fp7gf11zh5bbzehnb86FOK6hfNevvVVrTsPf+WbHFORkDydI/P/4
NUgduaNW0gAL8/J0LfGPyGoJQXq4u0ax7luHjg70IXxJhWS41Vu9G7h4iMjt4A6D0jdotnBUJ2GQ
CQRtlato5FUGoY0zpeYPX0qR9YbllHqvPRXYhNZlT1az0Yad8Nb/si4CQnsEpL6JvBBgDeVt1PfO
bMNZHPY4cq7JPw62jGl28M9VoLQmVrnsLrr5zZOa6XgHcCOGRl1nhX5oobl5htOFSrH2XRQbD/ci
SNQsV6XHVGmRfLKCWYV3z8aobcfALT0w5G9U2AvpOFpyaKDTz0gy29qUkhBOQOGnqxHhRKZ7B7b+
GDqPCQqZb3IUlJFw1Q1tJzKP4hh2yGpfAwzAI9r9V/66R8VAAQoxELNa6dflILExyi0BNwknb7U9
YJbItwmVz/mmbykuqGBMdUUCex4I2gZVEM0F0jEoEjRMVZEnTwP3tE0LDQhgKO/62j9hnQj8lwCV
l+GWn1iqssgQfueLH9aoBvHYRcylBSPDq6bCb4jbDWZKaXeOqRgHNGogTPyhtHh4xRZGePYrop+l
myL3bABs2+w0MzK03I2OiXfO/CsYgbsHsQDfOlzJjOcN4iULha+g03mpdhA5qvP9BrVUsrQqKozN
nkkWOFBXHMAzK5AAl+HSEhftR8t07Y9gYJH9J0EgdTVM2BbTEvm8ua9Fi+OCMRxQkIlAJAAn8rsT
eQspcUsfoooPSZ7llVvb+byyz6d3SSjA0OX9eJIjracNB68GdA2bSwa763SjqN6PL4Rtv0ACSzF+
YJO82dIHOl7lHpcSQZ3svLc09eSdQNdxaqZdrpi0+XfitE6X4f/VJFdONdVBK23ezzmrMZoir7L9
SWQ4TPy9koPLrRA9DmiNqU6ARmpn5upLqEhbkJcrphvq5yBraoReQRFk6gOXTvGNTVvWBl0hLCAr
jLJVgB1WrrKdmSoqMPaICEmJyVW86KW9p9DGJxiavyg/YjECpTSjTw9YsMUhOvPANZZvqhxE9XYM
qYNw38fkchrMnj8VLUP+tzENB6CSb1AlUvqTV+BZ8mZK+M3Pv6x/TRzcPIuA7UIcDqPvwkwexvfn
TqSiV20Oeprcg8t39nm4oB9BvS7lE+5VOkbDlAq25k+Sa8hMAiK1ZKaxk0+BOEmdtBuJTXnZe2SF
ZOaOTHIsFDFGEpFEvUrcIOYapSOttc9sfpNbR3+JW+rGmYRd7Tl9LuzcUDmcWit9OpipDig0WX3U
uPGHPZv0HT+ih7eMu0hAz2f7o1a2RAoynavAjjaUnwZwEz8tTlYkMCRzH57wwVnQguFyamWWaJFL
oSCP4R7Vz/hMtu7hogwHrqxHpxA5c0sQOYeLW3gvwneKK5CDl7j+krSqYkpxOG9SznEcSjlV2d+r
XVp54PvbZC0d/TDknPZJpdbIHBBeaWRLci+0hR7p3LkGIEVKulmbYxQD9mTm7+w0IbEiswbmWP+5
CJf/SQSqMatCNHy1s7M0dGp9fs1OYIOwVtp23v33c6FRTF4r99uNeNz2vr1hkOzsVfas2SCvR+fq
qpZMDHYOdzk3uHHvS2AqacJ6jFdqnZcbc0oTWNUOtwOyg9CjUowhPWi3J3FVDcMw3tr66koQJopj
g4HGDeNMFiF9mvW4ca7Ad+3rS31AGCuE/l+DMkzQ9VV+u5LtZE/hZC9Arj8Fb4dmQKbnWsV3AWLu
OVgOlJTmfhutKyPJ+IEjjDkzp4QniJmQiM/a+0C2R5ppa3BFbIH4ddu+l/NasTp0PwjTNsNqEZ4c
cqtVWb5WQ6jYYF6fADKikEfSl5aGPIpA/wcYPbldGK4YaZaPYe1Y++e7hXgY4IHT57p/JF6I+rZE
I8sv1aLexIEKkQTa/ppJPCVss5bqKKwDtY0sjAUsIg6sQUxV4yE+5Auvl4BGV7u8is/RROIQ4obk
+V6Xk7i9iWqfjd+CNIDZkns3ZRPcl6EdRWG5Rp5ckmR9LoM7E1mBYZpyihsTmpR3RoEiKSri5hRe
DP/MKYiPAL4aUIOvjcT+xyxK7qsKpbquikZ/XZXL6bFoeJGerZqhYFVGS/yqXaSZKREkNbJCCofm
l2iYV2Fg8T3P0m+gDh44sQ7v69h2vhWvXKfYhBFJ03K9h5dWnHLou7876rjauIo3METjd3V+/1H6
OkOWHaea+FG7D9bU2ePdpZIxOnV54MNaBg7BwpZkrjBi9FoFIFt9VbbZkncd9H+C8jgoOSvfKZ7H
v6okDp6f5rkTNhWYBQldBLLQDQOkdxbBBZdQjAqtGkKPRhjHHHZUjBvtPq7GoqKEezmpuBOk8KvF
AAYbwnsqT4o3vtWGE03KoRzGE/UmzuQ7BHy8/KnctlZxxBNFQfhbulSyLa0ohAIfP21BvHwueGtm
NaHkFTtemYm8T3gNdlgW+sbkE2gRggZGVBF2iO330hnuNY3hrOvXhwsc7SzEazsbUA5q3vQrKPJN
zByBlT31CN5mUiTMEag9C4LmPPh8Vep7I+bc85v1rMhJFcRPODL0Zxe8Vt8zby6vCNf4fF0Gu8pP
gAn5zAzCTb0RW/mThHsrVZY72LOdiiMuS/P8fC7A+GoMDv7BePfJOUM2UZpUzUjVLxdzi8Uuda2B
OecipPAS3ZZr6iPWN3aOEuZbl20qXe5KojfxfPtvhGt9BxrMw3JzImmgogvROataADBoYBeWePR6
IEIQhuufEq+HR9bAWXJZiYa2lGO6dUJT7fjQYO1qTwtN/tYp1+RAkiC7/DU8owiJ038iNaj7X4lX
jbwxkgRGC+eAW1EyjvAYf6Edkob+et3ZPMeQvBcUGqwE9Su/QhdcI8gH5vUyg1C808eWOIEvEcqp
QiDCCLPgMZCSNKs06aDRBQo60K4s8ritjO8dg2oOulDg7ZX+rBYacSTjtT0U4TJaAkjAyUIaxeYo
tv80p7Miq+thqrRa4LhBGZz/ekVo2LYqpRU9fxZJEqnzMLnWVwt15nsQ8S8tzE2sz3Mn9flgpmV3
wRhWkfaBvwozelkidhN1VXXrCfuQxUw/Ygux4ktjt61fRwTVef3a9+MTMEw5SVx/Q3wgGRaGH8OA
vKpkM0gkOKiuQm64M5I8PHYxPjSDs9I+PLyRa+qQmC2QWkOfRflm+8F548G/qE0xJsTh9BYKb5cg
vwN+g57kc2HDNFQ2tNyPx7HmRe7i86VGn4r0iTGDOa536iOqKRlpciJ2p+4IXHqmAuuzwgSU6olY
zbmkzAtZUkMiQB3lZNMtUdiLFAfrbsrZ5sFYu1DIE5+3HdvGfpD6eqw+o0NCaPDZKLbU9bIwhMkn
XCLlyHaA82dB6ihHdgg7z+6jpcxDgNYCQu+3tV0NbkJJ5OnzwTJyVmAPzilhrwI9PAkMe9RfZlWU
n8+t6M4hx4cmDZGhp0LpdjhtyKLDL96q8SJqcq/NojDPM8xg8SeQ9h+vkjYWN7QaH5nvQLfEYdMC
3qdRnHYP07FZRr89p27Qv0Dy+8uGjNcmM57d+Pqk4SL28WNnEF60UpMRbO37tnUfou4YfLYHxz0E
tm38w9Bz8KuNM6RTYH/w9oZuM5er920fiW2tD8/C2BFYnnxvJOMYwrVzUpiBrgWRpTIpCO9eqGHS
5ZCfki/HzFBQSuiZtjHiLqPfWOtNdg0spwIh8/Unjdnf/0k/X/X+cgId/rKE3VngprFIPqVExzB/
YWCSn2M+AEx4A3FXXMeQdtXciTmaDDibj1qYdRYuosIIaBkt0KjpnsO6MD8trA5Po0cVaXlxnZEQ
Y9Ah5Z5tiERP1N0wLqcB3a8QS6nADoMmUnty8OwWtJZo6osbaDLWlRU6AAT0y0vDgpxf/ay77kSb
cJk8ux7okNYZegy9sJxhl44rUwS4OpDje212HnvWGi9O6Wx6172NgOPEVp6TVjHgLhqcha9Urx/P
ureKOUKE7yqSR2fSaFrXzEhCvEsHUqwmNfYX5kfQzXbnzfL4fW1R6+DMRJYvYhRIQXHM/0qTRyma
K08iK0GUoI2nt+mJI/zgVyuztY4i5Csgq6kPV4fw++DND5NPd3vTObaKeTAIdAn4Dxr5EyCBurCC
a8QBRQCusizt3vVJg7Znhr1oyUx3qfXZOzIHk4QkwfjkEiMEaXZvr2Y6PxrJMGiN5E/Il5EIEK3e
1N5L+NpMaR/80upOqF7mWPFTqfXpPWYQAJNjnoStV2rmND0Mxs+Q8zWbR0cDvDAjemJ1LINM4Wip
BLZaSpeZDjpLg6FHXpICdBkZR70U8SsTFEr9GY0GrT8ena3ttsW0wTWIIwUKqTExqOaKrD2jnQBZ
5Y9vXDh2YeiEFhHEW4nXpMzCnJLh+pTZa2ZpGWQZuhDDjT0TL9+INaSl3TdhSb0TbKJPZZ11wRCR
1S/j3VWaIxjRqDFVGr7b7pPa1UQh+X4fmea0S7YRxSEy0Ue8jrJWb8/o6A6cnZ3QpEJ2QbSKIgRh
T3h+Q/qWRLuY+gdq+X9y2NFr1kfF9/UNPfBfU33A4aQCZQbvd9Re83s+/CdZWY73W+FCgc05Jkil
fl2AeonoqWpbi+sn8jf5O9JKz6JtqnGSA9YLRNRunal2m6IB15bZPxja9aQ8DHOzWhmAO1wTidHE
YVlasyNyafBrqb0nnSk6j2KHN1xH7UFzg6mlujTNU696s5Ji5VKYYCL9yaG9NJo1yEMXFu4DFG3l
bOdckVvOeQ6FrUAESv/daDYoTrcI1eH08duPixf2V7Fhz7iwadCrhOY+eTUbr761AifHS4iT7OKr
GvurCSC3XVeOMcYVE8hhty79JZAC22Hhg52Atf/lOq7wV7xDwkaRzRJSDkDt4oHwCmE0W5QsoVuj
vRmd+ux27IHDxcuU6CovSK7bltW+ImY6NnJ+3P17vz+JxHkeHV6jZXjM7pmYfGAZV8JhLkqmyE4V
925012bYt60pPmWKdAs2CAjvGg1QdAV5gUfWPFFAmD766+HXa4iK4JaQ5lOnSWUzNIs0s4YxlP1g
0ziwP2lq3OqBS08yWa+jMJzKfsp7K8e9CZrCOetdpIDJUDI0Ga9+XU6NoJRYL2Xeo7Gl1iiwK5vj
0kbDfcsucmRH4VQh9tcKoKp+jknTJMHSaFoLgq1SxtvTsn6G63nm99aZZBOfDpZ5kTu4OBhhwW5L
yJ9J4BaGZDeKisdPw7p29C69DvN+nl1tHW0b1OdMTaGvEPhxuT4IxTtsQaQBtszmv1Np5HiEFy8j
JKK3tv/aR6nhJVydYy5Zr+ClgfwH47K72N5sgJk6X3aQSMmh2HjkTGtUsJ0unLrldxeKxmVom+jh
YLWKEYNNQhecKK969lQbB9qVLoRAcLN70Ufx5DAYvtuyJ5aFfnPRq08IYQyz5hYYQGwrDTl+6tvk
+CikwNARC7Zj86J0li6bb1VsIWckCuXR5k6GRlO0KbOZxpdQIJGACnToishA3q+lEL2Y+UmqErrC
wZjQ7d3b3WMR7Vdupy5h1QmgQrepQppnOaOH7JBzVZM+/mi9lA64kwYkQpY6b1SphDJWsjZ5frCn
ju52uTzHBVmS/LA/7nvvBsrIyncN7YJgZEehNXVbGQqqRW2VGL5ilX4+M0mEEd2Y3lk0zZ1rbLU1
M+ydVKq1o76nQghDHljSPWTvVXpkITRcowB+KICfxvEOqiCf0ZwQ7aAxzgGnv2NBqbmiio3/iH1a
7UuUvfljgCD4xxNoNC5kILP0WQdsnFFPhFlBibBX8+4TlvS7Ks9hCCc5cG1TODbrNhmazkKE0u3u
ZxKwpWwbX4y+/KCt7bQ4JBGHTvotVUtRgKWLwT8nYAtQoHRvIGpL8wRQ8j5+rfiMtT3ECMaO48Td
l5ciqY34lZmGJjCRvAZ0aw7UnafZOoZl2qDI7xFZ8GpWpCBYWYbsmnRH26TmR3yJgTJdWgJOh/4S
eQ1fNgs4Q+nG4uatYHrpO8cBzB03qL1+1oSdmHdpXmb+tqygWjrp63Z/smKAlPsyyVKQ49Kz0uHB
MH0rBHZX9wvKvrlH2i43TJ+VG18IyVR1XvhEcJqb0JNkodhFXZOFbjNHuiH8G2V8n0vGNYqBTmd2
K7uAcr1nFOq3KcLoqrg0qcu96mSYizHRN2mmS4xkEZO0LxN4Y0skcgeVHExVErZdB4p6Hu/NUijA
QdSYY/PUiC7cFw599u7Y81otMU/R36aMukc0qkmxTvcwQ2ul1i7d3xN5HpPM177P2jDkQEsz3AdY
lIEbEreYmXA4nXWF+fQnL0mbpCbPD8Md58/ckstR4EkOxlFKvfwKnkuA/veEWNvYsAN35oCmdbZy
JSE8FvFGnD1PykFxMYLhNOjBn3f42cWZT9Tb/C5O/bQxY97BPVKo1h88FFyIlrOPFj86bRiztAzj
aUgsocytMuQQnM0rfJ923I5Wz20SwEOlxlaZBB4dSy2hZURfvO67PH6qHJrI6K5aphWZd+KwJCu0
rqTWyi4cBpUd0eJKP4nOJuNUJu40poujYou8w8qITERJpreUd1dt3D3YnoZqkloXxFvwQZ+GFOV+
SkluX2nJn2qfkdaL9E9gYYreMs1ZoByB6+32MTOcgOt8eI3G8VLgoIYQ+hIRqDawTtIGUeZVm+L8
6cApV+6I7XHr/qJXwfQnvDq1oOXPMx5TYxC7M8tY3Pmmgl+ObknQttCCyJlyBqPumN4SBHDU+pHG
e7qyu+uyvIcQ1aqCvGDtVP02/ycpw1lgdhFKSlxwcm2c/4cAOwuZ7rAODR/Ut0xs6BEIKONn/yUv
ZzsiqV/2WY4O71Ap3F1nXjGSD8Vh+x55GD5PuaXOOloF0B/loT6RL2czWknsG1SABfa4B6ykhBej
6uxKk8H25RDQBJ4obP4TM36pGk+de4KYkQm5f/z3J0OMOyaBXzdnMhawk3fol5uPHu1ANdPsNCZR
sopdxK5XHc3kI2lwKyBCRRuW+hgB0+Ht9TCFVw+Kao9487Wt9SLcvHX3WJWgvwRX4c/JqCitPxG2
RCXmFDxbeMUXx97vVhcTumvaIVRMqRIpFIY5x7JeU+xD48ULyXWZIcp/BY+3FnCxjk7eOm5O0wQQ
yk3eClG5/Mh0MyMBPWNdAt329JVlVaZcdPV+rgKo9oDk83oLVmL5MjgHsAhMnc9Hg0vSEVnj6dGq
KL47perqBHnzKtl1tA6iF10sfklPnOlYytbKQggsJpBwVDLCKgDEEYYKKEENHvCim0aTDzusUSk1
wTuHzSJr8fB0tA8I4To6EAX1+h2MOgy39M2gDLIcG5D9G9wAkBcNa1jNYuzje7mqqYOq4d5pYvXu
tnfPL8aEnNZu9+GGFhujTRS17/RhwwEiMZxcylEWe6DsTBmXsD7G+sbSoQmWi1sflskG2oOZPq/u
rHSbyGBKSuIc52NTr57DIgKMzFyAThG2cWPWN9ODD/P0KuUd5BEv4J6ms++PuQjXLSVm6jxuIBWr
yBLp5JWSbwdoBiDn5nQXdNVlNcguD517wYP+rGhXl2viGjnY8YDSLmAMGU88i7GWRsI80hYs0tOm
E4Y/E4ObWVXJA6Qden2H0JW9awrkDv7SxBTomT/LOQrN9+vdNLxKQb3uE2u8Np1Xh7QRobqmyhJs
qd93eJhj1mnqIl9R2pAVW3U1WlJeJ6krMyEurcXI3JdvPPnvPNoqAulDorRvvbI0xVwmyYjscY15
zR0gP96Zeu1/laBp0mT3o6+lSz+eiKQ3/SoMbMEq8Ry3Lt4woMTAoGnOut3h6wP4GQz+GhLbshZi
UX7H1A/D1LKhCiR5rVS1UxvbB82DX9Hh7ZuIdZqDSN9QfCYs+aZBZINZpk6vOT4NkZ5gsVRDnxWZ
ji/Foo1SSly1BLGLXvLs7n+zstELaR7pINsoO6ALsyLx2NZ1aF69HU0YL2vV8/quTevQls5gRFuI
mXcVAMKNICEg0IdjPP+e87aXgukpYhZOnFOHGvp95kycIWVpBKjpPgCZzMlZdAOtD3tM8Ja2FdES
e2htvEOmeoPiMAo5etSWllOcGjoq5hnwMB/M/dxGFDYO+Rvf1U36HBVmDl3w/O6O71+S5gBmzY47
UkwJx7RZESPmLCB79n0E37qBvENbetbUToXdSLpwLHReQ5ZezmcK/TTjbstJhSf9ebCp8uapnGx7
IY9ckyuWHRbH9tCH0wG/6/Txjq2qWqOlyQ/xs1Aac3CLoRqCHGfepv31oLNcyg05tib/YQri34p3
Geyvl6oXLYud1Oa+RqHo4DBWvRItqVTT3HGEOMtfFk+p/CCk7nNqnv3GO0lWEMtLoC7QYZRp+Zpr
WTuX9OsUfcjtsKfYtuDfmOeOQQJrIypmnThfPr6bPyNgE8MFcLVrNRwZrmdfT5QjP+qEJ5jbUGfw
23e9Sd2u7izxjgBHGaDPJriEs07HeQ+K4YFi1z9vYC0uitoxauKCrtD/SLhVWMP5vwbS3Xy/bLDd
u7G04bOctpKFjBCFZCT892wDRc/NlGm4tSbCBRDZ6e7YomYNH0uxTNUX+OGfBmHlWkdYLU4Vvmk6
wcW3ntNXTtPp3HFWn9xewLtumvtFFo31tj9mNAZt2Qa1SEStlbwDXroKpuVrS4nA2UZwUdn4SMfr
UxSQZEJ5I+0SjEKsqEVG/uiJN4m5blx1FZ2eQsySjKVFANH0gOn+KhTYeFSZD3vDN8V9E152yJZB
8lcmGmkwtlQW5O/52yF+5X2h8xpU8/IXbkQHiLPl27YTZFpv+Qw4g93BHgV/NqOtXf6HkvYNygr5
sL8F8bT95GpXSI34bz2pw1+hf1TpNIkU7Lk0YLkBWHngnIGX9xiyOvl7Fp9QUPzyCmORPvdX3wtk
Wdyr0Lgu9bD77ZUZlL8fvFETK7Mr1cVZ0lBafagpreRb0S+4WUIxiz+OOUJ8kcYOKfLHjG/CG4L6
5H0SEmn7TlQMM6JirnCw5dRlGB2o2qYqkRwu4fvpRMS2mjnLswQ3CX+ZdxyinHHz2x0wS+gGST9v
5u4XWPJathczdxBK0L1bj3p5sjxofZJOBobt4qVpZVIOPsmwwEZ46Fr6Rd8gKrlVBgSDjGjsqiEK
/d4lKBZ3IGVcZSqZQHM5DL7YpkSjwhVoiGmuw7/1aZFZv/bHMNpwIWAr9zYi5JhMPOuqIdh70Ml2
gZBnWUv2jlsrisIM8Giu98y3fKbMo+dFZPPGX6v1makpWSRdmAkwHXBxbCpAD6fNr/s7XRUQaqUr
rDGmkTVdv4T/wEHF/gmOb79Up5shdCEvMb2TMWNp0bX3EPnP8IFiYLi2cIV9F8bbKF6/k4zPQytD
U7TgR9+mfy5+Q9NxuUZVMOfcA0RiPUODx1ovHA/+/hcg2UG9C+0yYe7MDpW482sMiWp9K9hQw5VI
D1RIM/Vyw9hYtPx8/MTreG5B+Es/meof/yebRaSQqn1s8Zsud4DiNV/ae+ke5IBOb1Gf8DcEXco4
4KLr6LeMD28c0W/Rg4VYl/YliLoNawzfUSA8uwU9Us4XMdyOMOR21ga4eb88Kil3LhjkNJ5ReO31
04PuxqpLNoXFhr+QZsgMpR+LO6SpCD3G8U3qfm0j7CtT5KVkM1dC+BJxeSOlo/IdPwFPS55rrl9N
etS1wA6CQJlHqUVkGntKI7Yc5UJrkkdeivZMWveWQah8ugYSok8Gv6hfZvhPedV+ScHlz451tI23
guSCUIcJH7wHAqCq9PKwwaw2vZw0EbErbrQsRzOSBJNDf9+VutATMVcrbnkE+r8TPNgZ5iD+Nl1U
GzMOrTh0BDgTp2nC/Hmb2W43uL5HEl1phpfsPnAacNIv4YXSs4ZtsCUCIXfO0AQP7I4dZZSyne8r
GLBWRiNz35SqtsohX2C0aJ7LkiqyViUcBev21vajmC1F9U2+tgQ7UbW19Se7k5AotpJTbAAx1CaQ
2ANGGfOYSVkRghbnvJzoyaRROzjHIxHvYY7lJr0ureDqw2NaGWEB7v3lQYUAwJwdhj/mhOIKHruH
mooWQJBO5eDezdfeLqsJ0aQyXfgNli6LVAGgSqk52JKT9EmYdU0A+9GyyS4C2yIluE9dO42hDK+V
4pSHL4syDoBhKftepxud05v5wfTqb2rxXwm7Gb8xp+zqPFdbFwLHEykIylwAYwaaps2yPjlqK9Es
bGEw+WABiTYhBuTNEtzWyYJYSTPZr9TLchsTaOhlznwGcUupsIn41RLe1JPUPRDqXEZCZUkSxp2y
JXIfx3eImtq/nHbsO1BAhYXW67d1+RBhuRiw/MBMl8sPHj08BIUSbYrl50NzkGL5xsNWAi+L8h/5
y6mTNq4G4qDX8mePlCzFluRfbjTLeqC1q5VadG9390Fs/Y/YCC0N1cH1tydN5/ehsJtqY1QRVfwo
D4HPNIJIjHonKCGA9ATXi/xwusni0rX5CIrY+iutmRKIn2aF+6X6HWZdCfR9W9HY7KkVG3ljBklL
ZM4ZyhsDo3ZO/nbWW1dfUSSvJPgnJI26Gaz+NlD4AaCIMMLmSJWAEWgdvjUgrEAIWNh4y8Q9NTbv
CjDngNxzAh3pJAnCYzSDkznb1GY1Q+0x0yktWyXgNIKy9L62ZJbfQ0CLu5beaPGm3u9oDXM9Cg31
sp0I0te7yfodIVj/EtuTI9n6i/E1Apu77zhHPfRT5bk5St1AzbUYx97vEasOgpRl1U+ODPo5ZMPS
p/Sr7IwjMGMQUPxOsdgYK7xoSpoZRdO+DIkVR+YdU7k15Spwognz9rfx5IVvYgWKngAKNb8rPBza
UCQYMoEWdYGsNGh9eWOTrfazWRuLMnw1o1fEz6zQspo6bdNAc1TElYnZT6lldqy4UnDyr1Y557Mf
pw3Cax/y4SrHk6NfvDsVIUYmG7v67yqWMmiogFcDUACvlsL6CwshiapXZukx9kKBNx1GJ1l/esGg
JPreQM5TqsP56tgOrlJuyjjd+SMtUgfGlwYfpeuhye33e0OxM8YE+OfhGn4wEJiWc/49Ayp2CyvZ
YP4gdKW1CbFHvL5Ljrg4PUYQ3/VA2JKkSobLJCMvJlNNsbWO8BYVd3jNh9XR1JSVQTOu/2RlQ970
1+FXT/3QAgAFbrP9seEPjKJf1cyt6xYFWzfdfHCobyTGh+1OnMwG4P+c3jjljIhZ/SbE/yZVzg7s
M7Qcxg8EBsOvaqbYJl/WJH636rfaO2yBiqug/6P7JYmD/6XRH1rdtn3+vfNnG8cl9ze++3YtGzLe
euIuFhdsZYn7+x5J5UrXGK/X9xo7rQGEg9vHmykX71L/nnv1bzsuEuufa39hW5STkX8GYSvcFYid
i0eA0LZ0zoTgDNOky+gD/EP33tYqc1D4J0CUvbIpQDlVDc57FvkM7qpKu8uPA7uMaciazjIIFbj1
njljpJXWaP2eWN9+OOaJz9dsCKe3HNnNxzZvqKr/RaRlF7/inL+VrZbEo+hfNG9KA0+J5qlLLK8e
AJ0P55Q32HlyAVk47f3YutZhxRvu5IuQVfszzWUVFPiY6l96MJjZLeNeukZhaQYq3Lqx6Yti+ib3
GPK5PIae/5tD34VtRVWI2fyqI+5duCEF0W3Mhr6uy/zlUmIca5im4hlpu4ojrj1dBJTpvNr+5jYW
9o0AYzIzrI9F1liZ9nKIXKFV+9qxUGDU9MdLDgOWXd7LgGiJQmkW3cbR9Ypwaoxl/3uHKIMmgxkm
FAeVpXxzx4YcdqSxtONlKLP5rfvztle2kDfH8W1Cqw4s+9J/Ssfdh1DjL9dKsB/McZYZA12X0JxT
gmlX3r3FxyBgH+gvGDL9GEYD/qMxoE1Nd9wnV+SpMqOaV8dsE5QES9UWwHyJ6efP3UC+0gr7jl+N
PbAe477rdW6Y2fxKM/c7U8QOY5FZMFY1nKXIfTFXkO/qjReYnFf6p3ZQ2bgMnx6eQ01QRUeQxT3R
AmsuERwcK2ydWOQHFEFGwaEazj4Qz6q7NSejlSQH1XFsF3mn04GZHpa2GwvLe1QSA8iDORFQS07B
coe++7icG6Y9TxonVLWa6BI/R2a14vo9fZG9NeylwCEtcwk8tWx0Ew/FWxFlpSxVWHT0eDkimx2N
Zt86kwQwawXEsr8U75zTIckuh9iJ16P7Fs4It7Tq3z3A7YE3mOucvxoQdEZXISBfeEefCQjkszQw
/7EtU2KXMIFiEwvbrepWRNFFSRBvbqq6PrheTjqzg6P0TPbGJjNwFlAswsDsOUwKP9Gk3GwruX8E
1puAPImeqFK9DAdLhWCO5BVVth4bxFCXTxB2isdg4XgAzUWteaQxEUwzf4qLrrv/fekulwj1f6TO
EFP5kxJmAKVU+1zfZ/Q7Y+w5zVYY2mY6ox68dzHCj07XNx0bfU2AgTY/oBop57XC51qhFPC/xQTj
wzwRbyGE4iaEcPuswABv+bZie161Oq0th22du2Hf//Bphj8tIxGNY6mMgk5Q0g4zeiRI4DKZ71e0
5g827XFfjMkWT0UDLtq5yCNOSR2KFWkdYAKbU4q3lMyrL78n7MoUF4rT/PSd7InzihK607L44Y2/
JWghfx9J5tSfT1aTCGdEiY/Hg5wRhbMymgTHLgyhC3Zj93cEZ6OzjG5q4TaK5cJOJrJNIWe/zA5/
W8MaX+uK9yE3QWwrs2p/Z3h0dF9+Q/XCDjppbxq7SguVsvGd2empdvBTQHJKmf32ZZoFk9825ceG
XSUJnmcttRqqsbOse6lJ4QTpptY+YoIxiPxhnm7lugW9BhhjQlzHlUxCt7zVvtS/hkqfpO3Snun5
FZM2osS6e/O5S8tg7QevnaYz0K+u5Lkl3o3oahamId9Ms2jwIh15t7mFAGajS65PSK7af//TJWim
lBIMAuMkAg2sKVH0Xq0evxcA6HaK1MOJiTKQrnFIu45OYXJPSnHg7BWxa4CcvK57S38PGttTcDlQ
UrqYC4BA+waZDlCZmWIJT2bhFE/TBxOXHFqEbkK2aOVIvXfUYxzA0h3HbUIBigJ1w+YNaEGGNeXn
9qLmofvu5oXCEZ67U+cedqxdLfbUzPjb0KsOr2ts0ROCqLMFWmAOsvbId8YRENbNN7TBRQu0TnxX
0T097JV/dwfZ38ROQIHkaLGXYGK2reQFmcUMA4G/bDM4Rf5+zBv5/bw3YQ7vAjgP7ODv3Ch76uyH
XSb15b3Siwi45pTLpBFELVYgUKUMc/8ujpjW1dBv1a7wqEGqkJ4gukp2aV+lWiPtCuvrWPX/uYWc
0SAdnuKSOIAQJYy58iHBRzVJQP4YLDX6wO9wgxwzYhCG6IoTCEywZKoCJAwGJ398zn+v7vs8MwHa
0WO8HCYdQfCVPudgutm0kowvYMfHPkUBquBUevEo8XQaO/OlOAHQND55v5fUwovFbVJ5lFeSJkFg
xTAGhpeMybnoyiQTSL2e/dmU4Pi4vAG+Ghe7GkxmyPUxwhnd8PCi7/CIGiWROVudV8E1ggkaUpwW
1WsFlSR+bEkeR4cppqaqkhG46KUVhjYYXFVk3num9rkdLcQSiqWmKWELLfuU6ehX5mPOrGJgd5dT
D3inzpBy8a6ylvlWADMRpf8+a5YsmJvOLHcqG2pQl7DvPiF+SMaOcPdh+VNgmXugbycm0J14ZDp/
XBZ1Qprd6IfNC92QLUhzwENnfDd3HJkB5nFlOi6lQCS3HhvAe5KtMqdFzJhmoOMPg86ucSJ7q5YV
1yPvld2hajTpEaQdhUXCdOTpI1NaC/BALGj0IzmIwsBC+smm0QPy1CCtV/FKV68M/oW2sBlwhrPs
3qs51mqrRPgZ7Y2oC2b4WRFcFKWoRbPonknvoLQeGwywOUYAP7OzoKxHUZIqNt4NESMV8QhdPPCX
ZaHK4pBrF6SmQmq6UsNmQ0vZOmtjO04lBFAZaAwZw/EQF1AKcZcMzKI0x0hP9enC/+Mcnr7b3GqS
xDgEomuhAuRf7EQFukdRn3uWVHdiQcOTPq9Ndtj4hutzexJ/zKr09qj6XfQMBnCbx/1xX1lvVHHH
SraYkpxVMnuODnck4wGntyziIFrNKILjQkJ3ZkxuHxjGgcrydzZq/Eq7yUTOAYU6XZfXzXKBg0Ae
fv+Mca6oqrH+kzNBNdzOPd9lhQuoYftm0oaQfUQZNQdzTcsYkb20WUunhKrcvR24VXaUirSHnqes
TlOMQsRomtwplWAx+SlXmWZBeZLJwVTDaQhnubLm9aarG4PzM1uXtBvWlhhr1TwgBXjfDuNSa0lp
WQ9doX/J6v/EzR1Ohb3Tbkk/APdXpCbUplMUObj65ekx2SZSoO8/wig+BodtxFl/f2MC0jWyrwZ+
UT3gPg1xHc/LUGrgewnBw2kUhEMpHywg8/rugEN3XPjOXGUJ/SR/iqCDdjl4lwu6+Y8rWWGB21ZW
V1bKMH3Ugf2IZ8W45W6Nq7r0Lm+bzEmM3Q5dgjzklPcl9g+dUIcMezOCvvWBzMvRqzjCHgVXCoVo
yZn6IMg/qV1NTNEA499NbYqIhORaqIhNQ6fqnnPgHgDyQCw/QGHKLtMwcUSIn8J1HZ+Nre7us2kN
0mIKUSneNaPOEPciLG+b7l22MbdYLH9zPkvcGpZZwfxKfchNJ2UYL5zCi+nYK+eGxcDeguxruDkL
tBqr7P00ierLUfmK62Bnx/LUzkkvwPzZQPkz6uJEf9hY5InvHBQAuTqergmW11vVQZQlFF22Ez1b
XE8tH8I7DFUK50wAJWCRGrU3n83Ip4GwdAoK7OibkaZwiflORvtCvKPHp6vrcituiHIptZTvFwsP
CKjC7eVyttVsnodYyU8odoW1Ey3ltI5dU+ar/bAcpmcKCWb4au4xw+ZKJTlGLaz94JmU3zvDtDlh
+UnWp4qV+V0OuMErOaQNE2tqaK0BYi9IiV11LeL5k0G+mnNHrJcZ7a9eB3Jwz+QuY1QKo0JjtUvW
dZ0aKP/t6y4spfgDhNMgfW3YCl2OgRg1CT8JuKUVSniaOjw0D1HBscjV2KaN5QzuyJz2/foPQ5bR
XDKgrFz7v8Vl1fAFdbCYddSMBXdKooqmrzmwv3sf4zzQOOGg2PiaYY4IiMNo6ZEEYQv1r87RdlTp
wsrC0wjm8UTA2SYjjBk+5iM9L8+HuIHK4xEMdOkCukm71Zj6HcqweHlO+ycIHAXqbSOL9Uggln13
SwMQJDRcpM47e0bwByrvBZI4avScRutsgwAiWhA76HrRATLp+mi9yD+AK9A3xWn1Vq7j5Lnj75i5
uEw5iShGJcYePyUEZo9FyTMi/qsQLk46LPCrshI8k1VrBgSo649A9lphj1bEGnlbVjq0SmXhgvQB
VQbUuIDIuZ0pOY7mq8c2xx/XDeE/6gPSVpyAdi8op5eLfmosgjvT63OJ6E1yxvz/AtJwAG7akxNA
FgfbysAmIiZH8GKvVDpPzsZwmJspBuV5Puf4tvZa+U2QDOlD883kioNhhEvJnPaKbHksothPtnsY
PAkrzxII5vuiEtKqUO0yIjKughIwaXc2MOjbfagouL+wUH5OgLP8VDfC7zVc0HYi2UiEmADQUUMx
GlDRB6/ZXgnMWP2Nt/8LfXPW070OWM3s3PQE77fN3D4S7vJ7poS0bZPYT/okyz2JyL7RdioE1CFC
4INY5z2X9y73codlEhVWZpTL0TUBQNbmUJuG6vZnIPmpcunPFNi9VjWIaZZWsNbV9QZoH/jfjms2
y35QO2lkJ1w7qFJdoCp8bcqX+sH6CAMWUTvpTuUrseb/u0qBTYpvfFw6NaFn4LObJb7tMny2foCD
Fae+ecoLIBK1qZn96rDtYiyAUzEy5YJqxwGDO4JH4Pyf6xOPrEekih17eIGVx2M6CubcueHS8lyx
uiiZ4T026H+UXaAk+RqxR5ZhVFJSte7wiCitsnWU1CWkQtfrmr47OE4vkpVQNU/qG+yrOjXhs+j2
g3wrTlyr5H2bsnw7uWWPhL+wC6kfBsPUDANqscsPb3amk8ex/5tptF8kQZPvALhWX4TmBG1EyXD8
j8r6ty3n29tbd/5kn2tLMVpXk1uym4XkJ/gpVnLa5kMbTCSpWUEUWBH+ZhxRpgw/Tsggwk/Bt9qO
ZRagdizMLTzYGUedMvdeLI7KaeY9U1E5o8cvSLBIHbJLRQGa3KAZJ/h3rmy4lUDCcnqBvwAkRbT0
8MtLVV7HUuvzp8XY8Fv1sVHVHXo1YDzpd7sdqRSNk5N3YNanzdB5R8wNq6CSE/hjl9f3hfzzsTfu
8P0oS7au4YJvUE0XAzeKltUorEVs4wDrruLWnKnga6ZRSQeUdMIRWF98FY/bAw7II7CPAJlDWgUd
undrqxQ6L27MgkNPwHMF/WsgSwELdlH1cohxFTG7e8d4Mxh+UUnEJsjxj7aoYYnxjDF2DXCZDiPy
IqLBNSzrU/+AyNdxFemc7rdx8wFQnWfAzvRrYappAINO1pty11txME1FxbwDieb5PbU1zwIr5Ipz
MqZG76yZFGauivkmVvjJY0tUYYeZG5r1SdvPVsmoMnXCDwMCtzS1spsiLDEjcMNhGqbo9hFzeUVt
ZHCdh4k+fh1pn9sEFhfk8SuEb3NfGnDZvjfbWefDWvbVyupS05p4ecpC7eGwvVa7mbQhaMV6+w6X
55LvJN5YeW7XB7L/QehpG6jO1bJZ5q/LJkO/jwkv3J1qFNzulX83H2Ak/s8pYNCh1NFplXyIIoiF
wlq7KdIUbG3nzyzlapFbecZAfUfesF67tZVowKZlI2kNcCDrSi+7arTlU5rJ+guEv1aIxpsIYiKM
8BB7i2mQzXnIxQcfe4wWkJjLgE5c3RzzgFMQaOD2tasS9pmsq0HwahIA8DIz7YwLrc/d5nOLeuXO
ZONwAydGYaoeRJVUwFxDBrlHTEuclX+HB+mkU6JIhiJbhbvlDjTzkFOrUD9rGJTefKCYPguXjedf
ffHaUPn9q76wINdHZblBHX2RZbf7kNu6azyI0NHqcJ9BtyHpcMTn4rjCUD+t2EZ0SeTcAgZ1fwKq
82w0lR8O0AcXwA5PcS+OjAbPb18TkJo6ZGb7zy19cOLT+iSIzULkI9rhx1tkyVmMEpIXnA93/z4d
BfCTLZdTaEDwkR5tGNab2I1xbwjvpKuQoz1usdOO9+f9KOQWtPxVHb0Yqk/COpOe/Zdn2nbYFKt2
0HvmizpP1QNHDOvd3O1KpMI1RaiTPGsQaLsLB4ay02wqaB8sWtGTHU+mdDV6anTqcyaL0I41TRn4
5pxEX/zszUapBaG1Sb7zLli8b7NSV0mjcJSkY1719U50i9g70xTGz150fr+JPl+lQMTvYbA3UfXJ
+ak7MXIusvVgDQjvsxJ62X3gZI441sByFR4C4j69CLEFBP9wM3v53Gs/VZwV0qxorb84dZ797W5U
X/rBTvEdAFRpEsN1z8x1os9onEO4djcBrCeYBUbkFeqj+caEqXat0Tq/2RJ87SfKhuEFNGmOOw8E
fVXVQXFK1bEu6ibTdRCpRxDeHR3bktJP8C7tdHLlACw2VJxQHGtLqzhbPjFb9+5JRMJD+ubuiMpg
kPSNT5Njw9Ex+FUwB4ogL83z6iBiGvOw1nzPCNiFn05mLV63qBayD8S/4Omk9nl6G7z8dXi6AoJ8
/nIV58/voMyWtv0i7a6hcAczz2ghT0iUIBM8oiuLUaVOp0ZWkiqwSEpPSy+BJz4PKgjN8gO1bIW5
kvqVJkevSnFWb9BoRRTdPahmw6I3tiPxA8f/loo0auZn9WOXVzsVsr8/seiDJh8pV1xPczuieUzh
FIDBooAf8y9QZ2cGji4+Nib2GYSxcP9MQMTYSStNQpl7blXt6PBI3GjHbtp/X2hdGS2ayFugQgk2
nz9fWHYAdmbPOVFnmz3R14gO97Uq9i9KxiAZOxNhRS355caOMvcAff+KkWvMS5j4HsHBN7SvKK6f
om9yxUVnhsZ1+x5A6hqeFTOEfru87i7fee+KWpdmus6T+begEaLsgMDo9ZwVVURKhw0Hxuu4XIFP
E+1vThMRdGrrx1louQnr7krLf8NSesGmx1q9z0DvRZzkXtXqKgULWq2ifcRT7Al7bXXptjpoUKsP
aL5XyI1xxA3a9tH2gBLXHfJ42p1rY/0Foen7wR5EqisAwF3AkRuEKZd3CWB9CgNNvrZG/i9glJDq
UkDHxR8YAHv1nM0L53OnKLK+vFCEzgaKO0rTd7kOoeszHS4FaT+POWd6btCC3/lOXT08caiy52+C
g2PMn0MzzO841C4cJQ1R4PQnrhmOwtW1qRpI2yvNcM7PbjdNNX3Tb8YPiwpAYrTfG+eYxti6QsXo
ev0cj0kxLerzhx6Nw/7+spXiRawSv3dKOBIsysZqbD8g6Y0baSMrGLA/T8qHAkibRfpWyOzSckiB
YrZbfrBKs06katAXxOjGaLETYR/CjQ3xZcHZYu3z8dpM2TI5v2/Jo61f4Ofb5/qg5U7jgJe3JXf8
oXDm5zA9DuxwVgFOT1dIrV9TX7jp1QiNGYknHJ4nsaBnBE/dqAEzLiqEnb6dDC/nYbinh5pTUd1U
U4cFOkwrdFGJksCSMcLArrEdNhMQBlYOy6hiNJ/M+Wu6PA/FQ4BdLTf9zI2bi9CNtPdyifziRV/n
+RUt9zzvi5tNPpUAZAqu557/r7rZVSdLHC78JIImo4OFjzwhmekJtJql/L9SEuwEDcCzaDSFsMzR
1ELSvA76qDoi532spBmiIvr7Y4UJ3va6WBILMvLMxvzj6f8aw1XoKGW5g+swcKuliWyXt6qfO2Q5
EibNCX1VUfMSQj/zE2ATvRYrhQQkyseeyMwwbxP02nWMvPCkQbICf0zARRgSl5TwxRfSilWa54zo
sG45zaIXUnfBVmKBwD5UvEMwp6GJ9xyhKAHPdU/wBYK21syH5VtCJgxozFTn9I3piLwOR8ol5MEy
WfPKhnzUJfuZj/wJlDrePRmSr5HR/SuCno+fKeiNydlWmyZbduN5aGEOrl9T1WaJi40kNMVi+C7q
+RV4LOfsNdalX3qGcewo+fFzf1/apaPdAcwS/OqKA30aNlCJWhW1BB8z0OXfsIy1bSPaU1M4tqsr
i3tI77kdIFQHNTZY+vByX69gx6zFRzhtgK9KSk6x1HAr1RGrsMrZecsFBP176J3uThM0e13+EiYV
ir6TZmiTMWFJW/66EYw7YAWLAJeVkfflBqHvcExH487sdKEz93MNbUkvkFYePd8ZfM2oMr7pVJNi
4J4uWVUnwhOoB4nBCfUjmrHS5bUcdSM55vGb/CpxpFwt86aDfUwegg78r3NqHj6TNieqLGTiZ0sJ
Q20zWLjvIDwMdZ+cxtEC8yJZG126n85AEEHB+8n1qu6DQwmOTwFUnC5KvkRFiXA/3x4hKy2v81tc
ff0w/5KQLy2jclcfH0WH/kI1FPpgfZREQcZWOLF0B5V23Uj/rMD7KdeATB92ZqxV3mzyCic/kwLg
uBrY7zHKN/FxKI7oS9WOlelvlp3iBV9jB2r44fXye8qQIyvOPQgNd1EpwunquHVlCnjS4ClYeCid
uNj8/Juc/ki8iuJiAh5+NnZtRKFom0GOy3+Ai+SccjKqxuynqWNIVMGzP+kq0NXE/0bViMNSZyWy
etrqIwLFGnmkaBcv+YRM54icoZeeFiZrCpxRGTQOFzTcnysbrhpYlFlI3/u2PVVj+KTaUYXUh9da
wBKZJbwWICwoa3th4+sIZnoLflwWpQhca/ZPin9ja14yvQT9Dssn+Rh8GOa6cdRm7qOAHi1KvOMi
Avm79GqAg2reTir6kC5a9VNlPRgyJ7wOW5qewLbzTkCwjuKlJSdrlT4l/pUBhAFdcnHhwAdZxzNT
6bhVIOSz2Ch3mLkUnjlIvEwQSPwhT6oNes8gErMPpq36Zadbcn9I48vz6sywbhaSANyfhnNCq+le
F5FLCH8s0LkeVKDM/Newe13Jk5xAzej/rhK2imzZndr6ttSzzSgzp9Aqu8FCiAbbhfzxqN+T3YAU
MQHRILPemW3Q6uNSGFN6SyOK2RrlaZLlmVdllySjkP0p2yjXwpcggv43hkPPfJ62xy4Rsd4YqLKo
eKvHIsbDYNngf9sOzx8ETYNmxqI+ZdevLhnv6JhWZeIGZuqxFONMoZSdwFOnue1GNBybIyo7NfuT
113P2ktJoELtcprLnjuuAt9zhHrsB9BWNYlFX1/yY2RY7m/8QDaIpWwHXtM3D0Ir1DcmpN771zB7
Fhk8qjGuM8lO0AbmXHirRnOHCNhRfC6Zs5Xri2qgQMtvS07jl7slYFWzNOirhRTytYnk6vtoL1MN
83xK3rSkGoYLQOK31z38vjNky2rYkge3bYLAL/YQTg9Svuvj8fUO+yGzMPq+WQAHedcjcn+b4t/o
fyOby7uQ6p8VCwnh5FUB10HFBRID3uJuXog6bwoQh+otGWn1BKeJSJENP+6pac/S0Hi2V4vLzYir
bCYqy2TLWEKx6ho5qgmaBdQukK+DLX58IAigQkqJyTdrEH9EO+e1CjWEekkdZhBYXEsHSwYSuB1o
uL4LB17RXSYYwRxJnWFJTvD6zqXRYP32GsTxcFCewFBVk/02dn2UOkQvZHDfgjF0Ff8QszN9kyv8
+m3SEC2YF7+07bUTkJVKdDvSgAXdamayV+cIguc+zepiC16G4PsDgrip8PDA/E7K+1nytzo2UKUl
K+Nu1EjGm+UWOEg4ZtlTGkfdvEJ4nXIOw3fmPWqY9b5b9qCerRhSQMYy/PZ7IWm87sw8m7g/ituE
y3oeH2wYwtTdLAnBjbvYI9ODWcRHoZQKnnutqrI2GbrNL1wLVihdT9Xeh4NGwd8FKRNeUAjj3fEx
4ybGXDP2jHP9jQhZq4wXuqCbbaMlKt22dmKW+OOOjOsTsWvwHCUU5d3Nm5yk8HKMBGV5rR2vP9CG
fxy/PIU6mP9+VsdssyFzP8xBluQVqMwuK1+MT7VDjmVwMcXpiR6iQFMCYLUaBh7w9uVPCXTMKnqS
L/gWYF5lhuWVZUr+BmwIW69VGVqkA5dlCWBL7irj0GfzjVH5gTuSi/r7bPqJpp2NTTa9IjppoMKU
d1FPrqFd4GbcqeDjq5TcyjrlgXHSA99MyfD+yKkZ/AMHDnicYLxJ9bGyS9E/B8MRViMNt7mzKuLQ
RFUqvXeoonzBp0BwR4HpQcpAMy/KBoSZi+ZziR/DkXapmZfIyTnBwIuSPfPL1ICR7lC3dqzFm5p1
/PW6LD746LFM2ZLUq6raDl3D+hwIR6ZoqO3Q6yQn3Fh41xDkg5gqgA6TzYKh4D+FGf9kE8BfWMTj
Ion/4nXeDCTiULxexCQmLCVQWdCy7p277bRmBKXki9oiUrBrWQ7bvmvl4qMpzMxPQhEuhmhsgtiW
OF+CIk9NDnNEGbAv8xqT0m5A+J+F1aWL3bPpdr0hFa7wbdOgytjOL7wuEwH/JOGmtzczC7QILXGT
cIAfqKVk1fWdhfid0yOS24uupyUw2vduaZT1lK5pDzyB5q+Q1Wan/KkbjJSZkdB/yrVOD1rZrRgx
fRT5VXXXFfrjwJCiRJp7TRKHzUR7+hajcCwxdzSaMwuV3Gc5zf7NqJy+d1Se4wibQux+zR7zjziC
AAh/QvBoM+l223HuoACDpV7iws3XH0/PoNGtg6TBgeGcbID0FPTYL+HWC1kyfHWUXXWLAdnIRSxd
imAJila5PpPK3nTI+WBPV8hz1vFwejQr7PpxS9eR91zjClUe0xHFa3FPUqBFIdLZOq6EKnukcjI4
9jquOiW+KVUdNWEqYVln4O6M+Z23rMHgqlP3OhPHnsYQm+mf2pGxLXaz0McpZLXnkxEMsVvl9l/I
VvI+5rmlbfJQRnWG9RU65V2Pb86H7O3RUP8VopkklKgOQU/7zBi2DnWf9eSgc3G10LKm39UrPYtQ
sP5HBwMtBE6s14T0hN0sOYGsxZcG/Hl2hj3QdS75kNM4pFUrqkpFXo7TLgUVPKs/05ALy8r5V/UL
ZYOYIoLtSAutWI13sOY64NWHSpA+xucvTY6MoFDgXwOWE47TjSqoJqbAExQ5LxP33yoZpnrh2rO0
Rw0mZ6o+wbqm/7w8w1YyePmTZckz6OwlYVbxwvE9pf0Nk52h5wYZM/STF7FxXeyztmqFzfyxQL7F
7cl6YghRmTwfiVZYEsMQiFUkpQUdL2//M/zRhVtAtF3edFQNUJxKX1wGe5MWI3UAHe1D4neCwqqe
IUhRbsQS2wLd7l3SzJHk1sOML8LkHEd1gO55TLZqeVBuX7YELL0Mul3jc9EpaB0gafFjCn7h/mGv
60T+O/0o8ETABJxAWtE9/6w971rpbadRMFJCl0OOyi8263+Kfq/RFDKhIRnbkFIFFqAvMn36xa+A
JZCOsDvGhqu/5QO6A5F7Qh54iu79XvIXL1mC9tbXUs0bU17PjGlJVh/jJCr4r4uJQuzrJ8o3BmqO
yLklAgLa7UHHKoeDb2kdJ6dgTmiAULlRSFpJ/88bEiGIe/QSt6tHVCiuFaKgn29VMxSH+c4QdRuv
dpJ6tR+LUGWMT9fsmf35witGktzNTGukgwXa4bvNr/7p+ALXE6Zp3ltk6ZEbYuroMqqV9VYo5cRm
JR5dJRj7SSyYp/uCkDw5UsEu2yyDxeN5rlBZtDmOPGrw1E8kuvRxAON1jfmB3tOQ9hxPphPbSysp
VY6CmTLzsIhlti3xomdOv6jIJke4TaxCBlA/qQqtXtVzgwLCeEeB7swcAXMhyT8GTKLA4UNg8Ufx
vx3ZoyjFcd3mF7C3RtpSP8j6dcuycM2zZSjpca7z29cECDniZQuSLqfg6P26JcbMTLGqpK1ghAZJ
tDjw6PT0OCb0QVPNMYCfJLFoBQw/+1X9f8mtOisoPAxSuPgEuHbUx2TEOsepeQhaQbNczOzgK7J9
ukvIXc8dA1rvREHszLzxsS7e2bHz9ZYia5cPQc6otq1568G+l1P0zdtFutRSCRsejCNML4ToF+R5
hAHyvbMxZyawzSGGlIUDQDL0N91cfDaw/uxMVv5JLzgnay5irRP8/6iH6Kho6Wlvih4CiTZqN/rd
Jsz+eCNaVjnWMxX30Ez/19apowm0hHcpEDrZWfrpklRQ++d434JbvW5GINVTOumLRlbaoouEIOyz
zQXqxtNUC1jC3ALdjBfmf73cNYXr3kcp9QXZhK18aTg+hQFPmYBvx+JRtYQ4bGcZoIL040kRJQA2
JGuhOWKZ3PdkS5C4oWD0Qppi72AGodH4vyAuyUO7bsZ8pNKYlsdqaDYS6AIrybZbyMf6ghtu7tEm
reaHEJq9dBbiXoMOIYrITijUH2ogknNEng0uugwvN2RBThAVP90Ytt+IXj86efO/TLYVDTAzROCv
iLG7aoNdPODuLPSHGZthfsWZmY/Nwi0CoM0QWVWMRg5Ui7ab0PA5+JWRExY3+K1O9xgXBMEOKjfa
45xRMO6UXTxAOgE8nOVGOWkuv5+B3DDTybHg7aBmR5txH2XIhzKQ5rcp73576FVn3FW23twMIEsO
dqov7cHS/cZi2HuNyhQg7iWQkNWFb5NuDuSFwBUsLwCbSQhAa2CuDmnE+vGDiC/Zre+0OA3hS9CR
bkJui2lVi7jclMH3tBGYBguUCkuBQwTnYbW/qbZCcEFjBVnxJtgHgHd5W6h88sDR1NpFo380U/hM
A7dF0Rdm4sIZ+gMajBrG7C+xVaSkNd74NR4OSBKJ6LewNG5sz1/cvdWx3Db+UHDV1mzW5AGS06gc
ZlMZ0h+unfkn6FtLJVQKD/j0S/3lrMcoINKg3yA0wKi8mo2Ab7wI0jEv+tgvJINOo/ISAJIRtfzT
OJfUf9MUF+cICgzcye9fYCX5ftPNYe4qfGhw56Sg0qOSy0Hyxu/R6XJnZqmxzH6rREKHS/Jpsrj5
HKyQqjO9t+6nSARYyq/YI/6uMU53Oz2ulQVajdNuui5SZ7fKW/UAsYqTEOa1Y1KhlR4M2csmUADW
vA3qDIOcOJsZhW8QmV4Bp4RKFYlSnUno8UuEnObTTLzHPKzRoab3C1Z72BTm8JcYR2+u0HYvrJNB
8PhBILiL63DSr2l0qPxgm+J1c8JtnWCsrAqgl2BFGfjzV1Z7Uuw9Kgq0e/mSfCv/uxJfEh7RKj6S
7QmO4m6qffgEocAxGP+6UpH0tEKpYmInGxC+I6rtBQRFJJNTIq8jTOcvdiBGIFEeLdJn9Fx0/gxJ
dGvfM+Znmo5DyUKXMt6NUAwPdIhQWL+Gm7MzHKqaNsd1FAVS/9LTMVThJ+JYB/eix9i/oq2kvqih
PZHEbnLD/moobsBv4F/UYs1kpqV565TLfzzDp0Qga9pAMme5HMVmmQKPgaOzUBl9ozytejFUuH0z
WCjuB+dM13MtGriIwlsxUc49T79uDRUtFOPjwPLH2mKZsjIZOX36HIuA8QeV9kBtT6YtnCCvsC/Z
ZftAVLwYISYQEcDoAg6Ppzl/F/2P7WR+JibDNO2+1BctMhT4OozwuGmvUZf4kytPbhMruvehE54I
HriPEsbABBHQ35GvjXvnmK/dcEKnD3KHVLN/6MPsDbaBGN7RBBMt0/e4Z3/IlWAzs/MgbbDhTsEO
t0J3SQof5MHPC9kO0vIyrx4R51BeEp+5I5vc7vy619mxkk6aHC/rIA0nrmwmqllOaRuvGZg58maP
tBxzXl8Cy62c8EfonEhUOXfPGwUZrrt4qIkflFx+F/eSRNMJYc76yCuVej9LWgvhNBpqjRlrBNrK
Yv4tWHX3+BTxDJq67tO9KrTAZEparYRYwbxfYPG5xKb+DGUXJCliaE/0VJmVF6BN2EdMPG69FsvW
WhjdMoXmVhGZLIIseuIUtgLB9xXqXTqcJ6stAHg8/G38KsxcSCGuryJynSDUP+Wbti6bbod3abqx
/cB+opSUoSBR33B4A4UlMyIaCdKj0pf3yGsitzkea6qN48mloxmKp5zGAwjsNQD+Y+dc7L2uv9GR
dJnCQMn02uctvghIvHPzJFPeMTNw8Lktu+h6HNn3IElVRjg4u1w+oup1I03+yqtIymG8xSlrnCob
OdQE7uM3p3PzOeEvC3ruor259bdI3pZbxA2TarRmD3TQsPZmdSSg78faTXGRrP5nd676tWEuibRV
t+XMnVP0b+0GlZYc5BJdI09PaHaDaD+IGN1NZ0aJqlzKOf6P2P7+8kKbYOMKRztlOPNJJKoIbLST
LVrVwQW+4xqUu131G1bjc5ziAzZVq0APyYTSjH4VGadrGOhmo4U8P47jUYBRBCy5yVbIKm29WStP
QwrfXtZ9O2dMOJVbbd3HqugjGIaKRjakJSJNHec6dUsJG+mjEZxCQjguTzLVC37FzgX1Q7SeqHJH
NOhhtCklRZD7ov4gtO0AMFu7QOmFERGr6f/WiAykkJEqHljvRl1UdF163ihT/AGE/eTygjmVTniw
mWZiuGOZpSJH6IRR5uYmT9057e13ioJpmHcN6hERNng8PZATRnEu39jFAzjQftQefa5V/K+MzRkR
ZQ+kCE+cLawQjT6OMFdoyclzdEoKtyjD3//ScCBhi/ijpJlV61VqvBRZjpMA2M+AAH9S8b+w+47d
OgzFcXZyqMNcDbn9l+e9nu8ve42xGnFifcszcxV+RV2GS6PG0wi5iJIdS0MNJrJBn28iH97edyJM
PtpU36hXniLquqWyM8Mg/MpFaYVfrk4jI4E+lNcyMDhBMeBe3Fp+WFjKKrEjCoSgMc6GAxdac6BM
7EnyuJd6w5gNYob+VnMzpaylMoXxyPipL8Jz20UcQS89Po1vmV7QQKd/M59ZBRqcSyVyf/J5iH7O
f2xg1uAyQVXYpgnFijW+zTdhuS0gRk9O18lN1Y+32bHIwqKBixINEtu0d/4cLu7J7rw2Hn0p1mCp
5A+0vnpFCG6UNBBWMo4G3AVF6JzwAZlbtfGZfoIPsRYXGPXE13QctUBJcqGn1jRp4he7XbHe+bpS
Ax+QCHu7fRksivAldvkDMy6lWHiL7RKmAaYd+wdfhS1w5ix1YEb4m3AmrzYHd2Y71t26QG7BCXLN
JOhw0vvo/waAdi6xvddpW5oQW4sdPVY7iBQZP9cSaGy7BgSvUJmSi/R4ltucLFKsbnoFb40NNSiM
VI2p3IayZaCvPaHXFtRbJdzqiVreNRviBZ74Ae2mFZb01WGkH1JUW4ogYPqVY4acwPweadIoecSn
TyVXtkK84iRIhLOeOMLUd+0r0CPwjL6iz0YnHxvRKXkzYYhkpXkKXlMzOGflNVK5NF9mtuNmfnvR
bEYEE8S78/9bYiGfNwwZLAwYgafWk9/J9Ah7/+WSVTZvTX70CK12tIJt+5FwAhkcEoqz+ovUCHvx
HLkDB0ZNmPHx32jZHyn4o+gvjtKxr/75QE669GHIJl4BIHbClyfmFABr/njVO+NJ0cHzKVRz7XUP
8d7OTtbAQGi+SQkFGyo2vYoaoLzP8ulPEY3EIOsugJJ9UNoj27/YD7J7Bcv9NUCxuB0VjBELZaR9
1xR68/aFHdlxjBMJ1MsS6VWbDObtL/h0Gqq7TrrDjEGJlXMekmh9d24OHpaTQYO3RuPPOrFw7Aeo
ZXLlSivkGzlGnMfxNVWPFUI+4hG/vQBpDRtEHuHRJZd4jWm5Rdv2awyPfum46d3Xn/xghyYAQaYK
rfZNKwUJy1E0O9bmlb0dpn77n5rwCjYcSTySBneFP7/i2Si/8jJF3zXe4G/PRKevHD2Ezw7et2Xx
SZa7MOWkUzdY9b9GYurGvCbEIl/J0RtZ38jgLbi++nUFvdF42c2AGtbNgA06RyfbMsr6xf1dxNt0
Ygkrs3sq0F1TbXrToyxqhdMI4QwbT8KNTNxXoJqnp6xqNprxmcpZxeTlNjBh4ORpXaV1ti3gBWAN
1Pb3olDgAtDXgLABCUa+KTahaXaMccCThZTyf02priOu0W1GJYbE8XQRnN3dbiLeu1UZJhUfHPxQ
MLT7RCmJXp549kNk43+SFpOu1bezapT4KZo8F8IIUac6C5o+tTzANe5EfQMNxDkTDSnq/icaq7UZ
Qn3fWWvNKhlnw6qVb9bw6P9kgdSETG102GwKAJacqyEJaoWDLPOAyrl9oAMrGfXwptGzzBEn9Uep
XovTEWCfyo1n89xgywRmY02ayLhJT1kUGbDiIkMU0fVQn5qW688YI9rJiXucDLi+pSFk9ePC++0o
r7sw9oClqI0XgJCiTCicXa8m8bNntkqLr62YXSlLk7XojorCYycODS4yY6WxkDMR9TX4AWU5G2iN
GsWym4wkRiHRdtRZKDf6JmQeFuAtEycOzMA4WTtMvIP/0C+Uwy9ugXX3nnUU0V8NVZmMO9bJiGIL
Rwlsm21YDm1fEiwqEInPxdSjZCbAabMNot1tnJw0j2yDwbEyuQFoeWWhc+h9vAiZMw6txhvR/xF8
vSzScRnsddWWru0pln1OPdKHKdRtGbYNBA8InCXHxI8g4VRL+5aEAv2Ds0KBzs+miUe9os7yckYM
SwkV5ux42zBZcpQFu0XBSDd5NxyHO7DysvN/WXbP8dSrxw8h+wuZxkjybqjWVTr73V5i1s+dtqVn
VmwHCX65LBHn/KF+aKXm8PLE1bet4KvcfiODu4UiwTTxTaBUb8WJ45B7hpPLAcnXF+l1+ouexI9u
rBE1Q2QXK2XX6ITAkzgiTbMLr5izfUL6gXMLTzWAocR47oONgEHq7v7EeBaP7Qf3YC8UEIfyyVWy
5WJJLfQq5vOPfWqqhWnt635qjhxKswnyXPNNzYHU38XRp04arHV4U+oT+S/TFdsWk7L8Y6rALl4H
aL+InuUMR9WMtVE1TmimNimvT3KkgpsmvqucLmhKytQ16AfWNZU7olOcKrKFOmcQwklczsF3aFRW
n2mCYAcwGZl2IzPCzaAKZWIQgJe3T6+VgZMgQunKde1Tf+WLZlXZPMmLqnx3WMXsKDoP8KXAig4X
7/GTqo66nX+PHR4lGocsvvSdBWGcvk9bHMXJHdbzKHSSLkeSbU+IQ07ayt6pgEbO3j/A5CZvV+Rx
bgO71DSisey05Mmcn+ypcgte530cfhDFWbvXa5/Q5nGFCThpNWu5kRQv5Zm9QM+wi+ab8TQJNIMx
jJvPHwngclCESQ4nZpjxd0rHqPhuuHGnYqoDE6Z+Lz6woxQW4npzLKUNAwruza4zy5vpfAYeXiEI
JLU2iZXorMShopcmiAdJ8kxIOgneBCy2jDClyudj7wL053j5rQRhfpQaRt+9iAA5Rrra91GUc06r
aFVFEBP/Xz0eIP0yZpTpMsOvlM2/kZALXdZixJhO2xPpyw7cFTyF9q2OZ8mME0mOHrfSK4g/wDBc
BaHDSfrztUnb6gx1TPwgVMM1AgGMmrKlMz5RmjO22DxGAGDFbK5duD7wyPjM6j4t1dzpWrjyDH2v
0T8CeuCplaz4cyqQgy84dl5FT1EN8/Kn4S/5xVrMZ6igdStOyHufv5ALEjQgvr8yW24YFW16g6Qf
PU0/Z+KABacmL+iw6Yt66DK+3xxw2UWG8akSs2VV7XWmMIhgQtwPGPdaBpgBGfo5yL4pzlLu2DWj
3vzCsQ4ynmMP3eV630NswzDYvcRf4AwiTakWr1e3dz835Vo/t2EjJ1KbcxuZul0Qt/+xmiuPJhiE
VuQ2iQ/UJgkBbllegQlAUrRqsFRP+KjlVfksUOhoATGs3oEUf8lCFO+kwZk9hkIG4UPqdvEWi2gO
RCfuwPpzzq/7n2+u+w3QTaIBisfKbf2FML8xCd7tDOwSss5gcQ/iKL2axAHMww/aoxA63Cm+2C9A
t3i8y0pFx1ScBPXNNDPS2Lfqts+l6JUI7UplTJlZQYo2qgKDUiGnG5ki/IQ1nqtFrQH35FVAzHGL
fQNwkoOSlggFv1xALHRYFLphemB8Qpro3YkJjQQszeWc//RUiXZk+7SxjPDq3fACX4snbp91JmlR
IC0qN0fJn9nveyYW40VKUBzVo5+C2y5DBMiXP+sz9vUyT5fKEQdBsNBiBla+sFvk0PixPooYvwAU
HXVfuCJNgrDkSZ8urnvJfYzCkEhL4yg9JV13Uf0nl+XsMXnBt6vS4yI/KN0YXurqUsBv7gO0wUMx
2thPGaeNGOSU4fR8vAKt2AU/pKEb5K2AMVCU7LT5ss3u7jrRc3JkB+G+iIbbDqL4g8Rw7IC20jFr
H4VPfhTlkVIkVk5/6F+fIxvQ9BC/+Z7W5gSEynQ4iXteV6S2CIc+yFi6UhDLYF2h74sShkvANCSr
TH6e/6cfDYQUP9Mt3C500RdSmkg9m+XC0sIynQqA2giriGALoVLSjVhBOEygc+vTwevZLFA+f6PU
827hLYYJIPzFUO9YKWnq2T1DsXqxjIm9ljDGPpHuvwhsIaip4V0EqXoUfd/TkHax4ZuzvdlUqXrh
VTGfPs4cXDSS6V30ZPeEymNcYCjiwBxfpTN/IlnAs62rHMDchzFUAqfJwEIEnQnECSkeYl4BiC8c
AGsJjXDjIAq37aYfoT3QxtujD8CdIsg5PzghiUquI7y3O3RinnddeVqYoIjggw1MM7HFG3vSWA7u
CiRxvcRTAVnekXpruTtmToWtz3Y6Zp2K6kJD8eRYKjHKFUJb9hB7ZOwxz1bnchMdHiLBvKYLM9FV
m35rABawK8VZ1Zcwr4yq2lKLYQnWUmcepuk4AdEGedkiiU4nO6+g9PPOfz0fk47qdk+QXxrOtBoP
SvV40VbPh2q8aPcfM/+1jpncGqWuf5+EtK4tgHAI7Pje21/FO2pVDN5ATpXcbwkMA8W9jiDeQQE+
9LXig0l2ZcK7/rjpVCwgzGhqP8ofXPt1dxZCPq1ZKZrwNmJcqmF+fqhCC1+pLIeREntwjGOXqdIu
TDnmEEsDqJV3sGveEW0kharpKXiCXkmmag5EBWz/AgjreB0cn3ykEir4MoAqDkUy7Rs6Xmv6kbc3
LRC0Oq9bNNF9crgBCUnIJKrWdw3MaKQ+I5NjM+s5kI7SpZRt96NML0tO703/iOtYPgh42z17RLQu
SJJxeoUAJALlhD79F9MG1ITYb6jgZVUWjNSrTQWldDz9qB5THjBXV1tpXmA1f2BXOY8QLHVPqQTK
x2cF+5EfLyj+3dnjxeVK3O5CukAXyHvZZfmgIiS8e+r95zUpYXzvsTKkn/+3DHJqTaHiuQQ2YIy7
Crue+lGKo/DAoa1FE/V5BuTHGdP/+TvTQYUpWk5CDBqOfRSe83nSE4tdiFSs0b2kw5jbksmb/L0a
toPvWiHCPVr4mHcnxJ/oo4I3J8LzqagnjnaCjw7fAMEXAXQFmWehdtGQJKaT0+xWdH4qukqDN+gL
pdVAhEl9EA2IXHINr0hhaCMXb/VZx+uxnMEiReynpungWnd79lfFrX5unDtHTw/QVxuT08CNiBin
ipZIb7KaEdQusx2qP0VVCA8YpWXsSR2dD7NacLtNr4uBzxuxOmPlkNbhNgPnyKopbmcAT/uZ4tW+
w5fJvkyhM56OJ/+1PzqwvasLHzPvC6H1FhF0zwV/TEcZ5nb6q/T03nCa7igCjbBfeYrEKa/cXRi4
KgXt3MYUoOPQfTg9L2kXEvNoFu5HGJ0X5tuYWTV+c2hvlJYlSU+yEWlmLaMKq3NxW4Hav4I/ogvU
ckpEHGKRPJQ4u0uByb2t19g8nrBL8bwbX/HMrLBFiFK+J4sfMU+ELwtufu3aWLve0FxBHiu+ygpp
a7wZUmk8l0+XcHRy0bVS4fICfmGvJTpnj/OxzDhru1GadpJHEjYl3dIqQQ7UlTQu1hZHhHsqQii6
fdN7DP2sTBu5WxYJkmwvHvH0/yX0cbhRqxQaQBA3LCGL+2UL2B6KOYIdRJ02sk1+oXXtXhMu5zt9
mUCMHCnHNHUgzUUp6wB5s1UOQCxh7i9QOJzPHTDMH8d3uBTMMJS2YIJak6qu3PzZkP8mZ8NE984p
o5VDSKm/qnl1/m8fff1rX4EMwmFIKo+78XQIAcB+ZYxKZZsikZhTUAKVlRXBeskyL6MR6myPWMKU
TR4LIsMde6kdqTNyS9f0fAOybHpk5Cvq/HEgh5r3O0QSmlGJ26DFtbTGKG/XX7o4ohyJZ/AZc0wQ
lA8sdQAvSYBk/Fu6s6JAT5CCy+Febebkf8tJA4WdVrfefhGEdEcfP3UkJg/CbEQQAs1jkcPJCStw
ojx2XoxfvVeWLm5TaY16DDfWC7+M0s6wYa+eiR2Sn50pWbUGqT2zx9ShZ8mI2WsyvExQrF4IcO4n
xbTONk8vZpfy0PFPseh+0cDKc1vRRwz3b1042IUJbvB90MnBEkQWNVB4bF69fJ2BhU/MwFTX+fj3
GgQ8q0lSIS3JWLy4ZOSBZdiUwVdH6K4jAgMmK4GAC/rglFLrokIOQZULInzA3uukqnaZErbAY2n/
qJHJjv6ufa7ctK4Wo/0ncT0K9DrYhi7/7wtRBc9bi0A8lVdbAVJNJTU9N4pjaH34MXzVkvsQK+yw
xFcEqTmQ2QF2p+yYWGTLP/PFL1InSDEDnGLtB+zMKjvC52h5uSxsZ+D+qbblzH0Dim9R2wTZ+uCb
W8lbmV1YyPDAgX67bUrdfpGB85UePZe3B4NkipoiV7bJXAAbrXhQpu2LQ3qi9DVtkIsr5o2lDTfn
3/1NEvjtQti7mJNrqRLZMVo//np9F07HR1RuOpKO5Sj3uCn8XQDaWs1gr/s0oCkXYScjWyfpa82d
69LDtxY+blAKUDshG0nq4xcAOcOfukidyaE1A/JrDIAn0iz1fx3utHDISJgH6qrNZIs+9gpNSHtm
htuVUaI+n+bSKy/7brsE15y2/5xc9rzWLxwerirqCgeXey/+C8IOjAweIj+iUuP743741NpGSehc
CdR1ooc7jMvOKZVVJwCKrR8C404MyqcNNsUKLp4WDv3eWsAYPk0Md/42mBQf0hm2ASCpjysesFYP
kiwTP4WOeX2796Yov3gHt7/HRpGp7BrAIrVjuAtyB3zjV7dKK4EJ9TyeE8HqI2tTq0Mv3fGjfdrM
qEY3hqtfR8+qrexLp2ZFtYrNegX5t+6rnbr2Ah41xfCGLqERtozL9Qv7LCcVPSQDODVCTjQ1IbCw
oK99FuGi5TatQpfpL5/fL5QD3ld/gq7KaKuMSxoGLmNSDLH8/w0yBPqEkq6vbdt0xVmQkwkBnYCW
mmaFfahFz8nWKHnzMluk6PEBVk4sr4cwwYpW7XdOJ5QRwJITmbBZJUJDYuzUDUU0qKxo7zkoAZRb
HsuOj+IqJDkoprcoZQbYQ32zZQFDUBjkpz+3RmEVBLB08xp7ifSr5osm2YF2QjxV52uUzOIatbav
Sp/IUh6kXT2UK609LCfyEMjSw9cmnXqfdnSJAiLxBJ2hiWDR2XNJc/KIPWBwRfQp9K0olJeKmI5X
uT65GS+LYSzJViKPR2ZiSFsiWjDeld73q+Kh+LO69gWSZH7y9nqiskV/tljlAMCqnsPkrf6qNA7p
JtbUvRchV2iAtve/e7/sPXVDN5DAjta4o5iiPYkjGnFd1iX9MNWugJfPROFA8oDKbtGThQcJBJBs
bPLZTUgEr8CDR7k/cVUwsw4l70zqI+h1hvWA1ZP3RghZ6rpwqRfxBSDhXX0YRKjiTWi1Qi7eLLAW
4hKcTDJE6tcbrDxLjAKhHoKqbmkX2NGaiWjnWXFBgy+S+TTwVxcOMminI6CE37Nd4Zlu3LFnMblD
wCIS9t0JPRBSdRDlZzrsjK8pFOZb/XosnrpN7N9Yu6Rp6834+O2cOomoKy66k41B1g55biQjtyWc
Y0DSZyGHKAwsLtDdu9EgQMSxcHjZ/UB4b3EoyeJoqXfh7vs1zWad6Dy4MfBXiwtnQIu1FoMvD9MO
9Tv7KzUpnYZUuvsCUCO4uwm8JSM09637bRsofqFibhQcVGMBrJS3zGb/hh2GKxZ8cW/DwLZq/VoU
qzMhq4RVlf/cETsv+vWwYFEDHQi+mGj7OL+xXfIFeaF5pGU4aWGb9oqs1QSoqOkwQ1gjyTyP5QaN
ruFy37PakI50/HwKLSjqwSaTTGthZOrstjK2N1nojlQgyND0FufQIAeC6lPve9+YJdRTUaMUxFRK
XBJJkJOgkfqfEQFJRF9fBWyW6452T0Sw1I1MPZ7hY64usp0Z0N0/i1fbn8Vr8mCRNhDNSp6ETq6E
N1RatSmDEUnI1+gmAhcvVwymHkksFaAyU5d+WvdEYvkflZKZfDhhyT/i1N9O8DCRNYV8FvImJ+0J
h5UrLtwQabruaA+JXBqsCsI5Kx8F7Filcm5Q5y2DwV63wxkkqqERZYLDrr94BdWOBYgLi/LO+Y59
f88s0W70ui7DdZO/F44VFyHOPK8/8HUa6MtFRJgXWWse6FlFmBS8Qaw3WFTNNdJg6Qhf+K/FEKOI
pmXkVmcRLuiEUlEAZosp1wfOZCR+nhjs2C4n7Y5MCpUhf3d/NDANt4si61qqdEnJnbGGYc5Sux8M
rKr8RswNEBskaMTMIgU7Yo9+hmpe7EfD5+mNgfoq8cHSzyv5jdk3pLW3qd7pwQrUJeR0h/tDjMXm
OslzK+52opd8A+b682MMMX2F++WEthc/CjsptnLIzRDwovhmoMhTnnlGsqAz8WNMnVRc/BVcWe6Q
O+R1RM3X+gBRpFPPEG7pjWY7KtHWMhyNgoRAKMB7H0S1Bg7z+dcQ/gW7kbX8bSuvvp6PL+7IVh6/
OhJaHrPrQ4OMU+AGI+q4d3qDpAvRtePD6zbdWrUQir5FGV78QvQ+l4Ee6HO9iOhiKiWF3B85FhQU
74ZwWezjF05v/FhlY+wkWdSe6sZ5cI6JEj5B9mwa60y9Rg0UiUiIdVpk+jk+osMwKZpVayXn9dgG
qUdPiwjQiT2TsGnR/WTullp1u0J1TzDU9BYIJ2rIKNydIlZ+5GEZapvvJSWuFyyYu0AZLlpFzSPh
JlvC0ClfoFBm0nYO+2JE1j/C1gOANZnvvL62yaj7jc/QVUzosZ0a315vwgfIBn58vE4NmQuRb58Z
rHIK4cBGPMyntPmvLxPFWLDKQZIciSXomSehDl6UDrpEpvRIq6ViQSFymyfvA00+jn8/aTaQFLko
+rJ5BGGugioDP0aFq799AGp7wY8xo4stI5f4pXlPdUm/bGtxcK0quqW/0LGVU15UTVjPL0FYD8so
BNRn6jYjJ+x9ylAHjlyAFOGHp7DLrx/DxNOQwVJbDq3HRoZ67w1lLhjfEH8uSVwXgf3opQofnSi8
7O2L6Y1Jo/ECRlNKNGvu6D2b0rVz+hQDELZUvtGoczA9470QI5gbob/UK/2Hld0Nwu3zYFlBcEXe
XbdMSq4VpczJ5MCgPEx2ahObwfB58I2/bdTL6QBruQgreeJdTBb5hXnLH18iX8zJcXaGm+9am8aD
J9yZNF1p788I42VCC71UDLII0P386XqTu35IFs/IliZzk6wmQokHl46UovuXiFNsT4mRR036y5/V
MTIgWrid3KbjkoXjkO/F8i5Fhxy39iuIG65bsDzZmzdIZTflekMWwmA9XtxEWgRTK/puSSjRAGDi
v93H1nsJpiDx04bvkTYnqPQJpGhHMfknHKndtP+hXMQ+NmVnfLpjW6KpJNWgpElQ8w+bwL0GeKUH
MM1sFcfCiP971jGorGwVExjDL3yav1qSW4djaKyxTzkNVkLM0RJs2M/z2NI9pQoUu6EIQEyWR+4V
2Ilv5LNZK/5ZEE1mLzmfaAGA1MH2oGlyW2s6zul1APRTgdXfvJeJHMA/uEYjKUo7DN5O6NFWVK6N
HE1yZEXPTCh8qQfe10UkfNd6Quj3dZcKTq6uDH9Qw+QJqLh8JdAVtm/eRiQ1Q79OOP1iXGv8nblW
GoyHu551W/IJgmK46hJ2zhxNSmetA5QZxgOudFFeWBkAijElBwAP0QRLhzarAyHUrWA38KA+ZWra
YzgbmiPjTlgHFrGjwZG7bD+7t/JfLu/jyVGBt2yvO8t22JDXJAFcvz1uPuSAT4b7c+n0DmLrNjy9
w828xQPRwEd7dLwZJ2tV1+JZ/z4yFlybmi1AsaCPp2vrdqm90Gm5Mi7YhIepNnBZBs1f/kKA0931
RCQd5HLfD4mwex0rW5/s0faXc/YXdcAUAPOwXhtFWCI4pjRMIYlkuP9a4l8kizdHd9kW8Y7HhLw3
dci9JbvNwJsp1GAeOd6OroasCEJjxfAL+m3uM4culw0Ps0uPhy1rMY3BqfmvUoD7tv82fuGLW1DT
xDjD8p7q7l+0CLan8EftUVv2/h55hVmbdW1X39iMImSYS1Nxk945e5mi9nSbYy4+kbNe2FSZoUSD
OUoN0qjwDyVff5WroKUNn7ce6fRx2C8CxN4A2iHS5YLi9Nxin/IathcOoNsaw6xxLfy1Z6UnKwYC
2DH1rD2BH7R3UNI4HLHHAke5IAZ7XkAeVJWEYyK2NWlFaFAdC49ItchqXnmOqQ0uXrvfaY4lEuvI
rWbgxC/p+GQQFH2GQEM+4obRwFgxahYv2j/nFDikSv0IN5Yoj93feBxju5OK2xhOhjklvyKmocxS
OhU/6KjpA2q7bk7mVSQdT8ag+aGefVvMG5DNG6NFX4+NAR4W6gZIdzc1nQFX1ssJxgrSKh7duQT4
B9dKchLvPYbiEwBK9lVGW+wZMV3RBQD7GnEXBVpCuI1C4VXgsP63QoT18aiIQ6nrvd8VN8+QRzGh
mcI8D6MdBynTLV9EICAtcWYNqPDgVbTTtC07VF2UumSP1EYbk9cuh+00JdyPUC0mrhEfuQzDxQI4
6q/38qiWT543tDapibwn2R4ArbqAR94ikl1tkn+XEZHGcFUEEV4NQsSFFOvVqMy4DkpPnGj2Z+Ms
KPWJEY88+XNRY59l36HnwELMqKtqA1MTwUxru3qmkssibXFecvPqCLNFIAcDJEsfxq8AgWKhIc/z
GyOMGGv6tn4OPhQLoQrdscGxf2eBXITp2tdWvpo40y5xPvYbrU4Mhx4bq3R2SukKcaxC+/2Vduz0
QaUvOLrP/qJSBJUqC4Dc+/D8qKlUsnug8lYB4oWAnVaVJIzM/c9j/QkT9T9NMzZ0CLtuY/kxaJpA
bm1ln4HZh/quwX+06SbIH33rv67C5dXkHzwdkR5ILfH0M0HWVokxqrumR9XTWzZJ8WK+09CGsv9b
CH5neXYOrHxhytjoeNBl20OW0AgpfdvstSqipAPBJqaExVYU/7M1HWoMx4yqG1kCV7/bKOwap6FC
htySA9QSeYrkTZjArGXZkhXAwwFSUssAj1yu2RqQMO5Xjxv7vQrqCynHF0PgMg6RI+kFxm6HNv0D
z2KDYnFwWO4eTA1ac53sgMLwPHZVoYqfSBtwU2CNZo/q3A3vZRNxyOFDKIUnC7prWGiWydqmMerO
zttBZhsceQg9i7F7EyUAQkxFQ5V+dP44RJH4K8kCG4p71vcyHKc/nnhNeOVnRVgTDwWy9i0ox9Vd
4h4gTd844dg4BxKamFlQVGUPoAn5M3tyagtRhwdLUoX+w1KYjT8qqUQT7CUz0cicl9bvgYKWWgcU
K2wRz09m5Y3YiTWINBbH7x7yEBTf4ZxPvnSs5H+aj8dCBmWjFpE+E21dH20WXpnCxI1/oL8tZg1b
l+Jy55NorZKtiHYOO6+9t4Cn7d97E55+7H9UZLSr5f22VSQtov4DNBjgEDS0O/yyE18Ikg8E2jvv
FdoPQJLwap3CRWo8GYK/t23K5Difn2xJTidUr+RLXky3KKYP+/ULLx4khHGTaqoGu/Fhac3FHtYq
Qq70G/MGwXWhyHivcoqLSLX0dQaNg1nUO3b4src6D7fUt3ywIREfkDdZZ04evOk4/FtcNTAs8WzM
AEDEfNnImnUu1g7ojZHo2ALYTCRL41+l+eEUPRdVMp2bySJ2SkIRHAiorjg5GxhDpJKJ4A6JTXiD
fYB4Mb72Dfjb5VEbioobHzijZQNreasthNzpkDvOQfiXFMutuUbGPJy8Ihd2q96tEUe3GRbU6ehO
zRMp457WnKUBRAsb9DWObX33pLzIRl+dk5q0YGlvwxJHVVwNBTnEwy0ex84cKr3qlGPwfHV1a3d7
YHjWIqLKghVUOL/dUVnCYpcZIAHkVbe2QSu3Gt/uQsTc3T5RxBK7XWrSJiE/ruPheeVHyzxUQgek
DzMXzliVTgdi/lR6zY2WFGSEm/y3vZIWysIEmZ8/GmycLfnbNMGc9fNQrfuA/h5rn02tH7Sa3Yo0
WJNZcDOdPBmbMYSbvLjjUYlrJI2MoqQcO4cW01nhhmmiF+Cqm66ETp/EsPjkAYy/Fwb/xBkHEDYF
tX6lNi5C4xZCQX2NCPt711GnVD42mEyfYx/CwO84I8BjmuxYpecyz18F+hHlxFN8UtdpVcmUG4m5
cdTSl6zVtKQJt/OFT015nUFDlolGMEL12Feiaz+vSn0QGLV1ejjOTlyzxxVCizSgRwk7BwlyKWW6
5ixwhrYJpMBkjBI/9hGIPs9+iwZBCA0VvzteeNMSAnj6cXoRQQ/prfSH7oCDWLZnHBB0UxlugJPW
c8BOSc40/z4scZzIxBtUI5M6yLeWKi/vwFNcI3O7ITWl1uvp8oNkWQISOm80V/PQks4J6AZSOEk1
KTgwUNnS2GOIeKytYAK0ynUoA62o5CDv2kX1fmExHdkJ/7KSCp8ecsRKcu6hVrP2wqGg7ZZIFqn1
gEGitHs5PQhoAsubWDpxJL7LHldeQ3/3I9BgYpstlaHmQ4UwiTYv66ynmGMME3mKH0Legq78AWwr
hXf6U+vbAw27iG87p0xbcr90+QtglBrEYDXUZEK0XLEUMk27+wy6kJsT6+158wnzV0Im99TnPQ9s
MV3L2N5neAvoG+Iy8DalrhD+5yOJUKUsg7IZf+Vf/1gs3ClDFZu0PWu+nC5o4/YSPFmyf2pLjbdv
s+l7yZlxt0gX/znoD2sz5AFnW936CwApq3OTxUYF4lqi/RFPdzaq95G4pQiyUvoKqnV1mNTykLuF
lm4zgo30yh5VgY1/X71MQDNHEti6J2H7fsT9EoAFac8gnNE6jrTqeyQFPxft5qKkU5nsD43f1VJE
t/js8Rn9ZkKXB5s3LEHPDnZ/RxKYY7nRg8ajiXuDvJJM+9MquvNt6wIFTfqI9b0fjEC+9l4h5Z2C
lfRtQrDbkGB+weTNdnJr37zNsV1d7O4YgzBYpfNP/vOYehoaeuEgUD2UT7Z5kAjRmk4Ssl1a5hJh
iFPAjJInDglKWj3Xt/uFsDsbgeOAcJDG5A4TyrshviCBtsc5dXYTSI/95t04nofhzf15sDuGEE9A
l0D55bxN1dNCRdsKxgFQeVhzn4LPtCj0LUvR7VaF66XaHJvAAnwvYnnHUY40xmAWlRBkDH5LsakE
N3zyo+U0BUKDVM0xOa0T9/YoDwO8pDRd/AIMakPCQ24AeYn3zeafFxib4jqvvDyvbJ0pMUoiI0rg
6DZcPFqWcyQS25VXRaU+bnua5CMTlagv0CuKUPbvqQQFkZbSbhgh3W2TFygnw0FKdRLgG9Tkqyqk
loI/CceCisBIL+fzUZqkvIc+Q5c7248EOyxHR5tY8cpr8vlS76i/DJiCIho92GUhji37iVHYI4Oh
39mMWLmg/ZFcbfgHUdkeGWqN4ZDm6pa+I1jzou/ElT0CO19iFQUlpA5qdp73FbKd0V4yOCKRU1yi
M6biMiXSIgu7l5WiYTgjA4GzCSUYK76Qi5yHaJPhSsaJmhdRTDtXW1c7FQ1Y1e/D1zyAdivaocEl
cn4Dd//r2JSfy530kyPwuCELeZH3u03CLEoZj2SapAeGTjRWRCcR7UFqlNpMaMnjbHowBRrgPLzT
UstD5ZYQPjt5rKVM8NgMb21gCMaqHd0lRCS+pOdj7fXeyYLncHQG4qFnSc90+hpv0c1LY6I/nE+Y
QyDlpJskcB1mB8QwJdPlUdyzyEo/TP4MXCsYCFF5U0wIz09TLMuTSJcJeXhhTZopf0bV3rX49wB6
8pqwF5WAbDf5aCe6BYB/QuKO8+068SF76DwcoN0VhM0YxsUP4Lcb4yuRo/mTUQyaK5+L35OxwMnC
gyLAZjgia2UCyodvE8dsFbYMmaKr2rb6veCOwmvGjKvJLNoHBWF9H/aI5jmEHfpy/I31e8kHKwrL
33Z2vV6MWt+DiklPcTYZZ1SW6TALZGf5fnaK2kuL5rgt2rcuamydpWZDsBpBgODXcOAozgwnOCkW
7Zb4HKFQ1Qdi3zv2aV+Uqt5s7ngn7qK1uC68K14r7MRDxUphTmEI7NqqtqLqYCYfZMu4+/9p4z7t
F91U+zS0pce9cp6pKitedpDaRWGJVLT30xhqC4dHHT7xjtcUNE4pjNYJYkV/zKw1CXfr64Egykoh
eO4V9MHwenm2L8OMZFhUbI/5IkRJ6iDmpcHQzWh6R47Z96tKSdtp87yQpjO68RzgqQD5RC7zt+Bj
Wyo2edgyo3JnpFe0W/gYmKXeNVNgD16ZGE4m5anwih2n7LLoeENFShHdZS8aev+bIVdfK7LcbjLg
RMpQcxKPkA/bz/gReTKw1MRCd1DXWMJCagkpP35QjRuNPZMxpAJ9EZ5JSdSie4p6vTccOZLjkP6C
Tqx89CPQdhJSYui7h+mRnyXV2P9NTCn0AwxcENMAiFJcN8A7ry3LD3O5wZaMaIn7jxUAC1JKGhf5
tuwr+TermmQx8M8CWvWpWNLTVWk9oTkFdf8X4s3UaXxNnGge49xIPYGlPY4cD1ecomqNwDrrgyyK
iN9nvttEb3CtJLm9zZxI9Nu1IcRICp49xJSh7rZC6/VAd1s+mKNgq2Ss+NvDF4CKLqNWChHWMb5w
TJLxmtCFLaIUx2OEcT4fMiLU8l7yAIVroz+3MI7NN0YOQF/nbjLNU0DTetWeKcZx01tKA3h4lzph
XJgZWLyG2xEHseq6XAb4xeIuGS9EJkhAmpIkhtN7UO1jDHGU7JHGiPOYFetwPTgwwg12UP5fc6Cq
2WU8AQAlBsrN8hql0geOMKNGSqmm194cw/qXhf5/26KR6YNcz6Ost4h/NzAbQRHR5eXUNEXa6g+9
F/2EQPQRnsOEnZzcQR5QkprcFZ0jJLEHHV2w0CE/zyGX74+G6TW3cSuAJRQL29cpxApaWvTjvhst
K0ZdzOMqmFvuK1hHypnZO6AqYr+E0KZPQCLwWb1Ll53pepDum/6WicubwoQ0UKS2T5/LUXezQ8IW
IXtM3+h0d7fQXf53zy8G/IivuSSf2PfaBeRMchCsDnMhvQ56FBQHb5rM2CHW0CHAjw0MOnUkbaeZ
bBanbw+TYvxKYusQsrqsQD6+BoBoAMoI0ogIUKrnj+GHPd+NmZb/ZvUFh11fgfXImvE+5F4Z08nZ
fMW1LuBuRyT+sbek9yxgA3JXhCG+3Yv1/iO2bwj7VjXVPgLpC33j9Y1fAShauX97HwMDqcUFKxfT
0fZQhQuUA3PCuhGKUg/1+ng5QZCIW8oT2TNEqt8f4qQ+JPqqXzpQ7YNBC1/PrsB1etxLbfpvHxKN
3WEtsNFCFRq5vksfunPWRXG1RNONXsj3sekwVmdaQyA98Scd0Bbix4bh49TMaipjNyOSBvuNUK6q
IG0cFHwZ26VDxrbhGP+tATikWdSQxtf5rVpfbJa60hBAWRSYjINLivP+bCFhZxLAmdvke43CZw3l
cUqU4vJl/GTOhcF4JTmL2h0nowR6bgf9vfGBdrOXVVIrTEMP38Pja/gZcwZOs0qPNHnCCu8NfpgE
uR5b+8ZU698S/IahEQbzjEGBC9pR0mQwdSjYYqWGZUG2w5sx2XnxHGF64g6tOYJTaTfZGE9AdZDx
MBES2myQFKmRqN0a6+Lyi0Liok1zmEOqzsB8ruJjafZFVybLydPNzyYdT2bdP5Q1yIitjIi4YPkS
mFl5HqLlMdNoTKB3Bt/QmqgHMgMZQC9g5KowXPSZU6sA/Tl0Fc3IsGbHpukdNCBgZ6mJKYqWu7o4
FM/TO/TnYYeVqwaIiv8fGh5JZqabitzpNkL87Cn3l/3Gy8VsIW+P/1F780fHfXjAKXVuOIMWewhl
c4VJYdcHGCOWAr+cMT3rqf8HI+TmeyJwOX7aLo0KqaCd1dQ6Jhakvv2Rncf8sbUtQTqlmWvzWPI1
ziqH8NdKyqsnqMLu2t/0dO7SORrI2ZD1VDb0K9LOtACNjr2j/t0CVp2MdAVqzyVh+UZ7Q06noWt5
AfVR7ZulP6Fs72zDcj8/l04RKXwOqFifRGss3xHJGTClvXCS+8NrrQHoHKgMOLts4i1+ysVTwa5m
P49ZNJ0NFJM89AjgpiqHz+hX5IFPp0jckMkclsY0OdhZF4f1hO0je/sTaOnBAr0o1NxE+1+N3o2W
27w/SWhvZMyfTbik7I2RPR+9TPhcnDf5uNmTifr/v4CdbMwbMWvM3r212nRVh6udHvOgZcNVEywI
GCa1sR1sjmtO90c6SWzMiHYpNcwvWiJmro7edKOvjs6RYayrFy4oZuvWEl4PtgecuqBNxAaPpVG8
B1puM3ip8zJQsnkwHd26q29bXNoxfWj1AqJ6VceVucIViZ8NbudTOSghYwF+vG7w0d1P+AJm5R7m
5X5rGxaupPzGNNMMv265o5+D+ORDihiLxDo0A8nUl3tdnizoC6Xke5tWIbQLR2iZNqApfeDtym+Q
zL9PcDyuSyDb3IxjoJDSRXjdkb03jAu/1Bj2uySM97j5dWIWAsMI8LW8GPkbfWfx6m0iYnuLx3oi
E8q1EWgsHpjZYQp288usgMfkJbFkTo5rH1GohD4KlW914LCpmPnGXLtDt0dzFX8g/3H7pAR7c0Gf
b6QmUieG58bEk+yXPtI8tu3hKOcdlPCT7tGIUexMD2Dj9yzq6wP0/aK4NQ+2nTNezNJXSmCMIJYk
B8g8oCbEGx/XrjUVfT/ZLWWX2nVy94o/GiNaWIH/wyytKUA2F965wotziuTpNzZYZuTp2QMufq1v
n2WtZMe0ruzlLKG5mLKRRA2/9t+mj9Gc8k/xCK5bOZ9CEBJSlZiTH9Kom30YNMgUW2OtsDVI9MyX
t8jicGeBIM0/Pib7oSeL+aSYA3PZ4q3qdlYVu3GQGgbxMwATYOKU/yy6sn634b/y6Uxfc86So+4G
cudVyagXRG4uLCZHpD0tnqe5R8oMMUDcmiZoBtLwfpLJySWKzX/NaDwHGL1egECgchcw/AnNh/i/
pITE1epvL3LGBFCBK1FPYEjzmWsYrbxHeTe53joXvmEGqKoNwdA4BjYf+jdPAGr+tHdChntaCSEf
MXNnGhnVF/gJuV9X/o1rD0UTo67lkjUB7vajCwRVFAwun7exrBsuj2ut9tnNaTbXM3Nzl2XICw4y
/ul1jYpHMb021WVChK5ASMQ1Rbamn0nzP10ib5MdNZdynl9MLNef7Nn77H7h2B/RF2twqHgMUxlb
ofOBsEq+GUk6XU7S+aKCieefYWiDUwRqLzKjM0xz6aBegVOh2MRmmnm/f80E119YQhO38ow4KYWe
/xHfX3RyL0HmamZu3BWEvnohQ9at+iLZyXBJinPpWGMu7wG1ybuvs1ov/0cH73rGzoCoC6LDz+t1
hs5kVR3w82S5+HL6BBo035+m1dX9ht9hlQDkSD/zD/pnU7iYU3m4MIYqjqtoZ0mWs/AJU9JcHWCh
StWgSU/0OaPzwNw6VXl3/6Ob+25YnTDZQZ9yDxAV2c7sFeYAv594sLbQDHP8QfjB2ljO9x3dvfxE
Lxg9aB7uoRS2ggKvkNbr9/AQz1PfYtnLbA33/0lM0iI92yurKYlmc126paHA6dm3dRwSVP6XKwN8
BSe8hwMbPYFA8eqxXn5vRZr1GEfhb/06HjXqz6UHjobXR3wekgeK132hk0Q4ZMGlEwQGUoVvLq5+
z0fM8HybxERHdXorr3WkQ9XuQxgcwupUFPJ6auwj1rqvoArixnDzpxIbmFkvGxDGHV7uvO05ksTK
dfkSERVxpp46iFEmjvnhj4UMlSKo4WeyPV7WZNDK1ufVUtKSm9pS8Zk83s3pONWlQVvYGcTD1eU1
irVrvidA93e5JFzTzbJdQ1WNeqaFQZsEKVmxwQOtPPIkf1nh7jr5c4M2W8sBKJHlmtWlnr5Aj5G9
dRKKzP92h9s7v25gqcTin2rWb4FWDuMbB7AIkklyRB/NGKNo3eAr/wdb/jHvrueDaNAP5lXownbP
TTPeBGmnMdAWfhisbPVj/rSbovXpSAeV6VlZ2J8dkGLxi6Dx0fh094q9vgD9tYmTaD34iOdgStu1
b39MCy7sgpnaThrQfzNnPE7HSxcdLb6S108Cb2ZXd3+A7RNbQqz31Q31kbiOsz1sKl7nnwgYdQZc
EAwfPweTW7VlMQTzIxSyAEhIk5gfqA3c9NmRxdjVbVqlcFck10VH5In7cuXUNRfxUtTEIB6U3wmZ
Hd4ECqDssNw3/HurNxNwiE9ShKtJWaXBPRMstpAMv5KWcUFqZQfAPW3dN8zGJcDYK3Jrss25bPc+
m+peQQRIT3iV8/GDq7qYj8wOvZZ5sZzclM1i3Bdxy+NDK8ubYY0xOMUWIwpnF7Be/lsBzSQ65rpl
N2wOCWbBccycZGZg1KJdUc68NkIMgkROzNU8DdXhT9usUgbOcDFNAw6UUu4PVNBbEzLIs5hWIwgB
lB9BOgEe/o8L8d2lFUnIWmlEdXYCDXTW3YgZFWO/0hSoc3aY399SmJKuVbilCC2n3EyjdKNH91Rp
0Y7yUPWg5DQOI+JH2ezTz1WxZCXIzqo8ArhW9Hqdew3bR0mCBpKd7KzkM+xaH2fDPuov6zzmNVCz
ov7fowjdO1omFPpZ+9FTWnoDt7bROmeOe3hxih7/Nb27w+30di+auahzM9XsWTbvuEw82xf85X5k
DOYtsOaBzSVPPoSxE1ZA5E8XTV9G6DFCvaR6/KIoEE0zSlUxvGghasmaYzkkLSL0WvelqSlIuuac
HTjvtRXg7FiiQ1gYQmBonlh2YFF+KilwW12es1jR8RWweA2y7hoxB8VU3L7+9cHDK001jhqK7qcd
DK0K46haX1rZ0XPJOFBjvhdnUCaRgUv86UuJUqA3zfMcGeSCZpf1SaNyTKWJyDPG3ThIcrkUucuT
K/8ctYQSA0WLI/s2p7EYJMABfBBbKMkCWIIbRamnjyBUxApOzeyLk+9OKqsqgmAHM97hypHREa/t
C2IF2GF5intJ5brNKFzhRsSpbq/AQwikRIfql7dcNLIr4lRbK8ewKdyL3pz1fyfJCjjUNP4lTbHh
1SvSUUb4KdLpzFFdoaejH4lBX8iNFtPGIQOVRVOGBUlBoipX4d38I6ntK8+NoJyKsZ3RFFPa+p21
OdNCDDlbnd7xUd6AUf3gmSbmkbNTfd7Nhp2Ohb7sr5KoqpBjsPzBucz8FWTlvxO6af6cA7/C6UO+
G10qogKXgLU3dynz8dzkGan0M6EsiLd3hez2V/N2GE5x+PcNR4U8VuBa/34VrlRn1TWx5rAnfSRc
8vYrFrYv1N4Nomw6ELol2PkjtXahnYMaDgxe1u/9vkB50HCPcJRl0lqXhL/wn+fUfDfhpXjOKP3z
0zZb3xsUWvlO6o2PbyQZ4qn7mF1mE94WgGXiqJp4pV4SjA9OjTCkAHsaaVywtngwbsp4Cn+uqMRX
OXPOHdOB5zyKHvUmH8pS9Tr1Z+huDNEjina0NlgCV0TpG/L1PGmdI7J1fRgw46zfZrSxFm3JnIY4
J37j9ANcMh4spWzo73PyiCEjBUFkxeI2/2Hqpdo4vx/YJ2SWDgNP/Jk++sCA+fERNo5QN2rzCy7A
PL5vb0OV41hFsTFPsjNr4Edg1Qac16CfbSrToWFgT1Pm+yfXw8SdBZyjuvyZqZ1Cv2UREXcfAMFR
CkK/bTg2p/9LoFAJWl1QgtRbZ0DJdRis4SETEMsAvlFZCcKzzp7FxE9kG/smF9CJ6ZLARoPvdv4X
cG3FKPehEQ8gvw8ZSwWlkAcnlsVNoJ+eJUFjr5aMCZguibE6ChUdXVyJWkI0MdmlqsTdeoDVabsS
XO/p+YqWOcUbSHQca24iysdiPahv+M8FK2q50ehlXtrtzA1YmdiNM2QDC7B/QY6a3c8MyY3WeBDe
UrS+dlsuR0Dtsw4KPBn8J70je9+FboMcL42VPGl/yBnvFzTe+39/aHcopRqAlE4j/GldDscNveu4
a5BHrl+kZxpDHLmR6InLUs4dg3mpCMtdhyXV3wbbFRpZ3kqiXqIM2Y/Oy9vajdPMMTjCWI/rI2H/
ktIWDA+OLoHkveVpLep26us4sBChGbBEof0aWGwkOByPKJ8BG9SBTeJ+vmFXY4MIxwyPsleRxkgv
+6KzYy8hdiRoiSUzobF4jWdIVaIgs+dd/HQ0AL4tq11h58Bvue7u2mHpkNnFuo/HHS+ID/F7POj3
zCEXd1KYtBF3ApBI0tIPjjCRzmZUm8zMEXgDhPtkclTDEOr5MwMx5GIpVSLp33rS+B/V3wwRg/u5
y/ZhMA7Z6j8UR9I42v1WBoPSCGsFK6L73hBE2/DmwcbNLXXoMiU2X2g0VpBlNZzXuUOIr4/1D6Oc
coyvTh0oD94FChsz+EiTA/jhKrxJZ05TSIu4lP/0XhlDwhe2jYX3XLz/sc8SYNKCweHkfM1hVaDs
tyc0TYEYW5cDJSFu1C/fEi0mcnl4Kk9xuawYVuysvE0zod1h8KU/BEIYLYlPv5/Lu5rbl1Q6lNWo
inZfAxH1zOE7YQHooW3puZ5sg/H96VAAYvyYuiuuZKvW5ZOjqN3Khl9orpb6OumSBZ3a4380nFrk
REqMcvGaVbcJm3OxhJvWDcqyn0B4EUtg2trSUOelRRn+NJ4j3R40NMgBpJ2SyBHZB1As5HME3DS2
ljYc0yp0zoyHuQlkI6vv9d7Del6xf1STwVWj36Eg9kd7cYY/+kbxlcCNVeOFU3oHKCDpDEuegY1D
hph9fc21F0mQ22WJrZFEs9ErYRBzx/dozcZSYW2Ojxq93o8QMu+OtPKjuO/Mfy6WaRT6/5DohPqm
0Bhf87g4aYKvfCTNRrm6RsZyOuCISJnfR0+Pj8Zw2xUKrdqaoDp9ZRGbQ651RTk/juiq2bBeX2Kw
+kwaSIEDr0e+Xyq5OL1BX+6BCgd8w4w36adADvTcLXnNgGbfCzFYc0XbGaRdNn+/fIfms0hB87Yn
CImlZbkZUv11FhiHK+sEbWoSgglT9AaKIdRn8pSvTOCnNFr9EkfISztuNCJ6PgUgaFGtP3U6PEvn
eEIoKcUTWaRcIAAvBtC5HR6/MA9j8S+WYzMBGTI6HKJ0zx5nyc2X/6GEVxOY6+0YEPip9lb7vROK
WDPOzuz2algRQtq5jgcAIPfSOHD5yGK/1r3TC5Hi/dGhZTcDHLzakENkB5cl0biNJHX6dRak69/6
xVSR79CJ1M4msGuPJg3hgHeoGaLA0aH0QAO9y5UeXE2Ur/p7OToXMP7v0OA1/cCAnT/8ERwPDCkS
6qts8UHjvELJHg9CeUCaZ2kaK+blBEHPA31hv6Fso0TskvGtZnkx2D/gsccukVUJfPe6Q8SasY5m
QLeUodKFfO+mO1SFuROiGdhiV0c8hEcaC53mS++lTfZgODILzJ7wumUrqk8yRnN089lc5wHAce7f
8HTjM80jdXvXOo4u1E8O79zof/Ie8wLuAWeqlAbxYHHdJxnS/4OtG7RKwEQ1XhC+8IdzVPBnvlVo
Yz8R7/z9k8fgpFOhv03CHFMSif5hHjbN9qjurEyMo6gVNh76bn5NojseBvtne6Yx9tPm/H4rK3tj
4q8IQ5bGXH9rqUa8wv04Or0r8EBPqr+BuzOK/Ac0nrdWS/fqgpYnpAtrs/StPCHoLZ7hNm0OgNEz
HN7S9yuC+3R+JBeMKs0uzIf1fXptKDdgMDv2OCbLWruhpMqTHSmYbM4Fu+POCO5Q6ErxC5m01XOO
Yr9XnnuWJMUx4pxLyTfsbU7oS36KxPJ51h5ZRIjDDqp3jj76HvK3veC/nDCSEpFPnYYcg8qBDTmK
xDn0H9VuXVgvvaih8YlLK7xZuSRUCCFZUhbzFwANdOAAiO7XpIXqVbWmu2G9w7kUvXPX8t5EY03B
lon0h+gZU2oKYNGQNLMijn72woONGGDq3Y/4LNT81plBKagzLbrgk/LzeCfaiTDfIbPWX2zgLZDl
iZps4ZMwAWZ87Tw3WDlRGRld+qvocaKO3OD2csRbWZLbDzLw672tdsqISxqvsI0O57jkJ2O2LoTD
VDhq8BPvANMhgmBPG0m8j/uPkku8f5AYE53drfRUqGzUi2L/CBDzLL4XgTRK+REUzqHO99dp3UGZ
qAoeT0CWvajQmbxongg6/vz7KTF5bi0fJIAH//7RoekqRXmUGqCsWdFhyWjHirtVmrLcqFA/N/xA
E/CYlIJ8spG2ufJtuGvL3YwXzDVQCUICJI9qfYle2sKFOMbHpewzI+O7TttUyDzhAoqSKywoLCE+
Py6fjIXujyVNVaX5WtkLZnoHSiLvAxJvqBdzOUhcI1T2UHD/Wgxk5jJR2cjoSbgyakUKdq7doxPM
BKBYG8p77k5WMf3a67VlnF/S84qu4CwdD2ZvI/AKDYKNriqScRer3+KkI1Ct6OlyC7yxiPp18w1D
ld24E77JbwUD7vvSNoeFMZzflyXZSE0sanqHbHIQpLgC+3p5T3zCTR/X0th3/2qCpqhMVcCLqGGB
ixaS66NZlNiA8WAkdE2mgqKe/fJeiweuPojqeYUROtaapiBmT7Cc4nmD+4rMp5VzPL2AyzQwuYb6
N2Mhbu84NL9COuoqb5w6YmJ10rOe5Od+uVWEVyqIpaLvTtIH9SSgMMoZnuxsfEJ/s9hB/PScRtdJ
5EN/6jhoTXOg+69AKt9hZ+/w8ajoN09mQzqpzmwBX4uVQjIzlMGiMUOjlFWR7YFBBelgvjYUX75C
cwuqQbHn1a9ujMVRYgfupOVGQzk/akaY7r9c9B1rpskjwN9DC3BzEs1aVF09ExDt7gvdJ3STuJfS
kzgGElYMoymtWQ3Puq5SVpzXb9soxxFawaUu4D/zI/J+Kuva3TV4D0XCuHePCRLeBpq1RXF48pva
NLc0V7GqwRgloyc+S69aF0j7nnnMA5j1PB8zyYbc/eakmyJlXBE0vH5FDHqk8R6m9Eh41PaUQGcr
dbGtdOqjDGKcKSci1cd2HI15T6iT05ylVLARDRpB7lnUaxBSHAV7B5BtHG8hFUQAi/ntHVybaJlf
iFTQWa3AGlMja/vhfOcmb3ASMl72+B45NGozgw0Lk8BPSVBLvCjSs2vWwzM9x2CrQZCAGUl3qFWy
jdZdG9kre2k9FgDcrh0/jSUT8X2iU5Wi5sSKWhf+6h4LVTrWfQ0vGivCH7W0RFeiMxNWMMw8smM3
z5+7/qXCBXU3NCppmM+8J+42lxBV5+F+5MNgha+FUG7zy9ihka3zlwYum9goK2yX+rm3KuMR/VvQ
t95iIE91n3c3NNsFw0nLMxLIBk61wuSgv4bIfx0BlSnlB3J5aCSieCbtr5fwekVAf+AhJp/9vJMU
n5uZBTvKKAQ9tn1kbbTbsb+beb7w10PtJWdOBJT0YHPKF7tMZ1rVOY3sBGUrrEedwdMqaHJE/MA/
JagXDwyCdfmZy5TmXJHpJvgUrj5lbxXi23SL68gnPd5ZiXkDjdxyOmAGvDoUoPQ0ikuZFMjdwB3N
sIH+Ucud4pHiDcT4DQfuE3t6bOtF85YmcAA8FqMzGwn5/aoOiIw6qHUpypVCvNHIKhf9GgB+2Qlw
PYHL45I31DznumQu9OrWRcPSbun40cLZkou+aEFKQ71bgWRuPjUJXu3uk3YLyyjMLBItKZ4b8hUd
hPfbSqATFjyWYJw+nf404KaUVaqkQ42FiU8vxaq9IxAOPAEEK5SIailGLA0Y6Ij+/8149kUPi1oL
OkfH7QSS3oLVy3krxEH1fGoirdEgK6L5rm3vibnqpxzNLM82FtKr6fB11RvUVd5lmPEu6TYTox8f
sr3DZ5In7h6jMj72jegUOJ0XDVatu6on14RS05Oml6wlxv2H88L0XB08JmQzv3i+f7dk/8PeaxXx
yYPPehlYEU1R9rcykPn4ChHLvsG57twWFduq6R16IMdrYtG8M7XsL3rhnyJDB255EZlp3xJTAptU
5gs4VsltiuNrThWiwd1Thk6i4BhbVqHqJjiWmcBmZJ1PcxkoE0eDECublNX/fdIWTfASkqLzggG+
KXjWFytkVG8dDWZfG2ErS0SwL1IUw/8Vca6pQNDAcE0Ff+ZsicnxkZt8XEzZJDoDIVvBDcVG0+U2
JQm5r/QBbyd1xN9jVmuUAVo1lKYDQBlTvndUMKoy+Z6mgFz5pkL00GHf7N/g8EsBWBZhUo5odyfM
YUbnfrUeBnrm1GB75yfnhdl4v4z4FqJh/LYmfgYdrxOPsUqkpr5/8rgTCkpnESmPUzkqgSiexbCO
H3sE17O8Oarby1HFWRxEpc3xDztduk+NyfqLY3EVan5IUDyAhMDWuvG9PqGLbEA2El42hgeZyVwC
piQ/YZcWdGxesPPRZEZ0HLpvqEWpl3cGOqW81sy6t4CmupxeGyqmrd9g0C7VTCUbmig1r9kqEkpe
KbJcUQGKmiOi0dHEMzI8w1IGUmYOrVXCVbaSsSN4B416dMkCe+tvl6kpn6cUehVeGOCmtsPtIQ96
J0N9ZyZw+f4hHeStz17Pl1ylqq8RGFaeibIMJ+Pog95Q52zQDNPn/84hL6SQuovPLhvPvFKfFy7D
Vj3OCU3pLx8Ztr0xKPggNQeyJVU5SUPCRzCrwoGr5tAf8+m7azmF4SCQvOoq4fOxvq46YVCiUiNf
TYZrEubCM0hPVztLYD51tak67aombio2jVu3Ncd2c4Hw8L72hu1GmvA94dvF7ZcJ9Tgen/vCWVt4
RqWvzxdfMapm6uDeH4HatvKzxzvvBaYwxGMnPN/Ikhi9DkTx0ZXVsUkthbVTGuKBgJMosxIP4Kmn
p5epngHKtMa00+Yj2WNdQkhepTMU56SvPK/TptXAbGfYrKN6IgfSpUp1GFTuLhmGPIvCExJVNvI0
c9WeOxVcbSJjY5gyiVmraxww4WYoS8reHiS9cMoIi8fBTbEtc24lbvlnWy8tvSH8fJ07VGGM0Ais
fGeek8YprBgNCdzYZyxC0k1tFwKxPWuAaHuvOEHPdlz+rJtzliw1xGZmY9t/8pdsE5e4ROMFJb4S
45cGukv5u8jpJWlMJx3inoGjVJG/gNJwZbOaTlngzHnEJI1MSLuBQFDccWQtU0GWzaZNoHawVYq3
gvIR5z+YjLMyZZ0Jr2+/CF1e0buxGdHoiCFRVp+yZAqR6+bmVcF6OFpFfFkkKAbRnB7w1UQkeVt1
Eu7okcLH2mb6Rrmr2lXzfYxO4JaM2N5ch66en97iYI6xo/UeytGdwYuENgJ4kiRITRER+Xg9ohqg
5azY4Fl/o9OAGN+2TMGE8BpWzZDjQ348t34mnuS0EKYrMf7fvNrV+jK6HNn81yxL2IdrqetsldGu
jOIPOKV5Dp1U/naOmuenilqBb0w3amowpFDOYFg6VkLnPC9KMIMqGS6pgRIcmHNqMO5TZR9NcD3x
aoGMFdvwI5zc8eXoLNsP3WxfPugUSrOxBhV5/BBz8vLL1mFrZL1VHIEX0Vo339m0Wb+Y6Mm8smy7
s7a1rP0zBV5QU6z4D1Nslf1eGIVGVkGTXY2O4ynDyHy9e+fiSk3zo5PpF9ACbYrIMVd6iT2P7ule
2oVEugFAIZ0PCHcWit1L8ef2Ci50JtHpDi3U4JEpovgZnGGEkhZJG3jP+OKvqu0QHtXHVv5njjt3
emIBJZYSRFbg97W1xqSSzpg2cL3pdkrH55lGg0pbd02l97vpQPmE/Y0Oi1mR2zsMnssgu7gHl+Y0
G22OyWLDRa3/7O9t6wju0J8LNSzoRa4uPE01o9ls1Wtv5R0e4tYRWEN5eABLApjdgzol3ye9Yc0P
y3mlNTPwpYbZP7/heocpcYf0h46sKC7+HLqXbKdSKv37xQB0tcPABm/HGDEpKgeU1uvWVtXZbHik
v2XSd1Bxc7VeXP5rny6r6kNwPAzcFCyOo8RiVdIl4BKgZu9ZjnioogK7RV3rqvd8VDs0XAxLbILe
rDDvjZUL8hEOr/qS66yfjzlGZmAbCAwWLMhh0Zf5PsYTCHgKclDmeGPEgpSXm4SoVbipKPCDgsuU
y8tIC3y2ufur5QVFb9OcUO200xxPzHJRL4zfOUT5Vy0AIE/f87fMQ3Q4g5O6sDjx+WIrkjeIrIBl
kJl9arHEYalTaruutpoAGy6VcBdrnyAb8SzskSa/Tv5NwqNP6qtYg2p+U7QOIvwjaWOqqQUjs20j
/VAYWztn/FWGxN6dIJf3sLIaIrf4H9M9lTPvdf2dxuwBidcFYrldSPMNPgASp2XnSi3RLLpNbCB8
B+9Ufw4DO8W7/KuKlhZELSUH+M1pgcVILuNKxnbrh/ucmip7ooI4dJAzOx4HtVHm7m4lCOYc1sXf
qUCYf6zMrjKJrFpnlmy71MbJJvu4WovsltAdzttsfELEOLOQxOqiAfiD50ORSmKrcI0OLeVFRHzc
8ajkyQxB6NC+YjqMf2+b9jH8OFfi0DsH3/J6RL5T75HaPPlKxYhdttmsixafL84zpNIIY23lRd5e
gViveLpb0wVBe1PeWVVkYoiH/Hpijt8nDZH0t6SwEULXQ/2Ua2zVeFVDoasZnIvt0cjGwkBvwJpY
XhL50hGSQ9J6O+2/V45HEzH9sE1pU36vbfxeaWSe8s63ciB+Vsib0gp4gmeuEhYGxHbxfzaZWIx8
++GtMRyCFAWYO1UzTKjoC9E/yCmLGxkoNkmcTLNM/wj+nM2inEpBNJKQRmaoAaPDFGSOgYtvF1Qj
LGR85r857qEpHvKVtlX85lvBx4ZSu8wXqxcBRTJ0RJtNbdyhJOr7GRHJvmtXSjpDmuzF66vUfgAd
G/iPWc044N4NbgaqZ95PS8p52ymrSTdNHqWzXdaw1ao3OuvHsuYX023McuvcSrCcKaqQ8ZCaPmPk
y+4MoVp2JPSLqAKnUtPSeA4usxdQaOu+0DKFxH2p72n4eQpkiq73w2sJK7xsH/KFliyOx8bBmp+o
jU+MRB9leR0q+wWFoDJJN3XblO8pSTR70mk35am5vNLrfgwX60hEsS0GL15mSwcIBbK7FO2k1GZP
ZV+6OC3vohHODqkFiHho/LUBn9qOR6OhQLjlONQ6asg8+9/bLujXXGjCZywORPzpZ1t6DC82CGXa
BkcBmYiabpIUCRgS9m/dzkOwKfW1JHf4ql/TnI8VaYPUvFNm7aoC4ecElXfOjqjrh5K+jNgEVd5T
yisyrLvv7do4/LAYdB4Y+O9kjAEKDiIBX6C8xyA/nANW5w10lJDjyGw6w1bZ/XxuAt5YvqH8cXil
0IJlOB96wlb0t9+LD8wvJxI1fZfautPzQFlYBgfBTAqPLg/lRjvwSatqAd6KVw29jeFuSnYBL+kJ
vL3AC887PV1TOTG2MipVZiYt4rftDJsO7F6kyU1CaOBvjvezOzNCuKx1ovjLwT0xiRaq96/iWO57
+hUypp7UqtmDRL5yLyBwsG9AfI1EezsK7Wx6UEsYHYkCeBtVZskZLxyjUw0Q1LFMZdUGvT/V3RhD
me8U4nHbcMwKbH6NorAlwubmSAFzCPNa8NqQDDRxU3qHR0ctDz+dAUxetpwmoNqG3/T326q/+M9t
QLnS3ioA8MLUd9aPYZUTHHTnCyFlLsII4IgCLmJkT1X8+imBDhhLzT4dAKp8TRnyTMkXTNYnrFvq
85AnV1LGn3Nfl/e0/62SkRajXMGVIOatLqgtBNak1wH3hLTgdArI1C91QOmtnFgADl7ptnpJ5bAY
FMw6A6qdaj1Awq0yGOLRQzG74PQllybQxrEHv6WCdF6UCFq8qTxvVLspOCs3dbCd53Y3AKxJeXvW
Q+sJlGofOj2t+N8irJ6cSIReZfrnuiJefTLrIBXttZVMScf4us+3IEMvdiQ+kz14qhA0IUI4Fm9L
sTNreM6+oZnr7yQat/aE1SJkIoZ3LN+Eb1NB5KhFtFO8LSm8VvR6dk9WU0nR64DQUKtTHD0MHPov
BD/bMiEJs/8JGb/SrSOt1LHn8+PKqqdtHdpT2yzTpUzAkaY9cN9egE1GGDYnwwXUOFou/FckP5xO
DxgGnLdGaAePSibfxpIGjIhV9fUORAWx3gG0Gglq7Ud1aHgWaHQM83x4EE37D2V0E3r8nQoImszv
JvlQnTCrYb2Z6XncD7gCHDijwKvzHARcHDRz44iTey3d+r5ejzExhTX0FS3udv/IsahsdImn2JNF
CjR4pLVujSfksktm0fAZdu6lvh1v01d6iSUKIOgaz5uYk1t9i213Mqn4QEQSEaF1xdC71FmOR8gn
dyeRduVW64OkuKjntiyVuSnUtu2j5vggvXND+sPFYDHz/6qYvAK7XRSYbutPAzwLtOWdSCQWLjay
KQgPTcO3W9IOJwGFt4EJInDCEy8sNOE+QkW6JEeilu1AxzB398608EkUtrB6ILkPmjng4niocE2A
IAq7CvmUDSc9mAu9k92vK2ltvMI5Nl9fVR10AvTAagl1+7d2Btkog7E0tNYd7yPvbN2g65pD3PWf
V6f18k7grCZdzriMstBrJtIRhkhCTa/R4YuzC6JZ2FPfYf9TXhq9tB3qjpE7jghflYfcV9/V7lmu
CZwwSji2B0Q1jAEAIVUMPRH1h+58Wu5DFlEixx5uTnZt4T4+PKcdTMnq9Ydx1P6ea5NQbmlXfAqW
0ophEQDNyT5VWxu7mPoFJZNJ/iWPK5jtRBMMG2UmqfHO98V7xIcu9xyWXRebtE2SRwMXjwDnc03G
88SU5xRnncmqAFZUrA+fTcKwy6MGVNwjDSVB0vdrOOHnmu9IULvxpTz2W6OKdp1GwpXqbG5NTvy0
c6BKI6wvkWMeWDc8lRQO3iLNdZR/oWDmOvb1B3AKeHSA56abkhRxk9RzAA6GVt1Vtvp/QRkRKowy
ehDsJawM8pHim3/s6GVHL0DuoSepYGBAwMdvW7qVaKSD1MfPrFGjsLGIA/NUOpGNGMro21tKyyfw
priPMb0SHfXdcysGav4eQY7x7W2KymPk3IT4VGdxgmjp/UW9tjbR81zvBP7nknT9aC+GEfz5YLm1
CfGV6pMineK+Y9aFcy6Lv70/2yg0GAwJ1NvbF6P6SxKE3CpK7RXuIzCkZXmS9bh0X79OiEeUaOYf
nY+2nhI1OW2MzEqN2d5WFVKuvF9fa1nbdWxsk+ThaV1orujyzR9QFBy0pntl5xNe8HJdnEhjp13V
n3EpwVdF1YujqOsopMvcP6cT0BJgqWUGU9CwdlQy0wCeSqKJlgIsSNGOmulsoNY7igbfSKUg6JQZ
2XIpgWw38ZmCZcRZr/aq5BVRnqPTugva/Y2xhbaG6y2ER5kIPVRBsWCh+QFBv0IOhmGlZOQGp8S/
ii8GY/faQv0D8fUZtVTt/dQFqY4Ct00WuWqUvswaC8bwFmNT7LxsXt6o/BwO6Ozfz167P86amRax
vb4Bo0F550oNeY7b1X5EN5piGTP+gjmchJFiFW4sl7sf/1kAr6vuoSgWaZmPYiT4MBRwI0kov+ZE
d3mDgeqYQmIyfpIb8GkKUCuMFXNZ3LxkfBe4DcKKKU456ZyDOUAnVt4yqpn7aGpk9FfGIPWdiy21
c9EQXeLMRZT5lnGrSKijcWf18OdZWzM0VrpmenvAMKJgaKERksTHkt1PHXoom8F4my2BmWcKwMwF
SMlU8zCLLo7Du0O85hS27HMgKfkXjNzTaUFqJsOs30hnQ/Z7sTMWQAaDD8ZtcmY/Nb05ks9gTPCt
uDIMP4OrpTHlwB3Sz8dgG52b8YP+GUOSDw/dP5UmfRp7A2K2uJSUy/YfLaBKFnSHHAYYdTLZ9Gcv
+7Qve3YxD0C2MJva4gGePtxrk3j504gB77iiGR3QGp3dFTTsctNKW4/+NF9jwgEw5V0Ev9XkWyOR
DIeUV9y8652OFHjs4EuD6jfA3jW4U4UrlvWQyAg9Yg5bbesWzkDTdUNABibHaxz8Sv4TsgYtLwPN
8xS5acrjUWG4bTibPBmJzjHGRJm6WJrjIEeFKDZ7spL3RrymmD8ZwsNVYpkhtvssijbTEYsE9Ge7
OzaKGhrrDQDHauL1+/r9lcQfKt+IvHgcJP+5UJCXIm5pJQaVKYZbeELU2GcE/2YSb08t7IcpghIP
2Q+PEZxmeBL3kVHMKCo0Juhv8Q4h9z6TUKv8Ox9n13cCvERxG1PdsM7/LqqACvAxvM3CpruSJTs5
LCSVOASucSQBxPz7B2nRYe+LOWZB189FPVivj89kuscc9u2ovjMIZKs+5Mj8QAzDSaGx82QWK3dg
5Or143h7XNSLZ9Mj1AiFlowIaeGihBxXRE2TF/b35Vh3vR+AKclaS5+sQ+kL36z3WbKVuJPVIMj9
e3j1aCZzJc14DEfNKltLs0cZUfT/P7YK/5pkehRNUeKJscAUyN1BfFUv0KnZIXdi9xy7dMurqwFq
lciwjibAym7cNAC75WmPXFBy3c9aYQEU8BHqhhtjZJX8bh7B/BaQBWNSat/5M83MZW2ShAOKUktX
cDeqGjr8T27r3gVuRdhdyi2I7o9TW+4M3g0a+qsc57ekvUwAd/kFdlI4ZqIoXchrL7hBHj6zMOXv
0XiMXu1KnNsxn3QN6gjgZT5jQZUZwvMO+n1I3kv4M62DeOjS2NtKetDyzOh87qA2PhdqEaoGfCkX
rEii0ufxARzne7Gp8jqMGnk9M1Vu3fnHga1sVrkpO7TyG6bgqYV6SXz3xd2PCZ0sj1wrnGtTRmQG
4msMmtxEOZOAzNOZezvPNk1BI7z/D46211/wg2Xlhfhm8KpQgq6V7TAH8A6sq749LcwQDyli4sjH
vhmNS+8bATlnrseO82iUU37Hnvbj537/xnxJkWe4OLm/Zd/QpqbnTFcUpTJRKF859irNtHFAHUx/
b+Rfp36K+vvxAUxlz50Cduq/xeYmlCYjoCLjElg9tHMxpAvhX1WamflASxNeGz90ifoz+b5ju5q0
Z69fg+TQVhTYKqnaN38ArrdBkM1L6iGb0KASIyF9zJhJGLIEDkREhD7vQXzr6Qmq/fLoQ0ZPIYCY
0b3DeP9CEYLLfLNJXdjMDpQKAZ347i4OUzqlXNnR8/LfV8g83rSsVnHh1mBQnZGOA1ky4xi21Si8
/AUEsqjA5lpyftJNNx/mhwFaNUkM8yluR0aTdsSiwK2NZKkFuE3sJxnLL8AsqyjGUS8rV9niU/g1
QgjqjBvoubbcKN/49hw8vCFnSUVmp83wEtSOzz1OTJezzafWl7OZDSjmK7181tjjiDnwL2x53S/m
gXlVAUpURVbnp4Io+s/opu5ps/sBkVRxJXdqOoirPnluyXeuoHhgphV3+HpM5Lzcvz2oeBjWZmDg
D4g/wYlETecWnT7tr6Ysq2so+WSs26Xslx8vZ96p/5y1FuRrL8Jx8KbhVmBcU84/b6dp70iw5rmi
gap0lUQMbjIF7bLs8ZfgVBPJTfwgoqctqAYHcac+6IyoLO0oG9U51ZIb6cBKhbyEnGS42YW3GRRL
yATsWq5gLuLf6O+7ITcVo+lgOSXRb1EKH1UARPPMUuB0bymQtVQIUplrp5GXcYqv+BmenvEZj7a1
GmjWTwuV/CtROPnrUHeYFJn5QQkivGxx726CGDgwIxFO9Y3YgB1hEAU2JzSK8FiJ6VsSKYTmheDz
ZiIcYWT5A7SnbD8AeGp63w/OoSOvd01rmBvywBtRtd4BPe7pOPDblwcOKJ89tBXjvSKb1j0Jin5F
rTX6Yeeif9jgdDzETUE+iImBPFGAeFyMG6uQFYduhDHKp+MA6MjngN8sUTfLrCFaONmLkQOHDsRe
RDWdhX3roSGTmTOIuu4taa2Ae3A62XkvZw46z5nmfkdTx/KYdam4IhJnlHSaIgfUZrtSlB9Bvm6I
ey9BB12/I+qe5XJ04Hs5TSTceXqDf9PbzEOFTq0OO+XmqbJ88h9W/rGYf81TZraWnkQxF/OWNtsT
DsaFeBxoOMepkxJZgitYapycBBGtYU2h4HlB8UW3z3SBqjmiNgqnpascGSJ++wYQADcvu5OzaaxW
1XT1efj3WXCA0FCzXf3mvLyQzcKsdq8vQzlaBmLxA/Ik7z3/L5kB/Ww1sbo6iIAPqT1Ifv0k2Qz9
41VqNkLPL20U3/SLlQUEUlXZLmxM1KXB8fFvbwzYxyTdWJMszZQLW+5Knr6OgopmqPc3e1e+VbOz
gGf5Vi7wGlCso0k4LSgXeLsZGVcJLbO/J01JyK9wQ6X1wVpdPPDnfKCHfVfWzcgcYECNL+gWZBtm
2bOtiHDmDX6ilc1+US5Tnnt/n7PdIh6pvVatbztj2NbFcKh8OWffHxD4L0G3sFR60CzxhBvtGemU
P/5+IKsZScL9OKpGZF2ExJU+/CJEbd0KmAXgM8UD+hemxAaOOzoEAg5J8Phv2cCcGoZK84GU84LS
NoBJCU0uOdAuerZjpwBMwjYOHLblq8d8XUgBjA9rLJ7Rzofy/+r/zmoB/EtBgHg3BWnQgiVyTMWb
o+5M+TQKvnf0wUPk7vTMdPokcB/h+zGuudTA3nWMMwRu5mxjANLGzVH8nXffOoYt3fh7UsmQllr4
zQq3prpWxNq6YC0R1mQAa6Q6JW6HBUa/KJfu6fxSHmyIcHoUEuY3jZTGXmqKJUvhdrDGCODIlkut
HhjkVLI0/Jf3rHFXgEWvItpNqilLvazUDE16w76SBRJKNWuyhDwBPB139SNutOHWurgqLvnAicjX
ZCqudilZ38AuWAFuc6Nt4fAxNM25upxzFxPQcH8PYs76WQgHjfXAHegetE5QDco/zaSPomsQMr8N
ZGbayYO6z0ZeZgF/5mFeskojT8c4PMa6qKqcTWB1oBmWJiwnYUtZvofaq2ni2+m0FgrcKTqNCImd
hLVzMYCcOeNdrsV9Z+owcQQTRTYQdpxjrRv6SEghpSPam8A2B6AShllGverzM4LlJIbq/LvWaL8p
OtpNia7YSOnRRE0fYVHklGjbw832KXEvMHeCiueSJqBEyB5dYkCQPYV8xhVIg/AW9oTX/xZwUrrF
8crnZt4ic7cr5C5EbSgzDljJ3mX3o6FMIcRKxKa4DFpFAUsKoKOSYSlXCzE8mG87PJwr87tym+Fm
2fSlKmHkNzK73ODYB2WXvRdU+70NpUjOIBSuSPc+MO+FjqiFV6rlmsl/FmAFknogWEs5kXPzR4jx
Cc/Tfs+XtzL5zvvlWfsowgX1mBi4+23iJGkXEHH43CKp/hqWhnqKyqlk0BbSWNdVDaP4gC1ISw9M
WBHRNUTRkuTuR1yD7Kf2GL+Bjdvg9YYkMAt6oP68hFwkckWf1NGgRB7OpGwggPTO1Oy3TxJmZACY
gmj2q8BXWYsOuP82xbsE4/+Dk/dz+xXVI9u1JlylcW7GRTZAiGapt/geAPnu2brZyLzQCDxPcSQy
Jn1/p7H56RU593JZpvJlqQ2/wH5Gaoy+loRafoAjd1lYlEAVXk1KeYZyMDznjf3JGTkUZBbEE+zk
iabfWUiWry+UkqnpWfywPrdfPcEpWbS5q9yAg8RwR8IrozKCvmz+QPbx7mdb78VAx7X5SzmU1HO2
WPh9aQ3ny1I7Tr6zVxKuAruuxvRWOtfb9BoA6DJ7Bihbc1kvbb+UD2nQ37jToEA0lrg0tXe8b06F
9ZHcdB0NuoXSZYPnMQEShI0KDDAvKbe/hkpdAawZjmvq2ECTyftyyG1POyy7QRg3hlWY9/gA66M2
YQnCOydr8Zy2FJ1bDOrkeCOFq71Qx3pDeppaeMD09+8f09OGwTvFDOrMr4O+9rcPS2fM2DRL5ljI
ptIpOTfqKW5SinUiBtAduScaCyCu/s3uMspJFsdoRn5tzkcbq6N4965Av2b/t0jjcwZYqjil5/bp
OvixeQ22wW0TH5BgR0gct/GPINzALg1x2Ty2W39Q7iLDRLQIhWYM+FwcvgcVT3J9/M7EUDVoHdUw
6ABpiGiKYfvoEX1xzFDtbhwhtybNU/w5Nr7FVADrUJapWR/y5e9BlsKcONIJ8U53SNsjCvh1mx5V
iUYB9i0Jrkc0uT5kIaJxVvdOyCssSDSd2m4IaQEwAtAruKhmcVA0i7W3eocww+7wIaHqVz4liIyE
ctB5i8XoYoUdi54T5eLqPkZ8Tpex4xhMclbyro5dPb3key4V5y5bCHefhcJs2LOHjl6/JtwsBR9C
5HEGMyOj55m6r2ZBnJv9K66bhWHhA3qJzApagHPfyBmbOtICRATYBO83TpCW4XPc0J1Dw1r7lWfz
bZtHbBfN1YD26kqOyl8RQWXEYXKdfKacZ2yLWi5we6CO6YHrZKqYs8H6k0pfWu3M6dmT3dHi+ER6
LMe5Vp+wgAHMNt/H3hcGOPIbUkq+bo9/IDVu9kjSsj7aWYKw9/X1mvmyG3hRfyTkyON+OYO9walq
FEQn5+OF+eXeRt5fGPKmSPbn3co5TL7ZVg9VxICyNnDk/jDCHkBvGvE7X3PPXUSwVcpm+oIDRyUs
IaOoXidJejWeyqPg2CbWzBYnHI3lGnI+dIbNQJ9NMG5gxEtGCWxQ+KkCCukVaYdNlV1dzoNAomU9
e1ebhSERCTDdktDTH3MDPGiemA6bPNwZrA9bme3eMuIf9xRed5MrEUbP2Wx0zVqnnM6Butb9THtF
Hnb/zZFdJP8I8JseOo+4A9K5+7djogrjKNgAWGoUhsaGGVPxBKhA2IeAjo4WXkE8QmuCAKACRMI7
ffVHvwsMHkIYRb+BrzoiWorOaprhNalizyiu7vuEavbxfSWgu1u/Sf1rfMOx66Bj7Iq921Sgawdd
rZD6I4lPFhAoP0gePxnMVY0293CNTAGDuDVHvHTL4TlbAVzYqSb9CQ4XXY456OzbmZbo7xxVCell
Ayu84TUzKxClcLiLeIgkmf8la4Tjs4bvkO463CCHnQcWzA1tB9Sz2qmT7UHcUspLK238mUAZMAm6
9tLC5ckwMB/UotqoFs5mwYkqS62rz3Zsuty1EyWbHwP7MiASHTpkC4NhRujuMcMHK/OiWOCC46yZ
iMbLbpz523+7YWMMeva6b3cGOOzh60CwcG7hyCfq5HNk+vQ03iNm8TuDZ2X/ya8nU8EfvvIsjNYw
pwxrcpGWo4/2Y6rV4/mcVxHRCDB4Ogw3KKJ+n/UwQhkBnN2iJiL5KLamCOXnjla4jyjmf/YMvjeG
KKCLQKIaGxjvss+saf481K2NOEM/8w6A32XU0TEzYTqMXRQik2GaAEqRsNKX3BEykVDZybSOejLX
HhduoKyVpMLpQxKRzvtN64fNizocrPePbdKmsyCNyQpx/DILBKiV6dDxfu8NpfQC9xiVAc1zlmBl
tGgAIwmUzWTlbKgNqAP0eiq1mlSdj2Pto0Mfnto/m+UZSrAYmshCoAgE1qAzvcKsgyl+k7LQysxl
B4XnGsn+JZH3qp3U0F7FmjRaJF8AAGBO8n1bQ9c+jySOobg0ekxFLVE5xonEoF7jt6HaO58HGxBH
oc19SEukepBNIssdq/kuTjRhWTvTe2zlu9hQDwYk/aSIcxd/nX/jBNCq1BTKnJJ8hgDVHqEpBNqC
Zefn40Wud4zUZoKCbLep47ImwPP+7tMG6w/L8Q/d/t1SbUG1Uykz+nPnj6uW3FI3tyUzU1FOyN/1
Gy6n34HdnL4zRJjeK07kZulex6nB+XtGlOA9FB3+yCET39iGi6+pyudmDxjJq6jzaa3Y7atDSg2/
GA8KX+uFhu78YPNU0WMcA6/Zx1obEC3DuaD0NTFYxrRfERJ7B6PxaxC6mzYzzjbjSjTpZtqo8TJv
OOJI3NDFRECb29aUov/Ym9q29dUnwFrbS5ZI1LTrqgzEW5A39F3pu+ofpYh1EfvQoRdk/BhfH0/s
S3tVi9Ei3Ww7pgAiG/e7XoTuaqOFXuOuJapITXPWNn7Y1mxypzx3KsWlD2BpZeUeSPgsA+/PrGxl
aOwu8S9k4SfPc/wwRjWwxqNuaJ9/78E29pxeqrgzHoEz0v4YUllC4/IJTQfsTu0bJxmFuz56oUxQ
Vz3d1rsKPXMKH6KiKmSlR3Omu2DBKdkVDBUn/Msd1/ZL9MXawHCCgcSxywzriIficegPjK4SFvd4
1W6GvzY1Fj2E9Dxk9CJMTKLVLv062FYp9MO/ej80wDbd9oETbBrrY/Cw50MuqaEpR0FuKT4rv5x4
qWN0OBFGMLFGd3XHWbEx62LUOaZ1hY/8x3Xo9oYDCXG95uTO+SJBsBVGUmCYunijAUFIBaUPcm+o
AhYN36N3diKouvU1Avc4Nds0el7gehIkKdLIcVGL5ML1EDbIpgVx5C2QavCyPLNROJY/Mu5HY9Cs
AKPxna09OFLVkzEQxm/IdODedWi/n6Po49AD5vO8UZ/1F6DAX4tDiyChG8EkKjb0kdcID1//aw5V
PDCCSQCqjldESrZMj38Z2ay0pxXAZmERWK7fgLbxsXdhguYFWuEy3S9AMGQN4lmkUcdp07SRU+Mc
hTgbIlub42v2nL1Ql4zVvG7fTbEaaeVue5rtv252hVVTUx5VCNFne06odlD85mlJcxcnaUTtIZcJ
hqVpsA2crHqKCPIsCXKWQT/T3x55PdsdenwKjNspmUvPiRicqJnng99/ZjU6EF3v0g79sgmO/Ajr
G33ipD2Q9QMi3iOWjEOglVJB6FM5jdwXApQ3GeeUGth/pTIbdrS2VWQQCOTSOsq4VejkKxQNxvVf
Y8HwD0stJJ0wSj4YEINQX3g/RHn7u+7mm1b6ASO/fleSmFI7E+Nou0oMi+ZkukKagLsbLNJv/C42
FQGLCOF3fGG2yLLddomzDw0opUme+71lwn+KKR96KulxnLAH8OC/c4M/vtGzybci/RZpsC9VjTwx
ljOXRWzYQjExfJtCs0M5FLnCN8aOKZLEMoHpZENC4UypLAGOoKtupp+mucm9DzAR8tAKDNLIV5yt
1OTDyzJlcJpjKLE03T+vBBUr3G5cEE5ZXCIBGufjRhIUqmiWmanpa17nrGbx/NeufSuxCv0nL9ai
aAIW1jNJG8/ogezVTrHeLcLXXOA2ggxdGp6edadG++STH3ukUBJsvpCCiGy3AJDH+Bmf55405UeW
ATM/x8jDZpLy0SxBa2cdswkIB93vbQ+MoiE2LfDV6g7yRXrILZUz2pS6rBH/APlkkIECjhOW4C9M
gRFx8ZyBbQbV/z4/OQbe7a3FRz8JWFnKetxRrIb17PDvEYc/6H21xeubWNwZyMjIk0bJoIGVP2G2
n2kjkvc+HgUyu1k1D6vuBZ9zAEbDff+fFOyVjuVm5uipO8gEm3jGtS8jjGcr5v2c2GflNPUhHZoW
DGihsccchxFwDTm1z6emNfBnbViOG2Lq48g55n8RZRTOa4jcUzVESSIwZg3nf0Cz6U6mK7luNcvY
ctyL9tMq0XPe76N3rQyYjLC7Fb23/734O6dnTjIwGfVD0dHMYNuH7FD5qhHJq7ygz4SfahOmQXVR
ZAOtLQxnfYrA1GP0eqkW46xWCRen+9WmGXRA3RCW4b2KQhpFATFOe5tdrFAG4JeOR+erAk8Jfayv
LKYJFYh/eAFKW6JrTL31JOkjpNd3DfJ4OhccCwtjE5ODJQ8/Yn08qx37abgQGN9ZXpLKSFioDxJA
kzNM716/D/rBst+eWq+9anEny5YpSYl0oNrgDBMf9JcG/KdA4zVdqjlPYNMfx/DoZjJp2UYswg+O
iQj6eX7D9UbNpy2RDaTO8g621s31ykaTtC57UvTscAvCb9mY7MJgbCpAsg6LUli7KER1eN96oUkE
f8aKz9KIW/KYH6pZZxJicj/wzHlMjFDpZiATaC5K7E7ibvIMIKb5PMIT/PtPBWXnZhSOAY5BH5gp
/0zUu5mRaqoSTLxlUNHSGb7lqAks/crKjCS2BvZXnabXiF0IWQw4z2vp/pRKwgk2aYQbeAK8qU+d
FwEws8o5TgaJlARHXrOgnv3UoUfgMmG07lky4ETqT/JF5n4gmXjEfNErKnVzdLWGYmFGDZmeZavU
AI8WWg5xh/SgEoIHMG1zw54Kxfi47X/xG8S2aONyAKjkbYJf73OLyK9UQ5LS/erIMYu652rs+cFR
NQE2zE75Ix+r4m5iskCA286qP7yzrZNu3DOZ+1XbGqAbzrwPrq0gEws0jH8a5F/0CBYa+GnNGSXq
4Km83MoASEoysxq5y22MK5gZz1UyvUHGJWPwL08czdRc2Ko5QFgu9VXZi5AVin6tO2aYG4XV1c1P
0/82t+VpKMdp2e3oPCnXMjLcCj+jjKXM8lCVYImml2NvNvTxC2kSFnukxzdqJd3zdgHiewhPtzDJ
UCrjb5yulzm5e8/zNmW+i2S5Uy+7TjgsXXN7d9j0lH/UNrqwFDCOztUrCTFedVf6o1j2pVxH5IUJ
wimcOtpc6engRE8HY3ZrBoQzHQZiEqPworivRlRdsZxQ6TF910np6pJCzpyDd2lqeKYxFmimHZQU
7BVxnMZdvNsPsfz/tG2py1kYQe4xRb6IDybYFSpoVrzzeq3P1NmJbLTs4LoZcg0Ckr2MUITyt3tt
OHr4ZvOLF4wEsvWXK34x9eZMjJsbsUz3ag238GnYTpWk747NEsYZvl3T9DiKi30Lb6xWtvjY3pnN
Kejyuz8YILcpi9E9IYwCoqVbQ4QvvU1OttBA3MlSVpUX0Wbv5kPfNrIMwITlgFwHU5EIXCmGakCn
7RxVIbjuN1RnVk3SYBwaJSk1Ur8JGAGhsewxa2qrIXEc8pbS08jbyI6zfpA0+N0YcH8b07m0qEEj
hqWEO6341di2KtsJxgJ6d2dw2Bt/NrVwThbsNXZph/gBQ8+4tOPvv3s93ZlqO7V2VvjZ1ZLqL/3F
QIGlnKaI86WnozAnUV+qIVCxVdgPKHf7U+207QkCY9KdFLCuYSj+8DQNjLUEsbYwXA8l08JzAgT+
2JC7xSxGYgJNxwfZ5U5yR5Mdb8UWyl56LjGyWyVq2tsogiN4kNFsOuWdMuw9CA19yApRAQXJejcW
5WGkONtl6j+Iqz9w9xp18xU6Ru+Tji0nUfDOZcVJ/PqoUpTmiR6i1QBbrqL/Govz6L4uSYNSz7a+
iu1dZleaJOTnoxb1VWtf63SeWYF9MWC6FBFt5LMCgQQ2CVMa6oLZKvUe87QXk3lkrlLpRYn+PqNh
J+ZQitaqkGZBKL9xmKShGja1YegVj9rcB0dquXpm4aLcu1HY9PKBpv4NfcZrlSlH0x6ZXnIzucPi
osSaQzvZPECVL94RN9wExZ5nsr30GoPp1EJsDHnpP7eB/TmPQ5/2gOKDXvPUs5Wi5sinYHdPP7zC
tmEZsKe5C3K2/Z4mmb6L+xyww/7vxTVhrPcuFr7AcOQPFeSgmL8uSU2nhFp+7dbOGUshw90TzTFJ
5Ira2G3TOli9veSFwgjouRV5x1lAcIw2ui+B8DoRYQJcueFD5pZRNkaNVETc1fmu+a/AKioi98DH
DCaR8EgOLBQEnshbywBLj8yLNs90kdAxBJFUVDiVoLyg1C5uzEd51LSfN046mfbE0V/5t//PnVRL
8OrW8VsGG7kJXdxuKSKxWdIqfXk57AqXHMPgBHKjmjryN4lC86yGovQMuDBvFb/53V3CLjRxvbaV
KkwvERiJB5tQ/sf8+f0/eGhjgGIniXIA4y1sUb91AGOP5Lu7hmj8MO1XLf/msahQPRUG25fjmW4U
jzEEA9DKcahmdqS238w8D5LXr6ZWpTYgU/akv+SVGHGWqjZU1eh/pDgyVuzNNMNlLT02+9fUeii7
R81suh+OCsCKmRbOb8sN847DrIImmpSnZR1KKAahKTJYvjX+zdEFdWWUh1K9OrL5RJP7LSBGuqkp
ziK1r/ldxU7TgFdfY/jAvknhGZKbv4FSmvOOWbruG9JWOI/x/n4JJK1msCPJkNzaQQ00wlO6NMFg
FmprBQ78fkrhRJ4Lgbptg1Y+3UU6n8WSC5MmW8btzC6QuSepMLUeuYsr+RpXqtWielXWWF4Ehg5P
YewjLXgzwDKUjiDCvSIJbSINIqaYwuS2DFIMbTyUGPN1jFOERhuOQ6EpgCQFcPcZolUTJkTG6F3s
I4TkyNYT85tDDF/eUE135HVGwvYCgqmpoLfM95zPcgc/kOmUADxAd/Vfoq2yePRpxjgidJ0hqvmP
+zmfOtn8Y1GYbnKnspOaFKpMgUdbPByfvYLv4bkZlcvBN5Fh49Qt53sTyI9WoY84SvMyN/OKag0J
0/leUb8rQ0klpDL4IRHzDP8h5OugkTOOdcxsnIbfNSedDKcdXE0m/rCYbBLPrOVzTdG8ZKG9RCDd
bwGoIUSW+HNB856FjiZ+RgxOLlMYjJBUWGXZQp5wNK+aYgKcl75PB4PrYL1jDRt6H+MSQkLHad7S
XDk1pejxujnHKldDasCPeuuZf+TCC1wq776EJkbw0Mg0NLmPeh9cuXYUTRS0XyNgzhf+NiGciT7K
vEAyrcvtx4DgFoXkACyrEjT2DySw7dfAkfewyvVtlkZ+XUMg13WEMAOpII+74rLuoIxxAn2I29J6
lyqEXJCuhXbpTiDcE4rfYjAT7+bzyNobQyZIlEsNLfuuJHImOM+9KyRgEzNS4H0SxPI0KdkvW3Jw
GbUU4qXBhLujqPaO/S0PfTJ8TYSihwMWjh6DlccVO+B7mkJCH3pjttWUayBCH+QgMtpJOk603Hue
dcTb3TD6Q8gsqHvppfHeNXh59sEpzg0mWNsfVRT+z6YDo8uWgQkT4zVUOkss9vtHfN30DtErmyix
29m+NhAS3PV1aqKYACVCzTiDxFz2Hv+tTv/7QcvZq8cpaN6iBMJIUvdajAW2E/BW9pflnJMQSRfU
f72zNp04NGYtboG569l7rDi4extI7eNt+ZJ2Hqu0O2e6sPLzlNd/ROqb4H8VAnQI1ca+1uRAzTWO
mpcQOw9k9UVmkKMj24O5xFRn1lNciAvGYWFJuo2NexjT+RIjchix7ZjjPhY2eEuimOmpynFLg1l4
n6vVIN7r3Rwy+PrsSMu/+UgtnsZZWBEUOogusD2VWvGzu9hMnMb1R1wxA9Q5i1dbQAqryTyKM0Dh
A97BkpwvgwGlKEFymft69FrbnGJe2V3Fo2L503y0+suA935TRXE9o6F3qOZeQwu+iheffcpkKOuu
gvrACiqtUiFYuhLR9r2HZxfBxH3F1uYF7e6uIjtFypmldt0jv09cD80DstVz0lwsl222iKSBc6Lc
vAKa12R1aPHN2t1zfsqXGnGaLuxV6SNIYOZ0xJtJ1YyzOY0kPGkouq3fKnbG4c6RHqXhogw+u+Gb
PPoeS+r1pqPCj9mp4vc9HfF20+3ppSEMwzTk5urZqWwRONuk/Q60V7SeytFThzavVeU41aec89ai
Lkd23IvQAkQdsiTKlskRmCtrst1DKyPqTWSj+6KQbtVTLvZYoANVAVnD5AO6OBy1SCZ0IXIWAwic
KZqPsGnuuqAFtiv2/bxQJcoRdF4Qyh0WfqgAC8MjOa8IHYlFQSkYneAZrhmFW+pdRfSDBYGrm6z9
6FuSpWCJLIfyD+AwXpn2K0TkWeCSPvoelkLmEECVA8i2waZsa08kXMWM0ED8F2Z3Wk5S4RJoojgY
J95L3QpfXy96YxGkGQQvigRczoV8WxEpzkJGJM3g6+zdeTdh+2iJF7ELMPgeQD7R3uh2Dm3yU/a1
NcSkDnUIe6pUbsn9D0ioudWMTuw84Af/xJtHTjhtqbA27TCW62E2idnXYMd3pHGsUDl4nMXRlCyB
36zsUVdwq6BGMy+CphHsbjRn9Ouh41b9A15mSQhUl/WFbx5H1wuNnKBBPJNgfgj+mSbh+WjJdlkD
8boo9c9UG9+emTyK1USaDQn7TYa/xUIn+X33GH9vpkU/d3cmsD2Dt7+bcwpSknLCxFXibTXu8coG
PCBt40ZgZetVtGOcBTFIugm2Kgs60CARwAKg493NruLOT4ze5KhBwMCPSs5SyivilLRYxutwj8gu
tpuOyblgOwrs8UoV8AQL/wuuK9Yr/d3gyDL9eFjKLVDYwv0X4rJCAqwrVVuL3ghVY2EOgZ1cw4km
zjMsL0I0OSsSUnPR0QJ/qelpL3qrgcfdaLjQqRjh4m1919hlygoc6/+uQtEIjR2Y0XeZAnQxQnCk
hLLOILdlEOX0ZCVqv0j0I+baYetszrfd7+ufj/OZbjp5A6Hs+4XlIHkwFhQmIxvNcKygsApSbyKg
VRRxbqouwdGPBIoNQ43Ev9KtyXibxmZ7yYMM1rYc9NzbYeDBIDzRO1vyWLa+WyFJnnf4JVeCS6Sc
aEFGWU8ETpBMukjslmwYbkeb/TUdHssueuQRi45w2Eu/FeNJlv26RmJAqdaRlMkaDYBk++fCW2Dc
iRGY2+bWJfNC3GHvrE8hUjdh7HrAH9rR1V/Ps0tBkRQ7olDPv2gz8qmRQ4aDu0OqPuLA25OxPmN2
ULA8jjC09PtfBey9fdn3xFaq9NKvG6rHzBNlXVhDyGlJD2GoQRx91MXrBgJr0frw0J2SqH59dsNq
wFRuMj0opRZ4bjxKNfng5bG0JkHEWrkgtFKtt2lPhgxEeQ9JpxjMRoKoMIgOOl+/Qyy+7ULbyIK3
/m+GoF4cKmXoYV5isJTy2k7HKOicpoP9OTfK9DWta7ZsCq7RWho+XFOLeP2XjcsFQ9quAqmt1UPd
CUSP4U/DIFchB+M/ZXXWO8YB+NPZOfiaTJr9+Df/hAWtK7FECeVPrWLRONOrqZO6wlooGfjIo6fz
EivjhP9IaVncEXRCr/T1dqKKXQmmQlnm65l0P/eIq8hQcqHfB89ZEWa0khhqdYQukXe7pcO9E23e
qm7IKOdigLgIupg5FCtwRkmv+xS5x3JnlbOi5S3p67PUz3Yj3G2p5Kdk4npUxyLUMwfN39x3T/im
RDjA4uF2T4yoGzWr3fiQWTgD3YLTqy9J07Oj+XWjEzU6gvlmxWn18NGuGm9CQUs2Nw1VWMe0311l
qGAJmMsMP9O5dEP19JjWfen0a9VfBYclOoyhpcxp49CPMNl0nxELdPnL3p7eJqx/mjQHkXL82qjS
KsS/UX8w/PyrPpZoXBoLirQfmvRDGyiUdyttlwtUXydC8X+yMMrXSr4X+2ofdI/0T2PpvbGwfl6E
Dmw+cdEC+24McNyYra0jQL2FKanA0XQOU1mlh9ggFzHRJDiKeNn+tLONUW1L9d5FI8Cup82hbGOE
/znz+56uYeM01HUG1A01bu6rDV+p2z1L1AJROXeaq3nG03L+abPr6JtiaUwXXHPWM18ju6LiZijy
L4vNbPFlCFyKd/uBxqsRi2MyDpMU9zhvU5nYEFd+SxfOs2gTPY9h+h9haa9QZsyG3unFQgYAYOvS
YAh3FQbLLBxHoiIdcUbRM5dtW6ONqTCXEHUIvu6gNl8zVsuOgrTKdIhpO0d1hp1hc+3gCfoPStg4
1SW8xQpe6Fcs5NhZphevybDgYaBQ8yUKZatu7bmySKkNGNyHvfav0DlucAAIkCeU4rZx5wUWbmmh
41p618Y2BPjS5M8J6ZMlnMWqGRJkpTHuP6MWCclVYflgDnVJfq9X6BppEPrFgEr8FKq9mDVBriMD
t00mCNAp26plr3nk5uxlUvUcJMIpiM9gk7nzzoZL0x9Tgz2w5I8BAtdfQ+TSfds0f7d8/6htwM2y
19L04uoLlJTaPbgZ/BJl4lanGSLRej7A9vFuGKbWjUWu5EF9Ss/iayBCuraq26R4abA+mj1zV9/7
0PRG4rV0T2q6DiEb9FL/TBE5TDs3UAcnJXU6K9c9zkN1grP6JB3I4ryQ5CmtvB3ODeMquibPv63F
NlONHBBBRbc01jijdrW+F3cYOQDZvTsZu7lgLEWkjAAPL/OqwGl+su7kkUR8qod9lgzLdTa0ckfV
Qh2byBLse6GKcFTmDqiMHrrUItMormAMqbaPKJjIbtI5EOEVFKnuotTTU/aYFCzqEpk7+X8jlq46
i7YF7TAZuicHNd2FH7qRjb5/FJmLRXSG01O7M2dUQAFpbeGE5yTrgZDZ8eXPOlC3aoU+Mh9A9CUq
nFHWocZY2E2XBXyk4aBX5RlgTpZFUkPPHUFTd348NIeyoyVAUhhzj+4MOBLZ2PdkOJ54Lad2Eped
+q3qsJUch6VxVwzLzb/bjaDu4abQGWtOCDlLBe1BIdqVeM5hj9tlr1S20g8lcgNKQhVZhj9/bbMy
jAELg5GIjFL4tsmEQpLmcals2a0x13n/Er2lvJU3uonNFmL9BmoQqyA7SoxhiMArIuUDkBiDbdcx
8t2F2L9tNNdfGT1nrrrNp1Tq9Tw8h3lYjTdflZa7hAizoG0BZKpXhtrGqAoOq9chTispfOK2Fc95
Fhv7FIXEJeBH86Kub3SPqaUIbD8c/9G2VjI4vLsN0ZPsB8d16teRYUhpgAJ4A0S2v9m0b29tjzvN
DYbG4OmyYeKfhVCquBKbhne5cyi7mh8bYAD06e5q9wla2afshBb9JhVQrOqHbRjWWYc2J1DCRxNp
jzCSctRmjbZ5XKDUW0BAaVe0uzI8ecxZv496SEAzX0HI3EPojEAd/hpgPV8EvmFkZHNmStp46rUl
xcm+m2DiplRFYYvQF50I0Nj/Gefar04ELu3nZW8uSh5371XCa1ZqN7VOFpjDqrgm4Ax+t7bcLxGE
JJxFvrlgUp1WWGw2squC91YCGBFC/Vgc3VmtkGYbxbmwpvoLnOG+pOsAoFFI0ZFnos3vyT77/2ZY
BSihbZ5ywXDUquvHgi96cmLtsYuql+85wr3V3pZ/DpxMmEAPLBBgt9wO10V2yEcdqmoAKv+dhMx9
rO22qIOR0yV+jXeLKbSX1BABrOWkkp+GYs7WmWahUOuvn55iHk1q7Hl3c5HP8x/V2JwKaTVx7AVM
ccaxXKtO8G4nFxbQPXPSCXcQb4F+C5pWK6NK1Tl+R5CA3HmovccFD3Kwt8pXtSmxbq+Kzka8zqIY
pgi/jH/P2+q7jGZWY7ZCnhzzjdwDl0UABcEO6WyCZ3K3eC6cfVbHRQj7GMr4j6WhlCbtBrUuxWEG
nfSw0QskZqkpbUqlREEefxD+GYKeyL4/6i737jjiIafaF/0PXpmmJvK4tVrAjO0AphRU7T5OaQT5
y2tc19venKuYYK8jhD71slL09rY6mJNHzNkyZWxiKznAYDJNZiUPINsW84kQkkgq3hdIJMIQCx5o
wphTuSVyZknAtekqijIt+CPZl4XABjySdjF7BFslnT1dId3h4sLa/4MlY9tHh4FWVd6HXokYIv3z
+OvspClNHQCzS0TgFUtHMp47Ci6PiEhY1w9PzVsYPm5Ejfh7VJTe+sdyLxUHR5PFqfVXzcHqHGXE
OLVsKaejep3Pri6Oh9Reiw7qRbC8GVeLcFYQ2LRZwnxX7VUO2czTx//g6paoRyXRJG4wx348vAF5
z+7AsqhyH/Wqsn21apnwhfv8DzWlemUta/9Rb9SyX100yVXZph5EEVhu3bVoMuycBngkSAfFHJhs
qa7LYmVCcJ5PUVUQFvGdOxb0AW5MdbNyEMVJu34Vs2rRonUCjpP+t2zxMGfLk00WljDfP5HtvqU+
x5Wi3zqBtzTLpw3/LdjcnNJVZ4HxtRRxdJlZR0pXwql4fI9tlHn11mshPg5WG3CA1we+k4SK6drg
9pXeDvqlYZPTDeUp/F0U8u4N23YXMDSSVS1gGvWuBA+fCbHJ0yiDnXL+0Mnqb1G8JSMqK18F5KCc
PjQAYL7VbB5jVxVEnLqtZlssk6txv9ELZg/3nlwa5Xd2QSaZhYUwPHnMyZI0n5ub/tNE9DkgIfvY
CVzfKsEuAQBc7W5NQOMahGQJPv5m7q7QuSbrKtFfO8j8FUTQYCckhvudun2lD4DiEsmJ3rxdC0QZ
X8XR1HqXKX6WXctTRtFyIXqmbIHPv/ZMAEIIYQYXp1m1wuj2xxmI+jM3koL54f/TPbOrbf9sGuEV
xhxoLLcth9E1owSWmcm6MpgOmLwu0SX5FTVr02ieCG4aRV1r+EWhEblP7/gtj7pnAYFtSv+Yc/Pc
iscKmU9Ip/ahjgkeq4DhwXoK9OQsReP8O4McRxHl3d089/McbxjBGjdr8RZtFhoYXnypUbuska2K
VTFMhf8PpaURsufDySmlfQdI1wRWObnrNGCE6mq0/qnvCdCsZtUCLWodcEDGOZALxGil8BexUwNW
p7QnC4ExrIbZSTkkwe12kNiqNugATJ5uF6nk/HkTYGRe81WTU8qguIMEA9aRgKz4qj0eQSf5UKHJ
SYXXlEsr/0uJt9FYSjhnD9WvKK3qxoTNFSxmD/Nw+NHP0f6fSZnGQIpolO74N1vrDUlrJ0oVuhl1
a+pn0IiQ8Cr7BDGiUmBuVE/HNbPkRsPZFqMFRefzFdQ/Rq0EOyAn6zoADCJFzgiS+uxC88N7EK24
yCiZOL5/ZdA7CLlKrU7O756dqOBcedS1vI7RfvWu8D0RkSN96IGN7mmeYcPlR3e93eRW3/uLj7JA
cYVLR/LRkxNtcEbmsKvIGBgdSisZGOwb4povxmu+nq9L0KwPs686IbC4eVnIYBLmw0OOYLGsUAqy
9kqUyADFQP/6izWbThelv1ndnjP8W7LVpbgySvVtxkPQmUHtRgBbfQlpuo6fbPV+mmF+LbRkHarL
Vlp9cMXiPm4Bfb+zCSu0Ndw79Raw0AvZUEWZMGxE2xJl2mq+BQxi+7BNk1JlWt43rIQ3165sc9MV
GDvxoDu1tMd7eoBfjjrgOMJlxC9MzOmIZvG7vaeghc8WQDWSBVUK4FZ7V1RQkkAeq1nI4O5UwXdC
MN0vGlSqa3JqRz4egA+004t1v+1ClbuAs6SZFX/OEl8lnhjPI2xQzWa+7DCuwhsIOdHnNj9tYXAs
ZESejFutU6WdNvNz6FRcx4RVKy0ENE3fMB3JOdiypU0VDSreK2bRUr8Y6pCQM78aw8jqAqWCc87v
oQW6zIJ98ZQhVBGSWLLwSnds5kNKe7B5Q9aIv2IdRVpec6hkuNen74TpxxkPJF2Ps02Pqq2wF0YL
LgnFytDBAfoAhlTr1dus7vcMErG62cODylEP4amlJzqmyUEvkjmm8pzrMdKL30epAcenTnEw2+un
50A45NOSuJIWPk4lV/k57XggfBfneYEvIx1LIPvnGDZhVg5/IyfUXS87L84kL3Ii6NLHSa/NMsUz
7YImN7fGsCZhk6tAhpcmmGhtkzLCeEqbm02k1lLQNAzCJsdg4oRo2uQVBD+J42y3j19+U38ML3Qc
BN3oZy9FeovyI2/9V9LKFu3NChE0kjpAIuhKdP6HegiqpSRzNNgdfVKtdEst0PlZGmrXXkyDWtY/
uvznyNSc6KgLRdhYeL9ufqxpwe/sqGETSNKNWilWT0qrJAhvctWhxT6mEc0CGsQjdK49icyqbn/t
OZFy4sVCDycU7CeU6Yf0Z2eMGlh3hbqBh2XhfWJ93ORZXVaOI6IQzOW9k56zF7vl1KIKCUJWMvuR
2zpVryAQGMJP6eT9KKlKH3Y51qMxbdzhnEWI66aC1uyyjz60yT5/osVmB+J2+pHi52728QIafMFt
2l9MX0eUOsOsCeVQ/13EsDpJyY8zpbr3172nJK49vwiEobeTNeqkZZR+W9dbg3y7DPnWO77AJXjS
hsCT7lKnjqfL07OaYRSxQugqdi4j0MP+GW/p6GtlGrpo0xIdVP0dE4XyTUPdV62PnGMNarM9GQhV
eKwxompn61VkbCufnJkwhBAu2gg9aRNOrl4ldDQjHaUPYeQbx7R4Byy/hdTcL4ngfJjj7R0ELAwI
91tzFGQ74c2Qh7eZzzoudDj2JlsfeXsG2p6kuQVjne7IwxYlY4aJMDO5sN7wIyL1zq4FDYxgwURD
FkMHSwgf0b3F6qupyL0KWOW+5iT7EFTZFlu4T9JrYgxwg6OBSQS0LO0kQseoGlihhRo1sE/+bDFp
jUNnqFvvmPgnzvDO/FnV6ijb47DVry+g4OWzncGRUg+3mQ7BMy7tCGgOQ1zCPUjheSjRxVjFVWvv
z10stPmfRYPiSGwJCm5mBVkYqBpXJnwzLzwPyHwU+qB40Wy7Uyb46xK8hbKi2ofyDTQrO++k+Xwk
R0O65uk0LHJXgzMycqxWWtDRelpmWSJhgJEByr5XwG2NNunHIm8Z3V9BLZXKZ9WvosKaQG4SRQ9O
+17lLHZcqAYra1Q2YNz9+30VXVIpgRQ4eOMIZ5F9AKsFc6uDP0IZsEtAOg61rp90niV/6dPe7uWD
WtVkLpTBSQH1SBEy8Y08oNOHFgzz434k0lT3xp3sqKc2ludzsJSs4/hmz5dDdUlWs4umJQ8qXMfx
sgMfCZ7WdtwDzaYqC1jiVsTDybGe6JiMRTXyXh9/vUqBHNMcMBFvXt4R8Q5Q2SClu3vSNvyyRo3R
lZ6+FLRrRtjne6DyD/jYqBmtv/Y0yUsrcBSYqygWLx/0P1Mmu+Jtu1KNCxiB3sImVDafPR9EoPjx
uo7I2Q/l/RFcpwcKmoVWvBSrgK7yKPPMBrIKir9gz2JG4KaKU/g3q4RtJn//6p87aqRhaebcouhh
Yy1z5RXtkQcXZt59xqDWaU8Hgj/g5+ybvAlJ9Fb0dtjrtBc17opCwbhExZP+S67TRfVWKgw0HkE/
RUlRmyq9RW694zIAsLcQaAXi2nS5NITNibjoMeWp18icCGEGpdpOuN+TC9VzO3ge66kqzWvbpoNA
B/38JIqBhKCSO2FiQ32GOg93RCU+dgjKshy2Y2NbYHWnivP7tbrYDlHz3zy8sg4eDWtq6UlvpsY0
wr6jQRpwrxItS6Ac6aC7jFwyUWVsWIkMlbHQaF3UtKtvowzvO+7t/vbSTs3jsIylhlQ5anJ9j7ez
rcd84emtrXHRSKF/ctlgNmm2I1Vayui8bw962qgUVkYDbpy1TcOZ7V7K9275z2mAdJXnch1MP8NT
av0Xq3NRyqwY/2NpJO9LEI63uL3CUJ8X2zF8i+Xt8HRGaCeG34+t1OxxWY02RyBNDGvJz2J0jTj9
/Rw1/neweW9ovNsgWzemMQDE+4e3cqr+FDdPf9BDcc9jXmJPPoH46TOAM5YBnN1n0+atpjdDbAgF
uPvbMuJXidJeVQbRbUVV4mCENY2zjhvOyxWFNYmN+zRz82Ism6TdtwYka6Lgxvym7QSsKNbq+Z2U
9FaDpbAi3lCIEWBfUhDRaLL2ygIHywuXi3sSdxiCWwoX5Aur8OtOlf21WgDYyYscUaHJSSRZiYoi
41AVCg2462WqCvq3JrbNwbwrQeaQaoB0Vcd6FcnOQ2razKzNhRi83tG78Ym2naX/TSpaoaM1B/nx
d3rMciOfj4WmV2SXlKzApE6VV3CiECx668K8B34lyAwHOjguMCThJVKEii6FZynkjY2UKyDci/FO
A9MFdXsCfq5jRGHmjp45H4TsPNSAIVxZcb26U9mgsM6GfwqYOIqUhsdLUNJLaWUN8Oj6AGCJZd8a
fiBEixT7FV53TSEyzzKSuHijpMIgzpDbEggqHqK9OyKewUT+dJDxAQMMyahowkAPy7Qzi9REA036
DKzVU06650wFgImXCw7ssU8dxAr+e82UQLzK8p6WUnshHbWYc1kvVCEaf4MWHxvWxOVNG7BXsNXD
LeDhbfyWfSqdBhU8Zu0WH7TZS9uWvBOEfVNLB97iROXQiBGa4vUmUwX7gI9QnchRySgTAV6/iRS8
PXhdVbqgXL7XhSl7kv/EsR4J7Eb47Il7YjM2YhdjuuXBSzotTuz4NbUOblK+dMzQKh8GxRineznj
tINNiEHO5XfpOiENTyaS+Dc0C5mLS1qAlT4hETJ+KmEpEFVjOvRiwS9AcpxHLb9DVQFPhOVz6jq6
g6zEhCwyZdUxxszejOmWGu7nEaH6zp39TwaQYDIBjkbX488k+fVk2ylM/VMKLqazXsHagGba71a0
3TNsEtvAa6QhLlzYJSGiIrs2JFNSwMDgQdqn3MUoUja27Qke1LV5mxuzkHf94SrQ199rUDIIhMmq
NWXbt1vsTamTOvrCj44gIZPnEEFnv1AE+xnyysUpbueZAwLf0Iv37ApCEzf6mk/RrJleoAAMnlNx
q98SVr72yf/0Pdp+/AlqEQsIfrYP/KU36Qa+QVGqrs04gE3Jz8/7WATfyd0c8RHJp/xD/OosBjfD
6YTYdhHAmSdlw+e8q1bhS/uAt5KxqnDkJqAL83Nb18mtlFeRFzSuGEpNQHL7q8fSlIYazLxtcfEd
ZXVLzXca4LfQXT7Dm9ewQ1/ggF1w2Ad4R38NuN9ceEl6wXv42zHsYqZG7RrrSgWOHHFOI65tkmQD
IIvX55iqaWet8Gec1I7foIr+FLqBPDCBzBFpVEZxlF9f4eiAKGsIyRz+Np0h6fh30GBsPNNvnumo
9uJIWxqFSwmD8uvjgmw+4KqMKNkzlLDJWFXl3B2dEqp2+KEVIJg/PsxfkX/fqtlV8G7EXI+76hpk
K51m+VeFc1QMqtMXAfUjzsRSxm9CRULoISQ4NLOb5XZMkRZ+bDpv3I7AoT/qkTU8U7FaolubHGcN
/foJ0ssYx/jvXLRbizAnAgFNK+5ftUYF5FTknuYxJ8NPVm9flcGdxfUzBhCLHeaPDWj92dstuKZ6
ld0an6PTXj+x0hyFg0R6kdR8uP7FHSh3HiyUafBxHlkY4xP/003r5frEolCX9SPvquCVt+SDQb10
LGs44iIG0ZAFgEFc6P2LCff5aE/+2GSd8HuUSd+9MGX5rSmf3sjvL7+qdueRcrZn+R8NI5AWHu2O
DI6C9swog8+dy9QHZIJHevU5mMcNgJ3Sv/t6VJN95PxLuQoN1BSalYc926k9EdfdA8kXJscIvTlm
CSCdEPX3fxbB3U7oxJ5y1IFMNwuyyQehjBr6Jat5Kqabo5V/kaJUuxhh8fheK3ddEsZd0qqqKpLb
M+zcheyHSsQz9Z7/mIIa2rvcSn7jak9EcLOazUG2pmfELpgVNwem4Dc04HVTOZG2eTcVMPTR6t8O
8OMPwwbF4/b3ABun4wyRhKU6/LIiKj2MGwUr66X+F/UuhWn2aTf9u6AgKSMqOjfsqbqNJnq5BFDH
LilRIrqhamDp5CNo3dFY/gATscq6wYJ3vcix6MruFj2Geue/NKlv3Jd9FRxVYvDVSI6ssZVaTjHB
gdGLlZnBYDF5gO7xMSsGOZthdK3/ecIG1IYgC1R64OFp8jojfc9cfaum+N5Vq7aojYq9HrOBRDNf
K3ukhkmEzDsnAxVd1ODIed7QzSDI/9ZTfDLcTpIGczsXd7EgCP3kQGMJKRAudyRWqvGNcdEgYzvE
Ppf7fA4TAeZQiAWwZWzgYNVBIDX8rHB/U2vVT5uvikRZ6tudxPxzq8/d6NjT9zXihcCJkF9xsOgl
L+W+1tVlXRw7oBm4WJrW/xCmqo2req1lH+cUZUlz0GOeKyIx4c+OCgdpfYPQ2F3DxOcSoWHa4hCS
xs26nu+pmI84Yt3z/Q+iqyFGZVdR548OVryuuoZkHURV9z3kZNupW3Zz7sECv5DMFC0TDg5cWxxZ
dLa071e2u9afcgsqG7GJ/p9r7KnkUrRLeLwPhBGfHncNV8wpgY5K4dZUIA8vDZVcNhkJEKZxO4if
8gG7bXCmBI1OzaSD/C3+c3Nj3Do4HuHFhEIPv1YXUWtitzNvwS5tAKU1oWZxcXbl/OZXdM3ccTWw
3BnIRSsydPReGJxpKqkKVghJPwRR/Pi9ptb7hkXaNmQMXOac3mLXxNVtXuTJ96W23mldelKTZVwi
Pq1CzJjtGNGxVzzJi5LWAqotGTgMX2yt4A3nHS6eKu4rEitASO8+aI9i760b1clXwYI12YJL1kCC
TIsynx9cmej+toHTIORnPwt/WE9U+U2a5npmYGw9sVyPXlQ6XQKfflf1BObEZBKMhGNd+S7ZYD+b
bEBrwlfRF6LAOVbxIDdvOqCpsSPeZJ9xV+ebL/WZaufacqyaC0oPF/Cs1VNvCGyfJmNSO7W5h2Fc
VpBY2mPWtH/swK70pn7Zmb+ymK7gZ02Type+CCf0DU1vGaP2e1X1fgcseOlx6jSPq4Z0jRoU4E7V
SGRzAEWLHX5yzV3u22WLd+AxNagAmzIHcOzfTs6haT+hAuNLSO7L2n+XBBUc2zTrZPZ+YQsLbs7+
xEDSbAp/M3DClQq0/tMw82fpZvu2Gu6+Qf03smC1W26Gp/kqrPTrYWW7mcNR99tFd8kDTxoR+dCe
9q3pzv0rEgJ/Q86C0eVTr2BaG7hE+33bVdCIPF1N4bzke57XKzKYzxNBD54nYe41VE8MUeRLhIKz
yD14qEWmJljMQBqVFLJNtinknwHdMvlMWpY0axt/vRBIQdowAwmJwKxKMN8lvYQllepbaPr9ylNS
2JYzKCYLBp8RQfHymX+tQstfqOXWz5oJTSSLzVyvwpqXF8uu2wvcVqw5Jo/+ZOwjegN+B3GxYY0v
WOxSHNgK1j6p0sw3w0NJ7rU/HRcZgktktStrStuYRq4rRj8QmVy2m+kMf9b2vzvjoaSe/+aAXU4h
HHXDgDK4qPScqSlS5et5q0tJn7TwQp2DF8NpQD6AYeTm6oqnBiDKecnaqJUtI0XAu3NgTYNyCJKg
p0M3VIbrncaXi77ucVXDhf3gTWxCpOkySfX/ZB7vAIgzU/vS8wRoZ9/j0x/2RCeYMAfXllWf7f77
33O+mfx+cwFdNymNaHXZhPg4OQSIiPdrqHOJbgvbIxng0GO/PXo/yeRFHYSKYugo2AxRIPTBKaLp
W2xKcXFjfTTnnr4Hx/rV5zTnL8kKlwBWVXLyqc7kSDk3YwysvfeT05cW8AieID25UmI550S7PVoU
a03Kocviue3ItyNdejQdHkm4xHzO4HtJKfT8tFx2jbJFj+qqW086GHGfY61piKasO8KuTTHZJf4o
wdYH4+4nb24ehqUDHouNl0Eg5ZmTJhSCu26V2YlYKtsocGvGuxeGbujfuspI+VbLF8+rOkSrR8QK
eBo3stNbiyyI66611vojc3lYK6uSLgKssC7K/iAjgbOZDO01Es/9AJPp+Q3zR33xxUdr70gaROfK
QZC18AoM8RQQY8oIeSIe06vugGFOQy6VYcvxtbumKSNmtYRCp2aGReRa60pwNgTF7du7nC95vLSo
vz2tBDsN52L1hSW7qFqlgY0zAEGNA4/WPpWC5ijEQzIbr66nWVTsm/ZUz9oiUc18l1Aer3ekGp5r
AJueRR4ivVaT/HygSMxNfxqbQG8ep3fOexdpdYnjfWBO9PSyQCcdu03QE8oAuMTOv5GB4U6CFmSq
wMbbVSA3WucOL1gSaKg9q7uguFz5s+y/WArgYdK6hmqkwpAMu55+KRdSSLLTeogrIIkgZkHX7PWP
JSGxfWDQbGz5rT03Wd0J1stRCU9XEYBDearKj/2fGYbqUy9AOZXZWG8t1dgdbdtdAH8B5vrloGVU
Qw7hNJ67g4kTLh1Y3BWS6gEVHkXfxrO9cgAndZc1ng+SeldJ0UFDQ/3zVQ77Zn8Rf7OXIePC1lVj
TzqCJ/bnSJMZ/MyHsP9oYDrbXavwZ5/N7DxBFV0Ny38urvbHtWNS1RfBHHUIGT+1Y+YIITXv6mLL
ge5wJxYCssQ6s8mhGnAT5vr/BjoPlH7CA4ZY1ArUs3dyManWt9rQ44pklEGTFpogvFmfV0ZuLx+7
fRmZ568t9P6kh82MbWlyOsuypH9Lx3X3al8HDemQiTQzFjtVbP82JmtBlAwtPhkCh30tPyjMACl6
6gv9XsTYxGlRUEFkJVxLUvW0/l9TYiYJtHG025oFfcd9EAiOmWLt79f6oKY4dZsrWsbZQqi3JXHN
BpzyqQgob2Vbdp3NruPJZy6KIK2WM9M8IMP2dMKt/uwBDpTLL46XlUEBNquIJMpKx8uSEKXd/Zei
n5OmggC88ZbLvtWe9pj3tfJ0uOxEHebCO/PELlzUnHrLd1jwdyYEBbTQPoMlJur8RfXbod53Ygij
HBBPNNBS0+TSkF1hNv3rE0sSg7MN28FsAtTFYoE8qh3u68ZZyVNc16MDf2XwcLcT6Wd+jkedtQk4
yIrxL/0Qgaf2Y+AugqDOpv6rcfOpjQo+SjOpTGM6yQZK7lShTJ+V4Alh2Ks5ZmwHa6jPLK/pjwix
7aIV/W+KmprcTdCM/UqEkwTNNTKDhwVMqqS0VkFLrf1WixyN+sAl8t8i3wAM9rMPMyWyvO6Bsneg
h2eXcsDf3yirj8055SX+SEQJrGKXXRzhZ62Ckl6k+P78bZDVOjWHzvQ/LumduMbG4kkht1fTyFtJ
5rG5pI3RVgHgTdGeNFh721ubkC3Dt/U07zYBqkkCIwFlsNHv52ITroglkgShTPK5sDTioOuiVkAj
Iz6Fruc3iJcyQIYeC39SowxGKhTYuR9MbBZepGFyS7Tlg1e684zMJW7tloLc1vz9vwZzrBMpVCrO
m+Xv+V4pXMvwsj6MyS6wiQDAOJ3nPvaIBrC/jCQvdysui1NLCdISrwagIOENKobA+zHVV0TnOin7
e7FKhF2zknFg6pjjeFYb5dfLyKuoUnLcql3RmqUp2EoPqIaTYSdnmgiP1DtCtzzDvG6rTfMo9K34
h5DMdNbq+qloYTXbAEut24IkGXtztN2atO/F1EsPR2/WAfBqUTxMLS4/DOasYvg86C1xlKg2nKwq
8ibLq3fmRT2PuN1n3CSLPtqTAG1FGgKVq8bJQuy7xeBXmEFowPAIeqK2zUPs505nHSDwhv+FR+RS
XGoEmNyelPsiq6qDK6myHmUrXmHt/ZqU1oMuOBZZNF+ezACXt+p84qYgcWe0nSQMVirZFUpZLiGu
icY2/jeHimddmGbl7BDUIzrHBf/PlnMkYls1XkF696ckfEoOeAvujMlpU0S1Ve9L7ETu7eg1JDy8
Jc8oQez05Gcs0uLrWYenyEDxsP4XlEDBWEVR8k24bs8rahlIe/46m+e2e0lPrEF6ibHz/PDAjqnS
7Do/wrJ4mfqJlGiBbddqephGeY5a5BXKlDJL9xf33k/DmrlMz8DDF8Z8/1NPnURC0A4xC7Sr0a0e
e32M0/W7a+zPQTrQIRtBWZ6WetNleK6XN+am6/4fiG+a/HmscMtf9sG2W5Lagm/fcR0anSt6zz3Z
EtR6KPxpoT7xiEIMGlqe8FBUikYYNCHFfwHT3lxYrLq+NOaFXF8xdEKRphLQpgxLUvnG/g9I9evA
rIgFzCBDy26E/PJ7cGaUP/rP1GZ6suf7zqgpjq2Omv/FGET3W9rwCiNS8OO4fYsZEcPTWArsB7dN
NhQMGPW8I+34h4GoZQLd4+gLjHZejLp0wUCU68vb1DiVklWUbPrBkZ1mHZTrRomJPhoQ3csNhSmo
/SH6cC7xcjwkdWLwQuOmXoQhfHLDNg8MiGi4l7Omy4dudGnhBCt5WdWiq2Ygrp2LK40nWsK/fyCg
Ieq/Nj8RyhtB8duZr7oQ+SW9qPWFOuzsLlbivZw+cuHO+D086YLmuW1jOsz3pFUcDs1Br2HMjKJN
R7LpL7OkDyJNz4XL/r1ud3bnbXwB5JqRK6wl1xWs+lYMgWqQTc+3/h8oB+ntTMsgBUd4vYsjjYBQ
gqIBLbZnc/eEywTZDm6qc/YwLjUOriC/c59YhslBfqvHhSfdnFCqALwjoS+2aA/OrhBr3aJP16wC
QSSMqWF5pcEdbf4SrhM29Ha0wvgKXy6Tkzb6nS2GunAtJyezkMlotbgUIW/TqFbCO6XQAcQpFxix
oS4j4QiKmHs4EgK+wSeCWhae2yrCY+7jidJ1EfAUF740pEDIfuDQP2NOk4CddZnIYo02j0ARJQNQ
ErukPld/n3VqzCfCflDe2NMCT795J496dmLHCwC/HZxsb4BvTpd11Nx2Hwx5K+JrdpoJBPjlMjUO
+ZXO4DUL1N0C6LZ8GL9bFIoZ3FgNd65A6DW8nfU3WLrwWBSw3DSa+vRkYEyv0Km/ZWfkn+Dj8bX4
GPqPUe29+Rq56YBMo2YECCnreoc4IyqommFa7kKLNe3heVSdxk1ECNgoi0FCdeedWkbr3IGDohgm
29x6tLEvl03vVIrZ86tBeFU9B7HhmJd/2Hzm+TB3DOgr3bPKNDWgLYE28Qeaok7hRcB7YxgW9MmO
LZz8x00r3jYGjFDpuf6aEU+dPCDO0jzg2lFM9QPtrP7Be+/lBKjWIZOxqmVY2Q95nwvlHkJBQFop
sHkv2tZ2F9DtTDG5EMRGzlpceNLz11u/GlQr4/1gVAZzoeyuBh2HL1PxRoqEwJswxVS/d/1MYR0s
tMHCUUW9qpDQ6fYtyqbIH3GkSw0N9eV01l44P2r//LkP81xm+Ef2uW8qt4CIofRgISduTaioH5Zt
NpBAbDhBEbVsQLz1tZnXwdfLoNYCV+4pmky0Xd69mphwUApMIrPdCUqCojUg3nxOaYAjcr848P0b
mJLsQQha/30H8iBaNd6E50K36ywCfsFa+fa1Jsbl/jF+lmAyGLXYYPc/tZtoOHwYDXQ7w1DAgYyq
ZxEMd28uxh5fkWrQxPwvdaSAzr8FebS9qtizGJefmnI/2h47xXv+Wg12TwMo9ds25nyI0Cf/FvU7
DLhwmsPpLmFU5aNeFZi5mRAFRzr951pB/H245Tn4Wf8XVvdqWff3eqwR2UK/GYtdySLm56/SrPFh
nw8Ya4dbAVRdFqXQCR9BXP+gdCQAML3mUK+P4K3CjxDgK9WnPGJbH/tJwgT9H/RNQpWb3GKWkKb6
2hTmknh+FqUNQlRlmGYBCdojqNPR/qvO4wFhZoMa3eXJQlo3xM+zrbaU6nKixoMpE46vHIMwsiHg
bTJ4WnCv/WzaHNMmAxCj0mICllWmkqVZGG7Ynmy6pgCjiqw0z91Y9Edz2NscMc49rU/nM6D05WcJ
uvy7IfvnVdXnbeNyEHHmEWHYt1jyqmxgROW6n88GwKxIMOmrB8BJKysa6sGgMApTgZpLMYFCLqo3
c/3qFOAiLDVx5RmcJ0oWlY97KpC8a0YzrcnHnBOyhMUJsvth4d2boHDGrZRFB0vX+dvWgyrYEc/z
qPsg3Whr1u4erdjWeJtayc0iyfPAODI49kNFNJAZjPKO8av3KLHuZi6ML6wi2/T2BDyz/wK6Bq07
StorG0Si9V3JPGleFq6GuYKjJFxgv+8TTaZjb06wPQ+LQpa2nh8X1XXgZjDOe+zezDp/jDJ4OKei
S7ev6xgvJJag5r0tpq9RpGfyryOZsSY/wzbsawbv8p6y7l43RxWx7nmcwz7bXtSfSsGl6AZTB7S7
vfariuKf0wJ0VX3cegTJdGDtI+E3d+lwn3Aug26pPGTo3GDKGZZOX5XzXzFrRIee7oG8+EwxMGNk
Dp476e/QjMAXmqzBLkRwCXr4aM71PdIsE5BPZuSAscksM2NKIk+tJNvpNHsfknOX/pTHAiFJb8++
sr3QGEavQ22shStNEzkVAhgWuJi//H03e0quEMyOm/fUmJqERx/fAjx8TbMlUvZH6qgUFAZY3UWU
fMla3K5RMDvtD8xuLWA8EHoY6wMottphBPc2i1EYkbtRVeB0jAWKT3v8XiufjWoubBtenAibjAUJ
C0CvdtC3mVr7Z16qlVkmNRjCf5DRSptaZOEpHBNQpmFP8A1D+67F/kHOdzSMPTUYuDBWh21n/3hx
v3PcV/gYEnIBM5UEuQ8MFl7BImY0lvfTZ3cOtDnjLGtZDi2vwzPmj0q+jPUdVBGbNkYlthXFrUb9
F92q8MkYIhGyIysxG/ie3WO0OZ2qfP90gZimjLdbyNuH7yiSpgdgxrIuMzcb6AmNMQw+8hkde73k
H97S+CSzrxKXc+1jHerkgOPkWPcMbIxmQh+udCZanDy7z5/rWlBsphihNIxncQi2/9ifVpUgC0u9
uZR/NfbjPUOysXpjeql/+dMB+hE2HVVFMHkaE5DK75rnqcjPzH6Qozs+BfRfl93c21ZO6+77Yz/V
BwldhBetUG15vFif1HsxijaERevwsF7t6XOGCx+O7iCNDki3WkA9jaSshymKwVJuerMqBjkVJFuA
+iBvjJNhB8dGiU7I/yH9hotGelCTmPetWgt4NaEjw2bm9TjXb+gqcMhYBck669avQVO/5QSzUwsC
FCIvlnNEanYZjJ5Chn+EZ/pCgAGMl7komxVXn3FBH8hFVmpkdZ/KZ2150bqFvL15eXeyr8EWdWL/
EzYx+V4qKUJJdQ960pCsQe0YBAU2IfbxRgFYMH5hQEspDrSBIbDsTQCVU3rMMvGG8zJWHs80ffnu
gfWK5wEoY/Kb7zO6hwBxaQWMhaMSPr0XYDW/uKVxOBG34a9n0+Jqkkgkt5uNgIVERpDJtEvNPV7U
jAn32J751+KLacG2nrk0ilvQ2h7b2Dljggnmm9H8K5uajBbc89fEZjHqtTIERdFTNAi2yyzZLKIs
XzNLS1l4TSqNpvSm0rV9oL47buSvTfw32vBtH1peWrh6ZCq8iaUVQff/kMPxjylbljKVNcsi/NWB
UvsgPqpffrVgFUKuLDuawhh1DnSdv06jagJ/W0y9m5fn/AX0gAZtABGRMSYS+Y/ANXPW1GwdtpEU
Li3mDuVa1Dm0e5Tkgqly7B/1ubIDS5u8gsEF8oSUxi3sWxmk8DDX/8Rnc8WCPwD5hL7QgoVczJDJ
yiEFXiWgo23CwSpjkzU5pFbTumv9sbRnaVT3GJDMYLgIqKKNkzee/qlGWzl0J+yNUoouE4P11Eek
V4g6WhKH56g927N9CgLatgWX9A4HDMIsHCIfthPeiHHemDTQoDHQ4m6y/DvlWy/Wvvc6FxMEXw1m
/JZJWQYB1v3rCS740PVlCmvpWF39ruTXmyfH053/NunnFsTrlRAOFa+YYzdsFR7c7Qpfj4gmJl+D
TKIJWi4E0kHEKZbeyLib5nkuDtDrLW6aeuiitmgTgFDRkuC3YMuO3XRQ4ud0vVvAQOgBNwPFQ9Zn
29b1SfK7E3Zp+P2GJZk5XaoRjdN1pOBQfb3/rTPnHy524vZYCktPQqOs4W4b5ciukXSch6mtXxs2
V9GDpT1jKNPYZpbx9R+0z/0bqDgTBSC55A0aEniorDG1dUzIsTTZWEh7vwd/JSx3Hfuw5qkwHcmL
BWJH6wq1UC1GA+xL6AWZQRxAwVRBjyl7n2BK0YDKocp69ftAXvkM2VTZqlznKi/astMcY2eAO8AT
aKah28qxNscLNzf4pRSSk+R+YOukSXkfJdhNJ4kCMmrta2WczTHxYsHF4p8n3wA/VsPvUd68OnAP
9tsjFzTsmkadBjus9GOg7u6Sm1SE/K+B6e8RrqjDpgvdO0E/0rSkZ/LHB89etqr2tyYZOm+TEQSj
pxEMdOedWYWNffDQfJAp4WAcS/N6E+epWitrGw8OGexDX+rfL1BtbE73HdlldWbihuYvrVQzrZbj
1PiwdpoabKz8NN0zUaJBjSCBpz4AGk0M66bf7WdppNY1zVrr5ELcRm806aegMmrlz3niSQX7FmWS
kO+F0BwVSzrenY3jWySJbumrSvNu2WTwoecbT9EVIlPFjWgosqQ7qCyn2hMTX/6rHxEKgaXWJ1ek
NB/fOjHDEBlEkJoUOBK9VA8MC5jIuCskl+Uc0kLTa8mb39pP9mT+frPAThEPGXy+TYfm2NDWfVkL
ieAkLfzfKbZ7WG9PFWbOz0Gqf6ozEVRnfKxMGcQuY7TFw2CZyCvrV82j/AwalAZZJ+eskQBD7it7
t8+42YH7hd36uUlGK6YvcW/TMhjudV7o6njNJ1f9pVUjjIlKbcgUTelGCKYhwqaKIK0oKe2Idqmd
889yCgOOFwFr5Ww574kaX6JyQrW0f51/WSD9a/xMYwEn+q1FVXyf1NBsNVkzX+1MA+ESROG+Vdhi
NIu+n9pxZo/p0qhO6mR9nvSMu2deLw5WVj8Sw+jkIQavSA9rbjs3cZJekmoCNHjfmjNeatfMj2CL
8m1Vy0Eg/i6+XJ3Rrjxz2kS3XGRleaOfnetLqHypucX/tMzuclJ6n9gw9aAE6x2dMr+bIpB7KbHc
4xWToLshXHJ9Ds9h+9uVAUswCnznXKE8ngcn+7pzIH/31pyZrO1ypgc6W0SotIt0YedMk6gLU2LH
lEDSGZx4A3L3ij6BMEn/Hdzlsac37j+hIPSf/ePat4btGffQc7ga2pFtS9AHKZ4/96yXx3txvTma
EU/P0RZ5TGd72nVu8NxB1PDY4JyB6ML/3go9EdF24DVpbL5RGFQ5/+J7SfayGb0TLpKrWYsgFDp0
ACKyYmHWhF2uJQlh5Uj0zTXHHH9zB+nO4WBXG/5ZLjQr1S+szszdNQYCUhpmfgHb7AcxgJ82I95R
o4PYcOeTcJDjvLDsD/x0Ko4NwkmANSU57UJL50iWuQ5UygRV8TEd6IS1quzYL6m+1eSwZ9OfRZOw
YcpCOjfLswrBWpkA8SFN1fZJxTJaudDPAaf/qjwSGeT2UNryBImC6ZPU9CtpDMBodURte+8FyBTj
Avri98/mh0zvYDqTb/BlHdQoHd5M3817g7lLT+T3lBOR+/3bQye6b5ynJMqMUqI9cGcHHMdBxJKB
zRoT/R2gNA1MHAroABVUOouUKA7RtB576neNAhbZ4HRYCj5R9yNUqlGvu/oQtjgjTNEB4Qr0Ct5D
Q/Jx5Rx5/XSj51EqwrKvstBOWmaRiouReWMaYuTE6322Y5pJszBJISaTnLt759DH+i8POO/AmiEK
Qrn6XwiuvwEfSpjpcCoLKe72rd3s6MFeaj/MLgQ0YyRbuBWhWGo8spkOaptyeZVLNYJQNl2L71Gu
Degul6jxImxcZ/TAlp3+dHWnD6DUZYdghMUwa6cgxJxE9huJWL95aznwiQfC8KVhoHWcJvAHjnbn
qVymMN2znIgJoEFqZtTzn0ppjntp0IXbhXgQEY4afaW/R3EXrgW3ylm5KDKQiVj0/fuFgA9x/P1B
nu51P4DoGFBo6JsdDpYms1jFYlFYej8w1HMJBEVjZWPylp6t0I77dqxE5njjBQjjT7qZ6mVyQofK
yKqoJ4IdALUdoKrI49LJqfTowItrgSY5CsamYl1Ih1/vW2oPbGLffnVPRoIaOY97PrwomL7CGwDd
L1TxAZa135Sy1zS7ZLlIv61z7WcKJpVlaWAGCJcnQZ91kaHSnRJdFOXxBfM8iB1sQZZwU58xmGkf
g58K9usmPOz9AIVKhHkWhjWdqu3S8fDITfcjRHIw4CLqo4U1sky6cc2YhQDR2MmbDwbt9nhSGArW
lVJxtVyKgozgomPpGuRIfkjIJ6BAe18tH3ZqLc5Wl/R2T89glnAYnMVuwR+LlT3Qtj3IvE7XtO2x
3RXguMUDp4QPuTPPWw+lf64KvWgzHXgX5rV5icHvhI5vqB+UyJS+P3RKEMqQWetXaLWcXZ1eSbwD
X2mvE+CkIt3soxktrXxijh7IDEGd8hogo9x8IuHVzbNFOGOLDd3ke4g/xUvdd1m4RtwWQDswArNP
/VOhOdHtjmqZ+2pMRvJFmTB5uh0cs7ctKmRlgFBva+tZoxiIAualLVDaxU7Z457b0ZkhMuJAyHMf
g26tX1QjfVb69Aidmo/u4xvnA4UGq+L9tjUcmbDxlG5oRilgoIxRRxDFPCqoL9/C2i1608D4FcVq
CD3tVwjjdHUcPTUSjvlVT4vFrHgLxmcvcs4U9TTOH9smgEqZDWjXd7kE/yPItahBXhqbG59xQKH1
KVIKbva8u9NfSmh/Tv9PbjBImQqughjCMOcmroWrl1iu36pibZ+FTBMgnUvKDf/vnQ+64M7MZfK/
MUKJtCUjiEgk73nGHSJ/XwqMqV8Ler0E/kCGQegGpM7mx8+NIF6cp607ozCml3fICVMsNAh4opPJ
W0/NR+j/P9yvlD2O8antuRuEEZTxFeuzjW0c8mCNx3UDM556JYqZH2ecjQkaMOBTkjaA/sGMANl4
IzMuJJyXdaGDg875j7AZaJM8Vctv03zjD56Iq/yn0xnaJzp4wcHO1ReWbxFay5FxpiTlAw3R28Nb
scq+VSF5reRBI/8s1pddh1JJx7/W2ByGBYBZF/JkREo0D99TJx4vGr1PBz+8CTX/ymnlfQaM6dhe
xg3vZwI8X96oDvM5AmKRR1d1JpkPjE6lp+kBReSAU7P36ZGGD/MbsBxxX7WKJAB7/UCMAWpejPbD
566Ei7Q+arnoHPS2nGQRu4GZDiUlCuautrdtirOaJUjDMmo8tOaS5P5mSw7T1F1zRDyuOPGA2mrN
yWYLcrUuD2xBCOF7G6rtyjd2r7YJgcmX9Ho5Z8K6zwUqMB3DskTC0SHjR+oSxtJ9WAHU4IBV2gSE
MA/YDACGf1SL8ZSiAkdABMGB0B4Bk3j7OSiwzz/6aKeXeHY2i/04VSf2OoQztHhpoKFXlTOd77Dt
0+m5ud8V/kakumL5GyAX1ewgkTekVJnJFKt1uF0Iu3//yoyc3IQ90OJgyQDEzx97NEUf1OOkmCOp
VDEV55XlkfJLrmoD4SY3QX7Ufk9JzfkxrM/ftWxJAXdud7QiX7Jd75hDEVbkrRcC1OlHPD3gSwyW
SPqYA0QZuK5xlM9uq/Azqa3aywIs7NI4yfF0FtAdmj0UFNW3A3L8ru4zFmqu1gRzlpapw3JQ/Uqc
+xNXpa9QRDRDXDYMCCYmGNp8IpzhP3taod9blrWHuGRTuRLhCepTV7uj1IYVwF+Z/HLaFDOKaYep
i4vvO7fnEfl8pCUYtvHtqhpnYvXMwwceC6ykj8EpqR/k97mxCOs8mza4oFQd5dEyFcCxoQkBcGg9
z2SfgGFfRJG3BLpJIl1ZL5kUsLkd65C5A8LYq90h9Z2JllsCatfPpZeimw6eiz0qUAxiokBb1AO4
vuT6wfsfkFWM1218DT08g+FnmuQdFGeD3tcrjYXyj2FlTrrNgTShww+uo1sIPDHkbI7WHBf9ax2T
1Xrijxe+OvFSi+3lnNG5jvyUlzBeJn8ZNPdSwe3sJdyILnxnweBgVw8aDFJJHj6Fqk1Aaun3aGLq
2mspdMG6xGV5NWrRDMu+O6WTqqnC2jQJOmNBqmXoKArb6fHKHc05rQrKMMKGEWT6k0uLjKXbPDOG
Ovp2fyc0QD8RPdFvnwqYqd+3OeYLHQf8LWx+32zaRX78KVvN1IlDMU1dlajFxSALYqoRBk0fKi4e
fRr46dVm0zj+TrgmDR/9Ym6IPJfAZoEDFghtPOzsYIoA4YwJrdDuSPWM9lgvOnat6F6TvUS3uo4P
70UgadwAmKUvBSgNm8vcS08hSFWr3pOKoGDS4FIDEiCwzES3BDW4Tr6Q27yKidIwuvdyO/yhsD4Q
vJUZFbceo5yneMt5mD6up7k8G+/VgdlCoAXJtLY75zVznyv6oOH0u6/6btS0dZeaAkOXoEOp2VDB
3/F1z2R4khLGpg1FjJxwuH6Zp31+KvoATNoP0IYihGjcPZSces1EWzfgS5SQ2VaZXr/bIpBgSXBP
VNIzcAQbmByWDWJS1A4qZDir8CHgsDqplYgVc8G72dUWDx3qNreavvYTfhToAnbfvl4gjNmTP604
WeVQs1voZtkbP9wwmCXIOkVg4oKC1IdRP1SwK65+Lfl5TFHREwtlACuH3DOxEu/aPrRE8A9F+icu
E3r8xSoWuWsrATBEVnNIziyMREOVp1tN7Fp3GR0JpKhFugNYoffYG4M1n4sD6IrOlD4qgRIJLzpH
X5ZZozKBoQnmfUQGYQT3aeCAmjh5d8E2ibteCsQWqSJErFvW+jamsPchlWLfysY8oO4XyyGH5oXw
gOON2RFbWDPo72l0ybNORYLV5A1/RuJTGb7hQ42rJWcMINgGJn9NA/5L5l9Zskgaf28Rccotnc5H
tPspdB5FEMDpGVWWMNjt/910jSGi7wCf0esgmfi4Ys44nczpch6Q5tMnoWhhy6vvcFdy65RVRFDi
GAk/Y3lvAvSc+MhV2+oMnrHrY3zTgcuz5CbcZN2W0zEnVMuM+17PvAH3i3D85ZXmNQKozE4gPrzg
bdHRB0qDuoakk73THMF7wAbpu9PPHXmFSFfc8qhyBEoeoZA4lcW4bSaeXGX2AXeWYVr0P2WwFkXa
2Tm6DZdapEGto8F6GS/MjelSkXBPoPOR8r2gSebybRwj91MXqKqSr0QLnx/F0bi2JwCqV55nvKfE
9ALlMxOpSX2CJbjVyK70dC+a2nXYagpuM9vHiwP/Ae1AWtb2LmlmbggLVju3U+yT140xO00iUc5K
KRjOLnzGydhdoeVrfgPC0Zr1HTNJ/Zh6WH4qhGAOv17kRQSgGTGjfIwjw6tKhg0og+c44ZhvPqsw
AOce1l5QGGvw0No3LDG2U95JY53jGRKfM2wSwMIPmQ4L2k5TujO8Os6hKQToHb/pnbxObd08spHm
UEJp8xlKCoKOZdhqfX/J8dq4lvdpvPni8TywWOZHjZmrUZeJ1/6V6BxMajI62LlnniRC1kCBtcC2
MUxa+7XmSSF5B+6hiR+GQiSyZItgykPW9CDCNHZQ2nnasXr1YrWc+in6LAZUxdTs8mv/7GCM9KTz
IvdyD8SnkPDXqDtbQIyk4op97U4dO+TWIPf8NksMO6nIkfxl8TJtWCfPXaWZifSO7eiTSqKxudvW
gNApnsXiX4m0LaFWuJZxSIpba50Bo1arP9cKKkoyC6OpUywXOwN6GYYnePzb9REmOyOWs/6wrst3
WG5jw3dkBXYlHZkbLJynW8dy/pRJxru3gM6TrDxP+oi6Z0QWwn6mIinUDlB2Fx1Ofomo5Vz6itUA
zvjt6PwXNttM7BRk2nRJr7xwwUr8EXWBEPsTo0Az/rCdXED3KTbRjmWU4AePhcgK9+963mocaEMN
z+XHzg4Ogr4aVE51L9t/BMWuODeuBKxHJI/onDule6nho3Ae6eSmCUdCwc4N32VrVj3DvFTkEqxK
UrJvGexEZwn/6gIFleTSz7P9uDhjmMZbEDNJTPiQw5En9UndJyPZLwtGq23JOQUFI+dCjt7ntBM0
BWB1alrLRibLaQmHds824baLS0UTAtBiqnhU+aIJdbyY4pc469UMb53I4NK276V0AtaIiMFlKhZ8
3/7gr0hDWDihePETe6Lh+Np+6Aq9ZjpcuOWbQzHhWXynBD26WiqdzZysfpcqjo36vL7/RR/gK6nL
gbOxqWee1hwzVzSeZuL5q/8CbDZONH8pyPcy4DALrAqPro7UUJVUdB45Nv31Q9MLATVKjTOEpils
CG4KxhFPzi5Gusgm4NZM5uIwlUx+9WiHjNL4gI/Ykhkqk3m72vm8Z8GuuI2Q62uBcv6tMZFs7DX+
NWQCJc9iK2qsZSb53Ee0FQSBFXj7vt8hbLuTpp6VhBf8clduunAqMwlD3yFhwFjXMtu56nYG8Cmy
ldyc3HD/dlKDmQczpiKBrevdFysqomemWKVM6TnwhWZjdXE4MhtZ7NpGhCfypnT6Fiiz9ECdlD6i
L1Gfji0vpQ+pOSmeD/EAzDhxC7NHFp8b2qHjUuKkacKCw/q0iCARzqTY+F1f6R78YNbBL5bta+2Y
l4OC/vFNuNxVsO4boOlyFzXIX7FCfmmhLjOfvzeRefm8r2Mtf3d6MekEVsnXiRYTYhuXdnOf8Mo8
xGGGnXMwV+lq9vzNEs2QPjyPUnB7FuoHR5JOw+37SNWgfio8xz7ygaAIWKNwCjXd+mG2tnA2Yku7
37lm2KVsTFhryRzwvX06PAq9fTtJk8roJEKF6qSEJgf1FefMP90xuLVtd0wvResqd7nfbHWT3TYV
TWPURjjpcgrSJCVmDsKWND4AJjPZIwiTjR+H6ng9/AbPZbHZpsu0LLyM8DN9xHA36aWNh2HXvtmJ
tzaed+aL6fX+x7HzCrR8hQH0pwza0NIJo/wWpFqeXtFhAe3rOHHgmcmqAmnfrjyDu4bx1WAflH88
KY6E1gHYxuQZ5o5YcnEWANyz4+l8oEl7kpFAZ6rtCSTugdnYxfqpM1cLD1vtJKNe4X9exx2mhlHq
QF/4PzTfma000NzGTTB82/ILyWYHuHoSVpWpwQFnoLtcAXI2JJscA5PnFJTnRD4zF12F6X1yy/SL
iMN3rxx4/Ae/pkAvHE9l6+erAJD7lWhBe5XLbbl7VicLeHWVUErQCpvY6VZlKZLwwyaGqBRTxK3J
6I43zMdUiREzXtb5twQy+t+2GRf9KWzVuKUbmJ7iSVTMjdIFKkgAyEuiCcSA8YNJlpw/xm8veriT
h5hG6cxt758c7+WAH1GAiH9opH0V/bmbHAeh2/uOFzNov4ZTJESTrx4/M3LM0q28ceocxSjqQ1w3
8lLd72Ffyqc4EFUswKVnr81SSrLcxLfagvaTy4SAjHS1E5fLPXPTymhOLqpdNKBInRzvGNnipq4X
UKwQNDed7nE6XkpQ9cmDXegjybe06MNE7Ak+NUdBbYsPv1v5LBpr4V/DYyYsJGS3WpUu8rMrLCYe
5yIc608N9OZ+bzNP8ybgeFlsnJiKbyVGwxzgA18EQGPRwLwVih/U0JlmAVyosRXiJE4ZvOlNRKbi
RCsr3ATX0ukII26WLV5fjL7tu28L8s0RG4oJyWFO1Y75rKw6WPMXVqprD7zbC7S7eNqsIfO6MWgK
/Zka11SqXVJEvhMlQMX+D1RLf7a0MdgOmscMBCFI0s9cGA9JfRBx04Fa6aGO+Y7lSr85SHV2eIES
2NP4SyuOgZN0X+0XdwOIP3bSjn3FmMirNmy4jQeW+K+FuLi+ywQOr+C9jxtRtvljnpRRaHXmu8TJ
8GxVXm1RLCqtbah3I4pIf6xq8asZPftsCG0APdOB66GkeafYWzEabxlXNz2hOqTzQqwDvBxXI8+L
3RJaSOivxciMeeYqDY8vowuZ/26RiT8a0+u8YX4UxrVyIZreCALAsARQKW3wB6VSxU0r8DMF0CFs
ROHZTrNt/iijmFJgkAQqGmH2YIpauEJwxmBowgIrpz8pFGOV9Y7rYNNCqeomVP77lxmwI95E5fTP
f1OSrVOzYeay4hVNFUCON8t0cGDkVy6W68lnDwQM83rLmVuBlL6ZXaj8IVhmhP07KUEtxGamfY4D
g2vC14iXZ3nQZIfTcQDoMa/VdjkfYI3Y6ldqlG9yZcVf/Z8BISETGK29nzQ6P6USQJnY4qxEwXW0
7Leci8vMMM9WA4gooafgv/Tb2ZcyjBWQjoJrvJneBIy1eNSMy2hxgLbk8de9eAGnYBU/rv8SjuKQ
3K+3/36qDpYkLZysY8scVxr8Be094XdNYSMLVUzIsuSL/khjZWeAB07oA3yAGQbFQgBS/F+GO8oU
mD0avVKwhCiffx8B8+nvKILKaN3KopGJ4nWalCFHJ9KSsER2B3DwfKnyfYMLzUYQ7zEuW1pKT9J6
enhJQTY1wTk/61WqU1G7SpGhcIovy1Mm8xaIjTcgXT6yXrg2HHc0hLBa8FCs+EdZt4ULyMvzqwqU
wCNS6BSJUtmDImrDC/88jry8dc+lDbUD3dpxQhjpOaWYfa4K3iww71g+OxAE7FY3UCC1S6CyhUya
9RDon2HUuffeJGozNmPGtep7iyNYzPMvxYv6vb3uegLE4NJyJg2FyZx72qOW4coyednAtpzFZb8D
Vv0BIaTzi0zojfSZyFXo4itCHAtjrr2tbWOK1Fy9j9molSfA5r2hoQnodGiFvW1+0kw/byJ0rxJU
LHynCYUIpjmCXdure/CWxnzqXY59vPM4MZ1GCYWSJK8kGoxHfPQnzqq7CxPp74EdKC3FCc57drMT
Drs8ZCt2PzuWjxDe+J48baQksHI7rG1DNANYluUUJfBxI1o/7T2XWoQu0xPLhD7meN2aY478H+Nx
GXfXsOX14ozYfmGYkiVK/t3Atjk0Lyu59+nNGqn2ntHdUrw9xb34ggkV2X+LQHnGF9RvYNXJZOdB
QMGDfNNBZPCrWFKCWCuqdWGutDeLsFqrJQ9jTUwPLPJLUbWBemchmFoYK1LE+emHXPdaE+ROXE8d
xxiwm5t/9ip/n2geklbOq8VuX9g4ieyR6X1oqmkB+hwVYwcCBXqOV3Bo2NLQKVhOWlM5RQvqDGAF
0Pf2V1SddB1f6XGXUC2WC6Zxqb0gUfSRdGBBy3DeT+lt1SHEizQdaox7IbFiq9sx46x/+fj2aapa
4Y/x35zIpL0eysZgOtf0MtAPamCR5ZcKl7fD5pWfIVpuUo39Kn50Pg72+OsQfES7pacyVvu+aw0w
PKsw3eDgpTIEqYqt5re9k8JDvoHxouQrJcM3A0I5QSHNBDJ7PK0f6zt4GZiufmLRacQw8GF+x5jQ
E5+2aIcx7QK0DI/YYlXHUSeNx2tiWol8ngA3xnuO3is0mGYyGQqF3mRpuYzA4m+m/UxSntrlxYnu
X4FAQF+ZlEGakH7YklZbbeXaAhwEVY/Illb4WVhFreu5J4d5516GtB6uXRQnydLWLlJhPxA4kbRD
g8Tkirl9kUZkNh9imiE6u1ZTbRs1pq5gjHvAPyVulcBdLbUTs3j32AnLa0jeZQbJN+C17E0wbXxn
44K77Sm7x1pR0vbagwQofgtL+UfGY8AfrCXvmlGxPUxayCUrryYhJIJ1NnICc+8Q3emgBsaw+c1e
lhlnkl3mOIBII7EoMaXKNCpg2iMYlZQLKoY8Die07ScrIl59W1cMNHyEBasEuHjPJJWD68gfN/Iy
3+WUulRnV5E+Zdz1bZhUZlo+oZCXe2l+n1DBF4tIKhwOyJoPWp3a4K7tpfX/C/YOLfFbHdEJWEak
PbTXGYBQM01JHEiLPgLTdI7FyGOlGsio7gtikB4xpDOTpS5UyE6lDeifwgyJe2htahHoet+UeTrL
Ne7t0n91+6wjHyL6LLMNcwO1jH/OOuLt1469q8lQhw5Hwbuf6TWF32uPKXMdpkWPstmi6c/Z9rvU
WX3jXrZgY3J8LP4L/0FW4zDBOj+qPSvpGBD1k3ODRPXpcNrRBdVYUYdJIhTpgANMtAXKVQLD4XAZ
WgfiN/VYelZSLJv+lhMma9I7cBE1zzTa0T0SVYU2XRCDfUbXChOSO23Y9Gm/hZSUfsiQdCsMnHXE
gv6CRNOh1AwL8EcKi/kXOBV58CXXxsNRqv1780OaCSrpF2QUK2d3un6xCuendGWWxIS7YuTH852I
5S3ZdEnWXmqna4ThiZWpO2/3/YgUbs6rJ0KvXs/hZPzSGESRseZGSkf1pEfF2kxl4rvFdcoAINk+
+HR+v81/LeL+ES22GDQ79ZwFeOAUguFUxdRjrpPrX5rKHcxqY9WrVcDWLfG11gCZFPn17e8livEV
jtPBx+9yp4OdXZfh9IXUnAE01UtXg2/5ApT4i5v4CbHdE3db+puOsjKPs6TVMtxyJXXQex2io5F+
KBYQxKHF0AothgNCuyUvrVzYXrjrbELqs1OIB7Sqn7hZPJrNQ18ygh2cGwYiq2va+0pvwscutovd
qKD2zI/Uc/C64w+v6eeXnxLcqvj6StUOCEPBEWujcdATUsqm71K+JMLRowcGuZGWWvM4O98YCDkB
LVKLSoB7ferq80KXlFMwBW1Q2hAC1dI8ZV5NklTfKrzWFdjUrBkBF9dYt4ZV8SusgnJYnG3eb892
O1zr855N5ZU7YSSk5zfRQ0GHxFmNIZXvmYK9XXJNUYYxIbWA9L7nkPF/3yOVgSzUJnxerFgMKv7N
7H8C+pvs/AAUPJ+v68fQnl0J4//SvIWmtZnTtWZmGt90CPsSMu94JJ9GwW7apcbN4WVnPe9u0g+U
kMSAPWHXcWdnA13eQMhEIOqiTbUN+qUTKMA7Fn1jGyYjm1rCvyAT25XzI7zsGECCcFYsw7km5zcA
nKr7tY1UNkf086MeuTiYlCSIZ7NwGQLcjmQkZiTMbpkIRtQOZrHvzBEDf0uMlgu1vPEvPVZQ+e9/
cJL5xyjK/AggQ9kg/xLAR2YvSHZlJT59Xhn8gtf4brT0VRMHdEak5ABBAxOGSwabHdBKQleJQPlG
joAsvyE6Wpq5JD5U6nfOx/kZhDicMyDvg29KdFg1kvv3FmtIUqRqsLOT9qkn6vAtYPwD1PNv5Qd2
MQdbTtYycYlkIF2+gtf3FOEWpQjMtXin8DyJqywwkUGT4cBODouUL+UUIU73iuNYBWSQA84eYO8D
DNVDwH2rX+V9h95KB+pYnWjVNRsJg+8QMf33SPssicb28jIwqW+O4w4ZUs6J0S5zymiudcd50Yxk
SdxsV6lZP23m3oAhfrWxDCf6lXKaIdsoVcry+8SdquvkVY/f60R5wWdC374eMMYyLautEJHdqqLu
PmVRWZ99qd19ZS5qMDBsNY9js8E2andeuVcd2pU4swxy/IQvarZ5oWyP7MQVHL6ELAaXgDdctx5R
062eEnbYKypjzZ9aJ56IAEilF+R5tWapG3OFltdOLgPY+D69MOIWNM/QCTUKYCZTUNaM2iNS6P4V
3e0oyjnWQViMTwS24Nj4tBxTyenmq2wm/Sd56O/+jlon1nmasUpysuZkJ3uO94uLQLHMZ1nzG4az
3R6953QW78QEMcJemE4vOjIH/U1dTe93lSCeB8viBpJxuDhoGHMyG6pPzSCQ/L/9gMb+Q6au/fMQ
A3/ZlqijUSe6gwa4WL2Tr5UMLtFWk3nx8CO+jQwsHOzkDmZTiKD2A0jV3dIQ1DAjc2Wi5O0ArTMA
/Eh7urxYPLw82zhbYcSmKu+Wdo2HvGOygqqgOWzlOgXK36yK5W851T3WquypctlEPmStxvevdV4C
Vhst9n5iShqSINJBckzD33Oca0tFCYtnVE4jDrqLhc0Vdzrkp/GckE+UYI4DWC378l3rIjSAnGNC
w13V31gAwbqg5BPDhp5JPTHxedl17EgTJw2UNXOMrNru+QBJ7+wx8GvRf6r/PxG4eEpjq8XNY2ny
PmX7326s6MmhhHZJen7Ru/wuSNVXA5X1QE0JHfJ4U3HggeAdhHFoN+BlXFui9ler3MIjTk/KEE8k
5Ri2OfSEdX3mccP0SluwZLByTaVS6jyr0neWuOciAbaQF//UK+D2p2/2wThWuPkoXlda15F2HjTe
mlsKeJ4y7A0O8VxtsjKiteYafkD+yL8uuSI+xl+PY3uqw+yjjpJIucduqwcJCie3oJh7ZLrtzVdk
QIUtsaYLgvCwVk2+BmWYvKYWSQi3zmHJs8mgZsZc7SLKpyWfPgWnCjqoZ71VGUfSEBWy+Vs3wHxO
UDxsQZksXnag93hN06ae7FRyQPTdnfC23QXN+sL4QzBewpjXW3BHoa5pP4Z9R4tWJA5N1ZTTBn2q
sN9DpfRLEvAI2A4q+rpZuyEGvcULmrZPX7bTlg73Z6AHmdcChw7dGZodCMp+axpOyC8cpTIyby39
Ulr1cgu0DSXuhVWIQJ+JQ+MMmDRJbXcQCRHqFCNIZQf61eN3SWxY9Y1QIFRWCN5l9uKc+agBA5Nr
W3mrzvfDLNjOWpKMS5mm6lZzf0acSV/zklyICr0pitUUTzSG90tGFrR6ZmH+2Fguh9NoXfAA9k3r
8XEfBXYE5lQCKiATSvVy5tmpVeatogEpFmuQXBu4mxnhcqhsc0jAzyjP2t9+QRMgZziLqvHapnFK
u4/xeNPCHHfyyELwokTfZxxwmIH5YpxQT7QZr8dzeeRTMIjMDU6kJBOAigu39n75EGTKPzVhux5M
qWDLJrXHSyIWMAub58mt29hWAJf3AxHMS3o5mJKS3vgIxLz96DwjxqRXDLRRNg96lHj/Z0yCpWpn
qZvkiCPbDUSFSK2oCbSWMSRZRy1msD1QSf8NJD5xJyvNltD8D00ZtPeguj5/YbsXJ3/Ce++FmkfW
y0m8IZfTZh7V4hWybZI3mCTtXC5VotEWUe9tm3PX0flHZUnz3NtpW5Vi6TWtZyB6aUpHFdggt3Bv
hZugKnp1TKSC7orgkynivFPOBOy0tE6c4IyQDJOmp29G8zUDjvyzPTKkXt4BjqFslF4b4UQnKfkm
YPuzVZG6wu6rd2iBRwP1piTG48CkLTUOOG/o8TVYC4UqAxfdAMvDQmBR/wbO8YGsgU1QBmRwtowt
PYw+r21qjU4+97VUuoceXx6vi01wa7WzLk26mth0qFXfo9MSiFFPgT7gvBQlNNHJg6tTTSXcMehk
AO1RzEZdHL3kzL0AW+giEVK34o89uTU0pQxHEzOPKGiOVh3M0zdEp+kaJomi3SiSKn2qpNRdJE9g
tVYbBl7qFlj+YTY4fMfHSI+MBtaFhXaQGLnjPCldwxywF2X1ZdPEADAMZDnVClhLFMQrFIvpHyEQ
+O6Wrxwd/TrB+HKuRg4Xwmlshs07l/Aod7zqx+NdguCl8/zzbIGI7/ovppgeyHzV+hC7wXqW0VNb
OV6nhgV5HEu+J6CYlnaKjZJ4S/2Ncu8EIoMMfrv/ZE/KXwJAwuVx3RM75seIFMiOSfZvB1TyLYlG
yaUwHDXAWkQiqaYaFO1jBbpjjnhVE/MWCMZMU7vykpH022Co42foacM4mYCFKm6UQ3idF+tl+2Hd
A9WOI3TkjXg6/2A7zyd1F5TuObSXVXeXATcxJ0OgsiF0TinseWu1v4YBgsa/EJFiiZlyv7JdYMtI
fCA0xZ5tyBxSH4D+1LkwotACNQOTdeDpzPdgIoM4SUOxt5/8VEOeLAKS5fK6LIhzBQ9aebFMdn41
vFAu94Ye7rJRZK75cDHS1BxwIlkBCZGPMTzZxKeT41gyrjNKsDZcg7aiMDUmOgY/yMFVvkcHENHM
x6+ZeWxLK/BpTJ5ZTDXoiedEbvEVdhG2pSDJ7zSrAhD8s81iDxcAs/LLQNkSZd+jGc+VpwkbuVrn
+ibM9l6bdCXMQc4ll+7lID9TDttrMqRGekCvIVDmRyKb/JYSZOoQdVvbo3rxOe4ql4FGGTaxJIDZ
Jt+2piQA8p8upIx7hp4mRsCfOPtVh7kvuVmaW1+vox3bqxVWV9Iffx9pPBetSl9Dyq+eikGRPwke
kNSH5+vp9CN2cdcOwBmFszM8XHdHTWqGd4zCcSQflDtk5pZTDZXfB/H0MGU0lT0d/6iNIpxCnK3c
Bu9G+EG40F2G439dY1AZAJKRupRSu4cXQWyVaTbmskpM9fIKEnFKrlh+G1SkEFPsjvifLbYWSoU3
U5Z+aTAxLtDB5e/aAd1FxklrfMn4ltCyxlWLnb4VnwzVNK1aFgjJF1cZHWpmaj+E2c7//a4bbyzm
P6U563rz3iMPQy5NoS1fduaoBmd9vi7FXwUtAoxb9qtRxo58Wa3o1bS5vt+jZI4N++SwOSaoJoFm
5dbVdx2WUSe5nagJpW63FYv4wAnFhIXutOnsbKZ9uUiV7WTYddeBVsWSkz4kheqXeAlkPw20oS3U
B6iuoSA9suGphsclJQX1WIApkDjIunyO/n75JsuRkh0TgAdqgCED57O6AfdR4eOQSiXYIjw2PT4m
IHv3LlnCVZ3uAByr6WLBYldj7TG6ZDjl9719+5KiLPRlkJXi2edp8pFDhvcW+7Yzz2uwCV3f/rII
pJUbfqyYuQG1UAYRXQ/J/ObyezLk94zW5qnt9nQNNex6ogWG2XlGF9Izqoz3VOx8T0WUQw4FjRWq
oK5HGlXaGRs1SiB8qJaTc6idqYNUvR60rUsOfJYU10hUGalegyBJ3iVeUqheJbTH8eCw7g+n+jmd
jQlJ3yWClWNDN3wyn+cdQ7bwrSX5rEX0j0nRfUpt7KctzSh7dNVwqyU+D1WpywoWF2R5+t+12qaX
HqaMhOTmMpFnAEK43/GF2b3jvZTBw7Db4A6gFsFVS4PQiboj8ZQSp0BaCLtXOjW6ShKHWAAdPydB
7NddC1qDgNN11q+cFIQXWQuW6xWn92kHUaWOR+v5FvR8KyXmXmtGUxuecEmJo6gNdk9/e5UIYiSu
tnQ6WVEa3DTsIckfwn4OxkstR9KCFlXz8okZ1zLPPTas56ukT/vudgSRSGn+rwlBtHyYLwWZ7oZv
c4UzA8fgJa+28mu4shd2MffhYCnYtJIQ6cUgk+ar3eCng/9RxjYJzu1nn5CUmyOSr0HSx35aTe7d
HbnVeA/LypBDpGgda6tUniMDrk5TRE7mbFYAiSaGO1FJ93uipbdcltF09WQPRdyVcvEbvJcO4BAG
q/GvwtwmKwmhp4N1aUvJOZy7grEqjAnxbkNS6Q+ut1txaLA2Wl30nj2jn0FOGieQTyke6ERvDEn/
FzY/Kk6MuZR0BVBdfYXkkxH1wdDi1F3f578IfsUSxo2akc13ziI8jFXUMPBkDzEnfx+RJR9e1hLt
uBYDaIxQ1DSTzofR8rAzDW/oifHKfcpYwIPyj1KDup2xi078tnSJ0C2OYgPS7Wy15fnzsM9SnpBQ
FiuE4RY2Ut7uh3o0Jbl3g+l7bAU9jgza462ljUTNY5GF0f6lTp+yx7s+59VreDJuRydZIdcmWgz1
hT/DoCGdAwTyTFd9t7Q+PZ+fl/xic7xArU+UUYXm8kpTz0rBM2gmyIXXF7AatcXbieDLFTmB4r5o
lCz9QDsEweO1lD6SZOI/Gp6C0T+M3OGyA4x4zXFOPHUsX+fxiwiE9tH2fs14c641JwD7nkW/jeYB
+Wz0h2zm5tdluQEOWoTC33J/vef2Luz0i2wJ2ZAjhTQ1VW8LQIJLS7xD/GWjaJEB/q8HP9roIf4d
d9OEBX/pb+uCvlC4M7D5c7vm0/NfZVdGjvj4s+L1fXoBPnBSKUbZVQ5roMyvVo6dgcmvgKsvYa1A
/jH+rop1nFkdFDLqS/0DSZqNom0LlaaPT4HpfUmFqJJmqzlZqTEKwBNNmZVDtwb8SSM39PPxURQH
90FxfRdW9MJ/4v8ifPfkwa+h94JcdRPNGW9ujqxaMLVJEvu3VUsxZuyQJEx5O+rXMXwM8l4WDJGb
cwQ83eUzsse9DtKEdYptfFDkx+Hw08KTDGu86QY6pMYPjUK6siO4WsNqwDkACKwmPqBJ7niU9KBi
asi79r4qSUCyh3SRTUukbPLBpxxxaZx3whrNoAxsb0nUAJkMTuURAnTpYPr2CgG2ZL4H0VFL3/7V
iKb2rWSiwstSd08nVrfUqPZt+8A0+q5vPRm5druaZPsGOpL6XWAe1iBo4zDX+1+wK5PhihihKw11
5GUOPuHkkgIbEB4W2oBmWXi+PaV+xW7Z8OLUe5cMjwhhXL4PfNn9MoCcrq1n/xxUhcyCdAD97PCK
V7yxgUz6hgE2lB4v1X2XFnWmr2KeMmESjQUE4LXe5vKbxA42MrCt5s5KxWXZsHlxdG369RtHF5SJ
eJIG5nai6DoESrF/tsJ1mcGQ9VWxozFmnjoTOLt+gH5Z0hUkwFwRh/X69QPc6/DA87YXElMSi1JN
IapG+bbt8NFPeAgvw5QlWpSRx4+fil0yRFE95/xx+LT5jfMKstlQntLAjgO0zRMOdohDSVFS9R2F
YdvCH36BH4uDiee7EQGaL/43rNV5+6NLJTxCFSsf+awMd/5BZjM1pBQDS3pe4HUnd5usSLtz1Rli
ayYxjbsM9xjYXr6aJVVq8qUVuzeYEU155l2Qv54MucTqbQwOIwO6uJ+1CGMy41fBC8lyj0YSg7ms
ywlJbkRMB1E3Qt3/BHVk33sRZG2goEfd2cKexSzhoJ+sF8wr5nwvoUeVUfZNMDa+yFqJslYA4EEi
XuU8vvM9v9/iR9ulGXixCoBEL7sjdU9Xs3lRrtxk3Jb1duSNsjbqFwRqOxwe9FAoqodyVkQb3V07
CdKH+aFO5Xu2+vDnXCJH3JULNNiCuFbZbBIYsUqgjwRnVcfCqTeGha13/sLai1Hg5do/0zMH+/Db
FVEP77CR5YNcKAfhfczqDcmgxjI+vsCHhe4Gtw5lhJ8tEzsf78XVuNqVODlto/z3TSk8Q2uQmPZ0
uXK+btVIrUjZDJv67rzHJ6EdESp7p+A3MO7yS+Shm0JsWKcChXwS3vVGRCU83P3QeSGiSJ2nct+D
u50fPAEun8DxBt7XcWa5M4KJv1q4Kpg0wNqeRTcS8Tk6Drla3JqN/pNZEDqc9PqOvoQ//3rkeCVK
23lQmat2XoYaZSxg6q11v5pJP3qqKG3Yq44QhN2dx5EyD6aU8bibqNc+oweCWm38SFtIhTPnu9q/
S6TOtL3XqLTlsYxnQ6TT7tBkDedTs9Ybbwssva3bzDq4xn32FzzM1oDCj/Eo2G9wvbkKKPIOPsp/
AYEAa1jvfRCfCKxaT0xCkXtP9WlHXOIkNK12M/ugD5CfhJHFGh93PAkUJt2SPad1jRmjfjphvIA9
j3+epAdhLWcTwGeMSuwuYeTupVLNOMA57fe7YFBF33U427fhg8DVTI704zVB9FM4tPaBR/wiEuWJ
kJVdcXyGHSszTlPZCxfnSguknCsXH2CbBs0fciKsewazdVok3wR6SGjNjKvBg9J268Z4BZYOD2Hn
c1qWWyIF5HqJfFK8ZEe4jbhs1KX6wjvtxxcuuCRBRMSczrUr+l0RBM9BJEwrRFhw8UFFYgcjOWTC
HrQKJeH9xNewkqQ8+MBIgQRbsH+ndP1uYQgvD5RG1dGzYnepeTQZEQ7Y/4lXjVG43xiRcB10EWXz
LrUY2yBwMxXhjHwazDuf2hxQM7Od413ITKl1sgk0qdalSS0+I1YPzHpnS06W9tUyA3Fo4fupHUTF
NKbv44kYAFdVyE87n6ZUWH9LRteDkAfrkWs9Bdd+oGwcVwwfZDCr+aLPLVlO2mdQZ6kS/mvsdOeY
w7lqeV37l2PM/AaYg+eIeyTbiYRy5gxnZTH8qBBfXC44wSBIgJ1URmDFbKeQMek7HkurmLTFjlzS
tL/yrlHKltYDLPt0Mut5qu4Hsi75v58m8gye2nurDaLxiqK547KmO0zFEt4etSncdQkWqXhap/BR
nvb+HsuWCeB2BNelxRYc1rxrNlWJbMJALfPE94iDqH+y4Qkbxt57a+1cHYkxJ/2KuXPEG/50VRN8
8ZVzshCA76E3dezPD7HIjiSUKbw9HMETSi1mWhACK/gAd/nD1BIGJpRC3GgSq95owA3pBjKeyC4L
KP44gA8wWtiESuZvF/Jn/gKUe6d5P3fjv59Z0yB8lvxb819v8yKgkkGPeZvfkoEfrrPqgvKkRFOu
fu9zintSNJhXV2cZ9OmX1Pabr3xfsGNdfAlopMay/dAk8YErMociOEATT3Ru/H3FhLKxP6e91Sfg
AVDoD9lz6o+qcIjK7CcVzh21z8XC6tJkDnhWVZ0lu9P7id1XltWcSXCpcAN04mY9woBrs7UasU+u
CkvesdO1GY9s1vjXmayJfiEgi2h6kZjyesyyd9+gkYM9dcJNBkvHkQZOPtp2Zptmj7Y0bYQWmThC
SkdrmAnmO9/T44A1IT1DsAIcQYDKmnA4X1BQ3I//nfakq6PfOwEFWKfjolFuCgQxukpld1jU+HMW
OLmFF+Az+1CGMCemJSbO8ctLI6FrKTxJn/Wjt25Hss95ZjJXMwNBy8nKAm0rAFw6arc72gqb6O0a
yvP6W8URL+6uwf47oyUPFoNjaedA/i2hOdb1ST8R7D+lOG7tYLRzbH5rnwfdzvl3/rY+8L+rMSCo
Ht4U4CnZGFZZLwj9y1nyBxWT/1DmY+CLF2scbh8wdQedGnTidwNU4cMUaGY7dzfrepR9TypCVv81
ii1HiLa2JPQNnMiHOX7VgrqeOxbtUjG5la3TRfVByO6R1JgUdBQ2Tn7MA3TA0wrKEm/1P0ULCxkY
XnEOWZrWyg341Q2SId7xbPSGH9Mv4MlPIb4nNTpnGAxF4Fuo3mg6SD0TEXRgLgADuRZYb23O6uCm
EjNSVmleNXcrdGLJKlDToFozZUl/lFmfwJeb/5/e29604Ae0mA/uOvvJFKGF1FRwGn0zSUDCVm7Q
FaEvKJ+WvPuson0tXMuU68Fv/vaRdswEpNywUf6s/shtK7Kd6oW1Yv1Sg9a1uMgMQHukt04asBq7
TcFB1RNtDp7MV8A3Gv7waIchJoUAV+WWHIv0FgKQB1Wn0aR5XLPqWTy7JyZRK6kTq+uj6dQKIEEI
tTrDCHfVapKw58iqAB0dnjaDL3cmcK/c3xPubtuPVNAyiV5WvQ0vsP4ZHw0AprtCPGygb6zPK3rN
bZI55G1eHiVtgTCgq9h4erOaIIML7wEU2hJ5mVJnRLVEMCsZ31DK7M85G4A03dXjO8C20l02HNl9
6Q9GPY4ib7V2tv+vSZjyw1TuTxI9kvZfex0lEUu4L8IP7CDum2UhwIc2ymxh0F2RW1s20Kf4DFsb
9YgazAd7mlM6y/W0saLpalR6s3RPePb0CPdxG43RnhgViYFZfoCCf0eEDE/JJX86xZPfDpYcGBJP
ki/NadrQZvd3D/n83emg51Uz2zC+WMJ7Uiiw9YDvMa6mIwLBPz40tY09QawU/hoq4YMUfKTA5L+b
dV6QWseYV7DxGyo6udqV0g05S9xOv8umQkcEm4wF0sg4tzwDD43JGD0Kpi69GhYZ4wbOYs8iI3dY
Gl1x5Wy8Aa96497wDAilFgx5Sk9x4nCJW2bSCS/l503bNsqv2Lla/tlNWLn7oqTNfCKJnIwMkYNN
9p6Uy+evlJYCCRhdldZdG3e7qHXe+DjK7cy+d4wSL5lofkW//mc+t8ud+FyWa3+yTVdrYLJzcmJM
CU4kTx78ArGb/eZptxy3+B0Ix3NQqcKg/iAQbfv9xZ8Jn+b8MxSDkp6xiLrCahRs/MBGel/kbExO
HbY4idKvju829Rg4RfDQ9dyfZH3RvrPjduQdPMvL5USU9YfPpJOYwNexSauv+C+62LEowSn84P7f
XBxCZMs1njImf0LS9fzWw/MLzHD/DpEUfeXXHqAyTdzVKj1Fp+tQJ3Ru2R+iLEld0lcBUylqBKS1
HFw6PJb3L3kDdm521FWtSbMrZvDM9lQbHOjKf2foxkXfV9v8ZQdTDnbA+DqupZK2SdaLJhFJ4xSd
qYsIStw7iJIR6/5PlYqOIxceuacdZ6vUdNqb+lfchJ4bvmT9VgscJPTEwH8ipXkesBt+Z6Y/80Db
XLKXnkE4Lxwc915QJIwmj2YxebUtGqZb2OFhnztSQk2ZXywDeQcMngGMCvs0JDXivB7DKdEwEEyw
k4sWMHxgLoZKgTqdQuJ26FiIJvzsyRiP2gUlyaDZbT38lQjpZyECwl/CNOTq3rcTbqveE1Sys26c
wcBfHb3SLRYceyaNsu3CHb3o/scjFbXXAmJH05ToHD360HUIjQIOjtEqV19PZoBPNy0ssQ1zRBvL
3c3dTdK2Hn/9+9ZTirUFSURdB3j6JLAiA8DJrdR9FGeejDa9qkfh9HZ5iSkP/1TU4e3bydIRa88q
oMnlbdVwlMNuxJYZAxRVJVIPD5gkLweF52245wt1BE8pbWD6Ysg1+xV10P8+J540nP+ukgn8Ss8n
jR6yd2fU753IUL3Do5niMFMNr/Yl87jh8iquVRuk8wktNsryuVNHn1RJoiuM48w5i+TlWx106soC
3RjJpcZYSH15FjQMZef9sp60PsAK42904bkWHKrI0TKeXxd8VsLOTX+Z5xRj3BWZfZQ2Ehy94rUY
ZVUj7PKtyd1zIrdZLeu7u0aNepjtRfjl0GePMIwBGZywkDUPfJ0DQpZYJqDW+0MP1/mAu8DHa03F
xNermZFiGq9rIzDmqmyIFapmB5xS+fEAQT+LydXOeDIX3bPQfraXhirmxyycUJg9ObM7Yy3Mv4c/
w70O09NnTrYxGj9J2NEs7Ze/5p5DaqNOQlMYa8y5Ex3E+dZzzWjw9FEDCTbjQ+pEGp58JpMgnfD8
CgUS4lgRkPUzw+CJgL+j5rPzQXO3ZIc8ATgfUhATRMCQUDUd+0IGe6/h523S7d2Ci3JNrNxW4KA1
bCgT0Qq8CFQm0zXOPsBGduYFlSvKAwxwujxJ7LPizoAuGeGH4/mdjtaFdfYEf0gobh8xUrNdVfDx
nG03wKFfVNPZtVdpoowwF0uMH2hVonqXqiGmx6VjvUZ6gccZ7MLNZ96dy8UsWCft015n9/ne0Qas
yQZos+ZMITobQEUfHaII3GtSWgYl4hE/bESGmtJoHG0QLQKlZ4oVXDIzyAR+LarfVlJyF2CRE43k
Gv9X2rRuqALRPiuWetBHAHn0Xg7iU+hK6tgHbwjvD5XF3oeodEY+fDT7GGBCYrKMFnzO5CSe9O7S
+acCwDPz8B4ZTzIKj0eVd/Fbg67r7dh46XkT1c7fnbJNPCoqmu0EEheG7/r/VNjRwC4kp+i+4+U5
JGTzgbOzewPBdVW33a1kXWNbjuMJqVRyZa+HOrWqULJcDRt4ZifialbWjTtKKVMlvpsMYTvEXzn5
9QZqHKEStP5QG7zGAxwoK/3aXPquoJvvb5cE+PRRwN5KKkt97/AurEjnO+SNxmFU4Kav0saAV37C
675spksXytLn+mEvkiIsFa01g5UGtxyEOXdY1SKXOwNFlFqtnzgg7qzEBqvMxOXn+W1ikIHOqQY9
aNpdUHJTKZAFCcihmEIEKhOuBIoZpvvYQLCna4eNi//MEZEzWIFgQzuC9cWc1y6ZziV5arB6at+e
ehK1dM0Fr4beNj7H8Q8ig6vtzjTEh4NTAPhZ6gmoXU7gGNiyQPSL8WUpd2kX4En/328eUV+crPk1
3o/XpvexlOQgN1Gqef/iFWhIqE7Q+n3hAnMYDUnXI7DGD7FmChVHB7OJE8UVnXbo8hg1GZRQJWD2
+xmDm8SmkznBqfKWBLiAF0BdHjePqcx+LI/bXZ2FyudiE0BZY7SAYokxttdJMcIGp+ePc8xM7dpj
56vhYhyUhj0oqHD4xdVdpp98IRkz8NUpvO4jjOawSK3RhuXHB91oabBYLrfgOz1tEjktXZrszK1Q
trUIFTZUKLeVmZgSofi7fAtekV++pJJjIQ3qgKfpdVB0HxiiGG2r3khvjUz0IvnTaltU2l4MTWar
NAxVeVGv7nK6wkHH0suRNIoZBdm4sMAbmMcv+cTLao7Wh6oU5O4T9ucritoZJtJ92GJ7MCqhUJsz
5x27NotfmjEzMc0hNOE7CMYA8z6bC7E47w9RULW0TuC5xX3DYfnNPRmCr0pjlFjuMlYQRlURljr3
YQGJL6cGJFbdy7rMbfS7yHnXr+mn4MaTDIBUJ9e4cHNWn19VZBSQJVQvBvOaxxgFC9YvyuuqhyvL
M7HL/bP7h43FgQjMm1qzGqkdgIPhsrzcLkr4vBscn3eYv0yzFu/OVZzHC7NI74uMdLn39rxw1W+q
0k5N5wb3ckB+/aMFLJNuOWH3mPlgUyOhs1/wzkRrfyYShPPRGAXeKIPiUg9wwrWCa2Wo+4I8pjBN
AqGv+eCMoPL63DX/lZTud7uVRoBotM4P94k5+ySfQUpFzNHJlWJHqtmpF+Y7/kiCsjlamYjKYfUG
1A3x7A7l/oT3jf8iE1XRZqzR1rIqYTffAFL3lW7FWPOCuhM42pXrbUst0ciEPGPlwqTrRbBoDKRB
JoTMJYbUsVWIiz/3w0cJ/V9u6BUDDuidd12AXGgwLs4Ic4O5BpjmXNpEkGRsjJvEEJg+hDZkQO4S
+zDKiUr1wqIONGZjhmiszS0ZvVIerB4tKa4kygfpvjmhSP9IPkHE3KiaTmqhBwtgdrvDeNb7kzEJ
jmo3huBEzuObp2Gn1JBvefeK4hSYzc/djCSu71d8RJ6+OvqdgTm+sxawC4mn5WjSL9jbiUUIJThG
WqeTvFLSzcQA1bAD6ijKzUfzyfgLjlABznPE97EN1Jh4znpZQJTwFu1pNfGFJs9Q/uJ7FlfOkDot
UDNuY9jgwRaFB+UKB2LMTJOFZQlFOXGV+2hF2Wg2J3zxtXdhp2hIC3iWLLl4x2P3hDBY8ymnr3v2
aA7E/DGzqg3PAmdwXJJ/7ZjSKhHKZgPT+k2Fr+FcLs/MAhH6NxizktaDavACTp6vl/FhXyFXNEPn
yPHOkrRfVjSrNJ00b+MTncn73Zvxm1nfCPyA2v7ovh4D1WNYN6b+5UwVIxv5REoL4zXVvaGCyawr
OLQHK6wudnSDNtATnRRjfRQlC1Kv3TrPIVh8yXGwb3v1xSYP8XjzoVZF4D01RbqAiSU6AOO8p8ha
cK4oq0AFgaNo/Ikv31ApGoxU2fRd9/Nv9OhEcAIjpebXEgkcA1rV8PgvnM0yAVEdm8yXZZbs8Oqu
Slgan9nncV/AW9gMcvf9gyzq46mLm3npJOfWBdSOAg70rf/L2JDPrqkxATYrr61wilLpl2RPf1gQ
+R8HPietJMbvjTA4HUvp+khnhNuS5ODr2GiGvFtyhCER8w33iKvggp+w6bpD/eycsFVJU5CmGMwI
fVe8Pg783M5nfMAlADsgWz9UD3Dz4ULjE/Q66pgGTaTL9ZkFDL863/jYOP7BHIZw7zCaE9AWJiRH
I3jAgjZBmopUrH/mks85xrWJeMzMCE8C8DHVhpijBwCYmmOAonyNFMek1yjm2Fjc9iGWQud4Oe6R
1cvcrCKCS/wLG8xpX39Gn+RlkHb1HSCMURj/pUmGRT5lXlb8yyeWQ/sm7Nny8rdjYnqCAamkb9dJ
FcQbIyzJLCxIV4wD8g3getDWjtzQbhZpsgEqfhTwOnkg0wgdaEAMLPW7XR0Wzz1uuUKO3MxSJsvN
cTwkaHEfqK4c+F5KJGOOJYFxs3Hju7/OyNhWViqf9MgEkAFyebIW3WsPIIiX95L7HI3rUjg4shuO
Q2vPzQYuRN9eUdjVhR9MC83yZbZgJAWWLpIRDLUkCvz/093Vs4qTm5zRK/3kfkcyITRdAzalVH2c
d7uWWkwtL7sus2nqxq/JzFkmmjk50KimKD1JDYgt3NrfW328iwBX+vVJI3ti7FjgKn68yjLQd2ap
uBb13cxtCoLAsjzuKwNLOvzOo4wV8Qq/jbuaKSGbtL41fQtG3E2BadqFnvoE0HrIelgR5Kw+zBY5
gBVfuQtKpjFg0XvWYE6PZBDIsyUUn5zEAhBpKBT/yVz0pTQ75H/5IDBYt4dTc+zBmbOMD6Y90RVw
Z8lijPnVr/nF915z8QJqoBpJ7a8JalKWtifPFmnoWnrgiP8rqpyA5QycC1Nc5zb/2iQw6/NiDhcx
8JYeTxAM79c/z1QJiy0T2PvBNe0sUTXRruOkw6170t8DF5CGQiNddnB9pCwcuGO/7+LG9sbkN9UU
iGzW8JNBcrNSUKBR1XhTKTZSUW6bhdPBmCVQ9cuYvB5LKu3vPBYMVajfCwsPcT9Y0lCExKKLa++l
O63ZUvKQJxbxueoqUEQoe7hHEDWi2yp4WcoNkNc7L0IRZmnRVg5KTlBKXz5y7Jo8x1Kgcak9Euhc
zM064Qq2dWMmjecMRG+MxQnldvs1AT0IU2+w/qjMgJucKFlcggJCcUrEu+HG2bpzqp7zy2a+Usra
MsqgGPTQ0seE1AtPUdr6VTYXPmN0ORjdYQsZgSh75DU0RYSHT1yWIYqUfCFw2Vw1ICnOb2qkJwJ1
ZGtmXB3Jqa/nOmbAlZ9NX+58tSc2CH0n65XfLnb133TBrcTLzD3iJt0k3wN7TPQClLORj1nAVvpF
zLyAJ3llhJJRxBuzCWa0e+9aFWwUAJd5bzOuESaPEq8aShX/+ioZlv0C4katgPZWxhv+EwMqVs9x
wq0gSgsC8LALo0Uvg5c4+B0dMKU/+JMw/eAcXDQDyYTbbesnTDk5NOPHFuerjfWLk/bohxg7fS05
K8aR14IsFp2oNXQ3bDTTgkuUPep6rS78PQ8w7XFwuoi2hJdsBLAgwHLY3NwmniDNcR2uPyav/Dgh
lnu+hzdjEKJOn1S+lmYRHUTL/ejZH6w0mwEenlWv/GLin3HXU9IFErVxuUX2G8zaisq7zeHKmDRf
zCIii+GYY4BDjZbUqZzxlYyeobFwARm3jzHpmNFNibQq3ExeoRM2mywT4xf350ojRINJSpc4f+Qg
cGOHHfoxTRNBjnAy4xgDUS59rRwIBZB6Wx21JZx8Q1vT2Z5Pc0M0q6BKTLXUXnu36KkeUuH9eWx4
d+z2azZJMrnGQ4ZeUQnvVwl9zdqyuqbAYDSaJ6ZKb8eCbZuxNIdcYsZ4flStUL19ZSv5eCc4CRQC
Bvg+pupAzUc4Jcs5wkvYdl843LklTJZQlOCWhjNKRGmCX23qKAQRLPuF7Nb/dlO/L3Uia92IRb1O
fJ1gRQm4QevVgrx6kie+gh/++ypPA7ipTOnYJWNP8FfllYDUE3PMPktlEo4AOOjM6Df08ohUWr1g
bv+MKo4h9wixFgCLKL6NcBi+vtdJ6LYFGJFpzrxtSYiwv369yu2YPGawARL9eKLip2YbZcBJjqF4
xb195JuvhwpccZXcx8+SuWiktvCV90+db3z1J1Nnf8RjAWUN8xCvNb3eGHgFpOgNKDquLz2npm/F
WdDL0ZHkefcVwmq0r56XxTWnWRJlaeqGKWqb9u1x9zthr6h/Rsx6TIRJ1p2v3LAL2YKsHGBBeaX+
VSUf7Ce3skeGKNQ+Cnc7sl8BksJMRh+uLCK4tt3FeY1SASOPnEiu1D625ctLyHBnvIMBixpoA+of
WwZlocN+VV9hUBCjT3TWOIrMg2uVSh156GVAJupBuapwSKrGlrm/0As/3Ge0oEo2g6meQeDBao0Z
GsFkO7X9ub98VSdtjNcQLRBAhAH3DJPkVse+eBQeyW5ApaCdBA3ekPwLxiESGHZzq41Gg1yYybJ+
H0ST0BEpXLDv/cOK4frcBT2S66wkg2wuuZIADMGw1JwpGM8QFwZOXF5IIZ/MQXGyO22wirh4vrfw
oJKxh8y2cbr1ExnhxIYU3xEVdgbpYsMurqZfD0pSvdorpWjoOIKZHEXFL64ryE+IOQdhzQoJMYvB
Z6vxEr6dYJhBfhuvgsLriPjwGLnmSuG2Yg6n/nycfB7RAXJoTLbXS/WPX+/aWFVk8eZHd8jMFwya
RHckur+K/vS3Z7Ggdf3cnnY0vmdBqIxFOf0MssQHCMrbiUJJbaPO1HNM+zcGXFZt3k6/0ZRYtJwH
e1+OjxYYNYmkCG3kTXecbFUyL/htFbvAihi9inY3hLf5qMxsMegT03zf2V1FTLXQ9dF8zBSJqXQA
4J0vxFwi7u1ZL4Agf+qrY/QanIiIWixk7XxU98rATflko83aiSn9NCdTGutW6B+tDLkO/vpfnpzH
CO3voIwuU3dw6SZck4Lib9OK+gxaYemtxyGLJJd1LqyzqF6jR9riHlLqHJNm5SPmTYKSvPb/yOBM
rzWbYhfD+2WueoZfMKXRyxZTECqNdyeLlOAu3mb0V7HHFbcuYoHdGZhhqn13HYWI3beBpXc9YneM
b0m7GAQfad/K/PUWtLv/wXtwHHPT8s+/oRkky/iJQWlhvFInL2KFBcApBrXsULSoa1cFE4Jg2FAu
+MTMFHOXLmX/d10QMu1f5uM1NLjEdHycH3zagrKN1rMJb3Z8fqLd6Gl5RhSvOXY2roq5kzdj5Ydp
9c+/gbSuPDnuN8LZk0iwGQcrzQeo+wFOVMG9K6Bgn7/M2Ky3vb00tTDolS8zSjQuisQoXhWr8bGZ
5BBbDogiHXMIsOEN8EP4UA3Pnq4OhWTjyNiN5lJUihZSVeKVTA0iz//xsvmWO+OXBnPNwwX3anDB
MY1sSTvXn35/671RhlVglVa8Xv9Gk0W1v3b+6m1kx2rvWxxAX9dJ4HwQONyZKWUM3t/4cv2mxRmR
oqCKqP8QA5k96lJ0C36x30dWHZaXGZjJxikm5dDXFIxLMWKEl/VsgY0tgkMht6Rv4nlYbfqWdn+K
UyLjDkWEuug8KYtv8E+d2dNfsw4ftrYNlkSnhGrsfvhSg61Xe4Z/ilBL0xROVrOSPbB5PMtdIGR0
zsdnIwZYNktsK04P+KU1WC6neuOkmESLMx2rqH5369HzFCJjiH1lfA5yb4I7sAfIeIoihSVlZS6/
bWls6Unh2Y9YzavNHj4pLT0L/J4dZM5VY+0pke68WTCcS2xum4YFLDQHWU6xIXgw8U8ud8MyHe3T
xdrdKPxLAWWr/kwQmKDjj7mYYjAPL42v5MEJ5QG8EkgoPkAMVKplHZ2LF/FsUXIoTwc+VnRDFPqC
pJxLn6PNxks0bMB6ieaYMoyWOZT9ycXZfCJhHbplOU83pm867o12uVDZjWi9S+YLD/z3y+SGGMsg
UAhrDDv1VDm2eiJ7hGQzldqJdvuDyoEl6sSzVYGkAk2Kbht/8TkbDG+MZv4PAoLJ2sM3zPDXEajg
MkqVGI5ucvq8/jy6ffunCzxC7mKMsLCwca1jD8FQM8u7ENvFG7+aUEaT8LkHQdHhIgmxmF+x+S6C
1dWv+f64hvux48pWk5O8kFP8GP5XAcO7D+Z3UBEc4+bkWmPPY1m9XPwlsrd5rOCCTHx6Fv0QOV/c
6GHmd2s4mHW/htKgYI3EVMd1qwGGZYbgqpN1254hfpqF0wEIp4pVgQC9RAQENP2XLDC+SCApcEyW
iOXbZrDIVDExtovrgMiuG3VqGmaDF/W15YEJvVfJC5T5badYkihdEL2NbJBiKXMGfhEu6l4f92cg
X5p8RTLZEOgGaNhVwDTGR165w1k5kyer207eqo1xsqudoDMk32RXnmd9hY5pUv4JyK17GHRZdMYF
vwIm++mkh+WuJKkgmVYCqdT8IQGF6bZMEBoTGVaPrTjbympP3CwwF7eM/GLmVXeJY1S6cphF3yLg
WA/7r+TFW+rStCYm6xGhD6JLe9CUY9b1IImh1aT3bL7lG6EpGArQUDy/97lT3edSPuBiDlA/6tz5
o/6EN/eB2BlSrg53NbX7891Z8wiGVVnxAs1GVq853wIeFYerl0hThz5uoo3F8LOCqR/heold8be7
P/YjxBEk9+OCpXg3TR81A24Znvh6R3Faat4HHU34P3oCsFNMay79Ucn++ckzL14B9Od557bnpUIm
SI2mdFvB8eSM+m8oMIMX0GtmgxxG4ILJNWQcScBHHTfhnoXjYcg589WkpW/0aE8T4bT9PrMfFdDS
eQ6gNkYptV/nxwt1/j6BYfdOlqOiiVfoyJC4FCriF+/sTjtigZiAXsYqizYXFMkuDKigq7Q9xM21
KkNSuZ3CECumjdoO+t3hSb+vNG+nHJVpAcq4Ln8QScP9oQKXD09k1wCKotINrf6GTKnmxYUxgbfo
WoQJutR7PA4jE5GIPO4ACNZwT2WB2dwgQJyvYcbuRFTOhkQa81ZN4DJGqGVD8ZjP5BbJpQ/zU/bo
V8GvgjiN5enOTi77RgBerdrEJsWwDFCwdpz+MKRqFKVCe/whI7j3pT3VejxS4FroiJ5fNpHinXDu
fPiTm3pvjsPlF9towkXG2XVSCW/gmle1nXZ2HzTqbMvkUzWnq6LQopuIu6O+X8ShhLXFmrqqehXJ
VGY9/eO41EkcfMP6yCpIz3uWYyJULPjXcZ9Z9s2pMbO33zPfAQirOBjesIKZQgXWarbkJ7R0aWZA
rRnfQAbazmg0ouqcImOHFtPDFNye46OwnFJHeNWsl5NR7tjqC+YVmlend/E5q5ZL3O/wHdp0fqYB
SLhqHe1uS3slmwC0t2w9Zpp1NUz8k+Z9xwE2MpdK4ayukOBO44eKKyAxN1yEFjO3WkbLXXoB8PPA
FVE1SjoOhX0mRR7Jx4G3LRqOgFlaM7Ix1Ne6FdwPfO2RxcJAAPpjNHSZW0aBe92YoQmDQoxEXiao
sklrhI1JBdyi74gULlwYK6NKw9u0BXOkRYbXaPm76aITsyoVwkqWFvnBeS/wgP9XDkpzlTtHU02E
mXaybiAeuwiWmeouYHoLTtCtdoj7JI8txXAHlOfsYu7XHeWCTmfI82Oq9oE3u3V4XdnNgN9+c93X
6Sy0/DFkeaYstIXg6lXO5aVbHHOdvv5fgfPE/mKuiYojhZoJ++S8fL8liWjpNvpAkLvOhLaVC7eg
MKlZQbZibT3KeASDlSycI8ZwoLH8EHsTZLNf7CLEQ2rpW0Hcka6wBX8iPqYCk1AMAMbZ+Z0UswiR
tzNzhevzz6IBgj/R9I3KydrxRmpFfC1br/mVWbYZWqM9Npld689ex2mORpicjdguQ+sh1TZNom8O
yLWQAAhfrPZ86lpYG8qqOyiWYd+qEPbRRLMIcna+jexHkgDz2wIK1UeDbu0IzH/d6K0rYMhvlSlK
PyEO4AdysAHTzPJ0REdtgKC25ZQGit35EBwA/lLxzkgDkNiwoYDYfSN5xAENN19ArlE3wZoelQ0H
dI8rRd2BHoO4LYchkDjYGDC0Mg2i6yYUzndC8O6KVAz+7Mtx6ZSev8d9syEEz2fGWnN4FBvDgI6Q
+JikBEWQb5JZ+3iB19xIlwqF245uJfSvhMsc0MD9ItzK/Rq7I1JpJ/IECBLo1yaR2/1mIMvDSbnZ
PTm6InnFgUCtPQyOm9Ot+speG1qd34IyobWvCH0HQbLSHs7bbDDQHtK0DlvrRKZel+XoIv7qhMV/
HbduxJyu+cKV0p5zOee5tdaAv+R2/SM4+8wxcwRPBhHOxj32txUdQgnBQy80FXaecfY5p4jLzGTb
zBp4ff7HzofGX9iHF2dSO+SjfGTPIc7cuDqfIdT7Zrh3i+fAYSZ1yXMC8ifwpoVrD7m3F4HDxrnB
QwEcNKTboIcDAJkxTdUe/N7R61B68/p0g8/yPKpf/3CQJi4KnHZ1kFNOC7EE6h/J1mBSutIP8OV1
6wGaoedSSJaPghV0DkffHt6Z5lFv5Bjj1jqFnm1C9BgYWc9Vq6IEjtU2l7ngcFdqgZhgDo03yQ7D
2rtZaunKrQFMRkAoTXT4xakG7J3PBpRq43e/okQLEUMvDISfrhjbKJ8qymB8zaD294PM+6Dt71wG
JtdjHA5FljaMWDPmZr3XQOWzVgtNYaRlnRDFHDyRMigaUrB4QET9a+LqJsb9wRdW0K4L2fmrGAGw
YG5rLQkLwFWhcCSTanW8PwI5tX4AWOCNFpxdChiBzA8aAFVgzuQJLgfVKN2dHcr8ET2o3fh1KR6Q
OCaEuZyKLjAJOHGu6Y5wlnC5cMjyisPZpecJcYtelugJ/PeN8NdracQhCnG1P10w6FuVeWIJVbIU
REEg4K98W9tE3Cm8WGGDBjfyQEGHfTtlM9SIB8Ab5Men4rR4ntUfQbkC58u6Wx40SQLOjbfhCFnv
fOkb4Rd8Dvuk5uBo5QWPW1NQV7CaPc4C9djP616n3WGN9b0Ks7EMjVI0E/2b8bJlmjWBJmbgmZED
cN+pKSq37lk8QK74oZjUj09GZ+b5P7CYpWEvXUKmwfuePqXhmAC7pq/8zto1ESTqwdWMTQJgG9iH
i/+KRS8L69Nj9Pf8Gu0KHukYC6g8G75bh0Q0Rt4mD1hy9FYw1cYskyTSiYOFhCEzXt7i/V5tB3Lq
E33+wmQPDLPgj9mWmWIJ/ehpheMXFkuiRKu6StCvHvCKNUn7pjfHVmGvL6kNrG5Jedf544iR5Gvf
xxvcFytuzMcz5bzpB4so3GQCdO1vlATqG9WuoQIlWTZW81bYfyOAVI5C4D/QtO2WbsWbtvrlO/8H
FMseizdSFxUlpDI2fnEyGfeSgpf/DAzYTcmPV5jFp9CjAfA0xGlVBK0itKyY9W3h0TN/Y9ff3NpC
3J0FwiaVv0YQ9iflo8jfdh+eOao8zaueH6HPyn6IBGn6DAAU5XnCsIVORCNruSCbE6eU8r3A1lLU
yOWwNZFzTsMKeDBS5IGHDhRinaPaPdCfktqbVh+U8nA5KF5v44vF0w+/R2HtfVDKYG5npO6OChkO
OlsHH6wyyyXxuiSvFbwNj3qL5tPr4qDRF7NXFhNa/T+5s7fbeDosrOP7HaNWOwEQDNQxtcd0giCG
BEse+HPPEFeiYlptGUdWbFloKYNOAPDvOMKL6aSeCvQkrvAL6CzBWdUT9DZf93V5r79wdcU56OEx
ipZBxcd+jNSIxYVkH++Dh+jM5cj/fs8kc51zlhrd82AzPa3+Yr7M1i3BKjrUcdQrukhZYOww8K+r
uA2HnWbOT3o6eihoNJCDlUkqnqH6nRpwe49Ja4GjybaJcuh0r8lqbTk0yIsdg4ej8WwQVlH2oN3N
kCK3mPexz/rVkKjL+JkC5GQR80S28qLVH+kOhUMvXz+OfMRAe6B91TSWc7r8ZQlLvDkCb9pArzIt
pN3oOIdqRECwMtYax0sGhSLeyIeWHnSOPp8GUJ1vo/NL/lOHxH5ZhfQdZRoECyXIwhym0EVbL6Gz
L9P/8p4FRFZsA+XOxUUjwQamzVcaFsCB9gbZ2Xzl5xYLpWSYLjVm8UCPsYSfmHfrn9oZbPJDhU0f
C4iN+ttaM3J8A9aQpkBJHGiW/uEBPUR0gIsI53DjXMl5wushpe86c6OkCY7LZq/OxzkzA7thf+l4
nJfnOjynmlOpqQ04gcCUX6z0ix/Yis3RWlGG7n/AP8h8YIja8VmhbpeskhqXYAjadGYZFozScng/
oUMb0OtoLgH3GPSzj5s6WChvzol6OEtIbc3aUkH6ykb9oMkjDv4TbXzmZFDAwLDRyKQZoPtE43Cy
9QDNvvDsxxQ43hczF9psPB3kZl1yPDzPZ2lWSAqZ1SpTNMXWJA4kTxgcDaFIWwvRknVhjgX/iXv6
fcKw+dYwflxdVCCmfL5fphw3OT7DZ43hARjyQc+DyXf+xL5L4tQ4PAvAmbbKbTGumtXSw6dHQ+yL
RbBBzGfP8tvlVMJmZXipjQ5D8Fnxm/+sWJdP7jDL8ATnZEyzdlFHcbj5tiM5V0PD2sTx7VNHiNf1
iqQBYl9L111EbA4hsSN8EUGSVURekD9LragS9upPvTpGtxiY//VWI6F68wGVoECpHtgbOJr1ndoM
K2+iDL/hl19zcoZdjOy/SHc1qsZ9vbMpZ42Vhp2Ar3g39cDHSAfsQrkuca/iT3415kjZTyMoPEg6
80H1+OvnMT69e/XGRP1J41C5Nzun0fURsQvflXVKz8z0sBQRdmp7USaxdXj/X5Q0T+XTVW2a+NHB
PXLhGPzyw5FRzIiB5yacl+YWHiMDopRCN3aQweFQXLxNttQNmiCTq6TwTxZ18YciFsTQOzF2kMbE
U6l0+ZaI3/FIYQWZLouv8UoDcR7t57ZfPHv3tBPpxiYbjvfhf3osnN+rstyYrmB4WYarc2gmMC9H
nEr+iFWh3ASfA/TEWKoVByInh9m8Sw8+0vPpnPekHnnlXyI2N8oauhLJ3ik/LvXbWkFIA8aWhSAM
a1XMxLvj25UAyk1SyvBe7S072XT4QZT7jpCRZ/QiJ/q7bzXKwfte/J5UpW+/0B3OJidi24VdnRRA
I9tqioK1mICmaCzyWthja+SHeii0dr9t4z9rlDT8zjh0Y7+41QBxlsI8Q2TSjdq7i8aK9l9WdKKN
SORsaDekKOYcr06RRELfvp6V+AgN4to/+cOT2QH4+l+3p1ZrRAYl5YMohRJneiHPzD+CXFRB64aq
aHMyJh4IGilOmdpNG1dU8O4Pp8W1lzkrRLVRv7K5rUSyvI3YUimfzRmQHgvzf6MXJJ4tFCbexjrR
n6vss/NCYd8DXevwAhVwFumWYNv95tB61Z9QdWN3bknPoKFgqFi8sDBlscsxiHE5ph0FHAqmDUO7
Ag6YBt1fZ57wHWZTkcm/B9g6+rAiaYbdqhlTZ+2ChNqWazTZvNndiz2YyWmSE7y9MOD+u+NXTOF9
yw5/Cwh17OBz9Fj5jRpApJlgAX5PjDnGWtF6oD4RRdEZ7BGqGajxS0D+/6jn06t9vmTl0WQ+Q5qX
LgufnChB6FQDtyH6iLn4qdvdUrzjhJItMyJqWO3k7SsEUGBsYtICZDHwCLAyxLkAziZGOcaNfXBk
MZXeM+2wknznjItg3CSEBxlkvJOhaF/LA16KlHXWsAPU8NNHp3c1L5GrPlZI8r8wln9aQj4fsvRi
/qHVv8YX/VsQh15o99IVq/hzKw5hZSxFJqs/uVxDRrYAOtRwGDktn6r3/BIZb9kyD/qDbgVeXrNq
STSjadhr7aNqLakOtnDuNjze/sv9B+J5NT/DteCgXgUab6hA30vySdGZv72VW4p+g4qujLmOE5as
9TmJ6uVhg+YOCWcQeOmYzlduDP51ff/tuZsVWaclAbdwYXzY373sNdbPnP29QwpCdHTHvzRgMD3Z
nMQc2hVPwYQKHIvcLEYHcE8xjyF2zdR09APtM8IUUxXUp9npDjGEEASg1rmAmufhusjHQFvf0S0a
m+8+0h05R0A9naYAeU1BsBeiFa7FTaOs58IUu0fBK74LZXDKXu9PT9b7NAmdvwQ3APkqk5VhDASV
ImLpm6h4Z+UDcmyPi8Rp4teq16HNQkMaKuaCCd6biWRVtE/oGqpDc+otpSF40jvMuRS4VGj1LzR9
Q1J3czoIYBc+u69J9ofRgI1rikj7RTm4IfSR5p80jtAczwuK46X3/9O5ucqynlGx1Y/5CBAgA4Bd
rvXjWt9ZmiE9qVpSWmIVs/xPNBt/UOkhVznAVLSa2hmb0kycqMD7ZOglJGjnFL12Z66Lip24V1r+
UDfjnx9VBlx0xA3fjk9FGziGeyJYbc4OKFq7i1GimN4GWl1L7xpX+LaHzY0E3myAiXnZKZBO5xWb
WJ88IKJZAocSw0WR1onzHwzR2lbI689aUw0kaRF0REujIW//zcIukSFCEpWXrPDJIET5XAGroiCx
qQYAocmEOvEYO3rj+rWPGzS53sFAEGOmzs0kMl/OinWsny53F7THCfqQhDB/KjJAjxRqrvUCHQtm
tyDvEM6G2FN2hmOgSm76MiHCJ8vz5v7ZNSQFXvCRchwxjofEyiw/4IJRH1GgUrMHkHphY+jGhrHT
a0t+2IzD0hg9qkNe6c5VCZDLa7Z9fDITb9N9W4yidFAA4xFIntsJ3EZRRJZQOQaNntRRGBHruzG+
qxzRteIHHFeygwDESRjUHX8HQOGT6kHmntmLnKL5qHkOvWx7+nc5Xr5YYvkJZYoYoW0zlDGvhyqo
VmmZpe+5D9HL3Xx2zAHieoTSch/0Hv7g7GcpBG5Dus2PUJBJv9IFPkzKWNT1QDjOGw3G5rAjG4Wu
DvA1YqIdOuqAhuZ8mpuxV5iDEhRS4/LNvYMftDdDUkPLW0mGr9ycHdmb2HFztMHXNWOD1Rr0Zw9D
ql6a0zHT7A2nk9un8IaqLSW0Mtte3c0LOTmoPLaKwyxuvsVbS33ugJaVqJuZ5lnC5ssJddULvmXO
9fO10b/5myVLTjwOcQU1CzCqKM2yPjYIJVplQiiQ5WiDYtC1Y348rcWuUSodxNXeSmn3sd3LUVrk
ly3IbFmID1sztIsTgVFfcrOM/qNXBHDSnQTvy0/o8u+uHDzMLTr4dhH5mOsrSfWMcEAu7wMr4I9P
6kBd4HInltDncq8CgjyZnQ1N6rouxgSPfH2CYLiKdWKDqeYQarXUC4CsaQPXqXUFcMuFnXzwxLVA
a/6z6zH/RJZubh4kD6Y7wA8qZ0//6IHEkXfrQXmKSApOJtNS4W144CkgK9X0h6fLlDCXbB5mw05P
DjqhfeTZXXphfJneE68AC7Zo9nSycLY5ey8R8ZCpk8L24HGii7D04nKUCaLANDbV6oQmsC6qmKEf
Loubzw//2UR1txBKTZiY588pYB42WpD924UUa7y1AsPuft6SStm7EOeGSUZTU+ksdI7Rmni1tlkg
mwy07ViyQV7HStX1SS/gon7ihAQBrSg6V/vTScRyduSO7mMvTtXdLTYHbP5UKvXdsN6gLMG/miS4
toYycYQX4I8BisnpsxNo0lomFslaCOPayTpDJjrA7viIO+I1aKargtPskuO40oUxYoqeG0GAWt52
oPk+JgbUkCBAK7TsOX9FrdnYx5+KAUQz3RKi9/FjPBhms6yokaf+VucUVn3FcFN7d/UkEuatmNrw
DYaPyJpcDt4C+2Sy8jIk69IVhm3fBJPivUgdbmxbNRbFSLeVtzp/Fe1YWCoAEtfJFntz6w5nIeDT
jUlF+S4ybfyoX4umuIo73XQ2MIDMJvZWvl6PiOtsnuA9w6Yj+T54FhCHWDRTw036ChVOdnNJV7of
yF6TIxnjr7B1NKoMDY3lqE4iGTllm7VqhjUYs1gqjex2AU85xLMusznLmRUuO7Pkz+uBR7+tVdqh
mRBFJb/xC7/fZBfCv0KBp/MH3V/Sm1ctNCM3aBosSgm2h7Apd5qyywxHA7rH4Uh5ScQCVp58XdJo
K6M+ZVUkrABu1ZKkH5RcP/C9W1R2izC1c1/UAIXKtmYddie748htbpt1Nh44aIUbSaK1dJJO1GMX
pv/V2oaMIoI/c+wqIdxrbanjQO/GahweyI7ckDQHoOaM06hP0aWgxMJIFq5IAlpfON5M9Pr13rX3
rDyaaLjxp3rGZYz+R82vXNK2PKDeykPatEdBOxWo1bNxkd3HVvl+ahYtm1OOLJiCPe2mA3F2Flbe
e+mlomw6dg60zMmMnHl1JH+GWxg97in/HqQ+XYLxrfKwS7QnjAINKkkd88Pb02d/vfw3DkkkIBJF
A9R/MRPdjPHWczuQ2k4YYZX4L3J16JKdHOL4YnvqEs9swb9hebX/gGI9qjgUfvPOOXFY+jshb0Kh
jrMm7ieC3XiOFy2Q1j3SmYZaKLxa2eHjPjB4ULKYH2JH2pmAfO+fuKdr0i9ctiCoFlYNawfP661d
usAqLbOl0L73gqXEVgWFCFRKPmG5yVGFvUzS1xp+ucsrwV2Tnj84VcD0YCmZK37yckWbjR0sY5uB
ZMg+fXTRbWzxhVAqYvg4reLq6JlxAyG7pHErEzqM3giTJTywIYmcLJ5UatdVvcPyJzkvTDhZnwc4
upzQvN7ZlYBRrGLJBEXTRFNBX16uy79IqVH8oD0m4N4mVRjFZs58HOtmD/gS+OYwE6EVovvBn7+l
4B/5duH7GVn+HxYaoZ86qNvLcDpfbYqLOhTq8XgCVmRryxtxCJSZTe52TIZr/SuwXXkUmP3u2aFb
rUObW2l4vK29baD9m0MD6/FiwMOYK03lXgaUCZgD9ZTgHFJBa+YyAANCuMfaiXv39UvWgglOtuHd
VKVGAezn1GcFfRSkVnG0zw/KTCSl4cpV955VHpDDkXgB3b8zP/Rr+hYoYk/E7WgHi+5Mb6dkMdIw
oy4r+lMXg40lKZm/yosCytk5krNd9OWX1HhN9+ZuIgwibC3OgeGRnRmmYJGqYfHkMyYBBbEbLNNK
pGEa9EkjJiVQ4gpFk/3vfAq2NEdlesM8N3oopxYmAdnAFZLNAaQlfwwyI+YfsLtpbPAff6fUfBr5
PkKg3W7v77plhu2fo3VnvVd8QdVlj5Tbvkz0O88Dd7GRSz4dYTe91QZ55JcYk0VzJFxmr0o4w876
iRaDwXKpOGW+o4U3p+Ia5TZPRDHKtvQlhYyQsQ1mYMXJV7VbwqlC9qziZyPZ0Agg1XsDiqeXtOJs
ojaMUuiui/7DBqQKnANeJt5KSvHRt7/ySLBa/mgrkLulnPMgzTdvxGVmTB6ucZUPsZRReUpAHWEG
7InK6zesrRh8DdKqj8E4PxdCjEzEhFRpzgpIrUG8NeI7DVoLbMzuWJKPRB1LAAWbsuinFCkkJE/e
M149pWU5iSadd3DIubWkEeSYF+fR1K77p0vr5Jp2TjhcN6jSx2YberMHR2h/6jOPwLqSZIcqd9IO
lyY/EbGgEEr3mAUkXe2pZSYzkqF3K9eSEzroyEuOFyhrRO3q6hkvU4S3VVlZie+wdgHHiCIqMKU5
lqHBjs00Zkj+bT7BgpeYxozEKd1BzQ4m52/txxBQrfIQuZAm6pIJHJ7CvXMvTcbpvRYP0AgpWRnA
uolycj29LfrZu98/87AMSITE9efgeBwlHugOUrbySqhNpvdy859LTHmfrVelo8Zn7NdLCnpj4kNZ
a77XHoZoP60mgrWMvoNDzm3TWq6e/bvlH2n+z+ILd634NW/fZW5k9YsHz1e5oY6A3nd0+AA6pAUa
saqXbXPHPEDQuo5AjSP3ebhKe5w7W46lm0sax40dfJug1PP5eB6LB01YtGur73f7b2UJaN9IqDep
AXR0gyYQYiNXuE8rMYTLVhELessmggdiKeTis0xFnJj0eZMXaB4BNE8PRt3N2d9LpmrH6Gw4C5yR
QQkj5Unbd9nfrxyCkp9Cc/aDQSM+WUA1xX0OIUrNcKAvs9RF7TaQKRVoGQ0CIGFKcJI6ajaolfHo
vb3MGkHuVOXRcMgJyj02l9YY16FlVLoK1PGWFhzKYjGSnts+hw8Jy3dLKn9QThZTQD7rHM+Pnbe6
aHGV1RtBKzrzPvrPj6KQlHxSGp9iDLklvRMTpM5yhdsPqBPVdBMa9zVUyLagp+Sx+VKOPjCeNX7M
PK2CTQHmzab1V1NTQTFa+LAMjtarSoJXqRGN21nhTJzq1FPL5MTQv+ncLkxZMIBkwnv4sk9IFaxf
4u9LcC5u90VHFN8HLynMhiaixUC9ke4O+jDdQCOT+zP4drWTKBhge9htVM0Yxlv2tF1aS+fi1scN
aH+QP/asd/obRnatOvEPJFEL5Fngpu2QvdHNgKoO6hNF4pBYXntz2GdoPxGTkC/PHyLuBgLpVQ/H
sVg04Qx7q5nyfBlUPj8JGOGIfqI9amV2s81xpY397MxCZfrQcCRdSxbmV2hf7skYtl1HjweIUTgH
eU6ntYutS4qRIhpVp39aHdqXqp6Jdc8fz4uRzrERLNqOu9u23sQ79QaSLD4TW75CUBLeEnJyE/EK
wO0UbFF7dpnsrpsJ54RuEc3B2Fk4VJns8e9FQxYRI7hnQJylAQgO8XZ1iwFaZfptv5+RoKf3jGXl
T4cY1JBEjj0PnUCZUBWeaOwUDO7hmalBy+G8XIQ4r0qIMxDBJoxwtAw4jeWNsx9K0dJMP6WGfEqa
dZHuBU5siCy6ZAdGw4ofAnWRZHgCLQXJNTCgX8i70nNLnTP3gRZmJc8L5nw0FAEknx6rGzicCuZJ
XpJ/Nuh5TgcLT+DR4BCamZB/i6AZ6U0aHpNhmdjd1606VCbpuQ2cP+hJRPF3qebZb2yKLtVbDsz/
Af/DZFKHhB0nBYLOSZAo4L2HbjOtwvjaKB8PhW6YkFYazBLnjym3KNAcYa6Xv/0inpE2L0borMOc
E701LJfDb6faoA3ypqa4Hx/pEAQ7pf2RRcU6IhxzcZsvAq1JuMk/04PiSta9gqcYYvCnZ4cjzspO
oyWVWBFHPQ+rDbh4eo5xBTsQ90+VPEcr6j7jI50Y2VjaZyHTO3UQJmNbyWGMV6G4vGTSxpReHRQA
AQQkNm8g5kKPadIAZy0xOkTCUOYU7hrLflQ6EPAXumwrt7/UD63ofWOn/tb8ESfpd6sIp/Kj0Sch
rmR9wDezCRLQr/rUD8yJgdKxuG3TkXRoXEQVTPVxg/ormWqQkgsuQ3JGAXn6PAeCevaY8MMG9J+4
g0L1MgTbNPIIySU9uDyDRgIQx6klw+AX7x6YHaU2wSsKjDb3XL7lmzwaIuHrXbXqRmq33Fxyx5nR
fDiXh94OCfwmHk6PVe0cuK7CrRqFvg8g9i918pds4EGI8DYehdwgCQHqeMjXZCwYWMCU3/A/2HH2
KWmZD98vBMJGmC5bE4vLR4Qlo/vGvN7pNQwM2J/l/Hi3D1EStgjSsU9Rg2Z3RFo05JREte1D8x4w
eKLAAPiZtQxGnEwVXG5mwWeJIPVgoT8jqRAuM8LDqbeYV/BzouDO6dEk4pIgevniawIrb1quC+O6
kVFJxw6vutjLzZLs5FdaMIoeS1nTNi9agPpmmexqG443HZnVpOki21jEB3AhlOS8Aa1nwObTgjp6
evdg7zN8Y5GFhB1CZx0S7XhxtZMI1DTOF34oLXnQ8e2UIQT9A+30jXukvJPyGQUmod8fIhxxpdBS
bMbzdcO0EkDlW/MBI38gcdksew71QD+dn4sNbL5z3AvNJWZXnyMjxuVLR3Ly/tRCiFaN37vZVqjr
DX2y5u+CW8vwNLV+/VRQiMVyTGd5IlR4XbhMC5+mDzshf1GgZcI1njNdAfaV77bEcXr8blEKCgTR
7YpfLB9NpYbBIpSbOwbuMfSJTI7ozWTUvagLFVNl7ZVtb3zRWXww3gumqcBACLXAzJrk3Di4Gmd/
pPyGQXQBwBAQ17HOzItzGYPCN92IVa1pTrAqjfN9P7ArxC+DScOs8vkq2qehbil4wY6tM7Rj7kHX
lYZlsw5bapMDUgPQR1r19NlUBypDkxsn27n/CSE0kD8IxNB4ctIpSZgsZ2KtNFjfIpRwKENYEJAG
ITzQ7B5aDS2wjlT4BUa3o4h34GlPyvLwi+Y0KO2pn4p/hwU2o6U9j/46cHiKYyC9j7V507W2o1eT
4yakSbMY+IvI4OYxLHhQtiSXZxltjn9ZVZGWPsPeadbue3DGQkodI3fjalNDHzupsF8vPTjTz9vt
mh5xWuLcWb9tZh350Hq6OUiBNzRsSlQo6N29z6hrNLTG2ge7dbyXOvNd/uk1/iLH08Zbv9JXNJuo
0DOZZPX6JDfV1nW9x+XmRMq+uiRlE75MS9wqS7K5pvowP935IorQpSZbKmbHD9adylpEk5w4P0tV
FF+h9IYyIVlr4hQ+4BHjyux8PM8U+WkZzzfD9quxKpp9rOt/Jm70YrHFmhFhHfxv6bssm+j2Lu9t
wC5vr1wPO88FOBQn5X4dBZej9TCCpfoXlvnlhyWHRfHxS4AuV/MYHvXJ2q9ONqMK76EwyhGvdJEe
4FKDSBSwsbU/Kzc2iwPgFhsEumeioygr7+FIAqgvqT83l8/p+rmMUTHm2CmkGOWLd+lAS71oZmiD
MIg8iuyZ3wlxqW2iePq0/dR/F7wMK5cmdaTdM4IjY28E/eFjcFvX2xQcMN8Xh2dI4Vd3C0Rjqzwo
LdFhRQMiiPfypJH/lCnd22vG3p+9ZPIQF7iRVPbSzogg98MEWTdozEzgzJozuTto+JpHJhfEeNin
aPiQ51iAVZINKAYhBAd+b5XHBoFud7wETh6KF84Ss9pcVZk7FllBN0qiX9Oa3nVii2+iedFo30XY
Cf8irn+WGw/f8n1mV7IkYNTA8/TSsQuM9WOL9QyUgcRBXyBj0xKSL9CXF0uy1qpnXZ3/b+O/iJoO
T5Izha3iWkGsKipYK3Z8o3J/6BtTwAFV6Cwn74gvhdvQ68tzqd5d3ClMLcA6lc6KUmUYTDVOo6Y2
y7g75JmVPkzqt3mqbH5XIj2xo8/r6FAfaug4UCReg3uc5w/Hmovtve23lJufmcqwMxiorQ27vXCu
zZOq6qEP04UMcehadQcOsjcIrvHYmDZqMXJKWKwoCzVrzcv8ixePnDS/H9mhWki2ECAueWfUdMTW
Cw/YxzfAkBPFDpjugunEuZK3dMQVtjXRUlVirA8vXb7029sWaL4bg/eAl2xuuI7B78Bzr654oykt
wmqjiVKMG1wZ/6Y9RBn2nQrAs0ymN9VCWzK34sT2cU2hmmgg1SwIx9i5hXssQ8fREuwP5zj8SdLv
/42Aiil503DmHUoGfM+wHOCKV48BUSLie+znJXKe6bRGFN2sVFqycIMVpfNtAUE6yqr6bjvZsj/D
s3+DxN2aMu8YDK8+WF5SohWzYMMJP6jlXP3jp3r4QFk+Vq206tynLkdEeP+MkCGgi0ic9Z/xTZEj
kW2DcpMHkMvN7vMMt/cb4yAgECsaii85D+w8snF8eqT+sm9p3mjfZ5ZJKWqP00Mdvlf6gv+ZJhUA
REkKMRvU+oHcf/NOpGSUsmSP/QiahoCk4o63V0I5KgA3oEyO+0VdFyhUGzPZO5s+obT0fNGcy4BX
IWuVJwiQxSCsvVKKs4ouBo6pCY1k+vWH42K5HxlSnXuDHBlWru0MLqGIWw+fnAVfXHBsFYaP2/3p
lFYBK6VWnqopE7UW589LDtPw62by0xXeCEVRmP0udnjFVvoEEFScj0YP6o1XLPycxPvI8y4vgRK1
4yhZ3wsvmvsCLiBGwrtGAfkRYW+GtN2GCsiX06DeyqbcX8fYRHDHelwmEX3m6zeNFhPv97LWpL2g
7iWJOW+AiWgnDTyTmxQWdd+NYvtkOFKLJ5k1zIRaDX+NZhu4x0Ctyw3He37Qq2cH/gNznunnjAB5
g2lHvI45cdq8qVGXLtkBEUAV18mYNMQHvNpBb3SlnZvkofaomlka5+Ev+2I4Ds8Kiicjev1HJfb+
1rrua1QrSg74Yy1Dr2luTPgsF/XibsAQZUDmj057SHTlE64MfEcVAgSZOyH8R55+EissCubDtZj7
A23YwusZ2Vb8JNoxos6W4hymmfD/sz+A8pvvGnpHPbXhQ1DwBzuUwVlho/GsUs399jPys8Bxxlac
L+0yllBDGVWPd6YT5LNm9+Yjj/kN/6E8/AzNDITSDWUJBhN0xh2Fy8W4QTk6SvOUN3Zdssu/5IRM
3fVPw2yHaS8Wc8vrzNSv2NArtxUHlzatGYhfQxKlacHUm8C0yBptLCVVV6kh0qn0+mn2XlgLUtmx
3dL6PJl1BQ+kQ7bTmGkKs5tLEF1l45jB/PgyMszYlkS1HWUidYHBnbCshPIXKW/FpXH/n5Xw8eyb
7cdl4KOm6m/+c0qVzckBySpRmYYHPnxPuooxGUvbBZYnvlARn5D5pL0bMGpJQYSFOz9c8jvyaZeZ
CW4r/35M6NHYedQQ+kFmoY87PgcTuyAh5zt8BZICYy1ZZnYl2X8cutjez5wNkAG+GU90PGLGmpGT
fos/BxNfallhUFM2K83kIsGKXtpbhHoyOiM9YK16ZBW+Vz4nidm++5nqThhoB9oGxIb1KEP15iXZ
J0F4O1qU/YOrNoqShzUt26+HCEqhYkPI6kbfJz0vnPIsqEceNFVDM5JKGlj/LvyOLC2oHrzMopCE
/s0D4MiOxvJk3unin3AQ2g0/pltGzRIWPVEfdDEmmPNg97NXuhYZkZdBIH5cJ35DzJXM4iW0Xy4c
efrNsX3Reldn3xuOicr+CgjhUi3DCIZW4LCzUf1f9ruZ7YJc7W17LhZeu7bq5RruMau/I1XOlWPW
/Gl6RtBkyb1B4i9agH/aXKcfPVJiLgN9MAV0oA1hclz1DchoJOWzFhV8DbV2YwaOkU/HrmPUsQof
bThHZXGbCksestCvH5QnwTxEqDiIae9fny6lp/qOueTBHeXj0Atoryl+1e/dpHCwHtkBHhboEcHs
BAHkEimtcVLUf7XUey975Qyuxk2wVSaiyEIFBezOVkJk3NeAWlp2a2vM2NRg/OH9vMlI949BbGN2
pdobkb+10WNOfsbUleIk+pz6aLPO3cfD/nYuOc0qZB/kLl31ueMcTuqJE/YxxfQ7dRyvyZ0lbd/F
2MbBgcUv44fmkltEA0YINJoo7zya6FNdwnAL7zz4YJMd6apXrtKXXnfMQSN4GYzZS4p6DxrTvbuD
dosdu2c6jfVq8j1mW39lQxHaCFS1Bt9vsDtc1y7tQ73mCnHX8Dpps2yuswsj1N/kxIFkNREsB8g2
GmkyAjOtEwDq7RZNqX7s97kdV4maFxY/w735TQ9+50RcQ4Nqg6CYi3Ckgu1BIiHFmpUJRovLRPI3
SYY15pdGuk4fuxMw49SYRjJd90TbAjQ2NHlM/4MJCWceK8IyrCKeZw3bJbxou/njPDUi6lFfLRG1
ykpmw7wxQvZqmCXlCgylZ0kRPYKFKYiAY8azmswQfgfkLvX8x1qwduuPoDMJNSp07fiA5ToDnrY+
sNj192ZRgPCujrNZbSmkcqAdYh8qbtmiD6FfOB6ouGBNxK2iunLUSOVuvr1zE8TSHTYQpejJw3m7
A+5nCvYsh7sqHmSY4j8P9jU3NnFqMHESVQYR7iBYstcGyUDPrR9MtszzobXTOUoC16alWW+WYWJw
zbN6DzxXPlVfouUomblV3r45owUamucdRrZyVurtYo/yHm1kHWENNfO2q13Drk9jn6yzZxHtSrJV
irtt8GmJjVlQONqvmnW9uzGQRBm45hzq+dE5GmPQQynCkfrsG/gzkQGgguzME2kqvAqiMBmtZXrd
TCIiO/S/1mgrqEoq0LIebWjLJRLPnwO92tyVsOkUo+prRUq6smyIWx3mEB2ynhGaBtAv9EG5VD1L
YGuB0L4bk4Ye9COgYTz3Syrlkjf+eiR028suui8pHYIDuJ0+bqSonTo0qaLgtnDL1gpR+1EUTkLg
0SpDfZzd+evoY90VJvgJI3Mh4495lkEZaI8/oLba+lh46R9CePoLb/zi4dJv2pE8KTR1t5pGYHjO
5LBpaPF7V0ljh7nMZu9VftmglEeEMvq2BrCYB1oFwSRwCn0TpYOzzkW53NqnCh48sYiPmfmT/gQd
j6Yc+nOz1OwrwbMuRjCDNmEOcR0ZBQLKmGWvofxXaaG5PZ7bWB0mAI4LeIgOYkdvb1cVSV8silBO
5UqMZBxj6YO2zlTi1jIGy933JTGUnQomh+2Kzo/jGoF8i9q8hiAytLzljlKJ2CMg7Qa8QlOCg6hQ
M7dc3ibAsPGGNzbFoLUTst3nYmsFC0nOGiKXed1UKQs3YdaHMwAp7A0XyJpiiANHVg1kZTZ7tOZ5
P/DR6zpfQzM+fdJqT6tu9UjF8x2E8FVbAA7M+M+7Iuh1pVVSH6SplJbyieXpFwYtvnEyGfPqf9XR
24mrbP0tT02LUIcI/AYisEWjlbxsi9tzWe9fzHLbm46r9yVeY11knvXA97KGJU8P30CyUw2Rphll
zlnwlmvDb0kCUUjdaU03KkF+e11rN/xByAWhnwzcZGWBZRnRmIv3Y5dqcCI/qaX8AoqCsaDaj54Z
c19r59Dw6GAjQAidHntZZSkdAH8MnSa1iazfHth/1mAoKVIKJ68AjDgCQM5/wTGbxsr/LRyVboEk
ZVyRc7uWOCBmGOw/4AR72NdeE/s0tH+ZEQLoM64U6r/GtaLiURjYIP55h5b4TeRAKaU0Uar4Q44e
o06cgD1raqEQW6tg8KU2Xj25xNdyg1pJHVb9FFk19aYbhsoacoOtKWyqev5iLo0iomR6YM3SsEe+
hNh2qMptPSAqBuSNlm7ro/nxa3naUknPAyIV24E/SLLtnydi5NjnWMwLghz3it52enPciZFrrG4q
5XU086yFmnYaDE4mLWymChWiF39m5BfomTskMYHJz/NILHWTnJb44iPdYbStWTrKoo1RHfltK1De
vvgzaxynQ/1jl5q8j6iO18hqsygKPK453F3lr47NDu/qQhShI4J7EJvOeMWBUuHXVXuKtCVSrryi
k6Zhh/IB2pKFlDA38iY/K/ZbV44sWAUp0u4uUmdHrUOE8HO/o52o9xWyITIxV/qt74urh47QKLnq
cKi5aYgcUhPZSTY6EnMe2z1+SvEZ18s9y1Uk9tk9w4i1fnDtXdAfmwWclxxPqBCtgY/6CPQ3arlr
ZNBtTpZoCDL4MIqPr6Nk4SygSgzpw6sKJRcjSubNoPlRK4cNUSXikBrSwfMH8uxnKoqpmRwriCdd
l50b3K45RpvOkXag+oNq9uykwiS0vCvZL0MTduLQA3b1uhhFXwhyQJhbnsdEkpHmTTsQumCcwm4/
xys0qdawL5kbieG6mBwGtti0pXkerPYRQc6cd17T+O3NRuwaUQ46eEsx8R83k0hpZohUqL3PmbaA
HX8dWe7/GtT2IGW9EKGOB95CNsbC1zgYNQELQwkOxvIPjsvlY99pC5tBpUX15ErgNLW991ptqwDk
uWdfDO6HR3wvQbVTuZMLcUr6l8xm0d6d+6kWfYeq4S9NJWyCUKiU/pilQtZVqC48KB7T3b+YB21o
P0nqwXMeJhofNEIPKgs/kr+6cIPcKrXjWxT2L+zAPawWGkCLqgIh7XpDZyLU780x58so0lRAMxH9
2DWsvblh+d0ESNe8NQgEluGt7/ZFfyOuMP7q+x45Vef7PRt2/8p1SQ/RwtOHKr/0taxl5DSRrG83
oYGNoVUTzulcWn91BFI6Q5zS6IYT+U50iS15CA8BJK05pf1fvXVmFkDzTaP4znNrCc0UCeFUAVJf
mb8QRnd2gr8Gi4mZSPh+hgwCdRTrGSMkWGb9vJBeJFeTyyguTlxUgYSEFBo93MPdMBzhNxzN+phQ
ECaV4z7WMFqxB789uVVXBmWPRw2Hj7uhvRstgNleI366hjWmVfRQL8pCdiLnFEIwhxgSgs1r3Mrc
nyo/+aKsfKAfBU7b/7UrhCu22KigfYFEj2Hk2KWSGtrtCUfPWBCQ/xdTb/mPx1yhG+1znYVbQ0+3
Qf34iRQlGdz2bqXSpS9pyeZNxg4kMU0q4VacTgbxWTsz9gZp6/OhfO1da2I1f1puZb0DZQdHhFBg
zs3hepFChnBUWKnlr7hpVSNlVaa+utCXROq6yfDjawOYZstVz7UV8XXoAlxAHpewJ1ep/U0JrK6Q
yUbQTc1TmaO/YSXs0MVfQQJqH0DLUql0qanR6Wt9hoHNG5jibTW+FHtKzth+Gxy/vtY85sdmfJ6L
6D76bSuYeQI/mXBSZh53vqR5pARKIR87Q8vqtJ+z9MTOu45mfOeJYxkcBzTouoL57rnve9mNUuoF
FPrKtTyqywWgsQI5gOwVWiMUmUjboQBtJXdN3zRx3OS80IRrEuGTy7JZvKDZNc1Jsm08GNssmBVC
+CmLVORK2xrGejs6A1lwFZV+li3jNzAx6PjUbM5gCbVPATsMQizOeP40pFw5vqZb4K99SlU1KuUG
7e+fe1kkl0n7PMnZtI2/00MdxnfLBeLuXci2eQifBCdAG2mMDXKJs1nuEHcyrrUyg/Xq6+niUuVB
L79A6BzQNb+gZrPN45YqyFmr7VETV7ZMF6bpJTq0hNhkjT1bnOlSmcn0Ni5J2vU/oYJz6lnPDkS/
kNAgx7usn6Qx3MkFGjlfZq0nmNXc25iirWCzJDN987e6QTua0GNf10sHzuBTzRJPukR75TmktcD9
vQ4wBl6inagEeoq+BBkTuNrp4/3He5J6B+/aJ1/NFfsGaT5j0FUdw/WP/JTBedqQ0Ya3YSLSoVB2
rfxBZz14O54RBBswHcn+koeeugQJRZpxNvkkosnFAT8PYiBIrZcWvoUoFK5U/C6ykwyAzGrAazjQ
LYxlrQyFoawn/8ptzOlKc/iWT3asA925wrpr9Dl6oALroBU9Z9tonqqKshZiMiVtE9QkTLbawdMc
h1Eo89wySkhVti/VLAKyGmKaLm+2vw3wlpF3Ednsf4+kS0jXVxPeYIDZd6S53M/diX4oMTSDGZp3
V22EjID23vww8fUbHvuPgMLHRfyD7ViiCRl3h88H3RO57FtLGxwle+kKqKO45//TGkjkpRD34ixp
s6PGBnOiomYDDhwMFh0O60pcSCfdB9tdqE3jxvo5ByEmXNLq/hkP+eD5J8UZ9dRrKtIhMQFDmfbn
i3oE8EOhz3t/gnYYo9rCK/GllGidukCcTcMWwIi5T+LS0VTEc3H/B2sZDOIP1OsgM6yccS27CrL/
1Ft7YDtzKSizmE/sjapqlP9Ix95tU+RZ9PddcRxEaOENAxMORCNLHwL52bdORFviHpBeCu4Evl2p
yOIyJn0pGo49TZhsLywuvRBK31OKrVpwQSZp6q2cM7monVZEys5re0aBJZpQRcDZIyKRPTJVZqqn
f6CHoC866C5q+BBj98xO2YiVLbo0hMRUvixEkVLQ2dn8lrujWsJjLKZeaXJh0poVfFXkR5TrE6by
AUB87CcMjrHJ/bgFLnb8TYnDMI0vXp1F8qrqLbbsaOfvrVX225v4+A9pY8G4fDmp1ETquJ3yQOO6
j4rvyWGcYCBvSqdjYcbcxssO0sXTdKyWETPy85M4sslDxJNoSIr05lgGJabqEAJgWjgov+AA3oq1
UVJI2qyR42zr8zGp5w+6VZO4mibwrDlgCk0prs5D/IIWd34154zIFIRIeVC8YD6K24tY7EmCuICw
3H1tbxTzeY2DOMV/4h/9MY9Fybx0ft5nCtn6VJRgR4cxC2/n36PxMApIgvUA+5/YEq6jYCB+AQFP
/bUkeNZJsafy3KnEKkTsCjWxpE/89mNCtJY3GNsCopFp5KJTBVcY3LlPb2DQDlftdAGeqYchQgyX
BvOExQ5id6gMI4INZuH6Rw0SpwdojeexlnUK2N6vjwZdfc9iS944mScj7iygjqV2csL4NM5Q7vMo
EYZpsQCIb6/nRxF8P8eV7L6ssnVQ7CpiALIsenAm0ms4fQgQONCqP6EIRrWCQnCaIyDiRPbhKHUM
JXR0ka4jVSI/RD7KJz4jJLLVrqoWp30KCniJAZINXnDlkY8XtvPEF4QLBNU2lHiP7VEjdqYS/RDI
KgbsBVktni+VZYwQLXjM06bibWi7Hi2l6J5mj3evDkWugrxsHUd2YJ8W8/zmozFsQ8uJN+DGpK/Y
IhXit0Y0b3yXUZENbWMuyiTMTKSThlyuX/VOMcydUjbcrAo8hUZfGsBn+Zlsf0asyc8p4/85V+7l
tB4czSHxSaAw29NXroL7hkgn3wp70gviCxUT+9Wfyk30+YUJegOKy9hcvcFyFfAwYS0U95MAJ+1c
FGjc8rxsy1lo/in0dHOHQ4kD6vWljdA80FSDsbjdOQ1u9YYR39q5dCEdJiP0yTmeecNdtOd/varX
Jl8IW3qZqs9/RCQAWEudB0e+0MEPnfRUsaWNHFBYYi8UVoWHWNIvi3wWzupi9TO871KwTuYJyJZy
YVfcbcrjjALEdgN+ArrxqlOp7lOIT0K01buS//PGuB3JQOfz2GPCV+Mu6aCZfWWLJC8ZhRH/Luhv
FF7efD3K8JYMdtCbaYfJKw+arLM3vf9Zq1VDhgOpbhtrtlTMyzBl1VWZTfMZzshtCBfSdbtsRIj8
+PNoBOFjHcHhtUPJmcv3Q7BX4dwNzOz5SmyrbTr84kblMNYAg8brcGemManlul0m7mLlFKBVmCff
0g6dDsojF9FlaShcZN0lAUWT7YOQ2lHtxMjQ9ffXQddELGwi60vSScHzqS+qfaL3VqMGopD/17oP
Ny/xhhHw3DK0T3WLeKxc3ksXZJP2AKQIDI/I4vV3Yg59jy2w7/+lOvUu6ZTkhPv7ruCCeW6KMOWg
tZbMTJqvqv1B98MJI54+PON7w+lCI40m4SVI/eVGwdlVP+aKPHbCmagvk1UIYJIGMn0tUkB4uLLO
UVeTyjq39VYvAwkYAxAY04i09OC3eBfTzhKYUevN7n4Y6TkCaRyXGaQXLokOQGCK+iijxyexIHEk
7syms2TRPM2DQJadTVHDO70L1yo3PwLUzmEhCDo6erJsPrW9L9CuG1jP6Gigmo6hNw383whtAB0O
0kUGNMen/gQko+9Pu9Z+trOLPMcKy+kOQG0DO++qGj3SCeo8YNKU0yGhUwt+wdDOyiKwsSXo8xna
bIAJYvfCEkod+90PP/zhd3Xd+UaDqUMsH/0ALebczX8IpejrVajWH1hqVco6sNWhueh0+xMRL7yA
cSOXDaNucUDXHaoqfPeRVLDiZTOx5uodyMLMQVGpy3cll2XCh2OjoyBcACZAhR5/C+hsmHOWwtJR
Xtc23stqxKiUrX2oxuNQARWrKu5lyHGwiHFQOCRFcZABVxRAMPec4hkMKBQqGmLZEqOs7S2BEM/P
i8kGl0/UZmREjOtjNFQXLpdiy+JGhomM89aMnJfrnrfQBS6JVwArgxUvWlpdsMBssaDK5bjrS5TB
bFnbjbChi86VG73eTbGu4zbRZOlQyBZUnWzOuLuceBPGYd8Nzd4krvMEkzywfcorh3iupkWhPDau
fu36x7eEfhPHCERSLcKJkzrZIMKcDpUVK879WsBWSqAZ3pdJc3OXx/I4qN4AjxAVPiEWjlCqTHJm
IG+7CjF/4InhnRF/NQLBqskTH+xmtZNcNAqNlimIzpjDhDctxchG1lACkTxidmw2cTdpFOqx+lao
LAKNQadQdc3fwmsD+Y4SNpu/UaFUT9sBKO/3D7N1O5+PM3MHwALuvUqiXVn9Ef/ksaa3aYDrhXnw
4e96ERz1VsBlPnwSD4Emf3NPrQPI8YMEHYp/V7JOKW6HkAHJYcZZKZV5I8Y4ADlahEm5OhK16RWl
4A4mVTIX4rMdyUDhGbL2o9BqfnkyuwOvQAWl38S8nqIuD3l7DN16tFMoqYh3QKkkKt7MC3LvRdVx
JyNWI0UHAnIUFejcsoyX41yfhKKjKyp9jKaIX5m7XFGY9EB87UHS9fCcT2NlRHvu25nyMaLHletP
eTURVEXWwsNobgg3hrR5hT9lsc8Ry+FOEUgbv865wCPB+nX2vb/YeBwQ3qOlx7/djITQ+UarP4R1
y3tQTsgJRiLIsiA5EU9PjAx0Yc7ncJgS9iWtpQjegFOzmBqKsi5EsQP7MA652VYGhz1nBRgM7JDo
YLBWQwNowIfo6coxSS4QnEBO7VM3J4Pext0vJjzMt4a0LtuKuL7rg2gIwsnFLtkCxNt5loSZg4E2
5/e8Nnyh4FLoah0548VRmiBkYAxMBGwPEwVdIZaXtWxa1xdcy+XALrPug+O7bmrhrMPtpg6P5uS6
vU9ENobsivLHtZBVGGTji/I1JaSunOjKgCDfoQLrEseWOcK5iUikYa1nmDYQgDJWIwPVj4S4wLuq
9i1HkStK55N5dyvY5Id+UUdU9nsDURT28RIpuRI1gTd2f00Us/UsGWW4iH5Tj5NqkM0OPOWHQxfU
RKboyAGOZoJjnceFg6c+tGrQ5L2p+F0zO6mz6yLWfhkt7Jr85/wNfsnOORiH1S+7yg9bKiHKcKXy
jyh0/PKyy34EuoxlpdK8BE3tgob1Oc96qXnkIX7SPe8HRlFoDsDJQ3+15J3+rLLm0j7BCSKF8Ia7
wjKvEyrn/gdpyQ00SN60c2ZXgTJAvgU5i+ZgUTpkTasRHTBtqwFmh4f8yTKJdqFFLzycR0AnbyVG
QqcwsPiUHeF+YUb9bZ9u6GjUXw5tHP0xv+tpa0wOUBlXx27ILLUmabLODIYT42qNfKRiNBACcwPD
T3UzcMo64S4HAFJYzHQmbM7YUQZpiAIKsGG90LnsGlIN/dxyeivi4OQb4F6lkWRhH1iYvhlkMRiX
0FT+jkfhEPBN1S6gGvHOTq7x1/j+cO1fEcXhfv4GxtUmShOU6GR71/ippVfUsV62l/sjmuYUm1QR
7UcUmQxxm1H93stQ7J97y1MZ2N0jBuZvT4g3M2BugJjMDLNfEY/JJiBf8baJotacL9tIZGfjAlu1
mdzIsnynp+iVQA+0JmnnIO/q483ypq/TO0pwhWbKlTIW1k9IYf4lWLxr7iVKRlQdmVUomJ6aJzeg
YXCtnQUwDKpiFc6Zck+llV/3ODxp/AOK3kFTy0aCamGqIaisLvcYX6JXBx+SkqC09gw6w6cKTgV4
sEAJeyiqJ4TIFHemgxADYQNpQHcBh74jGLv8LDQ4UwVzuz8Dtlo5rpa6DFJaUUFGeaHxXPQkI9xF
UH7/uFndt3X3ZYFuihHGwuFw6pGLv63o9A4ZUf5PcxtP3ra/z/YP1Dyexie41PxuMd89iw+Pd9P5
GhMhovyRVDz63UYsSQUFAYPPMyRRksFV6AegE7h6GTY28KUKnZ7sJIap4LgAKCnAM71FEvYIZLwI
cxnh6sg9IMv/rzKRkRrMaJ+lUzsAfc9upZUkJNUyJgFdW7iG9jpsImJlxO1oA1vXa5KcXmpUHhwc
8iSK3rZ/eBXuf2FyUeYxCOR5NcAduxx+9idi+R1W8I0x6i75cmxwSHofl2NXJuJvgSPFFkEmulJH
ENMVQB1gbyTcax/HmXvbO2wmk5tr68LJiPcJ83og1cIlhbG2mZydTo3Dis7QmGtQe9m6RWI1UZ6Q
HuhgjAT+O5oIvTT1+CCWvGjItcLB2s2uTVo3aD8TIb45BhZ8uknZPI3m2Ca2CDFMVTz0N6ENW0bb
VTrTyhMrAy4DRIfW/ABSRrT4veImuUz9qc8qOwZjQbNPzZ9VZJLDovuVeg/Qko75P310+NwDgPpP
Vchze/EUYKxOGnnL0uEJ7nj5fzX1tZAbbL+fFDHwcuC6Fev4eeGtt/eS851fwTNe3izinxmBx/KK
124796KAkmaEvtNscKVBRVDy26JyS4KVber7Ujy13tXKPZKZmjhTvuUOEl71OQBl/0bevDoz80Dy
6bUcPM858p2atguePmnfycZWqGYjS0uxu9vsg06Be1VeP7wPtxNIeOEG4cLWRxb3/ERxz3f13v5f
4MV2LEjGfXeQl0dfIDsgr54WyW46WAfwyBNOHJStUa85NiPehq1gXNyEwvl/zABJvZ9VkyvNqBfS
k6TX+QKMv+sXe3w4DKjXPIiz5KMbC63UYYBzENlB5dHFfn6VOx3HKwF2YeROZpYVMaKLbQI1hnUa
EFU0o5zZqnFz4xCGrdKkGoKgvz5F4yvsV3lgFzPSFXblz9+uHO9I5mbT46UqT1d1tbMtngd1Cbnh
Ox07BpCeCOtoqaofQKkMMVIqqLnMQT74kA/8gE91zxgdkMU5c1t94TEF5Eez77Dl9OaNa98iO9SY
Xl2dhjLQYCNADfhS4HESHL2Uqa9LAf84Mwb/TYdMllOgcBMqca++l+Rld80DE3XOu5gBy47fjSIy
pb1aPoTY4QlUtHJReiIT6sStXvZkM4cZiw5TeEdtxEwRBn8M0iLqZgi19H/Ya61iP/MFS9VEEOg6
obpUs71xUSV2uwKS4Ogn7sGpRv1Jt0Z8DzKjNxBpSU5N6UpMDi6Fy0DyJuQmaYy4kkrFJYwStlv+
nzedAN4RjhZij3WvxZiiTMYWFMA6oRqmcJP3ZflK3inX9lwtWzVoKMabubl7hbYUs0J/vh2wds+a
QhucLuqttgXifLhZS2q6lYNmVe0BZcKEAIG/cfW0ccYYhNXdQqRaseaYR3TJPsUPEFLaHuv40Xd6
ir+5G4hD/DYxKuH60S4ihX+Lr0vPkdc5D7p1AY7mgrgXLSxum20t8+LqR3QDi+nhFfDxX9Rm5Fig
cXnZqoHW40CB85DKglQyAZ609xn0DhMfEcxK47i7IdzqK4Fy2EZ73EuUfLsjVlia+fC1/DY7cp+F
kH0DtmGHkv7Fk6P53JFQFooCeeXDzRF3s0GMw+c3tQYPA6O5cMPLYjC7nJr5+IkcUsatAw8RVpOk
hGx2fCcS+xI87F5CSJEZb1w8oltvw5F+IrKgXXv+q8Ce+OsMJmoTGZ+wUniDOJHJUf0hbce9z4IL
1WCQwWGwujZfETHOX++gudHsgmgc6iGu/u1rVCerjxcCLEirCn1XFmje/Wa/cSHJRzy6jBqOfZu8
3tPxHPy/goIehdN64uj0Q6R+UdEFUZzEkjOSZAG6Nj0HC39+nJyV+E9p67CXfaxYkfk1qTuqKmg5
hZM7d01+V7nJyqmA5z0JKCCWaAOJOSDQXCim5Upn1VKkWd0QgWR709D9X1LuxJY+ojwAKd63kh1b
vXWM6Whq6KZ6sRIGnYF6dZpz0Xt3e1xJ5v5kS8mgeknuSQYXhhAr2D5LGlXxUXUUxxvkE1kM+UeJ
w26rfJ3U7LuJiIuiJaWLkM1WDE7cdztzz1RNOQe43MdPFUe5eN83Y5o3T9r5qzLo9Mj0bVZbPgcV
Q5vKqdwo+oc7r5hW4SQHR8OK0llGd7dKkyjNFYnU1tywnhoR2kSbKUwbjSfm1kKCjrpHDuCKMUoS
d9C4f2LrQr6Twvgnr065Agg7YO1wbAnslCvl1wyVdhx1H8pfFvTpRv9vXJTsEX3hbvzvKl3cYk6n
pUZNxhHyJbehzWm2ojvjz48SIbElKODzOsVyY/uQ8RxWHjBSnUWuM1rAVD09cxPfdXvoMNg9xRKU
PttBRTq/tdmA1mCfoG7hNhUmYl3EU/bp+R/lHAop1q4eNA02MNydj48Csw+NcAR07LjmcVoLtKxM
Cc9ZegdTR31A5NlBl528mmZSkbUBxp/30f0O7jLdL7f3ED+omZIYYkvHPFEyC0vPI3fLotTE2XV7
dzKmkwZEXPP2F5uJ808ny1w5KCKi+pYPoxZlO7+KXhEi1iZlRHy1ZIzpSKgFJcmE1UJCrY7NQC3r
b8aa1BMA0X3OA4LWlL6KJxFhcMPXqUO1gh0BMtw02cwlrOVtiDGm2JbR5fwZ4KBG8qxVbxtaj/zr
HAAhFp2wEhuNCVyn8XnMs9EwrcdkbZq7xWDARHIiH2+ceOK8MwJT1H1T0hJD+cHZA3LjefjJobm6
FxYeVgBhRauTfx0J2SgoJPCfB9TgGIrJylA4g9HMyEhFQbfrQJKYQjO5HCxFrmObyGU6pcVln7hh
DMasWIKlhZRIskdc3zW3DTl6b4KGpw7Jelvz9UZnEqpO0cAWGNCDtp1fPZ4ldoIw+GqI1is/Yotu
WmkL9hFbGsLvzIVoQKoBZjCGKF/KVAyn4CaUPC7n0so4/0YRmLmLZlIXLhklJs0lNAK3jA7kXU9m
vGamUWPrEwBeLqOAEM9aBRlZcsSV5UMj8JklUKCzND+OZD99XFQWJpAHS3ocCs5H9Z9ffc0vkTaK
IjMo2AaD4Ve8NNVNf0p/T/gK0POhobUdIpKnfpY9wmpyYesW7FsC7jEaeeRO3U53geCSvrjg2MlO
w+C9MAMxJvI9PgU12QBTA1WC7dPffsafrTrgPs/qOUPFWNIKng+a+DCG6tVlZO7SX83ENQ/90BZ1
lFmX4Nva3/dBdbkrlEl3m6js2thmRzf3MxAzR0H4aOtaKhkTQhONjOkqx7MrkU4beTQh0jOXZxX/
jjuuWzfD1lHDbQQu5m4Z5Ok4x9DqrdWDJuzvg8ckcue+UTsEqXVni8s9SCfUwO9xhDQA85iebNjC
rkN8Ymk3y8QW+nb+4VKNlE0KVq0pTp/FqQhRhxF4QcObvg0fgjsmPXv+1xGfnUoWc5vsA77vTJUE
7H9chMPMN5T3ZH7eo7auzT60OOnJxDfl8grW0t28NQufb14mC9RrGhzll3exMQJttSTOoEe0yt8f
GHcQclYgUEkzi4N6Fha9M8RrEr0LtREbpgAZbJcm6xI7qHeNMXjBNceF7AQOyIsZXmVPmRJgkwHd
1SLruACM4z4qE/AgovL5lyZmKcrfOBOxmrJTiknYjC0cfDFIrGCOAdq0v8rF9kIX55qIZ35aeNez
YP9gWzOe4rNE1VRbHu4Ou6aFX0nNVADNs9icMMDhqKkkj7ns5FEcU5HIOxT7O0JBT/WXpvHJP5bI
9bZjcWUDR3xqQr154acY3IDGHDR0WQS6+GeW8u9NZo5LHWXdnopgECO96K917I5K2wvRyYT1GJD5
EDvtOd89934eBZ0XkZAogkE9ckC4Suu/T3jCk5Whuj0nwMbWaSJ7KKpLJmwQ8+ZKeOUVi+ofTPmg
86b5PVeVs8IccAiHz6bXIAgs214p1yuxUNsgedcLG/SofjyOs6jg7vUl3jutkMBt0n56eYFaG/oF
ewqAf0269y7mQ28D777I5FmtZ6g5eaZaIL2k1Je0B1vgQekQquGPPLQ2L0oHbYyEJFL4sQGQSHlQ
QQDWNJFtfbr5xOR4UAOEA9gWe7AeBXyRGyUox008azytkJi2Qwb7+9Pwh+jwqIchqlpr2uYrgTop
p1Qitcj37ZNcsis0CWlv+AcY3UGagU3fewMGB3fSLWvPUDnILXhfyILXRVnNR9CPJGVQWngi/ZHb
1KTUXnDiNnpmyzr7EMz15MqSP/h0XAi3qpCgc0tvvqGulYIFbBXsNWUBXDZUMCg0CaJCMGS7jLYf
CRFjezMEd/nUhi/fQiHps5uzF3/z6RFubSSBhyrSegA5DbBUljIeOMEW1tbHV3zrGBgF7UesvteG
vM5n1RCjpN/WqPk4r7ymBpWxurKzP+4DQDZ1+fs/lD2w39M4/sOjWx7VWpiNFKQ0oIwrKyz5jPNv
47lSn0ZidtvZR+n5L1W43yd7Ke5AagYA5drZEwnuy6qt0nRGgiOprZk+V2zyvgKAehXyc/LW4xKp
PZmvnlBgpswhPZdHJIH5sgQIwu3Ub+1qnLocSMakx07dwSSnJ/w2VCcWb/yBSGlps4KgMy8SrwK0
0S78Dii8a9y24cuaRGmc/eOCRs3CX6KTlUT1q9YSY/N2diYt7fTpqL6oGGkeS4XfFW/VKJP202A2
+vWAoeBOZOVBIuu7ROn7hd6HX7abjv+JeCO7ZSRt05L4r14MaKUiLgOEgodv3eMqesJy50Ma04sd
4/+8RRyu8Cgfl01DLZUBAMumqX5CQXgDeQmIJBvRc/BcIlaY8FRbfCOQeCQ3GF3LuR19fbXAhKOT
KBa3+34IVlT8m7eoejiOi38UI5ikwpvYj4FS3aBHIMYLJBZhPMJgpBzhT2cvS9ivn+xl1pvCJ7fy
Swc/tf/RlkM9AwTjxVMuydJKgULsCDi6LQLydGHRO1NQOiZzEKpU4PKed7ZNllDDL6VlG2J8c5Ip
pND19/8I03SRT1ejNRKqK0Z6fU/Cw8mdKUM4r0I0lBvmxsV/OKR9J0zMsDLRryIPsaaUmzvNqSWB
Ps3XUfqYBscCZAree05cKuY//KD2hO9kTzYlxB0d1nR+oBRqGQ5p7wxgoEgiBW0UYVmt1qfVZ/D8
Atn/U27gAMhVNaisKXovDqk9/couyJTgjSBWXmMQP+Im/3Ty5WXSyPc80FuQ8NCSnraKWdwr9TCm
ccy+48eBgONENKXfA5aAVjzlv8YxCuhHiTAlTjVi0p6M4SW6vWAt/EPzCdFQ+1MfpJZrqyAO5gq/
Z743XDkmyro7TdLNpZIyfomKw1nQJ/I7DqUJc+9k0Dc7tLRf4LeTJCBYU78N/t8O6juQzQ1igJnn
0gCmSPkSrQT3HmZJ85wgVehlRD1MWBX2MfNu7YR7YTA6N58fctuYakZstBWNuu3tWZwO+d4irO0K
rWmQjX1H+g6MaXUI7NqoJus52lEcmh6KFHTjOvfNfJR/QWpoG2lmkPQAwKk1KxmWJyuf8PdDNtNS
83MzDXiYcn9u+FNipO7+5OpFkn+QEHkQ0M9c6yG+XPY9XBhz8PP1SJfMNuOrxoArybtGQdVPvfgW
h3oKJ1DlYRrd5U74o+AHOutl1FBkuPEzOO/IhHODrcnqvuq8TojOqoRgVUclkZvF9mRbVmAKNl1H
nxgW//MV7Som2n0SAYA5F2sxTgg1+ZzTLo5CquAr1r9FNp+MBVURMaW5iydT3hHXykCk+G97vRPS
BBzlQfhPFDvKs73J5OZ0fFqE4ZJU3GOpchJT8lo7PpQ0oQ4U/q0J85IjwtlStfloL0FvCp+1rnGP
rKuuGlxMHMIHHEgocaQDleNQzjFGRqyeV+eMWH7/S08zaYLXzT5cZbK+HklZevhPpI+Y0YPFuBTb
ckeFNcbejNiWA6d1MgFUA3plY6lvUiy/zHx7xn+JNK/tODdgRURNbTohMgFLPHEnu1PDLxOAFtf4
KyDAqA6+BP7zR50huHkxmqRrQZlucD1ERr5zqfH02G14FuD+rWyAA6RAhSN7s8e2jBEv8ww7PC6V
kpMC1RJHJoqyYRbr+uOYN+YrgPiZ1WwVy2SYA6OvNtYBYwD5mtA31NivHPG5nYqBbf5hiBonCvAd
veYWD8BXr/oQrAdn9Ah5fhVqclywLSmdWGlY78a3vS5JhdiYi1bHxMP4J0nsA6Zhb6BJ23QfbC1E
7IdTde7neTwGorLKTaFOShAUmvvCl7nWFB4Zgp3SBitRdVkB3XGM87T1EwbytiOHjuSbOtughQQz
egHptAzbQR02rOW7UsR26/OfJeT0+SIxUqfqXF7pk1VtxUSLyNMlO7AEcu2zL2VKUt8f40DLw20y
dUWgMFBSq1v4nX3Z9irsEAsOglraSeKHPo9qp/As24QKKSf0zQtVGW/S5PvolM7RnBMbTrxv0gg8
vElmDGEDhdu604ZAGMV7wl95sVgSJVNoxHzq2C74IPwlUxRm6W9njECjvu9kgzR4uoG5OsPTmV4f
SzSPh8IO76+7s6WK7aMKH6C1lEbn8YpfCCmzAVaL0wuv/WPNxmSglV28Dnwxf5gI/y7nv9H8Rlk/
y7cPzuRY2rE98LYKaF08VJwzmmZjMxEPSA94P7g5sCbmqtd3Ptc60QfV8F/a2HfI+Y0EIv85oVXP
Y/z680KaMZz4MfVa/K+V3QMB9J8QKIDT0ZbM6sP4FCaI8rzPt3+5oPqzNW+ovJpWbttx4D81BD76
EqsepuOCU/5rfi1c4GE8kHEBY39VFYQdvCSfDn4JOT2urB+4Yw7qg2tB7wHIOAqzAIfTTAeqZQ3X
LR/LaXTXX7SHdcf1lT2STUu/5PBROp2hUN77PvY4NStYZTQZTo5QUc3PaaAFS0vASXSa61NMlXvd
lYoar7YdEgggMmwzqjoqS2hThFXF9jHZt/ZbSmkFQLlMPFUrFLT+LAsKtKfMc68cy6HyViw3WC2a
9lv7bs/4Y3WOceRabsqSqfbSxG1WrfUVcmnUHVI917tGjczA0RV1bbhHuJyASoxeOC0qznDRy1Fw
na7/DoMusesEKDVHrCD+CzJdi+Y8wf6jYCH9fkunm0S+yRtEEZfhwiD1ViZZag6NfPV6GxHYqdrb
gpAnb9x+OxdKMyPrK2tSLfPPtjM1yPXBI0S+TE9HooioaXnn6CG99ZwRRNV4DwICv7q1inSCfoAo
JWi0jZULbFTTWV0FTyiotspWxUfdezKgqwuVfzAuXg7BOsEqJWYxw4y0mU6q5PFLhfxSoPu3G7w3
uERl4UFLzZkdMPXqSfoLljV1ys+qIC0ET2ShICYFqYbiQEjLuN8rBnJ/iz57a2x+yysi/cz6Y9Yt
MilD8OaO+SliBMPZYr3WF7q3rYIDkC1t0Kq1gXr88FrE8zFegvjT/iNdAjNuOwdNLOgTZUwIZ134
jyILjSQkm3+B7GImzodW8mmygXE4Eds/of5TuNdnJzc8vkA0YW6bZDXaRWyO26uxPKPiMa/uTrMD
hYXPoJuqHqvNoM7N2gJ9vXL/o6wlOp+2TpFxKKwmIbHqgQVNknm3zCH7o/Wrsan/kmWDO1giKqWd
P0GcMINEzO/gldKPnh69htrIKtE51Xy6KBey30siQSh4KBOqcv6w+/zdEwVAqJR3lAXjcnLx/dWk
DSoz0vN2sWP89FRFVI3R3R4mEFn3OTkH3LaWr3+83DRaWlHBIRPARau3QZZKruCJ35epcyNNndSr
ldMBYGKKQ4otMwJqcDS+htTlqHhyBPfura8eyRGuU1YWPg5djMKdDGcSFF0UjoebWKTg8BZ2y0VG
HJHtJCiJdZtBFDZjbJr/CMbZbi4uxDb4ck43SLj03jjm+vcO9a1veEWmUygcDtbxB1lgP2rcHdCJ
YyjqL3nqQRFa1rrgclSoDKofZc1zU/WO42BwtayIgv0ZbQxHW6S+WJbVrQeEGtOvnqO+NxNEK1Ei
wsAWXlfuA/giMgqgqiZ7NARbWepgjHfALXaXBQ/1fzsB693TOXVmvxK3ZnRKvvosVsBBSmpR4Ww1
QHZTaupgbhXSIlf3LSbc2VrL6KUG6kJKsIP8lXcmuoGQep4LXq1D7kGjAeU5Jptr1H7EZfmzjJzd
KojKm8wra12dpzPy/+vKAEqMVM8wC7z3PjZJzMTyQZbpuIc6ITS8wEUoDCG+D/R4oy30QDGiGRvD
UD8USCEiMJZUhSUVt3DAx81qn5VoiqVhelJL5bU8slhdjcgxdNziN/3aa9gAn1jG3213Iu7Dw/o8
ex018Hu7sh9VH6I9nuSLdDuCxWU1tfkhPtuUnwZlTnSQSEoATsfo2KQGlnUJ4B3HAsKPXDBQRmI1
LGFI+LgA3f3BL0OaEnxzVUWXszzfXhoGICaqiuvR1mKbBiJx5fl6t58OCFUuOGYhebng7K0wcwyW
aQvqr1NiSJ5qhGDi7ALmKR+Dv7RHzwQvmP7J81os/qslN2OlvEva4gqyeuQRyzyhmt+unhCvbaVY
bvznLGbvvLajQaP6zV5DLHjXRYwxxquxlofd5fUmcRkDN0Kw+uAPD1nEjYjYUIgPQxbt+RzxHrAE
vrZmtePaAsIzXFmghy/OoeVTZrleoqFTpkIiC2AlEfcHOrEAhL0YOpzON4ZIuT6+5bnLwVON5yxQ
kwlCWZbhluGLBIkRJ8T+t7SlrE5e3795lkl0/4tBGdvMSAXzBXO8ET2/LJbcEuquotlLhEcnRH99
H/GMDebG4Og3YgsgQdAAS2Z3wBuPDycruLy7T8YxrUDoMyT3OgbyqPc3RqGjSRi105V5SHVQxWig
jU53izZM96GwH7zxJttRd4y5RVWb2V9iDyKGBDH78ujUmjYHUiIZ3fq5t8DwoTwHppEnuC2BXS1Y
HAU4/0sANd5q8M3n2cGyXArWPLP6AQMoU/+w23icwsjYX8/k4APaZUWL78+ikLiJScMmGH5j4GBh
XMalLfVZBd1u+H9oUvEanAFhySRyWGetrGqCn5EnYSIs5eUfHu3OdYy7tbFoZktCOTcyMBVV80bj
kMMvGWIDHZ9Oyk8nn05KMU3I9Ob5G/pDLcTqyqQHmkzfu2jgzqU7E7iLiENBnnuPabOQM0vlIMqt
6+j8AvSpOobOatC+qXXGusmxkbIdCZq3K1Y98ywGo1V6tY1mg1R2uNat6g3Zkno/+o2BRzzkUi/R
LhF6uwKE88tUvbaB8QY9YHzfIgkCFllCMmbqVFTv6tHjDvMd4WiF7L65Bzc5TOUGZXoHZId4LHhu
+WesDkNDeAPIjLEF2diOGO4+t0smTFsz7fCpAMq85nuA7rFlzO68E2gS1FQG1AXifQnf3/BZ3ksq
lEJWkltf11SCU9nzYQ+SdiROOsGtF2sx5FB5Sm0wazPDDT294Ef/sUGZAHIM1LzC8xBNmIBSEdWb
CrMGBCraWp1lgkJYjxH7nvM5di9em5Q2B6/iU9MrbVurVvzo1WivimvGpoBICRUO4dKVD/9IFdco
xz5//MzZHBG/ghTg56BH8Iejjb9Y+Z45loFUMJr3dIlYQS2Z0jLO7L6gOrUgL4Tha/rBO8c8z/+S
Pwq+ZMwt6so8KHvFUkB9b/qYBZnIZ+FLS/6qCWoT3d+UQI8ubgMSgdr38VAu9DfXhAJysKQOys/O
IEF/hC8BTfKObCZyOMVo2TzXAUaY3StVO5cT/jRl+6H8Uxg959hQm+YicQP9yYSyjCJC0asZ9s1E
jxs2fswPr7TCPeR1iym4SUcAFnDST66448/YpkoGhj3H8iYdwd/z8hUyQ7AXm9vTb8J6Rb1Rv20e
U0S0/oJc/qLtaoS0BDVLzu5l7i3Jnt+Uoi07Jo/78Ay4YvrPpKtD3BijkEK7a2d7aRcT1y8G7PNd
3MToatIdkrSa8/jp5O5FqFeSD9CA4McNEBP2dxrNOrIkEpdL7ANva9TR1Teu0BN30aWigQn4vkaB
KD43hiAJu7YKABF4mZxwEddjpCZRsGnZjq11TAvsd+DDQaWrcOTRinKhBS4iKxYsQU1QvFGF6Luy
SV3jTQX3275sC6KAabcluPUhvQevuEOpqGKgxE7MZZHHieoJJcNWHD78xQT6nWo0U0inXzxygyMq
Wj6RSmjjnkOkC+iVUzL+E+Qy/EmS9AxVfGwtInhRuWMBesYWM7vRsxkhpf+lZJc6eutH9CtneEC8
X315/dK34iTR7vSNPjGTumv9+aj3By7JgJWvJurqC5rP0ATt7JevrljKZbJp6O+2nUj6wzGqXXoh
66takmB/z69EnHMThSIwjEHpA5E3y2payAxKPnP9eoUL6Wog6aVS8R9RkQ9/dKRWXf4wLI1O74iP
zzMCIc7H0Ii2m9SnTt5IOa9b+XiFnArgVVv86qVNwL3VVt7c3w575Dnu23vVBCh9gpsLj+TInQMf
yhPi0Xsc3sjTyBaJlE2N9tGrStmv0d9MnMpsO42gwKT5f/yihNpOiGGoGZyLKyjPBcMF2h5wRQlc
Qh+CUssEBFuuymD8XcNRjTBJMyCrMhxqfxOE3VRaXgNulAez2ZGDfnzFS5o3PbDEAnWFvNngsN7V
1F0/kqS+/7meTy2pixHPJA5o5Bo7iIJBrhiaZfIcx+QVBh1NLoJ/QO2J/DQPYw9EPjX6z1qsS83w
2dV+wQDs0uGpm3sanlI7SzJ7KVKPiqrDDwhz/3Ujh5IOfXqECXMrdsDl08Re6UtfZP8/MPL6mQf8
93XEq225mGmshMor6/7jpefuOgqiNjbwulXNwsuik7MHibT8RgBFHfkgp1FuFrnIk7EyMIZo6izG
UkjpZ402F9Ls5wf5dBfa0iIbJGGrQCPmthbPl22jSEBzYEIcuCGe3VH0sO5TXRGAHZZeY241EY8i
cuZSVQoL22pcH1GIjwuioadklLv1BmohP/yXDgUnpeVFQHVmNXU4Le5xfwwssXyWuqG76hJOeoxi
lFGTX6H+Bobaee03hKnmCAfjjtv8uXlFhOz8wY9tw2j+G4mDZLG99SBAfu3pPh20r86UvSUZpFxb
zBxnsyRVSslUXnog7du202tzVGkAlc8gnHALQUd9AAdnOZJNNLvqESRBopH/en37cmDHVvRAL5n6
mfYGneia/7sduYrg41oTK9NCs57Fou1GSe5HS5+0DOQfPVQHDiYkw2VMxTe5CHNySyV1l8SMqzlN
UrRm9H1+YEV029ilORqdlXXZLokWvgXcl3+YW6bhbgJKgh/WmGJxDuRWHgZkrYUXgJZnmqCq5x8N
o6U/EtEOhqoj+O8Vr7FBvFG+uZWENOE1ZrRu0Da5e78Fep4o2gd4mE1TbZIdkXsgPY/GT6qkecnA
js85VHYU8Mez3EzxL2c+OuN71UsbVLWFyc8s2ft1Iwo1qF/xjKSGUXVCUN4h+jzG/yGjOmpr5jch
01ywn/AZlGGSflXa/tUnN5E7ljgHi5ZmymfQta5m4xo84i0+mbu5zlVRRXMel24moCOxFAGWa3NO
VSijaoDQ+eYGIxdtsE17rgLOWHNjtEDfMh6vlMXQyDygKFKXOOJ04IGb8Khp0bf2FPc0iPfaPq3O
sS6HfLjx0iq6XwHByMFvZzwIFUueiucquesA4W8/P9BZsTPkUUnF5nfBOShwzvZN8/fJbIzHTFcQ
6iRKxVOAAH2lEoJ1eV9+klipdUAiynw3F5neyhfwvwKCfJ76CG9LK1aPbm0cS72dlYL1UTdilZH2
xOrdkTnhZaTJMXs6WRSYpJkseWmfkeyT0y+xzAwvzip6gKjC93WsnIegafv0ekBWdunKrmE4Wn8F
uQRXnImseI4FRfR+uSznpI+BgeN3dPzJZIPhSRlSsE0ND7NXSYCLfPIpJvGJPSlBzb3IMwfB3kpu
iLfQwcrPCFqSyGKOI3aUTCbDWbzhoRCMvxxG7IXO6igW6NFMy/mJEek9BEuXmQ4UifHi27He7nr/
msYcxzqKuqqWyyNrnsTwypYsm1fXUclkSm84+GmtF9ZCk4WV4/X/CG3IXJx4ecF1+H/fIb11NPhU
I5048hQJEpSLSlyhjHLwja8SIvCgA4ONdi5SK1+kSRxioZyOD3VAGuTdJ6Kbx6jqYQDe0MvqSuCb
QNGX7ev6X1QW8nFVoI40AZcvm1GHADHlf2G6DzFFNoCgKPG6VVZIseXNFCwhXQm5hi08D1Ibv9vQ
enHH+gtr4IMxbWZccSuUJP3+iwMZq7RDATVpJKU515JN5l2lqS5cFpc7KlQTvDXojB07k+Ji9gzy
Id+5s8KnS4HP15CqFT5vU4u5b8r6sSgNax7v5AYSsgHSWSzFJYnZaf9x78gwvF7itpYlflgUi0jK
fcMAX/kXKsO3vG5y4YVuYX+gY4ptIdAFSy2QZiCiI2Kp3hcfLDWmeKW+pqD0XTO7avFTGsRie6+P
x5180susL7jZrLF7A0X67B9w65itcb6bpdA/L+xA73M9xugAUQoO4wZilOqI9f5diD4IX2UMAplJ
M52SWcco1lWp9hHZzrrCcI9lBA++QY1/EOYTu6dVP8km6kcSgMTYZAtDQbA40W2dfVwBQtvGaxkn
sOi5OkngOHtEOeLKhOdig5wHCr56hskoCVvUv4P/f1FYOizceWJByRgl7jM+/OGbVDC8ptvlfGe4
iEXkU/+q/2cIgh6+rkw22hnb6JVqfq+HBLlHV1PVr//iJJZPdVXy+po1uCKF5YxHEnvtugGSCpbr
ke2ACtqZLiCEvbISTmwAGiZadJJynOf9+XnIgVYUABYN3qEE8KI3vEd2hXWji/MnxTWQkEDvyf5H
odtv9A/D2vgHVGMO71KpVWKWZVJLG7fLdpPQ5gUcbS3G5FqXa3LM9afn0kCxCvvCVLJhBLj3qIAb
faX8yI71ORHDSf+ay+MWvjntEji3QJcurgh413yP5JDlRLUnc5Elw2xuTAaPiXGJghjLK4/nELNx
x90/8Rrsr/QrcVG4kkwzuk4W7JsFdpbOcLWArsvvEVgl3KSi17nTP7NE2Y7OJvQBKWFqiMbT/s5s
5D35aWz+j+RvgVrB1mZ7MCkK70vu3gVzUVJfEBDJHC9zh0YHw6rLkkz8UxsymOBFnWaI6rHonaEW
LvYbICoz/Qw5rzSdTR41M0PNz6cj+mxw4Dc18l9BDH2hz7WxolcY0mbcVSJh0J70J9UvtHqWdfAM
n8XLcP8BIw3IMnid7dl0/5eY1FjR6DUNjiFppUCW+n4JNqmeIk2rHDf5o92lU26sI9GiA3PdxKG2
ArDGxHdXz+ybYN+5pMQpDndQqpw7isxiD6H+TpmJsW5lSrslgzovX6RyzWzTeoLRWTGW0aSNNGk4
TJNfbcXuGdtsYh4GTf7gyydkWeRGwG1WQZMH8pfefW4e8YQC3Chv5DuKIoLs4cXaauQhmKetHCgA
HUBLjTwJQBqaIczh9bJMNW//Jk7g5V3We93unKn63iihQQUKRZBqUn5ttU1oH7N/fncXfn6FciVU
2+GcezRtmxsyN+9zf6wIroiwEeTJ+mB/bAyNpLvXtjET1H7MnNUTUV2jDPH4+DQdKqobKcJNA4lI
cg46/zPOwqPMuKoXov4J2OmIG2XcZGCwR0AZLhtaOztV3jUMO6kEGSOgwf1AIs33blRfgItXSAqE
mjVcwc//ePyY1D1IAQVKfTPLnwTVzBkjciob6QD14C0IQfVypvyx5vUXlVXLViRM84zolQ9f/y5H
J/EtaJBgcKgNqRX6D6IxUM/U6KoJdEmM8zdgmnRnlMlDRAroG744zGKHtreYTSsaZqC+pArb2A/v
osUfXvIROAQTT8+v5VMnNH+2iDl7ryvRhiY8+u2Wkngl2gZuAFzZw8pr2v5l6dc5qp1L8q1tKigK
7nZDhH0kcOratyJ7ucE8LU2Hzy8UCVVY2c3VD/OgqLQs7E90qBILhglY1+eiYdNxLFxlycbuVCFA
3X7QWxgXuBTdhaTfhe+KJnqTQNJL1J9A83jbYOkp9S49Ey2zPBF+yhvLK7BozDH8R0hu1BLUMlcA
i34YYXB9ZT04vJG3dfOBpQwMZLR0nAajXu5BCGUZwF9/c5g4vbNKvEsNzN0+C3ZmwypLuwqFy6e9
hK82SzBfvrrzItsI27Pp565p9Yev9xqIqhJZ+U5dKB0hSWvHKhWqtFYxuIiwTO0Q+eAtKAyz6f9+
sgz4LZ1zMkcxk1ny3rZ2w7lgkQVVzQ/sddCeHwp7zmi6dJAg1fxnbntaVBE0hg9gCNoz94/JGOn4
+c/w4btiuMkZQDEmZv842RL8dwZnJRv7VmJ6AaMSb5j5uqHswjGwChTVpsLmZyXp/hQLE4zaO7EM
ar35QteeCuWtdMVqGNZqc+PnLGsJyCUxltdD5hxmStfUsnqVkze0iPyRsD6l9EQQG7O7FS+t4NFG
BMpLQ98jzFZrzbsfC524Ik+7mVSpo9R3D9LzNhaO/HZUew53qY7bQPxRpzsn7e0+2eWFZl0lDJrx
LunZhiCFUh/GeIlnN7T38eaVNgt6IEBB8ZMpON7T/2+vxXeVxxQRauHkcdlFjff53jxLG8/oqSIb
aCKGhBBym+njfeFr8DJu5ndCrvmCDWF+Nhgpgyvv5Gn5MS+ldMrq+YBXdvLTx6d/M/L1djCC79hv
Gvm6APCn1ysBpSY/ExvaU/aV6Rblb81SkA7nQjakL7aRhAeEHXlvrIYTWdIX+U95I8IWULJPKUFD
PA37dteZzsb03Oyb1swfn2Gl4PRyznU6Xh5ZEpgwMz5Fbs4/wZsWjvBCO0gYwdwnsycFIiJwrdJS
0VIr3x0LKZ+h458U7N3g/baVXQCIWALqgkUS8D/lTFAZuFvEVaaq/7ENhFqHp5qNqxXREKDb6G88
wufklhirFOZieVxfbNoxd6KI0fh5I24nYucPA1SnDZ+Z8KiCMjoZ78gLL3RxMgI6iALr90xRZP9d
7GUgDCaTHWpYz4jq5Myt9Xq0mHoyVgYNL1rkWz54EGYKifo7q0zN+/RIp4CNlaXXqWO3HWoayqii
1TJO55ffEzY3ydf7J+KGLvnrYCT8HmO8b0V/MhJ223lcSPZt+2xN4zaAhVVfs6QXdODY1z2zllg2
6NSv4xJ2PRLNFdjIBbtJLBpkKzdcnHhgqQRSEnyr2dLFMLeB6SrYrjVwLZr/1u9XYVTwa7R+8QlL
tYWeEThyTL+W4RcYO+x8hI3HX40kPC+UgbIx2ONpSB1nnoEIvUPQ+fi6LdTMUa0HbK4CICUWSRY/
0wSd5fqa44jiAh8IpENdeOWbgqT0lWOo4fdejJRgPol4nCYzj3aooeuezWa4Nv1qyVJyR0LQcwrK
/R4EC/fhXVatJvKqPS5DZE7aPZZuNosiBcdQDQW5bQ3c5B37ZD6flEIlyDDyEH4GCrY4dQYEFlyu
tcnvgaC2KDwfAG0cd27rNaasEqKMITB/fhbOadr7XwP/gZL1Qxuo9x/iK4TE2/pOiRq0Xtj84tx8
F+y1C2dkl47Va7p3LwVaifcwp/s1+CorQk+Mb+rD9ICqAcMRuGqFTw8rnq+F0T3jCsgxgJ6P9JMi
Kzlt3OD9tWFh0J5ykPPjcy2t4via8Fwi236HaIXBJYoiUuSLMXXYYFDwPbS/EInh//VbOmbQYeE/
28Iy+eDCMM9pit9FhviF7580Med7CZJUbu7BPgBJPahfHA5Uuy95aCstq75vbIwq5s0fogahPD/1
1N8dQs2/1kYaqe9JSu5FxwYSJHt/A+tWGmY35NFpEpqpFwIavCJQKkPIk27Th3cnstfx7LgEmMIo
/r9wjPQoo0E/ImG/qTtLG6GGZFrieAwp2QzgC2AS5gdiAVapH2oVXwiGcumyJrjVDI9NOExccZIQ
bezVhAfc18cQGBH2oqzp6m+Dv4RVZNHPtSGHEDTcEzmKhHFKalGyNMoTBJvTz+faZxh4o4qxM0l7
RWJQQeiGk0C2FAHtsOCaKCuRn/RcT6N9dmBwV2fFW48l8VP5jsICNcwFn930hsExQeDd9Grgt5a9
s+hvRSaFIU2JhHPnmAWJLgPJTQBqM3FS6qlo3zF9166DmaJyTqpbQ8pljEfs1hlVtQ1NabYQNXKU
GnbD8VuTsoRtT3Z3Q55ouJDlC9jxsPfYMgW8eOef4TfQM65UJdagQ5qwTl1igio+5RGatq8jmXJx
8FzRSScX6LQ55PvnsjJk8LVAEBmpuPsllPfz2zXwVAc3QUiqEUyOiLYfRscLZAdn1mQ+qVqd9D9S
pQwIKEt8gkNWAJHrDJh5LZlxKJcDWfL76PEfaH4TmGV05UqRCr6Zb/lvPZJSOF6OwTdVQpZYduM7
KkWcIYToBiB29fjV+pt4vdprTDDkYr1jIyhzNUywRkFLFnGXPIe5SVVelmm9s4D7NVoLHf0xZvvM
XcJs1/mV5cICAlebSYgpm2fGunptf+3vxIOb2CwMEDrPZJ9zv+DC8+UMml86spe6Bnb1bwP3Pqr4
WPNvRHPaDvoOAcsG2rftAvXe8MOc93DNWDuIYRn5PkxqSRTQHeKrMyVU/l1U/YLa4YLsbqnCBd9v
OhD3dQbp4BPcDk7Ww4OoUNEuLSgj7zBL1914lvJLRhPGkaQddXDUT079GYcGVwzvH8ramAWgouG2
KxEFWIYfUcUTJLwu34zfa3UVjk9oWEnawUUdN0sWpA+5Fil2tFBuaIWOiz8rLQ+sh/YUGEiQNyvt
1Il9D3n3dkqxqJY2SIrP/z6ojHYkZwmovFp2iSow60ZCnZD6pgxjyy3yc7O5YPiVbSeUgHwIKpa8
WuoYvfJ7Qa2b0r/b+lUfB2DQwp8a44Nd4+sh0snRUrpRZU0KS1zl7No+5WD0VbydLSZOOahtulCI
G8IU5vPIvx93Qk8Lgq5UpPyphhJdyYUAdhjAz1I4Fe6Ks6/N7qOVmyyhGYGlY0LDVIdUzmon0eya
KOpBbomAxbKCt5Dt3F3bIFgRhGNMH38vj1ezGnfEgbJ3foGPAUVfwyNDH7YqBytw6VyemdZkgqYa
lG2akh5oIUAGSPWd8CIvtI2hCDaHbkquTj2CYqaGYUMJ+AmLDY0VgMkB43JmBJCzPA0mkIq5T9WJ
5MOR0pqq7gXuozTgTOFVuBdbOMmOP7hLPpdvsmsX/ZWuhLoQyWspyzUIB511NMPztv6T2IqgDJqI
eAiZRsIdhqv7LmdJj0C5KGXPlFxpXDgYERzoTeXDS1k8igP0t3Vs6Fus2GDQXwOadBAVIxnTwhNy
LlFQUw3nRK+2rMMPQY6dCplzBkcH5xphROcHsvis+VIsO1Oi1cdBr4dUVe/DlccchdARXNq9dOEG
JvSf4c1k5PqIQL70um1SDM+qXYveSt38nHx+/YfTEDlor5cOR9yYml4L0NuWVnUNfdHuQdze7Js3
QmCK4rmlkJ+64CvgGODKk4ETk33EXmbcJJCteT4N9Z99ONK1Qy12zPprq1cMyMZEZhm4V5bUQNuD
Oj4Lc1IqRKL8/QY5dO1r2gvKzN8sNngqyay02+xqXicJRREnfH3w3d18K6USM68LF8Alo5xvtzU2
hrU0dXirjnUIWB7Vw7RFqVxPMXT9hls4KAa4Mh1aS2VEdBemVefWUm6P4Rv3POf0oIx0up+7gKp3
DwcZGdv03VPSim7k/uK7Mqww9s3eGJJtqpIyTSiWIzgycnNWVaX7qr+Yqeva5lMau5WInCYoVChP
d36v+Eq2UPZl4/0xILxmExX3WdED9vlZacseHhJkCh59+DZSOPqy1z/6FPH6/Bxf9E6v6CinStFN
6sbAECaRoSIGxdoE9ZhJ11ezch9wZLkI+1zOz3ZgC9p4MQ4v6Zl5dJhaS8YjAHkjy6mr8XXr9yTp
fG38c7PsuFixpt/ZfBxGp6yZutve0sgSytMbgDpmVFIEOB/FV7oGM9yCv3uIL2ZUWLkqQI/X0eF0
ktlrAv0QSUOUsPCZcMtI/AsI10pafTnQjsVilxxKqKiRQqS6K3IoVVHHDz/5IZyzj6bFAIKfyt0n
/cbe16xiygom177T76YpVnqyZeE7CU+qMQ1KneziwvNd1EpxSwr01szzqr9u32ddhUCD5sTjNFav
Zc8I+KCg2WKaXBM4es2/TVJOXJxOzD4EsntHAiOSs+iR6y2bwlg1SXij7hnNGzfaqfVvSE5a9m4Q
Xx1yt0cE8jeBLIu0yV5dWzZiw+kfZIdnvH3wav0zdvqq9JsDB48TLN9IzvFu/adsfS3xCxWcjAHL
QWWWmxyNm97Gljt/2i10PSPiRjddrilt+6xZZA3Ynhnz+yMD2Uaksz46CQrxOtguNNP3fQbz6B+z
DdmCTu3R2NHKQthmLZOrswPIUXX+UeYIsFFzLFEShGDB5xqkfyvgMK2uaQAV7QMYMCaWaA9oMCQd
KMK/lygYD+41GwxD/KojBVondDoPVLBbktqQ4JVZvPJGbC2WCWCm5Y6lQvlxaai5Ux79e5H8ZtPL
6Qq+ljyx/RCAvGUFJywsYW5asDKTzcDruVeN5fvsy+kDBlLcO5scHjW2TIz8Cuz06Cz9xLg1nrSU
wZUdwa0/mOMZnfn8fXNqluUI/gRAWT7yL4RB+yuzAer+FrU3SzIfQQHzB0YxKfyt56SW8QVvu3Ey
m9c72pITv2vXlBWFZEwNp2Z9ULIaliH/Ia1JcFzgNqpRbHVp0y6urc7lJ5QQY9x0MPDfsAoHzeMW
A1lKIZxC+2wuEbVssgSOGooCSwTReEXc2l3/emZqK7bpqrCz8T+VCgi8MAQYA/D/fJP2b3HEk4vB
5zqDD2tAGW3BNUIsxI6xfLVIx+wR2NmPxOgxpVSaVF0AdFhBoXwPuLZ5k5h5Rllv8ePsYFTJp2s5
uzNJzq3Hpw2nfLb0aMRQ7GSBv3Z+R2OYbw19RWqzM2BkFMQAjGZITItkW100g6n4LTwdUCarYC4g
JH5IBbUopKAmv51d4OU0ZkVCficx51bMQCVMhw+hZgLdwPIuutUWAVwpHrZ6kc038XTRsyWu68j8
XisUiNqRUbukV8uMvFY7zsaL2kxC49weysfrqBYeYgbUFcVOrtVJi/wBEABkmslbJR6nY8iEYFRk
BfWn54jKtTqV821C3IsIaTxp7lXugN5W5Bw81/LRl/aL7hUUrVunxnIoR3BjVvMkL24Wwkxs5RTl
jPmlJoKDYnyL2401+t6k0HF2/+8TS9ZlXhVmxrrcUCY8yRHLfSnTAZA9C4WQO8SS3TToblpL5R4t
fD44tdCrtOwsjNsylj3lvxsg9WhBvp7LS64NwiJRXPr+qhBPow8dqzdPaWVkEe1J5LUglpgPz+E+
WP7YJGXlKKXEO5unpLfx6d+1IMiMZhl6JScWGV+4mIN1NTclGR6AElRimYFvixRShw7DrKbDMAgI
YoiXQYCw/7xpuqeQl3jxb6TY2q7mmCwpigdvN09uRGBJ9ufQa6G1bDv5gmrGbHxw8KJZN7XiYTVN
c3Ck1dQWKz6vM2ePSSjuDxYuKeSOr2F2p5etQoKNbw/2iOSWfmhu3PJEXWz/uvoA/WuNJEesiRJX
YwZgoqRgxY6K19A7M6Vg8nyoxerU1E6wj2ekODG7Ek4kLzbnBbBKIsRtFqrOmUbRmc8PV1ZP453p
kM1YW65beKUgmhW7dV/cXmxIYHRibZFvLDD+pcwTFlsbVeNvsm0hSb4n+j4q/Xtykwivc5JpWzJY
imivq1AV1jWWjC661ss5jzs7t0h7L8hT+ikKDO5qSepXdxK8rUMqFnkOslgzVhmCOc/uBzJYdBNz
1OLkpgLee6TskPOwdIwklqPQ8C6mxAFOs69hiFIDg94NWoBMNgA+ph80pZzqHfTtt4fwMTsslvlS
2AQ0SAXZgMvK7BAKnP3gfQR3owjLbb2h0Z8K8HUty7TC+Y1OdjEphMmLwBgx7Au+cbPygHFG5eUd
fyixWJ864dous7pGpjaPTJCAkw6bnLS/qE45cOV6XcFVmdQVKFSDTXg1B743sFE+bwKaaKWw4WWZ
LyFjCchTOGklqX0y6oIta64Cftumg2pos9dJ4vFnQXYqg3A90PBCjdTQ2E+SM6333+W751v0940E
pV5QrEypTJfCMnWjQMompp5F97lmFBDhp/dM0zXvCKVWutxzC8sMTpOnk6EPdBdts5bMQxK8oe2B
WLVoqBeemGAlgvi9s1WIcliBeWf4PGoPq6qozn7YfWYh6TlGiLHjWB9kIe0FWYJEKp/xeCny+6Gv
pfbvUMIBJ+iOnVMBiYraFrF5N8u/HSbaa1tze3uepG8leduFULi+fuP6t+B3Xotla1Xb5MDoRffW
VMv+XPA1myG0TWgsi0MZhV27yHBKBrfpWvLRxWLRJ8SYvyal9IxloKsEI1cPtXQeFDgUZrn4YL+C
SSBLeqiZD20JjUAv2QSa4QKcCKTDyso6/+BJOM2SET5JrUNp1uX7lKUFvuFa0IjVz3kQJkWFSzWR
m4AI+CYQjEugBFi6pToTCeff4kwXo9ejPTqhlb1qVe3WxVQCx5U503ij9X3XeR9gdl3v88H4vSya
++ZRMMHH/oZ4mIeUgZfYa06XvxrnGDWvby2YHYH8k1heyBuNySAN6GIFbpt7eMB1suEDrUnzy6f6
z434Gy9E8UOpsbCKp62oJlyy6FIht/Nk3MwNEhNlZxQqFxFxKX6e8/g3pzcmPFPNr0GPTzwI7mbz
fpmvnpG2wDQrymtu0BIHnawmyU1efmrjUaybypfDhZchQuFuuWNy9H07/4Xe41Er8oJ8rpLHOZzX
w+FVtAYwz+wWQBKS8ZiBjc2VWTwnEC0yk1TS1kkfVx1z8fEoYd85GAUJqVoR3qQxxSL1h2X6EyrN
8I4Eja7bYxSN2uSg0AvBeB+gknQ1YKEv2UPtQWPSLnWUuNYvaPXULGLRh+SXQtzVPPinNtyF6a6U
L5Udvrdez9v6/uHvroCxYRWP+50CkQ1Nvt2O1ujIfU+vzUnVSTF8kNr50OgOeLz+CvEa7zqjOISK
mWM2bUeNKkcTPPy4uYUG7mwLIDAaBpYMg6umeH8oXFSXgKLkd7sREqGoZiLyqyweUY5/kRhh6Vww
mUrWw1Dq5fdt5DGqUtx2z254PjDM3DfwgqpczgF3BOHvO5+W4U8Y+p1WJOt24AchS/BJMKCD7fSV
ZWDAkT1WXZOsV6VemX7SPpS71MH6EpqLQFAqCB0jP0OVN7hjsYchmxGDqB5VnnrgxkWZCVDx4Kah
TJBiJAHRvK5auHCurmcYtxZfZ4FqL+itSkH4hkO0Gbt60FGFNIyd65T+9CWc4HwA/WQBPNZ5bi1g
l8GjIS8fpYY7mGQ1RAzVIznmB+jfbaeVHeqRgfwyIw+KuL4Ty4/gM3kIUjzlBrM7ej5INu7NTXXR
MYZpREouvk0ebJc2Zo38W24MFjuIKNaWv2HPyoHvyGVmSGdYxyMnshk3HJOLVYnS5+wcUfc41+My
mZH8qFJgJQrTEwdyLXJvvqYF0Wij00Rn+TeK/BWCbw9vjpSq8JBdWDwuSHKS5xFTG91wMKfHE5Bd
ZEUbf2Nr4+GBdvjamo7nH80VBLfO/4BS2kJgUqWW8gq0Dixap18ywo7tNeZ5e6zx1ykCj91J6rJ7
YMMNuU2i67yBIi5fh4XIUPYi2uS//eJamLIN0jlrhp+cNsVbYhNHdq/ex7NZ5How87F24lts76W6
ZtCducCq4fnZlAmcZ8mJIkmI+eKhNs/QKKQ3Wthgy0cUf2gd5UwC8ITNZC9rqhm4zGQ+BD2bD0rk
bBUXN3iumi0BdVHj44xRLw+0XSeBxuRJs+Hi5WZnFVPboHnEYwnIotLAVBmUeK39QUabdLrmHyBJ
M/v5cSDtbv2QTt55CT6u8ORo3DAqx2hB+VAmGvC7bsXrQl59Goe4FBq4kDfufVfsIHMJjWXMOCjK
jzJvSNhmO+bFslCa4oMhFVLGB5EZuIBtvoX5aYS4dlqbOPJ5cKe9Aj3exlKWTW+HM9BtVKMmXugS
6K8POEcikkEndZQqKhwodkOuiZtQuXUp7VfErwKXIW0zTc4xycEv/ATlmk0MINdZWtQtjocQ76JC
s4beudP0dAX9FFFiuTRm4Qmi/BIHlK1MG1OcSGkJVIT+Y2Zxyjsg6uU21YttJdsL1OLDdObN1/NJ
nePiT/7OnG1eOhk5KyShev1ZuI9CDCxYBfxb62N6UxkM1bbbihiDTmKGNg+fmkF3YodcxOZyz/we
VXGNSwyTz6dMCe/EBhPp20bwQAUXP4OOUWyFxGsgUUthc6NYbka/wAPszr6JDQcY5UGz4A3zNcoN
7Ms23QlIUsuYG3iN095ASguhgkBULDURdFVO7+HyjTJ91vBbADNKmAZMgjfuBQIhpP7VTDB3ZsIu
xnU0hv4gIWskcjz26QAf3Z2or83DTA6WifWYErpxcGgjvK3rzRkohEZi4J70jMQUVty0SGJz1ibI
F3PmRaR4bNzQL6Focdk79PjRd+XVM0jQMDudzqApBhpEOCBtBw1nlpLivtMHPOOwV9OGJFD393hs
b5evkDfT83yBT1jM49s4a39myMAsSOu8kM4CckyzZ4sCOsC4GLTZt9Nt6NoyM3PdU0WsWR7g7R8I
fv1bFhsjAQETj8obE403hSgTuD2y2QGAdXF7NVCSjm7rPuBSK05nZNYilapgDrp0jlFxzAMveeK/
+fY1rRw1cvlpf/F0jaLvL3oiWOnBNvG4wCCEb9HS1TdK2KsAIEl7S0NYhROPDT8XBmp74SSvLUOQ
GS53/DVGlHNlA4ssh+ul3k5IdJs0xj8jTNtv1WlXNcutjP0uyvUdx42tO8lcqpoH+/pp4ApD5bh4
bhPY2SN36jym81JaNRmyLbUJvHjgsojPYgHKBtLA9DgQpHkbRGji+rNAWFIjt2JWa3/M+1kEUJXm
dUvxmk90iyhFguDBGjeBl7/O8EMUzWyM6g/4FcjA0ObvklJSNPh59Ffczq1147xexJPfxwG0GQqT
ft0BZM8KuXWnFxDNqtfl+2UVGvKHWv9mbcbJtBRObC/Gn69XOqXUBP7yM4VpX5+Rzc/A3AYqEpHb
jwEdi5AlxZykgz8wOhulTizfKk8wbDXavmFZIMdU80wm1gFGRwAPMy9Sgx+uZ5DviNl/QTC2VaD/
imj2MM6LC9UA9vN6cfSiUNMlSw9kCXX9lcvCoCGu5gr9DE2Z9LBELqyXmUDAl2D290nSMg7X1ZKX
NcMdBfeD2RvD2qtTYNjvlYXKTDhdKP/bC8jrgYvdAHsGIrAEYQnFY4jSD/2spYgmB+L9/g/KmTKt
HVoW6OjJp6HPiopsNPfa7flhEH3gJIGddGapaBCPE2qhlE+qPgS/lCnOyVjNVYmJZLeSHHXjaI76
51GvYqadZLcrT+qyyJfNNydEW/pIHaPLTiLgLd6Z6vUaG+cOcqu3w5GsnSh4pZj22vNUpaFUa1Gv
Jfy4RGCaxpmV36RkcRHsoJf5HUbpJgiKZLNB26P1g9c+1e7fnJgXb9szIWYJI9Fp9VmGHnH+ivPy
en/lBQfZWVd57THaKxPN+c2+i9LUypD+4Znx4fQWKWg5MW6ZWKknKicnQBUXvuRCy4CM8zXbVj5I
TqItJ4tFwtVXYPazWwOz42SK+HNkxZ9XLlQWEFMIP3j148Mi/4cDoCiaGBi0ejdxNVfUsByNET4f
sbfgpM6h6x2u5b33W4G4nZVshhbPsy72yGmK919IMYt8ysyDFo9pEt1FkLDtHI+iR/KBn5pEmlO9
wgsISHI1BTX9mCR/VYcyIuaXZWsvkOGUGPb23V/H1GqbC1/HR7ZjPzaSe5azR6HsDjRRuQ35Kw2E
feVBDtOYqFpZUTcNxJ6+KtN6GINGoPY6G/C8lvPIrD2JClf46IyJfqXB5KtrkBFiCmJ2pcqyrcP6
/HW/5ERDyQED+a7q13o3oiyK83r0VTT8OIEHTtts+wxZBfoyVCWxGT5uiz4M1hh0iryfO+XzSiFT
7uQL5UFZfukfhVDMb9X6XAtgtcjx0P4XOVKxnAW0S4C6DXWMCKvPjJcSP8hyKwUfxZWqxuDboL8U
zmPp4IG3RMRDhsNY8VuyFge9ykURoNuVCBMPq+6E8euD/aaRZcW1yYhdbryGKLzSgjUVie1DKERw
u7wB/ohMi+rlsKO/wAxHmk8hf4Z+5Nf32ZOTxNUSHOQ5fo2uU3HhBh3+M3gytRBO6mVMHNBVVykJ
6IfbB1XE7CrYutJYOI1WdPOULiLMIpEaj91IMz0zZLNTbFEWDtniZhR/dpHraEdRE9D4cLMTkGST
cxTbF4rduo78tBUwsKISz40KeYh/E+rvdJv4Vw4jx1xz8FgGnY89imRwVJk7mQWK3dr8NyI3Cm8j
hZBhmEbq7JQrhnFVnR5n77IFBPnYBoYZ1aYCMg7idaw7zppIsgAABHCvZmU9uhfpdpdzyZztYMrH
7CBTh16a9/Gtmc0ZPXqlodJYZ2pNivV+YlVcCBQlGb26DS6mGvKLUJkfNJ9ZGdIFh6gWZST1gSVV
WaN/mSGMZ9zBGUix6MOqOF1ORAt9YMHBLO4PwrrBAznawgQQuxi6qQ02qweA68yyPjXPFcmZYCGw
W5/SI7DO0mDlQTEiM7VymdHX8R9dEOBCwGYS9QKjEU+FKSzclMMeFa/SO5aeaX91DcBRJcehQc8M
Mpble1Fivh/gpgap4FFc+5/gsUHTJtJ8AXqp6OD3u1fzYSMewQm98bCMqTO7SsjziE9p27tm5jTL
fZCWEtBRMzmtm59k0vPAGHMleRniZb0gNGxipuGSJbtX+wXlFhfpPTumzGN7iy4dGBEXRItiih9v
Ep3WMzegiq9A1DtOpfbzI38M+MCIbnM2BDGR5fekFxXMjGx6Hv1vLsTUHGo/xQ9XB1PAqo5jIR7Q
cgDC8WL0md4IIFlg0YRQ77kgYUtLXlbht9ruo9zTpLoL1VlYlWkuuSoFXhb1i7bS6cHPNaCaG7Z9
wfrKlDd89F71zwP+O2aAiw3kDEDdhvZ6TVhZb/eE++YLN3aBGU+SOaaLcXFjZMvSISo1ZbBYwClU
UVkMbkzgYxyOZpSvsfH7gAKUZ865dGn+W9CaS417UScnwJu9tmitfp6VEXkI6qGX5FfYYjJBfC9s
mwXyzp67s3payBKQVuylR0wVG9mH9pasAuhOSQ1aeJ4EByjZ/kkTVM5nVG+55JdkQYUhYPanqm3v
cc+QrW44QHzmMtVgQDLPGXgGL08JslELAISwjlKi1OAGSc8Zv+MsRNLHHwnIdmm1UqNLoBdEhW5U
zYATnd2CBF6aTnsaxxG7YpPsFQ5Ch61JPD8fNuwhdbamaW7RdE4kIVbLVhV+MKXkyURlsZaztw0t
vwtzNyd0tmZPK+ymScbuAklan7sU5uVd2TaztjQ05KqAmJSFBhndzD4omsjKL3WIczKvu49KRP4Q
cNW+0J0k/VvZ62MDXZullGRlWgygAfaFOyitsUDp4XrIel2z6dkgb+ik6nzSS74U0xSa+00Xtma7
k27lGV2d1AFh3v+tQi2Qv/1SL5XwmJOgAaByFebLAs/Y3Vou/mOD17QPua9MDHk8+A79lvFf3MLL
O4XzPxc0UkjU62BssbLMJtULKmzHeoGNb/W8TrlRy/7lAp5O7Kz4YSuqdlEJh2/YyNJid5b6pvX5
r7ipapg0+LaFBFkmtYQsu0TW/ZZTMjVuxyX/Zo3+ajeHsnBLf4VqaVPk+tEe+Y+5CRa4qnn3ng1H
hG4VmPKrYAYWgtdnboi4M2LGyBrl9kz8RpW5eC5c0DaS/LPygf4u3rTamXseZ7JU44TG2rc8c078
BGnovDn7YrPDfAwl74Fc08wfefEjavyTlWtmrqhMbusnO5eJ+i7si1UbSs64LzX+3ysKNCttS8bG
V95e8Z99EFoH8j1ITIa9IxIqkFCQ2hVg/xkRvKpHEIIEHfQnl/rDfblWyhUzR3oYFofzyBNdeoI0
hvqVOEqxPF7szwdVKL8z2YEyPgoaXMIlNhzmGAr+euiZ5u1uQAe7dW3u1jJVQwTHobqbZZgirJ4Z
HJl3Zo7+sF9sBNPed9odeBM9sKz9TCqe6s8Ys+vXyQUyPziuAj5QErdmRCx+zemjPdo27+GdtJ89
48AHqDc0lglNA5JPCkI+sVA+TKjY3ZIBGJXR/VcRufoDrVSfHGndapNXJofPKQdB1i3rpCp9qJ+v
OIjMK2Xxj2Lyt7hIPmQG/GYESHNjV8jzixFTvuK1VeKHWOUsTMsxcP8LNsq70FMzxqni78m/4tMz
5QxBG1/kDouQB3QkUY3Zhnxbake2pP2CmGJHzyt9QHaYDaoUjZ4uORB7v7bfodWbjw1BkNuOaB9X
CKi3+swt388apjFiGXbSVnMnSMk/+2krQmBonnGznMFzfqIl18EkVKDwhN0sJK1AcbQLSLyLxkNV
Aao5nZ++2lP+dt67XAAhH/FZ+p3bFYIfdu9FvgEuIiGflejKXsk3h8/oZ/jFoaDXskzXvL6SQesr
7ODOviv/tiptYlDSCZq9U8b+Ox4DRQDqAoECN4jgT56ofzUOV38/dPddq019AF4wngsSvUQA7xTP
N/yEXpDENnGAZxtH/jM76T2MG9iFqI65YGdP877ACdGU89iI82LPMU0PwKcjAg2ZsDshBGGj7CoQ
9YyX5bNLitGQjgWH6+0rL9gVP7OSLDiQV16mxyvOTob2KwmC1nH6qZhjDbb11KcVEpZgJvx1tUzB
thILI03hFCoS6dCIdWiNJ3P0/i6OsRWXSkpt0QtBXT+Vs0W9C7fMdD9eFyRpx7gNs5/H/Ir8kdXl
gkhhZYGsmtEZK1w1adU8HjD8Kn0j1EQsmzfAOYiPzlswT0dqcQQcFqwNVWJc+iE/S4cRYNt5DZlw
QG1s0NRo+xRrid8b35oTHcTOCsuE8bvcy/VH2l7lfyGAS0NuVRme9PeT60U9e+GXZglW4RqLTQxo
tbKHfKLzhBvNdyBlCswcIhneU63NWO2ugkjZSokXMs7hhtWokoB6W74KkcqExSYca9YvxQzfoDGQ
p20lGHoEuVnpne2ueffE8OlxjeI17idkORq8ZZOW5hqZ6xKk4CR9zxK57VnASYjlYoxmnenD11DC
yr6T515AJ3TWAV97ag5hwleENHy3XElW98wmbOtn8aB436OfLQ0ZKKSd0w2oni0Ig1L3V5xIwbVa
URgzQflm2fSmYbVkOYzw4PvNTgc5klZuWMBAF4zYTi9hNJrZfV+gSPFtU6jSMhSLPGyKylZTf05n
KwCD9F9BCAGec8pIwXX9romdkNLhxd2GGyMz2rUOny9fkbb2lypekzBiTOVjY1l+GzZ+PCHJUXP/
ZVDgykLNjiHbCWMgEErxg/rf3r3RCnJcvrSVKjrTQp1c63f8th33X1xbsi5t9TkT3knjCxKxqt3k
F1FTn8MzfSG9dv8Dre7ZC1vEnxjf0PASWMI4HBvLjuO7tCuz9fjtWP4CpBg4Pif/Hvg/UaUvioSK
WQ8O84Lxe9TlUxLUnwVo+I5a2TAAKR0o8k/2ElRThxJeWTeA3CMWpwAk7DwgXOxXv++djcsFISp9
DYVv9KnK7hL4rAlGiVPhkyCNHVMT7MB5pK2LBTl3sQxnTIJRcM3CDlIuZi8US01cwQHvBVaffhJu
UMrUMoBMQyMIYsqbolV5DLka15DgB1ojKMb4ejJ6GJC96O0YabKuE0E17ZmPRhYBzr/cL+2BXN24
0TX7Ljb7H5O4XhCyUuqFu8HPf6qIw5pG7mLZqMsr8D1FAfwXXDL60tb3CsFYX8W8aMbLgE4wBP9f
aUFr4cgFJ9XGbBuGe9WDBJkz+6JjcJokC1RXUViWK/51DSroOYvD9AooyGz6p4KZ0u1sqvqqWeon
ep7f20WiSbNhJ6Qqbkr5Xtat+ycNYZjkx4lTa7FIxVcNTAzaHBg7i6ZAqlWEYOtMbHnoytAnrAyP
wXt5qfujBTL7vUEuJrUrM1dsZGyC+/Gg5+oCC/tm9/gNy+vxnjPej5YDZTWypGqSM7wa3dby2F/7
Kj5h0ioWjbemgCC/xgbBYqHo2pgmKcqQsu5XyaIVycSL/yVihGQdnIJ80Ve0Zu/1EAFvxDl40Vo/
fYfxDptLu5fRnWqmQKRuxEXoIpyhvFuCDHsEL+QtyzbruFhS0yvv7d09srFsbpJZfn7bX3gP8iX9
7UL6Uc+1Khp5m3BeSJ+T67NmS4efYqSZYiJFDR66nMySDq9cr7JpSk0Pk8sYLuEI2gaJanyDIv4b
C9A0R/B3ZT8dwcOtYT9Q58MmZ8bZvXioE24AeYfvdbSB6E1k5OF7o9cU3pnWgKbU8rsdqqLhZR77
vELappOdOur94CvnQ3lodCmcZIsrxPpnJ5oTgZFul8E5XlCdiSdEJAPp6F0pNp0gTdZqtL5XNEtA
hw5fTMwOVbho+MGbTT0vzBONQDZyfDGVGJXcGPrH6pngnRWLqidE4fHSrmNySykrUJ8bxo87YtOG
D+Xdj55uxNUCk2lp87pbTBsnmHdr7ztlCyEA1GRDG/twpis7NDSW9MW9e0Nl3FsG0OaO0TXUyMLj
ttaNuGXqUMO7BVE+jYfwkOXjbLCWEl3jGvgY3e57NBMbKfNXU0c6txrOBX2P7kj+05YKlZXz8Tie
FlAufA73aTPSuYJrrHat3yfiF2GmzWYKlh30QICGbGjViNK8UlDNacMzyUCAhe1JDxuwM3USx8m1
xg4gKRrR90wL3v9phnpdrwx65rH4iIdQe+b48RbrbLUHMdkAff+dPwM8YKIINluirafeh5Qx6RWx
UBZw5KBYRWspotxWPnpJ+youxcgAPXoxtgcrcEYK+tLsgk4wWFc5dYCFSWkOH2ZiR4gGEDB+dht7
lKyuPw/8JpFZgg1PL/pb9djdnmj/wzt3jSoHDLND5w/F23qXzz99OckfmQeHmtqw9UbFrxlXSTdw
EHv9lkwMk1oTXxnsYWsx8LPyUMbRHVWT8rXT7gKU/LxSN9HTYIhwU8ZQmzciN8mngElkxa/r+kkO
NDqigeY3vEeYV1NMVhqaYgG/5JRPhJD+r7yiMh96ff0VpW8LOt1Ra8zZcOof98IT0efUCEdydhrl
lCHXTtZhL3sPbv1aFwZbMOPBoVLYl8bgb3lHsTZEumJfn9lEOvY8VZaVkvdcAd2BM2UqNkYr4VPw
AE+1m4DMF2957cswotwo9UIaaTAel5U/ouooQwf1mppmNW92MgesEIpIRrnbLac4x01Zebcu2210
OqweIgCPvrJguoMwFPmfDibbWH+Z4/E/VZxDjcbJqMCrB4nUn/vOv7YhuiV/UrRibflLwiCtSTec
leMEu5QHN/zq04wL/mwIm1rs6Qf9qZV7N/20gji24QS/0X3u3e/XRxdza4UZCsJP5zjyU3Y31p0f
l9XUMKNJWQENDTIM5Iz8un3h8gSeL4E/dnu1gL5gMNkg+2ooNdcg61hkasOeY/UpwnpfWebJAQs/
m1XCH7OvwoO5KnfnW/YwbsUAs2pGYysj0EUs8LL8ZTNGmqNoeAyRc/H0MvCaLvYhQ3j2GyztH0EI
CkaE/4qR7SWr0WVsp5kGWXMOM6XG7i8SmKaz918qpuGlZQng3YrjfPKwOIiCzYdILybCFyeEpN1f
DmWH4z/ficUCColf9jOJFisx1Wzbu2XaVTAiUgImu1s7uYuT/PRTMtQbil4/uULLBM1dF/QFhiPa
1QI5qMpp7KjKxE0YddFKwiz7/D3pbXqEjQtpMP3JdvAhisoBuwCbVa+nUtCh8eHJ0ppPldhUjC4g
9axxd79w5NDx8LaCwrboWRdR0TCAh1UY5eAInxjPA5JmMIRMQp6SaIg8KqXzPzuBxvnx9/hvpdLH
nf5lbuxJDpIryHrkLZ/Ll2yWSySeNJ0MXu2Jj6pwEUhJ/qRZO2/zUmpYkN7HFtMHNhyxjWdYtALY
fbDH9dE/HmSHfoAfb4ARXMxWrZxchJY0USpQufFcciO9phbWCgXn4EduhdzEEJlqdnJvr9g/n84z
A6Oeo/18zeLWXWFMHxPyi6Fr/77CxL8W2DkNm+jTK4eBnrO8/KRrwYvY49qOAXRC/UejlWhYgdtm
+84RICig1ceY3nojlpRKOp4UOYoPbR7cBlqtZj5WspFO0mUkbvBti/bkj4l5qDxSbqcHQWAZbhSW
Az7yf/BNfGqx71wGGtlVuw9cUOSDi2o6PdG6CBmyZhMqaapRQGvDlXkUwOXeXbiLmdY9yfQdQyGR
zy+n/e3jFVJW5ap1mTuwa7dwHPyBMZi7RqNDOX8xklS1KbV5SXASM62s1W25l7kNGn2kscgLgKjf
FvU4FlW/k1FBXDGjncGwI1b/lqUN8qTmvjl5s8mLjyUKid/te1pV8AyBY6QJNvSyrl1L5E9dHuLN
1dFCYrBFtDwgnHpyTa4bcIlecVWU71K35grXWXgkv/etY1e12zNk2TYlVbPyxPtYEf1/me9cMLrj
d36kV9JkHI0D1SZUbl6FxTX3qsQHb3vdqWWD7PUZyxgtRPK++DNwnmyzn87OVs1Rzt+yrOm4BFF/
XzhvP14EMvrQK5Xd6Au7y0c+rsmGhwoomhx+vYMmajADJ4pelzzessVgTX/A9KO45nm6OApZraF+
R98muN774BX8sWcfPHCODnrgkkzKUpOkR5Xq0kQZzaaS5yi9Qm7NTl2j6hiROd5KT+J9T4ySObTp
++HJnhaDJOYuKJ0KP6BnIuKHOje3EgMxd19hZSPjTDgdq1YhU6XoXHKDwYIXXwOdHqLPx64qZMs5
FNjDDG2aWeBvDFcyqguiV7C2DgwdEcOmCaCDepHMorQsgN8Jt6qwdYCdkhAahRyatFYPLOL7NTYI
qx68yHep85qMoBnnVSeB3NGv4+ZDGjylivASwTtit052DQ5qaQk+GUoSVtBNjYUianEHgIvpKQJF
b0QghK9hoD7ILITbTPO5rwwRhOJ/hlMaGki9Lht8BV9yUxlxggGfKOS62yhXf7zB6G9M9gd08L90
QPl7LoG95XlFKFHGlQvCMhqhTag9X33ti12p4qWdq2Ht9ugF3eNZO5xlDVnc0HJ2hWBTU5MuUirw
Y5AKCichSWPG3sB83VD8fgPVPZooAcwZz/hkp4mpzL0Q0e72LTCkzFzqJxlPXe2UlGsm/lPl92zs
1xAr50E7rf9DFX/2hIDuTyMJ96ODeKbtM1JS/p++p5YWS69ZqxJ3bjjdhLC/DpM2LDB+ROVeZDaw
euuPpGO3Q5M4fYiiw4OopwwqdFxN9WGoygBDCO+OPMvT/z4R6aQx2S8VNNwY9aKtMmip8+rGjpk2
D7bsV9AoITtcg9mInf84Nis7PqU/7PISAR82O43q7TN7o1OA37XGCSH1CKYaPg9qZwhFuxag3HOF
WXmKD22UKnFMhXytGIlrYE2ZSiW1AQukoScM5N2zazEaijYCD/rsV4/v3cp+5j/DCdrVWzuBj7lW
MFg7UE5IqeFSWa008ycoHZNSJ9rdlXaZ94pJ2D5VYtog8YWU6DW3Dgpljntb/lSIuFiF22tcAgVT
S4CWvTS08Floq20g5Q7dbsGmLeEfTuhleOTpyUk2t2jlTxfXphTfTlePrCByP0lbl/7QHTFYh4h+
jQIdcbaL2xQIGbxzgT314ftuvITKdVxVdmhrq60nJFEkVszqclS0lis9A+hzV8jRLJf963XqV5bC
n7BV7LbZQiLFY0dQSxymKbdU2RVIUutyatQhBfqGOzPGZWzKyQvY75+0bk3D/JBkKoDphTxVyh5e
w7CoY4xM2xai3CW3sSo4BY5ONnZuvezn1eqPYqTTMt/QmU/+fuvNnhxhXeBwiJ1xKoD+5KV5uMpp
Nx1JkyKJ5lssh1+Tz2uxLKE5YesN3TR4v3v/Q4TM2PsaJtB7I94bo5W/+mmImwPeFROyxnRP2p6i
TheDfygM7zxVu9q01rbZz3MV8wCJQhOLYk9ow7hxBzO1zRDYyCrtS8sTbq+v0MAmOBmWNwqhHNm/
9If5VHGd+Ut+OnIV8sYV3lw67A8uFJ/80LkifTcjJQW2S6uQeVShE9ac63qRLe0TqhU3hvR2oY11
TySTZUSHay2z/6aO1zlnWr5421ZOD4tBLdpGrvyvH+s/UzFlUBbf50P/w63boGa4gCx2NEfeQfLt
khamrJZIfDrzMBZQlPPx8PcnOEM2CQQQdpnCmltJGgi3OCT+hR+/+wkM8YbYscwJRkWeSQugmyw9
4UcQ9+L9uIBiFMzURPRFuXgtYOKdpXiz4/Gj3wYdvsOxgeFXNFU4K4altKt9poWztYmea49venYx
1jIU6yY6R7hx33jg5eHv6kl/fr+5CO3uxWRhCEDYVHdrGQp7UoXH/b7iaf61rkzVDK/JYphYrlUt
M6F/311dhVHSD6bdij2bvUtFGJADZSRv7aoWuBCr31tRMJK3Vyg0myGQn7UU4hWv1idMFgJznN1R
I3zg76j17rQS/BLgPqTykVJbcYh4WBbSRMBQznKilYUhvWkD9pP0u4gQkcxm9Bn7hKPCRXjlYJkX
aA2hw5opbtWo6ar5HW/ftMbWjQx4A3r8nCwbjj46jgFDNHOmMoXIVYAibWbF9rC80Pewyj/WlszO
wMALOTVmT5LVe0MZ0kCKjOsSw10HwCEAT91kkkJYUkUwnSDOcgorLDx0+4jCgQUXOeF7XjUD+HST
P2gDJY44EHlrRSkWV73TW4Ze5WsLJ5JsgEfDjLWoxUJMxiRhx/xOPFmSoAqJS8bTjwCRXVas8/Dd
sdaSvngDVGn/b11bSiFYZXXhDJGykFEAtrjAhBLPNTDivIB7ydLnxroHe45qMt+o6Oq/f6kWnoKI
aH6YbUPqi5a5ARlLYdngby/U3XlSNBiUiH5Tio34Sun/DoWRbdnj4uI39Tt9TmHmU0J4SBZP5NEZ
mH/PXT4l5o6IXYrqzENFkSlL4L68d4Se9R84hev98r6WeFB/xOM1BDjAx/o6GbZGZABPcdCp+PAD
THSqcXF4Yz3wF6UcuTYxyrJmKZOuZu0pa/5E/Zwu2orFbXV8zY66bNo9LY0dqdOpMiVei+6kCrH9
FmSNIIdcD2V6B5Qao02PHydhY4qoaSNaRsiYgvD0fSTpd+6TXsj+mCIYrXKFS0aAwdvDyeMG8PUu
oP7hT824M1kdmOcwyZ89l8EA1vinvkk/oH24ygO8byMP4wCZot+hHPmYfwxvI3NCIe6nkFltOCGi
l2/zz6FHf0kEB7PGJAwQ5Of6MvxFEKR5NkAsT7En7jAUWoSsoIOXjU5o61KdxMZk6n/i/J4az87q
PXwsm/xMIrX9JqZFnYFGsg8X/7OhwyxIaS5VrLCQBjdxMVvP89h60VESz1oWYxcc1MyVeOEocwGf
h3gGPMGoHhekoWZK14VZ3irPe0rGQ5/qKa40mrTxdgWW0UQI5cfS5Wyt3UOCR56QR33Y8cc1S84z
nOFmBCnkfKTmn0XLZKJziHattN5BTVcQ4c1NrVVoKyryXL2dm/uiS/BjH2mR2uTwj4LCMk/X9GYy
vAU0A/uZ0HoFYigPnBP+1zXvLSOfZ6F2qiIAjB25AAEsDL+fE8Y6BWca+O8qODVxsv3GG0vpoFgL
CjHp8d9yLV8oG9D6Vynz3eOiOjZS8pdP80SFna0xkIerO7WGzDrIiqbwKb63KaCONt+suv+WPY3T
GjfnQRGdaXNIG7wf95MkaowAlOz0+z67seYJs0UbMbZ1Y71JeknHSsuTOCxl/9LxhNDNEG84MTcj
SW5ifn3szfCFkop6DzU4tsmFb/9VEPbBQ8hFzEUAKdhRH8/sqzrPwLNyrbGcr7VHvfAxUH/NZUGa
tACefQAplFPDVpCRnbvanO+q+VrLEkE+3BFkeZSXfpDqdLsUwX+WIqx424z7UzZykQ5eR3p70oXj
cqq04QCYm7NzxxYnxKkdLunmJLLGVDN2Zl7O8HsV/g5MZ6HR2x9rj15FnUSszs90FULBD8DtT6Ch
vP8K4fpOiZ8whGc/1tGGvIT9+d2YkAoWQ0B/GVZ6VL3z3nG/vp7Ay10agPzWqdFGy/D94ERXfol8
DdC7AybHYJGZL7BpGym5yTRW0KpUNN2jWk38rO+lRPl0AwkSArSWZwKDvaVEvr9f64sIT1tLy7Va
CuuiFZygll+iakwEaFcsT6kx5raMI5WwyNZSTU9w8quJKXxadw5RgcTCQKsKS/KV1fbtwG6tIP3p
Y1UqIjl5rZ4G+DJ691hJupleX1Kmu4K5JR2vTnMktP72NlkdUXCUTGKb2ad7troXzS6GIGylV+kF
Vf4RXKtuVUJAn1t+8dGGSLSIPz9T97fwHvpTZIQ9NzBXEcyTDYvEg3+Os+uADh1rz2pTyPc498T+
ZlvuyCK5ks86mH0qjEhA1oKGswAL9veBxndinj6DulFWu7mTPVjbQEGBGSKPvkn60epgklP4bG+m
rgDn5KG6Fh+krcXIvjm5jultKLBBfYwJ8fPAY9i1Y1bmcKaMcmrQH15MrB3jhB3b03st3/mEDDBj
n9I6/uWiy6pJYNOSGmBrkM1j8FxVH/R/LaQP5h0SqwI0nn1Ch8SYq+c8etRJAFene4dyf41MLT5O
SWTDUdfGgcgXc4z2nISJUsd2hXV2XjvvSvcUsSn5uIg90VcmO19hdiYolRpxB3h/9vDV+MkR7dSW
IN/6dQWnC/1AaRRltayQFFGsea5sDPLGtNVDCYbvnyb5kBkMnPztPvuQP+odPm7d2R62DkaTf8Pl
Y5yeIWG3zdTReHGdp0h9pWbuOt8xxMI2VBiiWzlG+W7ygLBpeQxC2bxg/2KUq1c+95GM+bI3efgX
dq99qTe2K5vUwQjunj554ruO9RmZHTV0OSRWWgc07q2JTwN8T9zr1EhfKt6sgcVMJCCog0YGzKRK
Tsdfj9PUwXoIKiN8GOhxvT077vii071ZEh1gwCE5oGsfgLT6AevFQ6H/yGUs893ZcVJCxIFMxmPs
llam8tWAdxY2jVlbDOqZvgMwSnjKAruU9nUxEpGIz9mfm6canZ06imSHpo75hnjJeec2u287B0pG
XCY5tVEjtfbc5oRBi9ZhV9lcvMr82AfoMWTQtcdV/G6OPXZedpirZygxDqqwDN1E1PlegRQhN6A4
9xUAF90HI9X9x7W/4Bv0dht0hY4wngDoH/a2H8dbOvfEHuscyqG4lET5Aidif1YurI+e3/2jx+DL
4pKRMQ0Vg+r2Rycg0fU85wLSEt8fukO5JaZBvxEkdr5dZJyoHaJ4oc/3Ql6pmmET9EZ40tsVBvlb
cEqt+yGk1U+i9epw50zlAi6jXppBNYfbZWp1rHNwWjDNB8kxNiIdPr+5ANfoOmrn2bko4fqFnJ4q
8QuJr3GMI4msWhGuw4ydSj2RpapDgDj3XfbH1qlGWqvBoxgBayWpEbcXXfwAsC7AR0vBu8P5UUuc
Snp9C/SbPL7yg4IpH0cr8q068LZB4Xgf2HTedlhioKwLEZErss2Ip+DKp8kzGY+6Ghil/oAU6bMr
yi0F8wOIX6zsdrl/7dgWlQl43T8W2qJBTbkv1ibO6b6M9Cxahz4OOJcUnHIIXcW41XwNK6hQP9Pd
V2vtv2KIWXV8frJHH+dZyYJHvRITX3OVxYJu2vqJMBnw5u0WjH/YuBiLVte+udK0ribtoNswwoz5
cNkTW+rKDxxJqcV6iqCj4Fi0fU4GHBmZLWm0H0qBwPKnbC4vFvux/q+n6SrBLBHtVD4x/IUtaiWW
m9kyh0x7JdGptasdSdEo/K/0ouNs2Wa1sJcs/1fLr3T+SHfFcNvu+pTSuP0trtyoP55p5/ZMLKcO
ZZk62LqupSof5IKvT4kX3f067BmJj7azNrmluv8ROk5nskPs3NigWYBSj4BZcd6KA1pATasGb33V
drcV4OE3KTScROgsyLfE0S07Ocegwob0hHuB4QQmecpos0NWJhM3LovGtXjdAc0iKPD8iEuDzWnO
8PIgLtI2sAQanieBpSj9644sWOjTJ4DAjo3xLwm7jIA8Mhf6cvEchQqQRi2HFDGDWkB42ICb2cIo
XBOdGWFnqRRiScg+HUldKWMkQa2SMqFdKuCUQgCy7Spid1N5Q+6ZI/DNT6b+LDTFrATHl87W2TfN
jQoy9Y5fYWvUaMPGnQ/8A8uKvwdBz+zX62fjXClv/dtUI8/ozvJtjfcB9qxecAzLxZlR3zSkRiA+
+N4MJED13t9zWIzbxTSTWkKoTzazhqfVDMcmomiVGk5fw8EO6G3BlqUclprsKvmHoYgluD+VEHYs
audHMhonYJDAUN7EW+9u8nuOhPe+sd5R4XLuJ/UyXPsFpx5Pgw5ufWMSAR3WX7v5PTKWH2jRfGkD
5gwdwlPnSrfPGcuhWKn2e6v/gXX3FolEYnX6QoUV08nwpshOmoLC37/0LiNKkEwJlcZ+tQaIiDFk
q2SIte2m7dbmRTm62QhiC+Eu2GgmtFKRLFKEFtEX/Zi3Kv4yLBKaMLL8hpzOEx+DRYbF92wvolLo
JVAsMrgS/HZ8JJewJwn36GmAW8HaUFWO3w1ZvScFoKJcyBrS22lC3rftUyfqQdXkLsFXrlWmrDxH
jj6q4x1397PXCvXGFYaLErxMla+fbsihOQPrxkZh4dLiVVtGp33xlJNHaTG5Buh7jyGXX7BsbDwq
nseZ3+/ER5AHqV3V5Ry9mPsE9vz8mN2oj4GB9NlmMC6nIwa12rO4IbInJsMfaBRw78zVHgnvfHnT
vWGiP0AXFqAHWfI2tos4nAaV/OQtizN2P3JDBDyfUZgXAv0h22bc0rIKonKNdR2DiHLePJZxRk/s
2zQkF/bZDmgecAX7Gbk7kfEaccWZLIhysTiVG7Eys+wfanqLwdJSSRhARCRO+KV0g5WnTx1bBarq
F8bQZBR4RFT3KcsVy04aWDf7yH5VwtqngLWDoTwYkWVEFJObnFlrAJ7g+7DX27fp+1EwPLDDH9qV
/mDZUh91bn/3gXWzpE+wgedbgykwXEHoaBxpLP54jDTphKIxMwQTSSgcWau8Fj5h2kCdJVKDW4xK
L/JCQyKNcfXFjwojSNua8Gzy76BAHVB6zeKvHwU2YdgkbgMVTD7NbpzwOTLjzaxglTnP210/Y3fR
QVBbNNnvXLzXtLdfl32fKqDvz8HOe7dQTpyuFDb3eq6lDL931hbS3bVmkDiwL+pQ1JaqfQPDPSsv
i3WtF3wvi/+F/DgrvywFe82eDezDQ/qSOaBntJ0nWjg+QxGbZWEIWSQajbmS7wV9epC4PvADafkg
lm6UH7x8QexwWuoS8ussPQegN1INXNp9CdMQjqDhJA05VPlytXLn2gEiJpnIZRZlgXk/edieCCWv
zZwFpcTGdj3sqx0VyKNFuAYXBd6pEzNHAUOJGphQlQ2NN50znVeQ7xwzu9IVEfySanUzCHWdYHzM
N9kElDlsMEp4WQlU7+TJq1KtLoO8KxIGKTF88o01kZfAI4eNkSnJUjR0fQMg/nlg35ZUELCZtGj6
yC6xAmRq0arDcdfpz9jri+OB1+iOYGPEa7E2My7dD6VYa+3eTHtZkQUygo6RbJwzld4JWEb5o+76
wbEXum9f+2FJygs3CnitIzke8Nafc5cuBTt5dZ4MKusJErMXvxbY2jGbQinNAuNJ60VnzwHtrFrd
/FGQ5Rb2OXvG59Wj992IiSmBdTU/pNZ1H8HTmp903xsvcuOPc0j+xvownH6NzIG6kgOzuIDDYNsx
moPftknOjlsgCoG2FmBGRrWqNUJ2cGTw2CzRGDttGDm/0V034ifmzRY8Cbhf7DSgY0liGfi7JhrV
75CKeEXajbEOtwTr/+kQULC3Raj5kyDYE6b1NuckZ7QQ9utSCCl2qeffv8ULHoYElwycbglfEajX
JkKSoC++rFMwJ+ef248dbJxKZtuDZ0vlB6BwsQH1Ev4/7Wq0fJ085mgSac//wBfYy1gKigXmdjJN
908kcsN/2AVk6674WGg77zpatybjOXJIMxxFOIYgOZEuhfomfNI/kxghNy5DW1KbYhVV45qamoF7
RomAlh5qZFV9awN1yjmxQXM3+asDCISCMLnulPm4l+h3LfgnDxq3ueaff+Qf5LqhA0tytjR4VfhO
57yx0IcfNY1xuWAys86QHv72jbO3uEcVxjjjnN+Cp2Z08Pr0gLhcoLG668/oShVSXvAvxbgwtOxM
1MzdFAnKP0/P9A6CHxSec5opG96gZ+obK9KEDvaczI0m8yhDczZ59mx1CKmzs9RyzvxFzi5zAWpB
37qwquT5c8+Cv4APalfZNka3FGoavZcnUjCKb6JiX8bIGlc9ZBC9cVCowV06YpKXB8O/+tEFZT70
19fjFMMaoJtaHUgTVtueY59GWQm/D71S6Hvm9yKDIrwLCNKF5K+1V5f6/Kn8pAbLrH3iLePb8HlG
w4n8YNIWWiVPmbYX78ftTCpzSPnXcL9kciAK2tEuAX4QWG2QRCxFYA6JeZvqHIar5izA0iHujr0r
w7xcMx++6Cntjx+asLX3UYA3gmrfOaMqPPO8uHaJlzmyHcq4awVoxje9ubojOtKx6lrIyeFLx5br
KKyScQULMNVJI2TctsPUKytPRShPouZrFw5wMSAUYOHEtlD/dNdRQ6X2AxFixc093g/XAbwf6ZD7
id9dtGYrrlx+RbGwTdsoqR77V//EBxTL+P7yqJzUorsJK8IF8f7JhB/2zLeBN9w0n95lLLCmRDFA
h+eIlfgyqayk3T4ZUu53xcvK8R2J48VvX+4Cg+11SXWIK90A3rRcT7ujUTkvGUGem00bZjpi5JcX
9AdlcMPcfmVzOv+BEhF6k7a8usyl7dgm55k0jbRzffp6/rLMmUPGHVUfRPbAPVc2kFXIFvNEHiKM
cIQ+uFKwXJxYG3R24q3/8Vm5RxQcIjdGutPvMyiSh5b7ppCXeLQS/A94o4eMlQqWh2tk9lOYpyOo
Z948INdmS2oWhShayg5at4i6QVK1oeccSo857ej1EjAdrArzsrKceDKhw9xXoFWIAgHptmKoDhP6
t6hgL4PpJGZ2T3dnGZ37dBk4Gk//QlBfGIz7ssePEhtCLWqB6YxLt1u5rpCLd6hA1m5GRpXDTq5g
HoCCBRDT6/YkxgRsxUawjwws703RDlmv9ra0JI4+aom0Sa8iunN+K3c3khPZNFWoPjls15HimzYU
3JmeKBki2DXXsfAXG1cbhjTTFSByWAa3NBIov/BVzt0LFo+X+JY8wNJrvGnFPJVShRzLYa5ZZTep
49cRYwFBbEK7JVaK2V/yTjfZMxLzdLQoEVLgyHnrGuVUuSx/pxfpXTw28hT34dmPZykXnJ/EJLxs
t48e1oRbSCCj7xtLBiOzg6YYDR2XDdvs6ZfDqdYozeW9m4BF6+j2BAr2SdK4SZplaeh4U7jBgmMX
GTLR7vt0Lv5tJuqxmP0mKBRdGVKDxj0pjzR52v/IIZX0MsxJ4ucE5fjufcwM73QO0z79zIGGqcCf
b+nmzxWngVBb4Ycb3VzuRLl8tqyu1/S1gHBbvtSTMNu+gKRVozBq/WTLmOIJcMmT+4Hs7vGJtxxn
2lIW7d8iGyO8dvFz1mZCnKw2NQsGv3XLEsiXyKimO162XKyhFcdveq1ljmtz3kdfYEWcJbnIMrOf
r8eo6JJlydCFLNwPrWQspsoWMcYzdQc0kGS+qBD8pU4GP2sIWXT3lFqL5R5ZqvI46bCtqDvzAAdJ
NX4fef+YK9CZ2dMjop47ec4I/onIwWrwZmLnlxXYs1FCCbXyUnO3rZEMrfVPSS33lSJuyc6cDl9P
LVLflGHyfm96WX+AS/gtPDjXqqO0PUXXmeOrYEE3SlOW3g27FBmrusvVFidZ+f2dbZiT3XZTBOAj
WnzgWiqfu7MxO4TnQd7yrtuKxGLgQ9a31K4F1kRaaWIpdmKrc6a4QsDBu+tc5IeAnY7yuxpCk46q
wD06CDM4hnqs4tzEGIQlRxRFJx8H7wdafMP26b4KeHyHvaxL7UUEPCzunJndnGDp0P08gcne+DcK
ZqwYOtHXo+QgDGEcaIWy0RtB1iWGrnzPBmchGIC89RWxbRGJ0xZ0PBjyVbPCm0Gj41obu1HRoSs4
Z0U2NU4a6eV/j0twu2sEOXVfPYzEktBGxjCr/FqHerIxUdzo1W/4CPLReZAmWIW66tBQ81B44vUG
u5fB15rZF4n9BWMhiu+WV7mlbIFnVpxJZ57Hqsr0qSYCuS1mbjZwFS/p/rcc1LxcEDMrAjh5pCEh
b06r+Iai3k7KJ95BXP1+R3V1RVA7VaGyduJwValQsHeBu7czTdseaZj2+Ayg25DxiIRm+E2FDu35
sKzL6rgN3Lx52iS4nWAiOcvfAebkNlWDkC9X5c5G9O7iIoyvLCnnfM45//ftyCefZ57U91wkxNkF
6q5pKdElnd7nPXbjERJpTRFt0qXwNwMETq4wJKlGXddbsZkZcFyxh9+JRI2LNbNaXbmyhdkXHM1U
dIAteKJXVzu7AxRiUQSQGtmqhNGMS+v6+sCMychrU/8uxF9EV2f0OL5hycRqOPQDzr5MjYtplirV
AVpLnkRGvfcYVR72w2+OWwMuD/l0DOJ0ijAwTV/pzvienHKPgqkPSZNRQck+YX+3D3G5fb6BuFAi
PBFYT37rkdFj/RgzaEwZBIatkrtlJJPr2iD56m+VUtr68eAWO4vpXHy1aeLE388pR7R0e13NayJb
izwX6gpokyZfJ6/hPFJ9BcJpKDIaGLo1JBXa+w+U1tJSv6S3tcMWfp3Ay4oASnWEohKucS++d/ES
7dSy8dFZPTld5Jh/RWEqn+AgqX9opEZTtFB/mmAWKrW45HDY2XyWGeS8diphoeCmPa5oiMAG0WMH
7T9Y2tFby/G9hmeIfkRV2CiV+7qJVLAXGIyKFxp8U3fCnl9g077uJDiUUsLrVKu8TjjI7J37e5dt
ed5xPGqhc5IpjDCxNJ/2qfE0cFzZ4lrcYppicWbvexNbA+6jodq/xowh9maX+vqromfdWuBVf2uQ
eYKDFOdcyWlN4+8HbqN3W6zl/oxfTRy95Zx4XwJkg0w6gu8XW7S/80M7Zq8i2PxMI0il3SG/mgBJ
AbHs0mS0aciH3cMWHA2yq+rDnXwrqhOVTBwfpeaZtsnM2IIobVOWxrPErTQJWJHxO6JAg33mP4di
14jJ6jswuktmagYAZQCNHl9rAsYFkC5DqlyS2fAk3yT3JaD9yDLZUlCj+BdCpujXlspESwKxZykt
dB/hkXEyXpL8nmH/Stkyw/8yMFREAo2p0hBCLwp35RkgbvxMrMxxUH8ziLmZ8nPdgn1iqb9DEb1U
XxRnP9vY4nVPLXo/aLkNrDhcCNL4iXcPxGB3X54SWADm2chEYo3lQJbJ/Yw/hZ79zz2VBKKBLPUa
vya4FEQMXpA1WbZoG2b65iIoIpIz2WTToPjvXxBNhXc98XG5R1fYmQGyPr/7uvoFxWRvrDr7WBbv
NDUkgCqfkWurKlhBd/6dXn1UF2R66vrwLZoHAXRppoeqa9LV+v6RhvcYtFNetljTIraQRsYl2NAt
DKanCvYXPKVqmCMdjxx83chGG/DX85kKJapkCiSI6ZUBJqgqsMYKI8/u9phKnYfuFn5Me3ZwSxWh
ecxvVrXG8HMntEWq3JVWrpkDg7RMZu3qcmh0xWfMBxAf5V0hGk4FzjHnTAplXq9bIzUq3P7DgZxQ
Ek0Tw/infnM5ZZEK9jYUghqEX87ELT4uC1krr3q+u2GBqrZ0u5bbdumgfgxMLSqgkxFTUDLlXZ1r
TkivXwdWRzb73+WuVRmokVrXhMJEkEZokHnN7m+qAnEySV0OWzcMfp2Bogj3REjQZJYmn1CKDN6s
psEihHyfxTt0EiTIc1f5tcYeiFv3x2X3uCZD4b5TuanV7UjaTrt9aRf9UMCI9iMm9NMrCmKPCK+b
SlnsRsqrP9M/qHMCvPqCco2g49q/VOyeB2esLxkR+8Bt+GNBD1w+jGY1iZR1AmYh1SN/HscsT8Vp
UqxhjzUwaoYazQyqbP38UC1FABZslhcHmJmxMQOUw9AIVzX+w6CjksEhwwUHLpTywuIyEbP5e4pR
Hncz1StMrOSqQrMOc/6D93mLCdD2XNwGbix2nFdF8SSrR3JXLH8X+x3IG9GunPlM9w6RWQdl1ogS
WZ83cA5f9LuRGJzC5e3ZvwqIRr0DkcZox/nydWuLdbMxjk4AHLJqfrjnvKJ0bQmB+TKNYlydayMI
muQkK9CIW1fAcuxI8vsjCoi8WssXeLpGx6lVfBTf+novr4Vu1r2KIJaP3fUIRGXJlWgL+E59SOiW
qvZiJhANVpDGAGXtPkTt6nOUPK/L89m2A3u7Js574/k/XqsXGdF6mi/bgg5Ho0y3maLd5mnzQz6a
kA9E0uJsoIdfxp6GH+W0fJT68dCB+YPExl+OiojIHuH9LIsxOK13M1QjMDMkRrjq4JhTOHvmQDVo
ECNbUBPvwzPnvvSvH/vFBn+u7ssXQtK8fkOa/2neB+t/3/vPzTP7anXC2FY+RI/py4O9cKp9ExNm
o4Nc8Z2eSMe1W/8IzpKPNatIRUTAZv/RyjjS/L6c7bPCBAcISiIuWqRua9NsZvmbin4DF4ilR3pE
KVm3t6IHIrzy1XDEXiYpyJ0Pxhy11sjZM6M5g4ZMhdApXfTOB5UfOn8lNRuWnTZlkfH+IxOBELgn
kdAPbuQAN5/a2zAwFEx6yEO9/NGfHW/CsSRZLTGfO1A8e8VStim8mUg3oD4uyl6Kxj2fLoa/Z8SY
kiWoURIWGREFQ3J/fB6HVviN8490gZ332aTEQ3wkx+ID/W++JLBQ+yrklRQ6EJJc2uwx+K519khU
k51I0+rEYFDeAHEyPwqQmr/T48zfgKU3npVYOqhXOISVBfVmvQSgEvkchZlfaxGmA1b4kBVD2YtX
PF2Ht6eUcK7//85b5v424joTF5USUoWZFarFXJ9A7izTHKpfxz+hzifFqCfi3m7iQ+PgzcvF06mi
RkYB1DILTrRdYSgtuOE0wtylnpAe34/FN5pYJlM+FwVbSb6AEcoK54YBV92fdR1pW/WbPycK5CgV
xdSP1r0nmuBmUXdKd172t8No3PgvQY+dnkXqCOwlXaJpU4fZ+zuG/hqSFh0eX4Z7qBQWmsGefin3
64f1GLJobYIjCHMGl28Srwiyz7C0BqIk6j3Q+1XbhPFdndCa4ntMkpZzyccQ2RQl/dP3oTLvwvyC
f3Tb9t/yYA0N7NwjcPbSBsE9ViAPxkSYyZbbFNgVw3njP+JiSJpBmA2gV4SnfwTNdKueYRRbJHko
U/xsNTFY7ZV7G/FtWUvr+oC37+QPEgl3g9Osb/9/MnAT1Ef6wEYj4nVuuK5lMkAVcfKK/3lPvGIf
hfYl/rJmOIKsHht+ZMecMii1QiEVvFbqWXgJAcm3EqCYDH6UpHE5q8JLwj4xFwAz7NxS3+deD1V/
LI0dF3ABXWk4fQojK94PNPBlVGb3g6p+D3OWEArdhvdnGfFtJ6LYv74z9RvFcyZ9UaTPtooKu+O0
7ueq/fWgXhKc518gjtsUU2cTz6O+sNjTMzqKWttG5bLQhPfSN9udmZTfmsPWZean/4SGsStx8C36
I1gns6BTdoiw/6cjsiqnt9UhLzWHjdquwy/B/T3y8rccn+KR0ZK4X7MfKIi5Q7o5X18poGhvsOjQ
TCih4tkDEdKlc5e9lpgeEXoJNmFOXc3+BaHE1Cbgf1iTHCBeaZd9AoACHdgWT06Lwi5iYBqvarBL
bxkMzv8rbrN5f1jZJydcu2PMrdtRrZoumG+DBkUdtTX7omYu2fSSHfQb7YyRbuCFrOoAZ/vVS+cw
JQrPivziaTTpJrChIKLMfXtFJcRsfPVKMmvUmZEJRaMqBEukUm5EwpNgK+w6OspHfjzzwwBl7Tq2
VZvod40J3db8IIC4VK/KNEe2OvzPoFU17HfvvgK55DZSr6DBFDsvdqs7vwb2fjDfiuEiAlboab/x
7MNcLksutdJ802ng9MHISLSsOEstuk3tkJUm1tuWgzjxEkAqIZobbPu/kOWjJ0HgulRIBS2feOO7
MmHH2GKsyk9M7eZ5zByqOcOTdoHGSMlEWliQaWId+qufV8rd6sJE6vqDmStMTqc84Q6GkvBtvJxO
n5nGwVbmM5teB9vvJLmINRGT9fNAjBkrUGeGbhJFxVf4UcBQg68eJK1wW8zuarYkC7TbVtDpnYet
O/zp3on039wp0nAHdGHo6CCqDfNUVdjlPizxikMPt9eN4scFNOlTLAvSRAHu/LPULJhV/KWIkpWZ
Y1LXuZZ4bW0LAb7/4sG0jXFDJH7zjtl7oD9ElR+av78TYNrr0BLJ9d4WUUi0A6cGcukiQWCUwSrQ
a1MPRGQgjYmlpNWX+pX1wqbzvpzVvaKeV3ChBGb+VtjChLCqcBAkANfbrJYlO7KDerOyp3YY979a
B4wBoHdw3CeQcyNwqdOEj8JtAWQvR+l7TzngClsJy3mijaBc2j/yuZL9Vxehsr0LkzKvfLgkjbl2
yYdqcI8v/Nkfyfhujys804B8dZELpN8audhLRux+dBT9coAL9v1Fivl63XDbhIKGxs5Ul1UekXQn
zxUyv0i17zP5gOD1uooC/ZUAnF8EHHa2P6jpWvDwHkxiIX6SDOWAp5IaVQk2aGySVBMz/1WCHRSg
rQvhSAxIdM4SIIIqaPri+kX+SujvYCQNBugKwdzXIT+W5i4nSP4p3wI3W0P/d/CjzXVyMommTohD
kULZbVL5WxObtCmtTukaXYDfB1iiAjByM7bbFMVyU0N95+WSvPPaq6WIiOUHF87Kju8rtub+5FH1
I20OgMvlsvlyEfaPzg1AkqPISBTaIbsa8UeXvaPeZJFCp5ZlkkBcxYEdQJHdn0Z7NoZqoczafKmj
TbSq75jd1QzlvzDT8ukwuQSU3PHUeky9j6tROEyCVQuaf7vgE35oc8l7mhGf7PWEXu5TLecaBKYH
z0FPneL5klPeQkWh7lMpo02fsv46vjIGIr1hP3qFtR3Tk8mb2hDVbm7WvEcbpF3Ym15druhDk3uQ
OFP1NLmhfz51Ggt+lIaLsvDwKcU5rEm7FeZC4gN0HdmIbBHNIL83J3HWZIS5E9T1YMCeS13y8NCf
2eS8kjt8OU9ak7lzs2XATaG9Zxf40LgjZmQRqvJi7h6ySyueV80Kyv48uknDcBdInz3tc/S7kr7G
zfC/JJ34FdeSXPjJkFILNHnJBGef+7tXHzZ3wSDSzGzJRx7EZMAEqcamKXbVjHHjdDj8/5WzZlc6
6XakdxpGyaBjQWoKQ5K4ZG+3W6Z2aOv377ns6eElIpYBnr7C1pVcI4Wfq/3G3u1HoYdPfICO+wwq
+grOUbmL9mdFXWMUZ93QgP6wl6r0GvNcCrSjfKXt6WsE4ifAdt/X/3/Kp4Lp1GUF6GdTqfh78Jw3
VmC0xLjqEb93LrlyHheQ2x7HZ5HopQMP/WCIE501HX2onc/swbXqKabEwagzoUrINzJxfzzkJP0p
vvKWbii5iPqIiyl4KJPiqZizI8Johr9gpMRpYkDB5frXix60D0fLEQ2HKKrgjzt1UZ42oAQNPc2X
bmJwv1Irc/YjGw4JtfmgD+IMGbwkKD/C2cKYmftbwNEMXH4+WqaIglvd1vspjO9SdqTLOGbD7C3C
c7Xd6RR90aDbuEiQGH4FhKLIgq7S7+5hj0e7y3mJjTidOxVUbGpUBCA3W8ziBkluivhHU4mM8N1L
0MrNPU8LMxIBqhXKnQULY0OgntIRpGC6rrEEB5AV7n6RRY+828Naz2TGXlMgNkodt/vTyrZk8aw9
rek3fAQDI+kcTjBFZilCVWGOwbrINv28OrRpD3b46775J00cftUJEIsNkd2RHyvnISIAs//clUN3
KcTS65mIGeyAFT33a5/5tIN3g0gTrl+otPPTSbCImnytQifNmCdsMGKKZlI5SOWcXMbNlwXgWqxh
vSyE7nXgOeVtmL7cR2p8jY6RIbMVO1E0GNEf8uPIkZtyxb3Kl6ntydSR/kksyP3sga5Vc+q1K3GW
hkdv6WLgTf3vl8E3+bqajtwa3Zb/UesaF55Vn9/jF8BPsDSbOBL30801IAMCT8KE2JpSyFXXYLrF
eT4GnrlhFtlEuTf6JUvIZUaq85KmzbSxwi0whlF6vc55IcPOic/AOKGthvnimKL889U6cc7JNQ60
mA9Gr7PT0A9bUYdAAXqiy75xWHjHIY0Z8MV5vyUaVeVHaA6G1JEpVWG0HqxyqWhlAL8VItuYFzjR
sv+0Gy2akhQAXYMHtRfyMffwP25aDw0T751JaL7aRAR4i/45Et67JVIyw6sxbOZPPGozJv7q9GxX
uxJmcblpEIKtvDTunvWPu+CnpyLmQcXvycK66msSJfmpMPcdS77cu6jwNnjfzIOsmqdsUVssY+x/
CT1+frIc9q06PTAd21urQmrERjvbfTkzsY81SptdAwa9TJi8lTcXt5Toy97Jfj46hEmuArKOStHp
c4Lugpxz+bPpxukqp/jz4Z+701d/Krw1nwY9Bdy4IDrcKWv+HEimpEQQnw3wfy2Ii8mlbxNMXhNi
ufVJYu4AHQzkyABg/7q9iEgFN8my/Y0BChLSW3MGGAIYD/7ods2eL5oEGwvKxNJiPxcF3MkasnX2
Ai2IVHxfXemtLeWkDXwZzQmhKorVj+0NZ4meH6+ZTwAIPv66bpXuiIWiIs4NIhHTJNCqfGuRwTMI
nl/VPkYyImZ+U+1Pk7SbllBNp/JFPHld4ZSEtYZARlMa3M6nel4h5IRv93wym7NV7VJSjNmW1zIT
p8QwK4wAH1k3elwaVN2X0S1YtKlXnJpYqVuD/VjfMbEcj8jDkKCZ0msQv8wBNOGi/xJUwtv0j3EZ
DTa0yEWF+0LRqwaXkoPLXZZOTBgLbD1oVF3GBVssWVJiP9/XTJMAqWQ8psFmTUcrZanOvOUqJX5B
Sl9ajKqRWI1rt8vi3rIl0NOrzfBkxXaCTOi1dDykOQuAzQakWKXnqy0cUuQ9NosqNpVpA35QkqH9
1zDWU1fV2GuGAB2sbrFE+XDQEXWeCavTjackaraRErGkKDU9pS2HjMUSQipTvqff+VTnvIuPcF9b
22VjoO1WTUcUoLNPRpWHAvAdA0qJmcLhQSdWebnclAA7X8orcziXJ/WY3e4kmhrxgaRRRzSmZl8I
QJ4FPpvkSXbZoaAWLwMK5bqXuGbmOacU2Fwy9K54h4LVeOvS0G2dbf+ZnekiBVAwcJsn31dakcsC
+IxlwghZa6VY4Sr3YybNUdGU8t7jDsAvZwNa65imVRdi5oOziw+kGrA3bfAW9JwqZzUZv6bwk/TH
pRer73mAVhkJMTsyEj1VuZy5lwctGwwLkoOJa3naX8Blz5B5zlzr5Bfnmfe6HgxBJKzTPqcnA8pX
qr0bKAef15AVZAKMbUCdCNZ8QK3dITOm/R4ey7oTBpaYKiPN44fxl45SIPpiKjc70l225rqGta5R
PhK+H28235D6TrNNBkQrlnQ86TvSz1ijzBzwinB/xlCaKBJ6Iqqc3JvRzEJgnP7FZGIbhoBVEyb/
e0vCOtRu7j84dZqHzX/PcWCpmRX4s5aQ7GO8jSWvmIi1gnWjYBY6Vs/2U5HrianZsfhbgmjDXCUP
VbtOH/I2ZjUSvVCvpmJbSgHQC2AVKF7ETuhVe4vGmD6OsIhNuhYXeeUx1MTCzqPm8KmJ1vZkeSuu
LrTFiQDjKPzGukl/2ekS0emaAfnY97Uq7xC3IZGSr9rAPnhzxJjuCuzPIXQu5o1zg8KUhBz2w9Zv
zVpOovzdbGbkH/1/ImJwF4RqHZeO5zBqdf/b+1dPoJ3Rq81Q7nD/aXjMx99FQRbHSh3A9M8peJUr
0qNFH+cX6ojVRq66I7h+6du1Ti78rfVJB96wjdpGlBsXsg+eFKf3x232xW0sTXenXCrIYU0cCx6Z
k3sZLvm9WnpnHvgF/zi2zrjv1DzjI8AnqgOiY8SdVwgQH5Iydg+vk6wGO5DvHw4l7fSqOsOIxhWI
HDU1v855WVJ3vlo6SPn+qAkpNW98mCeO3K3H0TTefO7z0LNmRIj6EQztI4TqrRkKoz+USChMiwwl
Y7htLqg5mCr5aAhRoZZu8WqHbHJJz5r2ZyTeQRGORxDBmC5rg7XXpMEz5xMTzdgH58+PLxY1QzK3
qec1iUKZwHBPJuKa+OIUEbsXzW4j5Nd+kuEsoYwlrAURS0wzVK0jGnRIeqluVtPOh3sYmdfcX+9N
m0cETpscFURxRx5ewRJEYcFN63IBxGSSMUNekBxQzE80n4pVOMH6g3Gj4T/CO50BOGkF7KW2tAkK
COt5CRZobtBRJC1OI5k5G9uzv80hsEJIU+t+010N7FBNiW7bVpefCjE1uMFA9NO5MIGIlH1d3SKg
XDWjTkXeb4Y6gGxgU5ysQEoEgGuN+Ezf3zzaujqRespfweRvDz43/62f+rrI3qIEm3wT2hxlpm1l
M3ZjfSCpVgVO80tSJDy3F5eLmXXfu0hcjIq9D/4XZudDlKi1LU09PSl03/qk6yyeVXpQHbuFBEaI
4bLINTKTZqrZmf607zwSNIkr2K1atbZdSIljNChPBSzmsG+1dqldwVU1dbeNtRUJ/YsR3fXMF9BC
yyxeovugDTtaRaD9/+f8xfUUZ4UE8HFGWf8q3rgvW9xkB7eFLNecxlxChdXyJed9S58QYJHeQOtu
ka30xaJU3sKiQV52Ta+HhaotW0V2MfzykA9HtD7NCZYGxcV/VNHlG5VC4siurcp3X0xEfdBMYbgZ
cZCkco9MBwG9vyGSKw2EsEx/hA+HiXrseqVdyUjiIoqvoNuEJumyRkhXm1QVyGEWONJMxwPdNDKK
91ctJpnQ3S0dltwnKoDtSRPn2t/Ysx16eTAZcFhpGNE7Wqbk5v/A7KIyE20S6AxobLPxmZEEhfjZ
hpa4pF4Y5AEihuXaJuh1Tg8ye1sSqC0T+Z75LG1vZV3/9URCXa4WjwGOGpqL2nribBL1Tk3Csn7w
YPlXNEvBa5lFv1bB3gmUezBr2kf+c8xQHr0F2qqMrqD80ViCdtcdDf67v498nZfdgSyHQ+zCcCVZ
9IC2uFuIMCFhIr5NiCc9++VkN+mBo/S8QzbqEbsdub4JZQ4AuTSDhyLxVw/MTQKEVT90fj9V5BBC
ha6QwmkZGWlbHLIEx8f2S4M8mudGNcknKhju6nW/iSZZxlQx9owVNPlgeI6rMVEWVPkCG5OrXU9j
27y9jB8InazfczMj2hhmZ/qtzyVUlrdwh8MPzVZ7ezItr7tNyp9JbZ6PJplpbI2w3gJ1m8rqZuM3
hCHoD1DbW0bgsiVrQ/YFvxMqmmBqu78aE/Gjru0jqY5gXb0cnuHDhcIpUSRODbLc8+LVW462zaAq
0vnrH3HLcjNJ475ONd1VvjQp475qJZnJgtpkRl37IbMaQsEfw8vAwUV7Rgdr/aRqJG9HkHCkEP85
jpKkt15P430hW5sfUxuuHNOoDXWUF7hJCBB96Y96zxD7g1c2JoQS7Hwdrw13Tpdmg+JOUygXUdmn
y3yut6oW7lkbP3i5I2HSqHTFvNWcGH3pXzneSFAgs2+JUSrnN7Qm1LxEczA2+tc8pE7l7gJI/1uL
XCfM/5WdxLORQrtnCHqcytk1/8D3FCfThYmrfUYsU+59T9BcjosRn9bnFxG4UXC2onXTWXSuLhl/
v2uE7mJDX/j47h2kINynnwjQNiJehNtLl/pH/Ff3dQPumCMcTrIpddXEWRI8w/a3WiewzoWT8W32
vVrQEbKMHcX8tXPiHtGTAyznRBRO2MAcbx+wkX77r1F2CBniN7GORMjomhp+mJMmsvwZBqSXv3iE
BZZS71FxzOxgXFYE2iC7J08n0BHz3YS4ztRmpTO5esyHbQl90xaFir4St6SEnHvuzDMfQVlc1EVW
QgGWpSVHHlqscphb6LuDFqLmFRge5Dlgg2IJnCWHdCL4ta1PPUwJlD86B3LhdJBFdQ7mcHy5LORh
EXCoh8HEC0JIm/5bVgV1aGrjbKIhfStV7WgeVBlCoFuo7l+e2i7QKunJCbupL55Z3ZCXlWFr47p/
WdKgONHPe2sd5Saw8hskxT3yf3oqXhqYI2wXv4+P7SMc2xKR8CuWITkYy0O4VN4QheAv1SRHjwJr
laeFXWO5o27nU/AinNFvv08GN2LabU9oOBwiPGXvs2bpxuXs4q/WLwqq7Hv8G9Ddxx1tsuSI5oB3
XHptj0uKRSwEPYNnR8CWbhUUhJiRdprL9pfPBMn7aCV9WJQVVd/mBRXsBN1ZPjbak9aWZbxY2tjn
UCoUJ57c/vkS8syNj9hCO2blm7XgXYs96H5kbHmAqZO2noUvEcVhmVgTPEtCtNR/Jzav7jinOxfg
bLLaoRJdOoZB6TEwBJzyMboYTvUk6+2llOfLQ0KTBr9CANvPkpQ8XJgSTkptLxJcSPwaaSNIsl9b
R6NpNHT4LoAnsEgSLyxdixTSpaAiZ7WMpNhPxt3JzLmpPilu8roM7SBh2WK6o5uWsq6iK7m2ZAhk
96J+NC1AFYhbZ3xuaetN5HrJYlLa7RokG5n5qKspbpldemu3kx0Z3TMAVy57USy4WbBRmQZHaQLg
abhnzPVkTAfOW+hZILtJRzdEbzLCNUtJBTqjF3tXvHX3J/yt462qSrA0PT5E4pyQWXLsBDpEGq08
a9wlSDSZw6ziQ9iWBuIImjGOTB6wK2Nw7+Rvjuod4SyV9DQnA+iLZbBv0CrIaiNSDvkZUlH2OdWc
53jFvdekuPdMbFECLfh0S9QIFFgiaGpxOetugSH754c12aPcQL4fzP+L1AwhSUpkNAShoutDkqNh
4ljSyMCxrjk3VgeeDoDPqCcj6GnawJ/nvR7byf8Jo/1ceZxrYyJJcVqYF63VOTLK+QknJJHZhUr9
mAGBDgt8O6JPnJCDsXSArQCz9besKwVs3Lp7tEwqDuP/UCFoD6kNNqQW+Tt1Nan+CAhyMIDvPSKR
/FkMMSM95N4J9JNG6t/VvP5RKLHjJKMp3ckRvD49hMgJNILqprPFq+O80XcSSuAfsM1KrPYzdBtB
WRxlIBEgMF94rOrCFQeJ6LbFS22cOCIxOHQ4YBGdUmVSDT1bUQ0ZM8/ll/ioqxnRTEoeAATT2u3X
wVMSKBPoWqskHlZfcM0XoOrK91Ds646VXJWY3McpJiQlBp6+ry5XQVAaYQH4iK+/um09IsVEIX1u
itK5n/hreYGKfU0XXbhLS2r1WHb2f6oaKsUv/Arr3nLQOhvEI2y1jZmNCyLuSJ5hZ9KriA6BYZsC
qq1gg1C6hDIsbEE0FaFWGm99MmxBfIPgFO8elwO7kLVBmPfRXaC9cvP2YQOJUnyhYJVt4bMpojyG
R4mZYHgXkBNJlm3FMIvoPiR6zSglciPUpMRP0yWJGuCuijRc7iaVtBs8v9/dbEofjyq3pxX0g2Ua
zRihmJb9z9XM1qypkfJP40LQBXZLRM/cSu/+Ewnkcy4W+jSQycC2jVsS1NLI0fy1pRz/3bkeeVOC
3ZxktKXYdlmvkX+xN304Cjsffyesjuc0hCza6Eoaqp/qsyfxrujgIHVFEm0ppwn/BX2w3HTY8CYN
DIGeD0KtLyS+CTXtxiuC/pE33ix9XJCWE6iKdwo+ETonO8yZIs1tUznP4Gh2Y17sv/TzMT3Ej3sT
24OEZyttaTpNheeyitiV9LzqtW83lMRO+g6LACznW3DtmRa38u9jgFVKzYf4xiEQ7Zo388VJ5AQo
a3GeyFfA4K1zCJndMRqIBQQTkF6vNflvh9ille+eccXD606nN8HbEtPpuwVnDZFYnuloLJBKShIx
G5Kq6c2OcabEq45Pdb76QrDiYUhGl0xxCmrbOFwCCXpO04+5C9wQxERHAeg8PQ+Rus9/SEcOa8IL
JeVHvfCy42IIyi2DK6ZgKMjTNc45C6JkGmL1d3XBr9I8HWzeb9+uhWMtMv6AieaXXEDy7v8zOW6q
27dETQ4C2fJuAAQXqJTPcZW8wZK/wLbcO52qN+DE2hKb+ZEGv5ht9AZGerLeaMkvnWzqquJE+BSg
8VzmugRovIma0l7N5bhLYWOKK0ZJscnkM0/YMROcAlpbOQYfPqj0tww2Omqdv/0ytTWGyNo+UZn0
hCbqAjzJr8Y5SzPj/5ffLfhsW3Vm4vxMLME0Zs8LqGIntOycvR25FEgdbpe21eK85/uLOf0FasTE
YKa1X57PY73q6IqG03Lb6btewg/AteZ/LDAFtajcfpuKO05wFxnjBShSYb5xewOX0e4yvyb/KJof
5uZO0DtQenHv02xl1g26WJvgRxSff3Rc48vYYwvsAg1+JhpIQlRV/Uu0PLh7nqJ15tPQU01Lx/0V
+pm0hTkMNdg3GAhxT93ZN7s3QZYS6u8AUjeUQIuUkjZWQg8V9ICOBoBiP2igNnH1TCAawludTbPt
MPKOUg4DOoeLqE9oqMPaEg1wUTx3uHx1ivknSJ/0HxYECO4dzY0PI0KXPWy8fuVAeIPhi72nkJHE
K2oQ4FVgStIcAlWfTHTBSV5yT/2l4jiwjKtB3kIhtm9nTLwc7f1S1Gahhhj2JWnolkolAO1MCDz3
+g3LS6GQ6p+y34O0QvL9PIAit65W/flTGNeEF0OCu5rdhtlRcdBd2CyHtSOGqtq3jfn4DyMy4U2D
zenvAVIFkEBDuoGSYgaZk8VoQTrif4LWuc2CehkJTDw3XiG7aw1g9a8NnJbt3k5nsLIhqdeuZy+J
5bGzg3q3E1fa8VweWmEnSruWrTHHSXPKyP8gs+EDl+fmyyMn5XXSRR6+Co9buXBRP+YXxjpH0JfA
+tx6yCyxvq6GyL9yXoFU/Y93N4sAae7LzeDvPbH/XPPfr/7LMoNfAI1AOLYHX6ZCI9wXHL3DfbYQ
GOFo2Bfg1+k+toC0ZB0UvP6t6meilcPI2hIGZEGqRz+4sPIymLCm6zjm8/4dXLt48D24cjBozzAp
Jl0R3HjbWp8MwE11JPz8h6+H5d4mB09MtntaJnnGSRF0suk8P+kL0Ypq8fdPLMgNk8X4IRgwGMmS
YRNsLSLZo7quRLVzqiDNU3oeZyIipyxcQ/ZmUG2Fl96V1EFUSMBY5bs+MS6PiKqLlUXudaKzws6l
WxQELhWjH2lYc5ysB5xKFVD5eF0hHmP6nVRMD3nB65sf/KDvWjeDBY1nLL3MxaXZfHPCcACUhNDQ
GcT/emb8yv2UNe/lktciGWnvuCs8x9W/wQjxyA9B4Y9+CTW8rESl49xqv8OOeiuxcEK5CtTkhQ+e
2bO+va7/hdGJVe2bOq3lX71xxQ/ZpkhDbSf4qRbRz0hPqm0FYma7MxQhtRQu+aNH53ZtyCHTFGmE
IVt5XMauKwkHzN3ZB0pMMUByM5iFdTA230kxC4V6v9cQ87DKzDp/2ovwE6DiiGsCfnK/jna5GGro
nROwBl87my0sVDeUTj6R3h4CTiNCdZrHGIDcE4TwD1D3kuuTOjWDlDG1U7mBcO6mc8hFnvEJgkOY
4HMGdfxURs3nFTIf+M3i8wkVN0zIpSj/uWheIPekrPqDho3EnFVfyWPA3QSCM/g25j3fM3RYC3NB
yT6aQ858tygWGuGN/tecyH4wH0z7OnepMnT3XgnasS9ZOnuZyBtR9ju912OH3/dXGJDOVwl05wQK
tHhfEt5mPhK6V0uU1jWlVZLUZwuYa1WOBgUZdFCZbtgEFx/ev7qGDSav0rwwlsEg5XK+8P19nM8n
mS04ttMnPV1oCdSPHn5toNr5Xyj/ythIFgbiAClVd07OhSn69FwwHYTp3ITVdLItAM1jUF/tZSLs
WdX6Jd0NtTBo/D3ZJKKdKTM9eJO4UC2/XVq3AGkeOoUMeh1M4gNw1krvC19YKJl42cMx+lhcsOQI
9FGDg76YnE4FR7eYAmMtBg2gjHyplOzfcX97372KzybMNTPyMYljRzLom/Ks9UVul/s8Mp2CjEyg
JqW+wh0JpmQ14fFdFbw3rHIAdWQ+dGnlPLrdO9uPH9JUk0yu9WgDTRbRMV8zq3nApjmW9eqLY1tC
WYqmn8ckpAkZBgJsco7ClqsvTc2m2UlpSzXPiVMNOAxE3vAm8Ne6Kip/UD5kKoiwWu1G+rRdsIw7
wt8RhdQ48C5Eqa/FDrh0B/k/P3vIxSISqBLB/+waOQRyeB+cPG08XQzgFoUixdsO0vHNSxBqD0By
2BXZrFOdk3H4kwnDnLsEABCMcU7+0CMOpgmmQIjcjIXGOmogsatVSAAuwY+yI57i45MWNU2KhhyY
duRhMTrhNYvG1i9npY31G2YYS+B3u2ZGNaYeZwCwAK/DgmNMtgBNwSn0+xPDZJlvTyhsl5bTfDL0
ER7MZA4QNsEYIPf6YqfLoa16a6r8Wu4JoCGTgLlXrMqkx4gBWoKURej8oR7O+Jarmhf/agXqJta7
frQJjgLClgrlkd99RMj4JQWBHnd3HjBctVDsXQHzqEVpv0rkyEOI8x/YrYrLQYdxuxFRmvVkyhzI
ucMXBuJX1rALmsa6JJDqgCQ2nFDb4EFY2Fzu9h2S3YhWJGs9I2X3iNGz1MnEPsjrexhR/Y4tNdFL
gq0ytxO+oWV4G1CtTCKN4YPRdOqRW57xMQTy8s2vL+gL7lJ1WNHtYWmy2FgQjeokAK4hIvT0qjxH
MKEEZEq7zqtXLJBJ3rN+/mQB+cdPutnA5cdx+rG472V0GO5kcc1jiGcKjQozQJQ8sYwXVGnQg1fr
MuNgrD53ckPyN6U/ATlp8yrq/cyMz3/1MOCS93pIyBgbKTV67i72dGWAtSkONXqLY1FXDMyKRMlQ
tSY8E73K071grWtVR2jbp/J5OMc0+wgNjEIWnUGbn223uTkJJbtOiQt54hzG7p0UDMikV5J+sWzh
4tgXJIEV2QyaTjzUxtfklU+dAhC3IiW66gwwM9y96ZhHRIA4SckT6qpomj0EI9IaePqMUAJypiFp
uxwdtcrjJnQMkVu3b5BEINSaTWtg8oFpEghhnEC0c6A4I8nuAA6rpWQA3X7p0Z8IrWsE9GMsl+p/
ByvA+UAn7u6OEGavCep9SnbHZey8KKXwOO3sPYk+3Yi+Z0zpMNCTuk3rBcAE1K9y21F7mpnEeAVO
/7+W3CUvdRg4dNEZqaHBvHLfFm3dG2iiPy0Bj7Pe43QtlzpY94gYqgcXjTfqGfcDh7qU4TQ4bXu8
fwDuBM89Gnlwf9Uwd4xYqXFn47VicLsbj5+CD6WRBh+0nRhVaRrvf1FOGZSF6qdLXXJEpGhlELKx
zDWqkNvt/lrCgcGqAap/sHPHQH7nzwWxNC5tdGTrGZYCIaCzJYIVtaZGi2zjVK8c4HQRbWgL1H9J
06FVtVurQ9FdOdqBbJc0XIX0e2mK+111I//AkbmG6VT6tPCv+JFLpXSmDkyUQqfPuUXbutlCL2IJ
6a+ISMnxxT8v0Kk36nTnd2o9bVUmkITP+bmp4ItUbRXVlIFCK0IRAC91HSfYP+EAogaH+i0/aYz1
B67FareSPMW/+rjEtwnscqRMyCRIG8Nr1KUlY2H8YM5pPKnfORD0uDNgD7tsKNRvVXiFZOwUEcZ5
h81a+NzmOcqnxOhFw1ZuZiEEPqupiACvNiWify1AEqkZJ6psrBgf/HSBtRdMT/Ok6llE19WPOKxN
pFM2JBl8XHTbVaDaDEK+qFmqvzoUZoFx6ZZro/3M8zpe36uYA3+PF1LtEU6hUQn32qXe1STXBvLD
2ikDRPtkG83MgJ/mojHpra3fLUBNmZY7SUGIv4RJ+rp47JMDd2W7mhj4tmw15+NoAMtzjg/E2Zcp
t7bFauwXkNUlbnuTWXz1dbLiRV8yND1MadZjNb83NaBefmPU57TZh5CsGQ+euQjokHmxwH42B1hv
qj0hYm6k74onVzL2WZZsFvAoPX5Nx8b2LvKhbV99jrdbGJ5rJOFYBjLcltUxtnZvw/CBhrHZDMfh
3BOJg/YQKX/cOhKCdHKSOIWPfKcikYWEne02gCxeiDXs8IvBZjsD7tGhKl+KKyWjLhqkTru5JBxH
MX0mImRqmKfRrHUEhgPETmN1UOLBZvVA+trpsDJHRfCJvsc9sJ6vv79hhOID4qNt7h2/baEHPj+m
PURxZJtoRLnpwUO/NptG5fmZsqo5MstCoLzh+o0HLal7rn7AQCQX0/6P1wRtsDT6o0Fj6S9ZOBbC
z9mzw53d5FS98NeGP2sT6IwjM3EBUxR1vH238waqNih7xsHEdUnoZWYrmZ7/MITtM3N5I8N+4NSY
R5mY/3OtYNQTbhNQ9scL0SXw6uyN/RGEYUqMBXeCx9LEhsz07EaRFxhu3zKyLVY5fi4vSCOx0gYB
rmRyOV0eyhQPljJTIgtg1kTKRGVKA2gZ83cjOq8EHYvS6H/cYc5z/QcUMeWSdRrl4b2454hEjbi8
/A7Znr5HH3yhDIiVoEdHU0RXfBR2AgM8JJ9l4uNMfNDGJYl/y4EhzFsJpmIXu/+Ah3QDMu5jpAbS
wv5elDgvgZhvym9ISkyrxqwUe3EC20FSYlWQLaEYGsYJjINjW0n/X4gEPasZOZt4k4H/vB6lmgww
9zT2S+a+Pb3QTeYlowihyez979j2l6X/+d0gLH3vpinDuJDlTCxV+jdbln8vZLytTR2/590H1c2z
Ve3+IvTH+gsKow9DUJRvlm2faxNvGfMhL3eo9YJuqfVZUUUw58pQDFcvS0t3kA0SBh0/WGniGPdv
4HjI5UPNesr4bNPGGKNd8j/SnZ9ZGeuLJY3Z/HHgisHGwCRpvJf6yYx1IDZWPU64L6PTFulwWEAT
VMhYFBnXZuMmn2ihKgumEFtlvIuSrlgZhb3Grdpijzppz6z0IfwNznclbdW3OrpMhLm7lVhqNBaw
k6O1pODkr90cRFY82NsPJD6UjgGd8AEeh325F99zCcZRP/CfKLrS66diNWC6pszwkkOzQJ9ZQ7iC
u7ybsX0D5E4/q0UDk5HluLLxjEr+qzETu5D9sIrFpXAHSJZ9QPlhLpg6IyxVTJv0xKKM8GkputyN
L31bgkTT4MF6D3vWRTMDnE+DsJKfjRQuh25BAhkFtRdBr0vqVPd43jCh9tFzhJanAKrvr87ikC8D
cvLgnl1XxLOuQG4jYCfvfp9NZE71I5GG4Xu+bf8Zma7nfzRqRSd/e4tgJWU03nrYp8nVK9rka4NI
sVJnzLy/9AyIPP9o2xQGR5sOEYPlOwYsarB68McUlWuVeGp4aoReyf3RzXUn1ftTRQAWJi6gcGmR
11oXnYDLR9Wlx0hiwxy7/qBsbL5jrxlru23xMxh9zDn8QRfTt52m/PQ7SlGB+TScj1E4HsVm/aJZ
X+1ZhW76rWp+uoA7J1EMKRoMAmXCcwpPX/KUWkN3B4i4lpCUmH70g0wcLbbcIRZDG2hvUisXch0m
gG3as0ntYe+Mu4ViQfwJFwh1Me/QVHv00fcceTsjlmRmbe9DTwUtFpHo8T9+dwGTdlFw+aeYo/2b
2THqbPmLtvG/3iGKBYpjEXKBzK2pEqzSRQH02PGdIAEfS9f7Ubw+vdAqrVJ+ndffbaU8TEG0XRtn
pcTNEp01gK6msnzAzdp6Covnti20I4acDgPrXGrtkRRo9DtaE0jpaIqI8rx0b0SzhExMzLQl2h9m
00r5Otv4SzaS/au8hQ1F+asQu6KSybqm+mIsGcXXzAwKS7rB14H5OVQEthzgPHjrZSoZcXm16HWL
oh0pmWBi60ua1R2H8IGlqfAFTW+Qs7TODM5rHIlM+b6VtjB+wVF/N2AE8UAbQtvRH3WYouDIn9Do
VtHMZMYI3otD1RaY2iNYcXIBsovZ6Qy4gX6hXOVhrQ3EK/a4EpOJ7nJDMkSDuQvgc97YdcwsNFf+
tbJeRPYiPpPjGBRRq1pHBxrp6ah2XuEfKoliftdhXeprgYeO2DkLUk5Lta8X1IXL3Q9oj2EyXyeB
BhOKRNpx3wgd/MGvorCxjbjUx8P+vkTSQqy+YVsXC5mZjf1c1Jf3Z6IDpMQ34Fh7uDPS0dc9sM00
QRFZDH5M0MbhQQFzv79DpcYlrOyQoOgz2QD6g4ilzaIKEGq0J/qa03zZNCBGKaZcWbHGKk1UynPH
561k2zOREbp/E82gmefizD/9OFdGyHo8g56G68RQfJaZa1SLN+Unty7DAHcwpEeneCZB+PY6FiPI
YxFfCH1+3D+6xLj17w13GyEtarBklaFWPJAjeYysJuHhgriZdGRG8ZQQ9VQK7vXJnrbCbOS5dTNK
m0TJMCSGyXTS9DCTHcaIjABiE0viE3M9EC6VC0Qh9T/xHvt5iIi5yZB+CFamsWjliraQ6eIXSn3k
zA4Q4sx2WFl1vFWc3Hni2jaSh9zO1LEa6n6GetLK9i/VYVpAGF98VdZ+TrDyGB+tGvoHuR2bdc/s
dp6AHvr89iMw5DYH4FtuN8kzbbxV/+oAqI243jwC3k4sxnpDtZeH4+n0m2n1Ektxe53RhXX9TZYh
YqHcTUiSC0jSNxOstolOJUItInQd/2Y5ouWUScqOWMvQ96DiVVCpJson7KmuzB7iOxtK0Wa0noAI
0tiLWVbcFCg9crA4GEMTwGag5gZBKJTTcob9WMlHraTYEItbEDEGD9PT2c6vrsgEZznPuCZS525Q
GDt0KIbtfYp38T5fve9aKVZdi2qfDcIe5GtuW8wPRkLeDDEGtKsaJ0gWKXy2iV3AdrkzzNEMc7qr
jDMU8KFhc655U+Yd6+mbhae3/IM2Fh0tiTKoAuH6XVSYwNeKQnayYUtH7FOrdQOXkq7nJFBfuoP7
Tyhz3czyWyuLLv+jef8lTEs8XPXFXd3vDfahbNP8jIzLNfU+z2LHIM7X/Be903cjeQaU3ZCNhEk2
DUFIbLvhVTwHiTDnn9qQ6DWBGjrs0mxAdn9bfLgc6t1VRQx1lngbrWZ41CM4a4Kfj/gBaLOIawN5
ofuw/3DF59Q8bUYN7GExA2uM0pncFOkZLhbE6/CjO0xqdbFiztxA2JU7+cVmNCdFlgqlHDaLgi04
RaC9iPRNTt6DBUSZtwlRculXwCspr81kR93VhjV15QbosobaxK/po4bf5TLuCZLaTu1XIpUjWMxx
zoPeOAcgI2pAkx5Dv4CmgaU2tPKKm0RxMect5Zb5Ar5lG4ZYEETcnlIAZvft33V+6nfEsimL50jM
tZAkUq13MD918eauH3lGKKicv/6WBqanpwu+ybn3zBt6w8gWfBJPaABcQu68tn2J2n4xyszQa+vS
mAHptsaHVVn3uYBGdHO3A/ZAXiUE9y1FuzlgnncT/d7/DET5qE9Zx+RVK9NqK0sTXYUm1/nyi9gJ
Zyuayey4oEK5/GgxzBKN//SLiJ8LNnc2CC4XDWYpTfdyYdQJcGDTMiKaTw3elCOYr8Wnw+eTrPby
fOz1e229D1Z6EB86SFYA0XFDrpTvl508J1qa7OfDi2+xp1BRT2nOY6zGE945PHd7GzTwVQStO9zx
xz7P+6YBFkBg6CI7fBJ1gb+IRA7JEs8C+XK7Xclh+A/JCxY53iq/Cno6x/aekZRKTOkNZdhTDQkw
QQsUNCS4P6jfdLoZrZjtAXdMT/qU+akRnMAzEUYs9LByKpvmYmS4bvHix5sprJD224r1izKupYqI
Nj1Pi0JIlkTxddy+OYDfZjTp92e2QpiGBW6eTT1JUU/HqhKSA9WALoTuU3uTevMWK/aZi7BRUWKt
jrv8+cG679I/qJdXnr/5LPphCceYe3uQWAA2AqFmTJdL/cLz6cdDMWwm4hKxUi2vi4lylIhL1sGw
hBuHoQfIG7fJe4Pelf3U+laNh2Z8gKATcgMQQ+w9AcWi10QzrG1Y5mHsn+Ua97cR5cIKD5zs+Wj8
iRZqqd2dqlZJ6PfheV1ywhCJjZlp9ChsNL7MNHsVFEhHVs6/qi6BO3foKPPxS1I8lQkfhxtGd4r1
cxy+KQizjR94uU/+y/YeFk3soMebXUh3k6y8VEXDNKOwOeJzXhaFfbkMJYHMjtLT9/rL/mFeebaZ
GxD6OQmxDkLWEg46k+Wg653BCnCTyTTLUgWuLVkYzl5lIyBUPthTNjzoCgd0GYZHMh0J4b5VttVN
Ln8+KHuIzkX/U2HI6m7P8D5m2Tg7je9RxYu5SXzP1oQia+SkPDIe/u4EBA3+mHFPCBYUMmVYr3EQ
mAX7nstspQmcT69NgERWH8/g+KSG/wFFAllv1uOtMHDXvqKuEtmN6/zJnzWXCimQwZl82wSEIDpb
wjqi/QQfsPlDeS2IGPc19WNnH91Uip9fnXWZOxehqkIuBOH4hM20pT6ucdSWxw0XSrxoEVt222kY
J2vomaUjKgEuvuR57f3MJKXHaVd+vAJpBbKXNVZg2EJw7616ii/rUereiL1LD5twCkXIM5qMl/Mv
bFcYDyyLOvZJYaGMLsdxlsbQ45PAUiN6aQJ+Q305wCTJ7UYScwujfAxzWxAXrxQ211IUsJ3SiVZZ
7OBtgBpC75iOkTvlHb0/umm7D7zp3BGuPo3CMuZi7gm0Fh/O4mSGsekqCs5EtTYIGnU/FhPQRzEu
7Dp6iTXOg2RnHe5Xje2oZudhe8avqzWk/WkVo2ngI+P3/BXj+Qa3Ow65xL4dQEET9s42QW/8enD8
T3SQyWgGFyF8mEqLKNrS63Rc5gvD0427z8fRfKRQDIYT0WjdEN50sMz3nKTj6rkEgBRgKYkcRS90
P7L7AMFQ9W0+EXFPri14Hz5zsK3ujhJPQFNMTEmHrEliuDKqsSCFVaN0GUdja7iahBA1arwDeVfR
XG2Bl92m+XDnK7A+egWs1rNpmFH7oPVEZ1LJ+YXb2oeBb0GrVMAP2kUtWIhE2HwgeOtuoZGmu8jb
QfD2XLs17MLpQKkNR6m8IBXdRnlzopkkLSGuhzRHk4hvroPeOMfQC3dqIKI+1GWUjp3Sp9CGG+ed
PvMGO1g3CXKllKfQAVxxmTQyU0zCwWPiXeDui0EdpBRGdmGP0n/zqB4PpQfU9JTxFVQvSuBLJ/br
FFDgxFa090C3MWF7KV6I+CqW3qyZfWHRoWI5s/SQedg0m8FYlpF01PJQf9D8F+kgrv0bw7TXkeDu
HwblFVsfwKDlyKumTQO2HvWZ9RjEBQmvYaYEx/RekfaD76J2Ir1c4ULcOqM5vhjm3yAvRGKeD/ZX
49FUTrRPPuQqLhL2lHb+w9OgIwZZx1GAPFHvbCY0a1H93IObG/RkeD0lIendKTvi9QCrGCxSEWti
HdzE/00Vr99NYUmNfIsTgtobanh0rN+rL5GMqgP6Z34cafmdZtbpxwgLFvsxfFPN0BPJ+3Dm9wQD
tj6y/a5XRTstJ/CXlUq5aicAe3Gjug/Mn4D/oPEgRL23xjznOMzfI3wR2M/TtgELTDWH+FldrRtP
WS0lwQIWyQ62a42XTzTjDlZePTdlrUuIj5b3nTpEiXKE4AcGlFoxgQS8B9S7GYpPs9N5TCS9bWX7
vYnPrzruEln8hxAfcyybU50qpQ8zCZ+n5qyMjYHk2uNufXxFmIC6BXyaCF/R4GAjoUyGh1jPLDyB
+ErvidixuXzVIaJeeS2PnZ+QO5ngJsvQVmLXCKACou1ZyXheIzJFodrW72Y58jU2vd8milHj3EN3
47r/k9BNfzRd5yCf96neMj5VEMBomIP8GqfqDZ/A7dHyERD81c5qBl3pS9Fde62yVcOXckbMvfEj
2BUkd1iXiGuHZpVag3abgfj17kMk9bge7HCGzZfixhWK6c0eJGFXifK/cdk0ydsvBoAMNPx+LBpT
MoyQunwPxL0YxysO3kts7TZgrkdbebA0mBkyiemuspPRrVR7DoVIcznefOXWYRzdO/c3GqcXqz8A
Oh6CAqjRvC+sHi7jJhlLjFoULjuojk8cDqYyVT65jfEKyGTCbpWYVwF0DwKvYo/Hf7bNwmfbwhMZ
uo9TC2Kp7NNeiOzdadyrTCvHWD8Tphwt0EbCbsa2Uzc0WSVwTa5yZK2uChDEW0HHFQCYiKoAK+aH
rQa6V963AUwQjwKN6WtXR9f39q2l56KwHyYwvdw5IoiJLWiUKebhGeWjt1V4B1e/ODVz0Fmy19lH
E7FbGdvnisfAfcC7BzdDrh2ZbZjf9fR6U/ikBOJXDXi5GLR46owMuJVvUIU9AM6oQxeJX9aMe2us
ua5VusTUXgemi6D/y2J/ZZuBRWbtcC+ShwUlTuzdcSM4bDVMpXn4Yo+PAyrPebJAHB5/nzyWMMJa
P/mov0OFlRN4NwjW9LGsCocPhfEzWvS11kyH1ZZtyFXcthBreEEWy+cVwBFY6itTc9uVB0/CCz9d
QrDE9Nx3QuiBE4bL+P626HeefMPz1nEbJUo3fhY5a8p8xM97eq4wS+qB3iPHZ5josTBLMA6IA/vD
aiWAiyNFFB9UW9n9MSFFLtrl5H75N3X6trHl++jPVu7dd+biUBQEwUGzUJf7byppsyNTIHdN2Z4d
6mVuxUMVtB1lxTh/AKAOYaewl/Tf/4yU1etQWSpE2j5sUX/7mX+eyD78m1MjnbTB51nfpKzUNdOT
lgXb9SIN8b/kRULPUadVepBAJPUWCkqL8D3SFqVfDp9ltqMXSACr5E6heXwqxtocwBtLBNTAtXdj
KIMrjwwsfhZ1qLh5Ae/DoYpAQt/87o14VoTytfjfzloN+T2rgMJUoSWzyofwFL6uiTAxd3phTFfA
KHIGCe6e/+/MFtLPW0CRqFZKc/VpcjB52dqS5wxEhjUMGvZuD9rzOFvL05sekbDpYaOm15VBLiXM
AHdL9j0Y2Vrzm9WSjk6D5G+okoAvGhK7+O4gC9g4XpN8LSQdAs8xsmTbXssPMDHKHA7j5J9fxW05
s926ANJnxgfWFxiv7UFVR+FMKrMX+qD1Ech/bH93JJhuCGd/J8vB6Fv5zjfhPMdMMKmJxvz4xWod
4EAWnNWEvck0ftAMLnaJeEC6a1POgCv3BjGAnpVogOCtYdpPdalUNP3mArfhxpj4hY2m7vQ+tM75
lP9cNS6sjIJtHlP67DdOtg4yN7a68NN1poGUvXnMWG5kmByWOjL2calfYGTDNHw43hphk17LqIf8
RJq5jMoCrAO62rwN5E+ys9QXVZyjkYWjD40oQrhQyN9T1wP1INlerWGynr2vA9zekXYYXAq1Hmpq
HenQCcAxEl+s7+JPIOZjTx4VHwq2I5RslDS1pG4sAaBNrUd2aLhaMk9h9GpxNRG0tFjQDFV3yBzO
rVzp5ZnN4UHVMjRFzx6bt6sgPend2lI9OIEIHs8sqSmGAKJlB8DGueNEjikAHuqkiSuG1tqcw96p
qM8cq5ODwpYk7Py6vpRgDqf3s0gCPYWvzRbHXt8AI6SpU9ur2buO5wzlDGH8f5ZzN+PjDNi8n2AE
u6irbtoJZXgIqRR22HNwO2ZO/arSO+0xxmOBEiYf2y5loxaC6mh9aUxPyGwQYMPwMO805gtejMoh
82rDewK3yTQZcdgZIDIXrERgYoDWDi/Cy+A0NFeNfDiFa5kOz7gxuaTuG5HD8gjv/omqWrqaiQW+
qlylWqWLW2Xb9Oanyh/6wmLFWyCCAKBkWjLMR1pBP8O0JIWUolMzY4O1C9NV+gMwU9AamBWUUelI
AfKQ6jniF/QcUQZXb66S1LtMHPjAXB78NysUxE4fSDlti77aOjlh1vYO/PLrAex3rCX0elnlyj7b
D2yGQNAwNYYXgKMVGS8A2AwPjgol3Amsq3NMahzAQ2kW/FRwLIOP+vs7lghaj9UHVQU7FzfkF4Wo
nGiwDJ8k44WaywMKp6lQ5a3qZ9HZGvsGr9qsjogPAsK50wiK3sWDjp7YONB5vSepkwDjEUTXM+rb
vDHsUowPX4AwKMbyWCp/Epi+EFBLoXpryieObVuSXe1PuwuoIrq5gZChOGxRXr/Rl+FCtwF8aFu2
bAP/qdyV28S8A/AXzyrfY3K376WT9plXF9kNKcKfGCAHJy819mmtym/HoQ1COdtbzCLLGrhwLB4L
sH6ob8AeR7QJ76YBinwXKqX9KsBYeYbaANArK+XxuSS8WHih1cC5Ps/3X7HFmfvGZOcdY5LyAVAP
ez3S2w+tlda/A6cImDC9rjPNDAK5+3xGQFEiJLQZngsEA+x1sJN0rA7ADL+jCzdpnSWYYUvtITHd
8b3RHFdyG/15EGSavSPpl1tCm3MpYmDb5tRzGtnXELK/0uQacYIUKv42DjLF6ljcg/xe1GePnb+l
9IMu8E9i8b4i2H0UQMs4fIz9oDMQZjdOMrmTUVMxy9bLbba0PNttC+3Wq0IKp1fl4jmw4bxfIaGE
gLrQXJTUgMIhlKIgmeIx9zYfufZU5TCx84Ve0uCuynY4tzs49YzBt6gvsEuLPx7A/oTDKk0jtny+
OFl3BhJth7xaIoBknOiwwNU0/uFU25xbTCdu6Eza7ifsXuzh0l14gEqoMlq4mv8qtsP1qwBwj20i
ZWdV/rY3g7+JclbwWdp3WTjRS+udH0rVcU18+uX7+C2hWQx280yzAWbiNK/CnUtbCvCc40bN1BYi
tSKIkCAW9e9Vx3ucgruRBNFcDnI7WcUwJqfQqeus6/Ziqd75hGMOjMGeYjPHbcL8cAKOrBK8PXtL
o7WDpI3zm1ZLxWEoewKtONj0mH/AT6xJvqdT0f060/Yc54BnkL9pnTYwMgq5uo7bKVAFU7Yqn8U8
umxZ0bId4nyOrkeWwvOlcZ97IoS28bwUtR6kpSiGVBL7phUzMqdbJ0sLTI8pLSx2mtgWHyTlyDpw
n8/yKg4PVY4ZWY6Qpd6wcqpbTU1m0s4tlsrsgwlG1dA/efHAszVPGRAz8DxFO9yZw0oq0qI5tNfi
1WR6vocpx1wFAIUmglIgEB2KngAhPAugzyhp+On0KCDvc2NixUR/EIsA70Li+LKT4rfK+n8huXka
dFWq1RAHToV3vqQSw4+8+SHijpY2hV+u18yZqYpfQYuP7XJt0IqdbBCSuMNsVzsbu8ZTb9IvOed4
VG98E/ajXSGGoMeO0uHMiAJSILq03ITP9i1IQcuL9cv4+uVQMDhtGF955m6QyIi+Wy3YNqw/I076
nlhnbvOgLg1oSG22qCRwuKTw78kdKBuBlB9lOjg5/NybKHGohsYdgT4wAhU+VxCV0TwA5G0xo1gW
c/xeD1k00IGXe6kAQSHPiPsnHP+KNMoFsxhisbD/bf+ut6nj/S62K3dMVQ7aD7+6hSEhTl+3n3/f
5Y5knEdJ+xeswFxpQO8nWpUgQb2bQNKyQ+EtJ6EvqqGU4FOdJGBo17RMHOwvC3yuCvf3MkGiCPyO
/RO/8UBlo6OKxV7ffaU1/Qm0kkwVR0QSHB84EIxzyd3ffLlqS6liPiotEot+Trk2qIyrzE11GUl2
kiL1OPMF6LFRHs+CSfHnHPJ6Dlr+8aqUU0+k+9aRvavpCKKxCajRAeVefnPgFqHa7FtdUxdqF6Dd
VKPbOaaReNi/qQxwwqvXoW8YotqhJt5+0C8f/IcRTqmgWzURDH7pEIxzJCMeYtbvSkXS2/GBk4AV
+/ZPJOXMTnh2mXxqgbcXzPXyoQ84a7yEY9g7TJTvf4mmvROnNkMcVe4Gida7EeU0Jl4s5s4E9OTv
9BXsCe1bDH6rw5QjrqcElyQQ9offdbDmbB6bCiQbUsR5SINp9CWugExWu/TD33bO+3H0K2MHQqeC
HPssQZQA6Om/qB6ip/4IsGtBTBz8trja4c23Asds94SKTjfv+EbFj0rtse0Y7eU4fpkbkIaXUVY6
44Kb/DsT3jTqqjHT/cIvwjTEN6mz7H/NPYefWMSMasSv0oNOppRgt8Tu/c9UwoIVIzD1PKijF8Ka
QlBm5rICNTwoOA6ZUxS7wqMFtI5yw0PHWBlT0HNIlhbqYusdkT7BmBeSNp3QcT8aXjG40fJZkt8o
fF6JAE4SmseQvb/aOBkbQPd/6JsRmLePT48XdNM5HwVMkrUVauhFGRHwCC7EALZrXXObqeuLF1zG
OLzMpaQBwG8IeW9M/A7AAesHqZbAt9ltn0SH2snKUUbKPKUYsEQQ5/vN/OcHsYg0fOArsfYuiWhf
OUCP2Vw5fF7u6NI+JB9DNW19nZZXQGfi2RWJMKVW5ru7lGALAgx3q8JqSzSTS1EQWr5H8FJHNNXI
0CNN/GkadwVLQioiq5noGLFmLogMZezxNbvbQFY0E/CllBPjHzyBQa2laufDLIH7EQdRMI+L0AGY
hBZfm2DSko1Mogsbs3etfEvzSAHepUNbhZMB0pkOJjwSZ3idEQnxB3r5mXV/CGm7nV+KcHKrc2vH
PFdo5I4NZ6Aov4CjK7iKCtPT7Bb1PZUDk61c+GAqoazuv2tMgdhrivJyaSdpPpWHQEFtEJ2PXg16
mVfX9yywVTI20Hh/dWLd1EyRLtGmLq46BWb9ddu3SqBrCT9I/FiF+nKaJY5isDw+C/EDVTg3VPjx
eyrdW34sRIPf+Rm41utgUvzGW1cPxxc9ojs5rl2Trg8tsq3QD9EaHbHcK2eYw1JgS4YRGqQoRCJl
ZrtBYDhbMg4vfuQ+tyByeUwBC4rPqzS7oaaFV27Z/54Ik8z35P8oEsvgmOFGRSZy0iKBb9/p0GHV
98Vjm3zmYUir58C+Mx/yQpobDDMDsiiF10OErmuLZqzBMG8AHhQNDHkMa/NgBvvtXikq+dJ0VnG9
ZO9fCqn3mIiuaVOZP10YIMGV7M/g0nBWuA8gs8ZjUfkhRpI39f3FrT5ADR9MUGXesFyq8fvwgz1u
i88oobSAe1JHB84sTFO1AuqBZSHZoT+lGfZVDbF21u6xI+GuLG3ouH0TTFm+wLig+oackppJ946t
oZKBseyXsFOtbA3SnGhVJBrYnLV7QYhEP2RXRKFhDTwfLsL2WjiqpdoyUAokHe+EXvvHTebkwCIY
sKHtrKvaEKKif3pO0xI0AngwtV8Z6v4o4ia8m62odBaJ9Pxu8j/0SLbNn83ZhciaWpughUIcJE41
HoMz7UG2VfYVqS0ylkNeDjuUL+x/Aypfmh37848jbdVBNo85pBPDSeGftjNKDY3Bl0pYpFGM9uTy
MpFX4mWELWIzWkDyT+7RBHDjBfdifZjMqwYafMjE7ytoGhUhOSHURLONUrSjvIp+YjqXhA9QAWXx
UIffEKkB/iiLGea49hPBlcR1Y6C5zaRbJCHbC8EvGQh4C5b0dapXJLeA5gKCIcl8u6J56iMzUgg/
KB99d3sAV58MwkWIXyTwt62lgmsFzdnBpMKWx7Xi2Qci3Naa57QNZGRZPDYGTd3uR5eT/r1NxGue
qR8leKJkCBaIY7+j0IkxXaOxeQXOf88IBLpwEfM5NayPqggRt7J5sbkpKqzQ4MLgUoxd8/5KGtPE
AW+CJRx43X7+JjiOFnOLWre7je1cDsLjvc6A9jcfq4oJQCXN+WEGiEZ/95CZB7ZalhjFfDletBQ3
Rveph2SpU5tiE4j0LZSUKg6CN+O6DbCM5Azh4Y4pB1W4GS7C9k8TsOlBZHYtgBq6OjSoWgoRVasU
PJxih1U3GqUmAi4hY8Qmw+/pBhV5/zoN2qUn5AEW7R21iFAaeDURqHIH74gP3uniuLz6AL3KtvVP
ct/mUWImLvD0ROiGqOUgv++OkWlYuC7usRSerKawgkDQf9c5alyEc2ZQz8QdMYGUISzcgfH0GjbY
spew/RREvYLzw2bak/npOWk9xXImqcSauoZNcqOyAfLBowYrrwNi4sYpd9gaSpWby7Pq7CiYTmqM
CRTcwCQD3UyN7bsQITmChb+BHhkyhJxVVFlhTWUrqLqvmaEL4HQPi13vy/g2gP0HGgT3DURuzT1n
wdiTCDURzwuY2HA+5VtA1KSAQBm9n8HUjuPo2WrcZ7mCCxgmho2chb5d0qylYtSSAeIDdea0wBoG
M2+Qd7QxUGjDHiDtggiUBF4ipUPDBtptWohM0T8ygesHZBHgaiyWETWVv9VkBBF3Y7u855mZJ4ns
eUQAjN9XxqYCnGYNh1dYVTvF3mC7iYX0ER6pTzClYgrPdcml2ooIm6w/1BJQet6Xsb4LKq1Mzqgt
C63/m+HfjCXSoRIbyIv9lr6UdUwGbPjqSuk+/E13YVm9HKH42UQNsZdQVlytXOe2w/nP1g3jaQ5i
+ON7my1qZUhHK66ojyUiyQe5z2R2UMCf2Qhj7XDyiiJ6nazPQKYWp9QMl4DCiCB5BG/M1rfAUKnK
1MGWmjVgCaAMwJ25cd61kNy2iEtbaBp1CR+XKePfUniRk1eqkcTXMjUeLyF1zDam21px/4QpWe65
2kqyvyBleVKWLw4XLWC07/D07Ij193qhkNBn2ArDyFoBkOEsMHTHu2g5KIVRKpWbBvJmghYp0GJQ
oN3J0sX5X8epab1JEXyKeROWrwlyoaSOJohTUUDR8hxjuOf4G9Oz0u7S97iW1D/5HmHEZuAAcJTB
8yecHo0tDgD75GKQJxQlFFpu7ev4foouKk0mvkFTnPgPvlYB00nz7sCDPzYqrbU8VW7V5bxgyru8
5UUp69n6Uezfa0dhHb01clTiS7f50hEyIyMb0DZhG8JtbvJOb1g7AbQZSYS4lEXBy7hEYOlUEUda
nFJtK940pqnevkKjP8JVp+GxWQZ4K9FR8YG5r4qwKLXy+cwZvXjbXIeSwIyUMK4VPbqDz6RpFFuk
yzilP8EkaKbYiax9GY0YhfYkMwbCdAxt2uQBjwKhOTDzjargrfFRrMHQGX84jv36J/P9rpyJd1p/
nHPGwPmN5uN+hPJjbKTZaGET+fXOe86ZrWm3+8Xv3aaPfkOp09hIWURYt3HHCXORgYTTRd+uRtmz
CdiqNm2RGSzoRouLzu9hxQCoV9920nRXHthNr4mB54fKXJHMDSL/6avUTqMqlyRt0P0R414IGKqa
0LXIw2tp6F2HRIcXtnkXSBqCOsnsW9KlfUwg7Q7Z2B9ccq6xooKh8hRP5LWp1UIXL/qOJtQ1DcYJ
ikl/uYJvggMN4WDgcl1SN4pAm9Dvtt9xVU4RH64Tm3SrFW2lCUfEPhdXjGzY7aM0Tfd4FtOxBgtO
8ilZhbCx9UVD46VyCAHnujZgGaDr3bCGo0ErsX2YbZRqOIiLigipVZjzDn9o2ZC9efs85J5TZVG4
zN1UMp69kSBpfg0DvznRHBZS2oPv8KirpaiRmB1Jpjpf9i+LEeRb+4HIgi7CeSTwwUfImInMIew1
TQe9ljmqf6Uj3AF2m4kDl2+WF6zF2gMgvgtrmDFrQlIbgbSacZrjLmuAjl6EYSUw3XiglNzmvBJd
t4iZb90hubQxaNrGLWJftNrAuMQK5bCLc+ohCVWbtebRIPxzMAhZhfh84CNd/z7OJBGhfcx2au9J
SHhK+I9cgJ0GJjXuPpY4a7chi0vzveiL20HQiJ2paUh1dO0h09I83yxQuRfmDowRQ2lIMnHIhAMz
SgUmk1/HpZQP25n97sgmfJ1cu1tUlGy/NJD0wlGhOrOZ2GvFyoSN01cLTqa0MwtW+ieikchCaN6o
E3GzI4a7EWYWJn99+VgHWCyogNpzOjsygIlxu9J2SXjJdfwfu/8YI0BHy6XGmGRhqY45lJQG258r
zMBvhG4lmqYfaKRD/evzk8/oacGMrktIHB6KomzlSrhpjq0B7ySU24lWXCKrI+ZwQY0APfRLhsLH
UfosjaSSCIx1ajDdJ2Mx+VKuPX2X0ukFbxr/WjrQ/GcmYcD3LCu1+A1pUmDUGG9fVqyP47IObTO+
Ryd1vFhXYJZ+Xmo/e3dzYJ1qgNLJNvFtgAA3AAj4ANNbaQPniQt9ZpozOZ6qY925HtFNDkyqul9U
Jur+6xht6QpM6ejOGFoxt0qtxyZlEw+ia4Mvm51v0/amILGxZQGMAKTsNqAUzCpNVhTZqfC9RHMT
mVj/+Or6Y+9LPKVGmRDiPLPc+gLKwxFjqWJm2pkALMGMbciq8mGHpyJzJL2Yai3oNXyFp6X99SrS
5MkXpqKHw2wHRkLf+CAr6D16QRvH6cS+RUJu/lpKcV+9HRGsGu1K2QcIJZE7AzqkbtqclplkBH2J
OJTDXnJg7AqxwcM1L3hn6nxURjWun3gCdQJlk4gecx4VuKnL/kViAlyCT/bJxvPl74JzuhwW3QKq
2McaElWeZ4RJQsQNHQvQAbYeOLIrKSYBn1osjqmBFze6s8MJ6YOP//LnMweuLpPXCNJzixL+s/ff
3U7esKpU6LcYOV8ZU1Qx6phywjQAIxUjlj6crZddSPPghguQiukKDUFDVue+rIUZKrZ08ZyhZ8lC
hpdVrGeJ/YFPmhh2vCdDtrY4wityzioMQwUBRy7DsT0F3Su487PyWzahkzJb7Wh08EkbljMPbgUe
A1gYMLWUVKVkpKngrgtOU1lQJA/WzLJPntb5Bj3GDE+fvea9nqiyFxxQrlpL7zUYUwM/IzGqoDt6
ZfT6LlZ9B8BVz7pK1Z91U3v7ttHo6Tqs+4kYJDkL5VHyn4FVsOk4Zf+qXkRdH0KaHFRbBrP0KYCa
Ktb++QJKAQEGr7AIlglTxdvW7qTJADf0bifHMBw85z3ogoOihHtUnT8H8q6IFWzsff/9UdLIppP3
9xijiU+1BEGLWDrr6+V3bvllF8lPPhxjmu2t5a+LQ4ylIAgeLv9QDoXXgADgslDw8Gfbu69yTz8g
M7e3+6IfDF+YeS9DWZ7j5rSa7AulkUnwmXgj7Po1Y+8lJFUfqFwU+96WyXhIIx2m9Ms9wn3Yj6pq
tWCtXCjNUpSgHAu0MZQBK11chiL2opAMD+J7DNk4Z/LDdRHY42cGEa5GOkHj1gZUoXuRTDbY8oMy
lj3HhqW2+OoxyloV3+f68e6I+g1dLC60TJoPL/hxOooWkmruW5rL/v9Jm9PwBS2wnnNCgS3cu7GT
FZuVSvORPVtgQLxu3z6QfeNrxcpfdC5CL2vz+JLkxlQdzYOr73RN3T5leuF6NTSUq2g5FMknl2lV
ICMNKZowavHGg7ibmVKfyjhH68HWrLq7NZE6xbYHnr2ibFkc3+IDo80fr0EC4BjfdGp1V9r8G+HM
DTdPq4114XLsfQqchGNyPjx8hVUtrp1JTia1/2lUX8v1ifCHINYXNe3gOYc4amzsXK2hfRsYcDFa
VZGtIw4GG9Kp0I4QlZFevmIDTucKnDm3HgSmehY542mY0JcGHVIkrE7XRG3Z2Dbt5AMv8ydHfnPe
T06CgIU8l+zTDvkf34/UX6lNbHyEbPBZbQv6fHYtkm34ea/hRmfuhF/xL+hwCQB7ZdMmEf5GWvz2
WAUEHAyUiUAEmatQ7iWe4hmYx8GqtSOMj6xJtvd9LGqJ244YEnxGYT400g9WrTv6s3ODjnoQzyNS
c8kCIq8Zu+gpXPOOUIVuFgYV+k++B0Bh/tOp49A/1eoSvCPlBWJXt3c/LkldOB0FbdZ/q9Hc+thQ
jd8HrdVITFpeuDLZEji0xWu6ncth1hzL8kFhm/a5dpZgZvhQPOwxiIsgoeSR4d4tSDEh0G70TLUE
2WTbAsbmsY6J2yVWrO0b9MnmH/bmIn+6MArYPL+j6GWus0Qz3XH059GOhv/75Qniph+goVcktNsX
9ApkaptoKWe1tjziNazcjpf3HbJbfU+WkAVZ1uli6n2XpHdzJQJK8MK2D/8ZRJY0HbcMS4P3w/fx
xD9JelG55Vf+Kv9k+sGIgRFjFgWFM1AFZI5km0kvocjimNjUAS63hyVbkYgqoiUBuJc8iK6ijFyQ
XnFQev3P2taEieeDv2lLh08ifj77xeipqNRYQz0gTnwlDPFdmzqNHnM2J+QiS+wsXvAnBU+7Okey
ku/EQyGwcefw8JsARaI8XPDjRd3JileL3U3WN3AU9/YauFrHkEnpDg1DjUO2SrO87kz4Be2Rhk0b
yJ+4pQ3n3yn3sd2tqmZkR76+WPvFpVlEQ4ooS6j3iY8JrFnIgWyY2GddOWfi7Ujv5WN+cIiZy7Av
HHw5j/1KJfJpe5eijfuc1PtTxtvTIV58KCDzbpV0S4pzgKu7pXI6HY220Ogbh2f+Oc/FkrbYYaiU
p2RtILgYn3ki9Rm52iRb3ZNdPeutUTGeJwPaQlCu6JZ1bJ/Q6Gt8N3PKGkz/4b5i/1dZf6ym3feJ
x39nRCTcpTnmD49UwE4+J+XkA1e1fAtSMxCqO1cjMKopJ2K0uATievB/sYpBYV3G8rEfjahJWtKP
5vo7M+hHaOqxAjW/e/FtLjpksb87uMhcAjlU8P9U/UWOdei7sBMFlzQ2i52fIjUe3Ja62LzpzpOA
diErAd5oZ6TgyGGo8kt8qukvXNfRvSuBA3m/BmspfDqplLX4Y6pVUgt5593EizTXvWNW61b/c8Cp
zBoK8aZgIy6gyOgdupd6/j0dRpkFrzB+FftbON0QnpTldO/8QJTeN2Sc0QMKodaSfLixyDvHp0UX
hmVmDyMqBm0Jv9+iiX6UjcrQXzU9qIpZAIG+Juib8cl15RT3Bz9XyhdTcIm7MGrH4w/c+1U67eb8
tJbxZDineKRswaqrfqYtNcXBCBriSS319HmP2B1e/O9nbDn75XBS4RuppHtTuXoQMWvBe2yv2w1s
S6S3Px+xLyigMgEmT6Zw32W+s4Oz/vXbPMNzdZ6pA+Q2SxE2LQPe8GtPEUSd6KhOp7cqU8eynHgM
1MCbsRKGegni7BgpIXblIuAe6mQBNgkCPrCQaQEeqJqFkVAYBzTCHrcIcCm88KZ0AoTDblKbLjP5
JOhi+3lKRW3cgLgaBF1Ng462piEajbfyaU0cMZjJ+JPpKyp9tzoaTba9+TEaBWivv9NeOa7J/S/z
pqbqbyCAy7fl//sYrWfQ9Q1NnL7uWGFcjwNHNRuCNPiy2PDdLciCpjuqMof7/68V2NS3Bp8rZE0R
gnKrtzq3NRJGL5PB6nbDXnNI+G4Oydf6Jwm/aypPkPjKAKMbohL0rx4B2a/3vKodME/tRz7hFva2
vTXNdsynhxzuNxOiK/sP+kBRoDKISrffmrT93bYTrZ91wXW6txnX+x837NddC1rraGOm23A4CjZU
AQSdNnAmY9W/ZwbAmxV8nFd0+1YQqQc8bUlOCLD5wEUNBgZflc3eCSX/lFSpW+qxxwR0PpPqF1qe
5459kqrn1BOYvlKL8qRDOxJXF4bA3z8GzBw6IMgVUGYKLyZZPSpJNk5z1oDCYLQk0vklgDMH1fbM
z9T9+0ua/ynLScft3XaE53zVd1knhBlewv16wbtX1x9Vb0O4iLyn35r47rz7y1tJGtG6jomoP2g1
LPN6qJ5536CtpAGyc8nswY7rh8Mb1hBMZ2YlvERPqgabj+X6TSAazJkiwxCko9Oz54hMiHzpM3aM
7zPcc3ikQJeNDRO0xgEgIKJ7yUS3MHw4TimYtHu9JlFPaopbpu6rqPGsK39rR9GtR39yvCn6z4cb
4v0/22x/SoxtyQ0SmPJZSTsmvyMGRStxc5lXzz99HA0WPR5y4HiCPakLT+KZV/mrDwwA8l+wVBlb
hyJim8a6OUhXqE+5mg+UhCytNhZtYlT7bCiiF3AENeSgrMaTV1hNWFBikekUcSixY9nZjHZCOGuj
pYaYw7YPR2yleH8ZGqCRy5g05ihGb5G19usWF6ihdmx7UxKrDl+lQLcePterQRuhuqVFCHaAMgo4
gUEV/b0RaT5t8cwxft+i17M+c3xMgUv//iAWJ3xVBBZa8KE/qa4AElCOmJQpGe4KI7wMgP3K20Gc
SqQZG/T7RjiXXoBhnX/Zit+Qf0i5xCAquK11gyqG9Lzw8aufF6zdGAHBylAqtVZaqZ8gZpI3xiNj
LLQ2paQw1I3Vs3G1lkYMMa6FdjwuGSddEZkDZb1dvusOJ2pd1PvBmEUeqNbIOGv7fiudZx4chFLz
JQV9qTJhjIgE1+1kVDLBjlYouZGXPGKoFIRJaVtGRzELs+q+k6lAufftzwn+eOYj1kaHaDlTaYNU
7oYxjvmkVYQoRd6QVc1S/r62poeeuxT/j9bJdmE7oBzbLQ8z6cGmPeR431o9CKhV8Sv9K9EmSFWe
kGPkSqWHdPfWmWIBXqwefelem7DXTKhJfjX0MGtTn+ETD1yukpcjKl2cw9YaetTw23up2gX1hUvb
BrJDU+M5z+ph+0Alf6OEi1OR7CV7gPpu91LQiYXk8jejTRypy1iaPOFoS7sKxdTNzDbONAXDl2Ia
0pZdJLk3PPJB9TfzNE+J4fhV8/Dfk4G7leUzJmNdZbK1/iLjq967j2Umagg8Ilm1iLmDy0Ruy0HH
eAfukDB7RiRjWQDd9kNhe8bD8OIf/yEqj8jSnlMiLeURP1cHbR6AAMSNI6s2v+DgotUvc8lpEXN4
TShPbXURV5AUtB43m3q/ip5ORaQOkzbvNgjXQf86eKtNRCOLfgRrrihCu6JVdzPEiE5df5TI2NCQ
AkeZVYWKjmYpJIlSLZzJ4ZoiztD7m3w14gFJAIqBN6BiN3qjrgyf8Ezet/EnNYZ27zppBkexjct4
vbfMABaW02R+NcCz8VaU/+2kl+O06tmxNnCj1hk5NSI8YZnprP2SOBWTm5K23ezAL/rTjEqI/Cf/
51rwOJFXiWWwZRE0JIIS6wEenjSZPPOIFIXwp1RH71fYWqmEtryJBZhLfbDPn8c2ByHTt8PnrfCz
xSCPlEro9HTdtWwOGWxbgmC6bMw9SfrTLIz8dM5z3MN2Jm0za/a2nYDTOYgtpxIB7V65BFnQaKso
7WjI90wvmwLAbrpoameA/k4AEHOBF1FY6A+XVfIU9nMSzqN4TA5BpbsmoKTTdTX7fJ0zzS5i+Too
54ux2t0DAsCSTCGHeEMXZ6g7UcUnSibhaz7zEW6+dm2LkMwfREtgoFtl+jjHSLRFUjIQmzk427UR
rylDm05EHhXXIdq9qiIWun0NoeSC09R76cytdQlc2IFtLEjF+XxnIKXRaTX7dYyGKcy5ao68qoF/
r238dPZd2X08ZFTGnodKCuOf95ZKJxFnrmQ53Rm7kRG8vxI1H0/IfFRpKk5s0VtkfcFjl1+eaDG0
reTb1pWclbIdYoCcRh5KCCLKoQrJEGbaO1g6gm0P8TWpUD+HPvbe2bIZLKQmyq3YhQmhOlqftd0a
rlvZojkMoJExH2gwTBC2IjFsfeczuj5qkUq4P2qLSlnD4LErhzVoGmgqw1HeaYTDkCV4DKPIQ8Cj
zHnVu9Kb2qzx/riaQ76uh0uXHCptH7zd4o/9b+j21xWKHuZ7Ey/XR/fVIzRLjCklB0YP1jJDbCh+
20G6u9K8Zpk6MtU/WFtovNi533T/DDDRoe9JcLIqv6BGfpRnq5Obi1WAukTDNSvS2W+wZrgqSGz7
K5DkNwIWpux3deNPJppIDvEL91LEpNzMwEoZNeXMe6H3h6iJB5pA0QaEj+wQtW81ax7CDD5IHcCa
FQeiwFm7St4Fti+iQ6R+KlgPC2eMf3fnVIYTQTmMXw4Rj+LRFJjIzixkuVzuLJM7TJPEK1Wqnl4j
wduJVaHDfgdZC57jiNtujHD84NehR2XkJdnL4Fct47Q/Bg6nHu93kdjXmMldFC573L6SgjGUv9+8
XcknPDkWZEAYQ3QLC8YxSUISnK6L31q/VRRApLvhipZVW+tBduRir/qspRa3qBE5JG5XueyldSUI
De/dORvsdVu8jj91WCJjIf9YI7LI7un4ID/yRSa1vtz+qaET3Mre+nmueR105QEPezxJZJG3b5aD
pnYXCPPfkTijad9rgrOprScDUSCpNYQP7aA20gBZKBITIN7rQMcQAs6tOugYxmAmHal+MgmNJ8h0
euYqWVu3YwSaXDXOHCJrwNDYf6ZHNxjkxdwhOPj14tQGJ2TzYGu4xnzH1hpdYzuKCZJNQ/Iaji/m
mDIeYcYTXs7idO4yoZ0ROjpLoZdMEOwRZPLgMNahuIaepm6AMtU5l/X23HB9n9t2/p6knXKNfkZr
Ax9sVHLJFji19jgQjjNyHrKV5f691dJ+ALh5CUiwCZGPHLVAl/yjPygTI/bbnCLK1+CQYjnYKyKv
yTRUU6dPEX5PcCGrTsaHpAltg8leBpCNzUQWU0slBJzYfs89ZlweWpLmvjV6vP8O77lvAOMdaaTI
7nA1u2xur8iZdAwoCYfdREA0NT9Jso99sECOi5v6t5DBXsYPxTC5sUiGKScjyGaqDcpfozt9hNKv
heUk0fXlJxVTyt8U8ooHPa/9b+77I12a+qj0r7pZP8kTkrgmoEVZDc6zVEsQyckhXxHrfgzmOA4t
Ph+ByLenfmA7NclQ72+ATtNoWRMdJawi5MWS+WuDIw/4XUdn50z/9CJrNxYlkpBj3BQCTDV0wliY
zWg6qX3nXnB8t2iqrdfclfo+0K0ngXDe6MIP4btcUO2kV8iaQef3jGV5k5Mxhmf8DoeKE+BEAOFe
gxKma26BfRuowNbvX8vrtdQtXY7uxuBw7UgkCICKNA89TIdzJvqyf4ZnbJ28LvgAhYf5uE4+Y7Ry
JQ/xKRIhG1KoOFrkNQhWA0ZWAjQUJPXW2nLLvtFF0OEYX+7OF52YPu/sPm78cxYxjOUKMrc5naWL
3IBDzklrHr3H19VI7+A1K/LzGRY2qytL3AIelMBpFx+LzD9+ZimRPjT8+iqj50O5UvZ22zvpERQA
dXSlR+w8TWkl2iO4K0OB4S9frGWEFOFI00v04ed8mpqsy3jdNfCd+YQBpdygZhfsB6eGoT0J4wEB
mkxuwXNz/LG8t/6RuJr/WNq16gGAvdbSdtHix5zO8b88TLnqBoZ+mpb32IE6iZfTcUuG6ghNZ7Yu
WNJGg1fXAqfhb5hst1s1NY4zlNt/mFAcYvawhjKbEZP3WUAc/KKqPApVRuJIf04b/A5ySHOCabhj
w42GFm+js/l6/m3DfZRTYYwSR7GZSn0iYxtKGHvzB89Jzor4/9k1M5wYzXNUBYs5xN+XhVJhCVui
L04qb5SPFhF8RRfhjPUJoOFgIruBgUDlqyhhCwkszj7w4atVRZmQg1XCQuyHh0X8ZvbL4s/4JAPW
V80I/XnjRjvBQBA2sLd+nuASVCB15/Zj8RFFsiEZZtX1APS3AcQozdm79IlM9MuOKR26fs+8pQc/
OfY7MQhiYWWWWz2BEFzFYP5jsXkkV70SwY2zddj77s7czTTSWx4sesLa3w9/Cq5fy8qLEfTmcM7N
dMFl4wMV1sHLwiyrOW0e8y+srIEDXYSZzJcphfF6J8ldmEjNuJPBiHLXlkKSJxiasonvlaUHot2l
pYfNXd8+8T9Vn9bdv3zGNBulIrJaF9AVA0Y4XmNEdxyv9tJt51qAZMWrY1q93l3Gxl5vtCRxDhLP
vT/Jhbxl+8xqc+qmTk/pMv+wi881+OzyjirtyVJSRvQ/ihcDt+575+NcmYwXI3pg/vSc8GerajRJ
UcJ1i6Lh7tVeetEUnTWOZWl0LjMpummEWwpkxgRIg2B8lLoVSBUrsnUUz8pRtrQwqAssRQ09rjsa
ipIC7TQHZ6OgoeupGOLUTGjqWRFfgQuQwbVczcEIzXyK9LsMraOaONUjONKY1hoRmzMV7HkWYnw0
H3YQ/KV23qlgitUHVryHpwWa5PytzcDf2URjnZ4ts3OLQNsGMTBBVfYmKn18kltpYNW5tSp6xTno
OqHivV4g1piGUXRYBTM8/3r5wd2qHqxBRMefu2G6FyBv2Clx4ZDQgoltBnHnjlwi+hjB/36WRA1b
qYVAEpYgwlC1YCxQU0xMbwf7h5V/j8pREzC+zC6nr4HVaqYxPZr6XDO0gH1qgEKRZkzV/3rRA3hj
5sUJ4uRR7bFGTFlTs0C0cUomhHJkDFoTInpFjWO0gMVrnrlK+SDvoKKUsP55j0EkzfhjRl+9Mf5C
DgWGTHD72SKkofg23QsVCb5fN/OHla33e9XTnA5dhUZLKgdeIZSqzxHz2Hrao8WycdRqEmaNY1oy
Lp7J6uXMOiMPfRBeG6H5yJrmUppjtb6YodyKtuTf9joLBoKhl2+wcDtr6slNRpcx+eSPecYLg7BF
Httit+PHFtLuhKeHgnKDB15EbnrQIhxBHdN8UYWjJ5Pd2rbI+e9QOY2gNjKGG1GcHwE/gCtjQ7QP
flvvHXhq6w9nbSXTfRoNOyGKruMmKzNzglbdcnVjHgiM91FnVsMb2WZMIbJ52D6Fl8rU0WO1x9jP
+N9zsn7a1KCsHKafeqm9ElrON2O3jnhDcghZn4ti4XFRI1sekDOaMAoKQZO//VQf9XCrqwTDPGvv
lF0vJpfhB4IjrU2Tn51mRLeVpLR3dlSQAiF0kmlofY6QdnM51C5xBpUcvn5G18KUNbPKonfF0Qz+
JL2CJHmbEZXqjlBIkPkyWrFiVgtRhqm5yKaOuj88TsxIgDQmszov6/+OLAQWaHIPetovepUynLGD
5ATigUU18Sn+txeB28Dd9G0+fUcB8oFsPx3yzmOXaybgSdyrzsZNAEwmJBQJPZx23HPGiC1va4wJ
gR5nwFdOL35gOFLcg1jXW3Bqg6iJZmcfmdHViENjAAXvdr4fQOxrlmBwW6NgVvK0C7VPUCnd+WPj
F1bq+WWsliRAkUkH/AWhBvfkL+YBfAjzihc9tFhmQ2MxUj/QgS96akNlCQAfWty0XfnfZXxeSTMx
ggQlbXzJy2twoIGB039ChKOeAnw3gPor52+jZCKxZHq1puXRqEG5wLAxk3x700RGrjivDn35nj1u
Fx65K9n81gOycJEO9wnpoj2R3Y8w4SaumqMgZB55bZicESLlQ27xCpgkbjkhtdBmc+0Mw7p8sXyD
fUAMXHSXs7xY3a+DkiiULpgk92Zlwx04rdidSnSXjzInzfLOrJB2+2mHgajh05WQ55nF4L7Ry/K/
SEUZls5TNRhI7nM8ve1ForkPDZK4RV+FYVwXCLu7rKjkIb+hGE2oUnE4L83Ix7XUqXhE+sLegi3i
lstBHKjccr7O4M3c9og2lP7PlKkXHegoCNh03oIqJplKOMEsfSdTDjUuTVswlqBiOhBuEWMAwhdu
wdZKMoK7N49/idIoBf90blN8hbirnZP4TuFJ3uln1xsvBbaBtb9TVEllHe8zZouWXzDs7q7YbLK1
MS0UPdPdN8WhiEx1geFKoNRRjs8LK0KYsJQhcthL4q2Kd3B4QFtIZEQ+HZGnlwCvv+iw2b3TpqJV
T4fG+HyM5ilPTGPcq3TRNuilcYI3RrEVpCkfEfS+M0yVIpyyIxai6zRl1hWfVLWSA+cILjz+KrSa
saaSg7ZmBQyNdcPNJfhDnAp03j0wkN/ebbDAliy5ghWKbH8opjL/CuJ4mbIROOeQSrgAftk/AqWB
JKSdFHfLvi3ZpQt0kcDoWMAPPzK2PPnJbXXGjZ20+btfkIgvbsb1HmQboLhUve6JqtZXyXg30yrS
efipiPHv1T1a35BYkb8UTKHYtrZHw+uPXA1fhT6l3Ssh763w5O1g5yVObFmOohckaVVfqL7gZuya
TzLtkkQY19+2OqNYnq+Do3jF3PrHjwj1ZjfuFHKCReVTB9d25r+uomGcMeru2TIvjnl9CNEkaXfW
wgXeHFI6fbNAdc6hOfRRrgbcxbwOjwAGw6GwAONSYqCdiYJXIDVx3kYZyt6VS1dgerd+5opffsOO
kpEeIWF9F96W86JhzKXUhVt2nUAA+9ClarLk2IXPcv6PAMHpYFPd0IrDXLxT8uBviGh5On3+8aig
hp8XaGo26VzyyyJNDapg7dkZBB9hYuHMOTdhvI3jrMtPl5s0FWsFNYyYoZam2fW41EsQJRN9AgAh
WfTDF6fzvGYmtmH7/ZglYDRSgT1DtTyIBPy9BD3JWNEN+8eRrFN7b8rg9fiDO47HVRwIwDMpcZo/
+mf+3LJG2b/lEulqsPeGzKwN/H+E6dATzTx/0odk0obht7Emr2zrA+F5R5LzQ7gsHBKVYubm7Vxo
IU7ilJDlqiMaKDC81a+yVOSepygQ9edwAp40YaIJ+i9wHlsX3dp1nj/YLeYcInK42WVsywgsPGYe
4pSpBwBMubs0g+b2RQ06iSgkEZKZv59GZ4oigDE8UY5YAA/u+eksFbe6izSfh+hpSgGw+jsrUY6o
cTUM3i23UZ6tsUd1nOuLRbzAYe/dvZ5ZMCQBCCz6tQrkN6FiCmqqgZCftRGO16QihPbFVjVop8Wp
Ksh+DTdhovX5OC7q9+rFR82LytaGVRO4whfOFPs7YGvv2atmBlKjIfycjkPXCB9viI17Y+W/oc5L
BKd/N2qcJMwbKC2GpZ/5hRAAC+668FQjQxTJCfib6GGJzfaZXnDTYoFEYad8weH/7gq0an3MP43A
R0sWsVBXdlgjvAtQbcb9fq6JXaHGtQh3S1JWfmpE7SjYlHHDLW3sdlyzSUwFK0zmP/Sv14cmL1vX
0B+5nZquhp2sRqpccQcsewlkKhUkCgOydNkILJGGOu3ikDoNLzYd4eXjHX63YGzFL7EXn+YKgq20
DnU5xlrvzyh5uYE5kzTbAjW6xDBhyU2bN0vbkr7wGN5q7Aor3pkAZ2zmK2Yz7JgBEw9AIeUqEySC
9LZyNUB8LPmMCGSA/gqgL1HMgK9hUNNEI71QaxH5ASh277WJ/DubTjRah4YI2ScU6cIjV9YQTOrk
uQIFue0szB4oAvk4vY7ge5wiCxfFAEuxtt+CFIkTPozMa1FUkJcE+Qs+bqM98Gzjv6X899mQHyox
+uSeYkxvEE5pf32/y7KxEpfxV9xBD0cWJkhb8b7b/4b3wgD6YpIXYJ9A6NMSjlos/LF0EXwO0mKJ
eE3wOD4urXTJ9KnPrvFPxTyRMiBYQwX+gJZUOdTwJAI9BxF4pDmm0fUzYDIuCiIsg3X659tEdWXI
5i6ebOfSJaMjeAog0lT1W6MXmjc3qQ5c96WhVx79MkCBApp4Lm20wW4v2dri+eWu7jOUG0xx6OTA
O/z7+H6vPzUvAxxjK4V9KwpgyTaLZ754cFZZx7H4UPBYAJOlV2nWHmd2t08a+Mq+u/0eoz8yb0BP
6YWxoLG8TOKaqymmNWmG/DBl08puzxR4wCUDoSjzUIfluSO/ZKCmmcpiaTQMbQmfE7ateFgDRpRH
JVO6FVtHoI8JUuRq+kp6QVsnjuaZQSgg4k+HTnZ9BHM83+15x5/cG0sRfIHltevDuuLfQgINWopr
tvtCDO6IPpWVoEFNTHpaY2rzBHYlGfloYHO2yyMADNKiNP+geEXerxihm7h9tEQrV9VH8oBRdcfh
tCop3/me5elNSqnoSlTBbiWIEGfueHnC7uceqnjJ/mIbZq0kEBt3LfVbkrRD32k0MVs0Z6131+O3
jcX4FePqq0K+PTiqjZ7MNoScko79mTRJ81YekK5PBEiE0hWzymb9UrVsN96R28eHK61537skRErt
uJHaYVAxN6v7ohnlE9UoofdYnrJnq8KUPtJccJC99cwjJdlOrXHnW4EtCSeF2KvF87WKJsXHC6vZ
gFFhmRh78VXeiNf9sENvXdTaknN/ENMGihIiuqS4Tfp2UmaN7RmUybQDPjC/orfmMk1nfbIhnYAv
Z7YEj3bXQdVbMTkMeYDZJahItb1+tDF1iqjzXJEqTfGUQKd89bnDnkEsGpoL5Jt3LCXU/Rg/0Zbf
y9cuw74fw1Iju3nhG/dNYlrc8eR+6EWlWToFd9nP3OM6FtPX+JBlSc5ydKgXMQH64imRd4B6rqNL
UHRWqiqEJ2TjYY9ZOTXEm+0w2b3Keo9P4gsfv+4t9ZhEm2uVcYhDripCI/aoDC1NvREx0dTpseiK
zRqMl4N8s1NFqYJIBybHTsIs0QKrk7BCka2RZNU9/vFGupP32Oo9wkLM08CLM4edI3r8Gu2ZEM0y
+uCmE+8Mr8Dnhih8wMU3BWAGND5L8oyZfNrm6fGVPdPi3a8YsMqH4en+RPlR+RYZ0WZ2Ui2HNq3Z
ZCw0wx6Eb11RluCCk8Wd9/9JGXM7kvJQSxe/VTRnboYsuasjs0cfrbOpWCc7Lsgyfkme3HX+hoI3
lwSVprf5dNd6EZjtkLxm1aFZupG04n4g33C5dVPWKQvuQMOTqHTS5oeImAxR1jtm4Zm5muUhE9Hx
JjLuUR146KMsiULHikl0JrXojX4d9I+9NKLE++Hhx/8Sn/oMfEXVLXW3Sdvp08haBk94CsyKGjEs
rCFcebmrIuttXXtEvA6nwcVjJ3OYgBxhHLiCEIFdZcE9MUPn+sH5HFiL368mX6pQpyR4bE4BE/RW
gGlmNFbX8v6LmwbqKxSn/okZTsw7AwZnKT4I+DbQBpxNtFsx16D/iQXrGutWpTK7KX1qC0oLOFco
/+edW9cGKgbKvzVHnlYHHPVUdFPhdXr6J/bEPpnO6/WVvntKsFjPkhsfLxmHNh8S2vXCoaSFu/mj
kjt5V7BtdmJ5mogtCPZE3/egK1tSEopVkBSuvub/EQCV6XDiE34hI/EgwKeXJR9iAjS0N8ZvRJbn
g/nSLjO4XcLCftEKhPg985kNmgBDdyHOlCz5+DiUKZ/QY20yRcPSxzqk2QKA5DTb2IFv0X2pU1Wf
e41MBAPl4G4+tzcCwsSvscletTLmP2EdhmylKrhiYrXdQhU1BpOAZZe7mCPVAgN6uLj2r5wcPLUH
yTnnkTNvlrg1/NVgruFTwfOq7DQ6vFGnA0Kg71IauidUqO8a3UiBBEIAR3kRSooKyYgoty36O/Nm
bWnIFDi5orsFf5JqS98UukAkcEBsywa6jiDE0b5OUKduNYJitY9SuvQ8Ksmdl5UPq7Fw3seTGxA7
EMAIDnGxSLdvfreYbHM4UV71+4MrfwPehmUaUayCJIfQyvLYt9ODS3TQon+cu++jjEfSnyMVouE0
+7jTv3CXRAjP+Sd4KXx0mA+XPbfjC9chppze3nxU9zV/TwVkEJ9PENaR54mxRj3HGCcuRYyt+Cu0
RSWFmqQzq0C8YRo6mTunJyk/RGT6nlBCVkObclhheuYCLiaCruohEI98gow8TlKUJhgmQHrLEeu+
AA51NJ4pGs+g0yBxwORHDIfabX4NA2Vu4nwBVMxzM5DOEXgsO+472sEuAJ5ROK6rHVDvnelGlUFi
oSZKaybAk3eJZqArQgDbbAbnrL8FkuMgbul231RFuW6K8qBJx8wSQwc2wXXnCnXEvII7wtPZULsx
75dzzAx4kBArKVQdxKyrKMUqVRY4n/mA4DGcXGbjCGUkgNCd/bj1g19F1T3whHG/sBFuWB+rryO6
XQ4vbjZxOLnPdbuN39NXFjNG0EkPxx3IvutADgIcmDhquE8drzE+4WrAcomipVZ/z9oodG76ED6I
/NCfb2teVE0acIqXhZhH99P0hfh7q9zHHOF/SaCwSSwlIRBNhl3xZwnYB59g3TwkzljfGk1DrQAT
K8cRfyd82QUbhcd0OnwUj/nhmHhDqgY1zFMq451xjbF0ACrqQM7D+/PTmzCFYzY4LGrPM0ioR7ce
S51KhrtARnuIu8IGbAWAZxSqVa0gOMo1Roub+qnkMPFdrMRNwHdGuwOLQ5g4Zm8BckVlFFQYZ5qv
i/CujjOH5Oyv6zRBITer37AFAVUC6F7l6BqLv+ei1KrBJjFo+9v/cOcSLbf/hUqcLnyuhf3kFUYO
gc82PE3UQFD+xYRvxsetH4v3NqASpjSHoYGcdg/H7fq0OQmzNQRB9LluXwhuBf8u9oh59MqNUwo8
cp/TysE6GepUd2sCrdAILLkRprFlVufVPrzboPz7qKnGFIDoM3lkmKZe7gclqmQ7vtaUYIhbqcWa
u9snVbzu5UEKzbNcmslRHAIlgkHm8YGT+JeWF/3WmKRhKyx4z5ZHQrKPJeVZV4p3zpc+d6juMZDH
X3aK1iNyCUKaMUplLBu64qUxny0MJ/Km+toiIcpGg0Pi3MB0RWMNfc4fvTuTrhEJOBE4ZMX4RP4G
4xmAj9qgfGM/VSCn6IaEQrFhJTZHwJM190PzNuO97kJdml0Al7aHrvmMPvloYbF8z5xfgEXKnwhJ
7U6I9TRhCrnpOyFt01iGcPr2Y8VI/ohilN6UMYsrUW2WZKxuNRQc7xMEq0lS1bP0mpAI/uYsCqKJ
fxBlziZtn+fqUvAmSYv8iWJslozbgwmFEGjCzMDjJ3KSOetsKKaocsZOfq0/btshRaQ7kzFSli0p
oHXElnyp77DcNb6BVPIGoLjqF9qD2BU1UxOC0zn+80eIH7mvy4crTtFPqK5oZcwZ1gyPcjxv8pjQ
yrWm8KIinW96jeui8kUsQY9HtoYsSYDmqYz7RjlH44yuQY8QiGuWAsMPbPZSCwMx4BZAxYjl9wBb
33Ri7YVW34SAJaMIxFWq33mfQZ+tQfSQmnzmTMr/5RD7YPZXBKf6v5AaGZRYPeaGXI1B+ajWczaF
QZG9uLZbS/6fUEZh0jUZUDbkejiuPYy2Ip+BKYBzkUGWgO2LrDJDrtfJ2FHAoVAPYbhZC/uk53kW
EQMx4qKnkLinQg6/3HlAjxlgK5oHWR9c/VfPGnaDINX1maUjc4fEM+LE+L987mDeBkFMUv4TAgoX
tJfzoZTcYL3he+qNDZmFDgP4pte2hzB9qxgfepIjpjeQbj9oCC6aEskfQc+egZrwFgZjR75quSmf
KC/wuHvtrJkZ4g7Ol6tM1uY4LreM0/MbOdVw/dJCWc/Jhk5o7albgZesGHvbcvTKCQOCfFmKzd61
wRsYFQbMMb0UFEx+m09N58aR4qyGvApX6pF3yi94m4sCOtd34YlrH45+fd1ysf+HfvzSpg/HkZjs
4UEDqB5V4NoDrVvHNDwIxSOsZXQ2apCss2yZfQm2n1ziHPcHWSqjL6JzNSniLvD71o4DEWu6MYth
7wXhaWqZKAkfUbXV1AHZV3nMB8uch0VyHgOLFKwH6boMKlIUkBTudaHJvZUBtBQD0ZgnXOyQa5Q1
1Nh1V930enaw3RvTjh2rL0FTmfd2TekvEN0qmljfWmL/gGXI0oAWvJqBHh2ld6hnYMXtUEhnMptV
Q7Z6CgAbGSAeoZpMBuhnQr3zakmai3RUvNfZSA01r0nldfU7Xqftdv85WP4lZW+PAQ8v25W00+D4
nRTHulN8naqi/qvVrXQhgQOzzYBC0YhxeIVwLVOUtet/g/knpvvR2DKxU7zB0IAUmrPDzkS4IueR
dCer8SfhyGyObFwSF1v+cHZBU2Y7yKERxe5475cwHZahiD+D5lsX2R2juGRYalL69aQ3SeiEy2IT
b7g3sXzMG+4agLaW2D427KGA7ZkZG81g0OgZpc08rZuOhNWsFeKGknrbXFr2/STE1lj64Nn2W0Vk
LYbaLcuB19yvw5R+5UD2LePEPRgTgmMuhDuQ946xBwMxRMnkpLp1b5CE/es6AtkhnB1Qs58gCqqV
pouaL6PiO11hqjJO1raeF0rGTUkAlg8ULhOCDJcQFG6ENeRNfoygBgtjyHgJDVzNw3u1wl8tyaDp
etXnTUUWb8wT0tzp8X2ixzr7NS18HZmXquXlOK82evzFs+Miza4ZxPxRJK7GuoElbwud6f+P0hYk
phgYOknp3LaJaXrq6UMd6OnS5Ae0mZb0Ps/sVRKl7p6kvLTc23ePGq9neZUDDLhg/DlIAq8vNBzH
QHKVzb6StJT16TyAYi31F5PjV9pBtxsitvcNjRzg9mDEPn8fzc2AjaSfwjyWMezqiSlMKTnwARjk
kpqLZ5J3zWes2gE/WkL8YGpf/5zLsiiOQ+FuYh+IYaTlcDTdwb0MNL4NRYu8YtmlleXgfVJVkMAF
oTSIznSS1s2vC8d++xtFINNxYAWoN+YgjrH0C4lDlflLSo1HS3cOQKZerIZd+doXt5z5jxUr4rKC
z+tmpXJmw2WrCa+PALcuaC+8g5pmUUGLfIW9DeZ7VRMADXR+IdnpSQiaLLxrpSjiRQmAxzgLSH3I
awcam4+C7VyRGTk6gq6Jo98LuuhjV7D744QyJoqoVhE7FguncnCto9RwhxToqfoWddJITp/OB9xY
KVnF/HbqQECh+5RFwVk50lsYUlt5b+fUZfjptMYOjeLpX9Wpu/cW6bu6OmEaQhli/5nVrzOslNgq
2van11rwSc+s2cedBS2JRMfSH3rxa3WDbWzjzPgLBJmyqQU+7IUiVwQDmxm/ScdvyigrWhEiX/pL
QbZfIURqYLgjEkOpU9xms00IdZllu1s1Abs8Yz6W5cSgAtyTuOCb6mc9x2TTckKOVvTbCgr6PeIO
HguZt/m/Pkd18/ocUD5hUwMmlwUxlbdkz6IzyhbaPRye9JpRlkx+rKae2UeAR9vigwrQDaSd/AGB
z8vtjQt7Kkn+Gd9RUeIkZQKI9KMjt0pqS2de9VXB68dXtz7eS46F69xHt4XCedXZTq2ChtfxIaJP
Izgu+EDpiz051G3Y9459EyjF5WMPYCmczGaH9b8AGZPTcOdvsVyWYIh54IP3l3pCZ1nAkN7lqtEh
eZJ0HbAnz/ocDCJgYL0UjqZrukrPpmPLBx/0zaBUY3eIYMGW191fpJPpqOmuXpZLVLTQjqN2kDqO
88GHESLehxSD1ngTekq1XoZdOgy28lxzT2gYN8DyxG5EVHSbUgVN7KgnZujCCvqhCEMLUfZPmGzo
kqGd8f8oCsfhCESpY9DGTEGq06NRiNSbqU2mJtx2Cz95ug2zJV5LpzpYPbmxVgXE0WkM0N3Le7Ov
FNAAjO2ZbmPmSI/SE16pvx4FgY8Q1KK+Rg2iAWXKvfqenJmAFWS5eECFwgaFP7OiAraRhbfDKDWy
CbcDhgtWxhSPJow1NNgSM7FcuWj8ZYWDFqaszd/gvvhkouWyunfuP0jfku+f1pYtw/oUAu3nXF+h
h2xHkwj9bppKJIfzP1Jj7gLR5nr8rNOrMckIJa5b5YJ7sZOiTri5zIzVhfn96aJrZD7WNAuDXZto
GqBM8mk5O9TLfHSsufWW5pfyYiFqXZpxfLQM5XtDZp1C4sDXUVAycGCmGeJZttptLp5vJqk2wDeG
TNvDli3sxJ3KTtgxNCjoxbSyq2s5BF+eQX2RmefTZXdrFQOmdr2N/HmICNZoDrwIfk9pw8MwW4nn
9Dr7ltKN4b6+GIOpocMufdRS4CC9sY99W1TgV51BBydt8xbbdMbW7AjdLaFRcSLPu0mfvVxkmpXG
akUVEGKJXqwN8fuIQwoyTtBDSBScNs2vUL33SEC2zQNR9ZMMThW8DcBkPGU9WabJdkZ/7B70Eck/
Q6V7pJ3C+BZbgFy1X6qze1NX6i56Y98X3F+w9RGKo0xN/5+gspcwC1IewuiW2bDObwb0Ob9MjNVf
+zlkJVqPXaGuWU5IA5SUR+3XVAzngF9APmkLYeOhueqGuI7M6nuY21TsbsHzCjpYs6EDoIwyPLGN
aq5tbsq5IoIDqOFVAPmhpoitTZXEDhFmhDmi3DklE5FfFpTPAaTQ7Q7h3k/0knfGRF2cue6xxx66
m9h+pIquLckoOeHxk/dtzQLaKdTaQAKOJm1f3rl6tp9F54iVADkH3EV/jUMr1T5Zg1qbQx6lKiPR
yvCcFDBxMKUKyPBQqfQ3sGBdM3OO6nOW+/oQyMm+S2V/09xcfTXX/Sy/9W+1sf53HVIBT/nW4n3S
EMwPPllN0w0uod4a0KJPO/OlhTtV6rCt6fPDyTbXLMmqkyH20nLjZ81PodNn67RvzFe231R8OdBI
rj/MmBL6SQIPIABB7WxmNqYV6wYZiigUqYoOUG70lRGPc+oYJciuWg29vDcXrKg+2wXUY9XNkSUk
sK5pEkzJTSGRLEd+XYLJnRgpQq8VbvYoL+JfauLc8WVbeEb/SplFbyEu2FZ6YRNMNDfIjfrCiEyW
ZAjqypZQqifvvtp0ZAdOpjiCnBuAD3sUXF/L9lnvraR0rnnhxoH2ZNyWsFAy3+aKDaa6KQCe6Bye
QuB5O4/NERgaLlfo8vRICOUMkTQcEMy+qGV2RQyDe1ASpRMLPkrwGlNe9Yl90/lKnhQ1Aom4etn/
o9JW0vbVaaJxrWYco/3NNh+Skpbwr0SisW3oayopgZl3uJEJTqBk+RL9L64S6IEi/HyPQEjj1u+d
JIHmJkbdB+h7d2vQNtTScts9vKGkTfTrGdKPnT0yVBar43UGwTbCRaqNwG7SjXyokxcYcQ0Mh5f1
vZgGh/sIp4TOesv5R3uvdrjAkb4WruFlUrSOTc3cvsnpLJKULzZlPqBRIaARqjzMpLzSwvkz6h8t
Ju4LxeT5hW501bVSkas9xAGb22YJDDZHNSVxsQj6kFq8h0ZRlrO0ytv9sgug3xbhl9yfCD9uNtqO
A0HJGN5RoPmPcWUaTjDe5Fn+oYNkU8T91o2DP0fFwtr5dv+s88cnYy3iBPDKQjIQZsE3/UMVDLeW
YkbzJGnvRbzBq3Q4+h+MT3660j0Lb1hYjilOOQ2zZT9CV1MBuxFz4xUyjSQurColbOXYXx5lWjfP
yCX8zn9Y40SPPFE146R5t4U9UmKzSUQFCCElk1RADQkfeAWyD+6a5yl27w90JqtXq/ZOhdhruis5
NsHZ3ssJH97GY9+ZQF0g0Ee9kA/B8dw3UbEimazGK8rZzBw9IxTILzdB8HI3NWS6LyPyG7gCL7OB
G0vcyXr4RZUyiYk9hTRCGqyoXmbDlAiTC3eRK6AvZid2CuJ5OWLqsJMmL69rMcbBF8+voNYCRlY1
0s+M8w0KJvVnL1NuTxcgaBOLxYgWhJzt6lSQJDiQ7c3wXLdgnvhKLVeov8ykeqgLW7vOhOa62iHm
JBQVq/y4qjnitKFSwUJFGp6krHG5mpji6Ud3c3bP6A+D8uAHFe/LQiNDiHXGlxmU6rw4S4vUp/cp
rGt3Wx4waj7ge/f+5pus68JMckonEbWokLu45st9TjJOdYadCXdWIvGXp+W54RtMAqy5pkwxQ6VE
giKAKd6u+6dr3IyS16HiOcjNoesReuAPaeeu+nO/tqhELOEhLeN69LzsnBB1ecAYTMJ81oHIxAN9
4ORjNV/O2dYgZwMVuxpbjH6PWS1Dds6dt2JkO1E2vPop6UcncnUPBjVEWqrvkphGGKp52TMe87vi
7s0Edw+8TDL9hnTWWEGyF3eReT9uBvbiV5Z69byF2rrcBx5ywiNAVK6fcm410kxBLfmH+rMgfzbj
C5pHT34EqupmMpDzkZWloJxC3TssjcSqNFOWYhBe70oSgQFBbZzBJoejijTGplytSpfJUTsEvOev
L32YR+p7fM1/WhquraRntfCArCfDMBM00sB7ujM7GWraKFO8yqiSlO+KE/Iry0vWNRWnTGpbEXjE
Ghwd8WBU2FMashYc2RsiUCT1/vznUvqL//rJ7cd6AuJSYuc5dSf//9pRA7Q0/CM4ql10iolXnOmT
q/N1hE8+kTYlwdw4RsNs5anaQIzRWR9OZzV1+Qf6c5I1l+lTOaNq0jNntVdWTzt1g8xc6zdImkV8
ysS+AG8nHKn2wRsazooq/wlPcWVLuddtI+OQiF9L0DITcFDtLlxGh5vRg8tN+ysWLGFmO/2n7SDp
coUDO0sPH1G0VaDmoTEUwpwR5bkAfeVxMO6Cd8ehsWFQKsFhTlHQNiEAYeBjgDdjafkmIgUsq5/8
Lxuhj1mr0oREXnZfZtWME90pcJgKtHXZULQa+ovzEx/LVY6JdzUgdiN+1dN0F1WzxQiwsgnnVy6k
7HbwwH9juLwzhEeQhfr2ud9ufLg2v/SQ9QibO4plyGQdmBfr0DyBkTZouVfkPsouN7P1Wd+jRXQd
8ygnKXy0N+PGB2WJ8h2CgnXs3vxyefbuJ3innMOsvOdlz8o9mEB1fOiNF/1ZzVMUD7+W/K6RZT9S
DQ2lcnVP8Cd9j/0hSxW7Flxna90ekYUsCQjjWJ+14DDslyLXPBHEqUf563sz6ABl0cJlAXF7RQLM
jmfDYXsJleW8zBHToZzVakWHzhuvo1xR102EQpVLbxtNKdAOlFSBnBqAcwrr7JrXruVWEcjIaeK+
V+Xp79CaTK6dmrQtJyrlaFtOM+V/NWY8OqTK3wN8tSF1qtknCanDXbX038eEmVuUvm+9Am+GYW1L
YGvwpcea4MocCkxte4iULmeXGKbWGVi3tFJzWLLy438yvV5CPI87fsdz2Ds3TEipwgDEuANohQsb
gS8HJ3yn+DHSeVDhXXdW88gZRkFoTF67BpQ2SZVMfpdObGuCNkKzhlWmxqVWxRlDe1f9gsRjRKsf
+FU339hLqM98YX1bmeJuXClG7pvrtEt7IVgqLKrrDNyeXVf0ae3+61X5xcOnbpugDwveyJ85KZXH
vIXA+LD+mEx1gSmhnGNve3lUNrLjvDTf+z5XFOrmUW/oXRpa1i+tANJzKtpfCZ26VlyS7jmCNMF1
A07tC2KV1SnuXKpfkiTy3iMUcH9ed8tv4QUq0aN7XaSr1A/0McK0OV55ZvIvMolL3w/PKUoxrNXk
LOj+cLuTTmJmX40kBx4cWzrzbTW1hT+GUHiTbMVXBBb9HnPo4oj/Ht/2wTdDEK1+ZFUxOBBK8RKU
wDlax38HQuL89jV+P/6YDlSFhXwaQp1kaAs4aPdFzrbd3RekZUNLfMFM3Rha09fJVZTB/UcpTA2T
fk1QbUz98hbczNjx4FFNZabJ260B1wivTosKR3OPPy328pTHvB4yCTnXmyEeRm++DrwBELXGWdQ6
ubLFCKzVVjPVbVHZUiKRkqEm1NAZ7MjBct5tgrSZVHgEHllRmiFT4syqpVIeqW+LuLAa/Q78cyh5
9Q8CqQqwtvz+fY7VG6hdnoaYQ4Rg0A5NcA1LIQiiv4nrPPwgURjGm1BiU2OppwLuIEzT+PXbNsrp
XcafkVNlCU6j2tiXodOZHKkhePEmcqnlmC8dBAmVheI/FjZjAtF1jAo/ygTaRRA7IG/jN1OIpPlZ
ggpjsgmR+A91v56HSmY/h22Vv6ATRaQu5FJf7jLdFffyCmSTzR/nBW99iKGYPGVlMdAGf+LYcVPH
TNMEcZZCFdbdt3jhq3w1X/uQeI/qAY7JmMxKALsp6n6+A6vHsUR1GKdvD7jeznSklg/z/HhppH2S
JASV8KyhoHTwdVLko9ZBKCZduSdGKAWVXykid2JKW2h+Uuh5MYXoxZR5JXaFazq24wbfSUd8Zh6D
NoUCZ+nhCV9HB+JtodX4dgY2zrJ35kXCN6GhS+V/XGrrAglVfcHB20obQB2ncwXzzlL3gp97sqjN
aHE1N0w+nkQglOuvIJqT//BpkVEp3ehKwNRd0B8FMgJ+2Loa5w/Jum3HBKPlowtT4tyk7ZZywXh8
1suknBLqM39jxcnq16BndoDIPgP6cC6H6ILyeo4Yo5M8LWurqde1PDxa46RhpjPkmk6zD2i0Ih7+
wc/smJyIA3qBRHuX5VWrwZQZdDyy2phO51udk9EUTjUBjdnTUG0QqMiQZFI7bS4o4N+jTutVtv4o
Hh1/1Cy1uYyWvQNJ3Yrv5/72M1eXTYI+dK7nyDAV0One8XmmM1wKbSIrb+yzNIxlQBwbvhX2iN90
SSYrcx/hMkIEc3N7406evy3cAGvnDxAYuWTRG0wt0SSV3lzL2K4HbN0QhLy7WMawWfOjbMbYwyMu
6klogBwjc3cwy8+9iE6ShGzGRsaj3VdQ51MVDW/fXafpqhwSDCLtII99BmUjhMOv3edCvXT8V7a7
/DKhBwUUkaX1nYxAppDCtzKd8jyY2GMfQfVhAPduotRRw0dapU0pcyYdk9ltdbRHbHP+F92PV0+F
ZLpF8FsX02HzJuH+rg5H0NTREbqfZaMMX0dBQu1TUoMrTub85jYeMlV9N98mi9MDrHrTECpLfgaf
gU7LQy34/QibPs1bjX8wgBiMXT2lT0jmlrvaGc8LEemvanXTGoJlHzhC5oJwVtzyqMpQlITxI9ar
vhUPMM8XLgKA5VgXIFiJSVFLHbf76OpEX9/5CMRm1X7B1fLRfPEdrna5RSgkl3lVZo3Qsh2mfgBh
C2fT2LHoVCGAEKD8c2vidc9lUxT/MaCgo9TD2FifctfuN8d29W4+AhB7qpV9TG6BNxGA1jwqvz1J
fLTwOgMvWA4bnDzjxSnigNhIjJjwLNc32Bzb1FP/rcq1lxjydesDWgAjdVhlGQOtNtWXVpZS1chs
n219umIsgkzNcZxHNUyzjM6nVAXsYAraMbqR6aO1zjSHg6HTCUeTy7CBW6I7AzQvcyxpEcz2M6Sh
RZOcro9JF2dzfmA5XUxlto7+CY1E5nqDmTQxq6+ioqdMTlNC1IWOPAjw69aS92xD5tsGlVp3kAXS
uUPv5HhNNtQzWbpcuuM8Vt7euL4TEzkelOhcJqNnymg5OHze55fY8eALnOEpUIm/fFVy06wobEte
ulf6SWxk/s3HJ2Kuf0m53Xx3jous9glek4LcKpkD6OzTfpIg0hxBGRSo8yi6ZIn3O1V96l6Yntn/
XybIm6+Jz7mEW4rUteKRNNMLWly3IYoKhOWF6Yn/dkHU7U7JHn/WezA6MCTXpvAHYba8i6HEak3h
itW2YIO3GR6bfkJf6FmlvQ/sktj2o5jEusR3IQF+IhnNanG/HN/Ve11hAkBz5a706HriFiz0Xeit
waRzoOGkbovznVYGcYtAMt4ZkNvz/u7zdZCNpRVz4r0/GF7UMzlHPH228dY+0q1PjPzzmSOEhgrj
x8vFoOiB8xctq6XNzRnOzLNHX3jrun6FabtmDZ05rrZm3PhZdSlJ0d0xhA22g0ExKnkezCo6Tb7I
NQFLhogAMlSo/j/FOwkTjmCJ2I01Hq/c90rcZveeK1wyZ/LhZEAa1MCViNdRkFxXQFb3G3NXLHwA
9kqHCwq9uevJ4se2tOXgvck3bvemSrHLIDAGLdmaJ+2Vx8BefIkAgATrmVNp2gO0EdlhJUsbyczd
Omz7ndLBKwaSugpxdVsImdjq1CuLGGVU0mWRgx3jBLF2hEHZGzTrV+LwEmg3g2wtQN97ZjCk4NUn
E3EfVoPUr3UetH0Iy6QeXAt5/m2rgtfC9WxC5RG8muWxErAcJ7mOv62OyjH9zO/GyaOtqfGLbGAr
AKlYxCoQx73D6LsFAggIIqzDzuz3u/yvFXLD/evxWn+ebYljHmUwieYsZRkWucd07CInMPAK1JdY
+bQI1pZeSgMAmJ3QdBDt3PDvKaYKH3bNLfgsoWMKzNxjumZvIHWE+UFA6/JmtEwcVMtykhikZzV9
EWBJmQVbKtpTqfNPcKaYX73cESI6p6Qd6EJrYfhQcZGfWQearAtuf2/VIBj0SBeShUA1tqUT7k43
1OPbbyja5aexl+DRsPhFfCBtX8l9HLcJKypioiTszaIPoadFCaRz5FicgKdBra1JlVYGBrQlQx99
BaG/aI9CCt1sAw7sboymfUvRt4W/pFUTsjUjPuENiJHJXl87ytTmRomkoN/KE4yQukmg0S8oYutv
YVqQ8GKJRu1q81LtE3uWBlGpwRRlBCtmsV2tSl5fTlex3SOXveUOwTIXAaxrAwHaMM5tF8iLM9Fm
496jSYVjPIDOHUIA6yXrrwFLxjbqOQ/sJMqBS9218yuDlhlgM56s98DQehOZBYslzqotbJZyPsKj
GBlAnM78UHxhv3ufO4yBILHIjNoHD/LHkHKRNHx9/Krq6DdDAhSKcqBdbMQGFjfoMTjLgd2ykoF9
YWERkynNi4r453qhFfgGmGUW3yyYiLJgPglss6i/lxpiMjn2YmjitRLWFyYZN9P96jRSuTVGFijc
rzVXFAsutu1UAqx/2MtmxRaEPSqtMqzYo1JdDWepw0U1bR4DYWaipyBMdg7/e9xHUcXZ6e5m8JvW
nYkSB5XDFQlLQLLeA7S2eOX8+lMq9GrujZaUycmNhJTo2M58BCuDYqpRVURO4pEyxrQ4x7Zupswg
esUDD37Zn1p/a50GfHrZ9oqWBEOZ8qgn7a2P9RuGqLebsHy/mgJIrSor5qwujQQfC6v/ZL5tJY1M
rmmMNE0HMJbylulz0JFhp3L+JbuEN/fD7CMWNxAmv+Y+X4OJmR7zxQFQLl0wvP7YubbvSkXQCnqj
3SOkpvBBR/lJep8lZF58MQoqCE7r2T3L7Ef0Vei+aEr2406JLOqE8jCi+kQvLn6+hz4Z/Jce14of
JBuhZlGhWRexdZFJRlQCR4FOX5tNHrayHmY9bhOuwY08YvNH2b2311qoTBM2y1x+1/OduWtAIOK8
fduHbFFvfIggGEonFIC5R/s0+cudJSsS4i2NDIS15aUv0s1kFEZba3U7AZGAV/gtdPqQs5r6tMly
DuXKlHN5d9Kp3+op+jx574Ygu/wI1ZSfHtuYuVdhCle7HWJYXcl3i4EctZboxPHjKubUcn7qo7K9
4FmCNQ9zxiQgYw7K33Ngdbhbv75Frtegm9SVLP9bdr9YBlHVP1K7EjpXLW7ZV9d3vrbjyu64MJ5R
Nr1OpoCIjxlQWd00NUzJ4qzpUOdfjDF/3COQyc/doA/V0FuvvGRwJOeVxwwaUKRYVW7zGa6GeQFW
ebquVKeZugGUuy+GAJV6DGPPIO7SKSeQ+V5ZQi92zrQfw5uRNDcD6MtH13w3f2YCUITaO2PGEN6I
jawH6ujVM9ryR5jdGS6h3HNTsK7Haxa3uQuSYWDwwk+3YuUcVxJTxBaOi9ygX4l1MrtCXMQjNbCO
lUMiu5HKBSGmQAikLur3z8dFt3uPCNtkpjYg/wUqQa9PyaKQTjPA9pTCNVrRZiEHeGQgZL/A8mBx
Mw2jIQ8PYiU0fGV2XFhtEFtDgCYQpucVI1MMWrDWRe1jYLd24TRuRe1hBvNHX8QCucgok56k39og
3Ws9fnLOFWyXvUEa37SsPw+xTnV/ARyc/DOokj73ymNXkdktGpRWc/qU1uPcy8oc1TYHVeiWcHGc
/Cnes45q+mIUhoLJjdYwnSUKgWScDCkX76eHUr6WubbJoPBOh0WHxXSeC+PAVEYym5h3x/tb5zKn
1SrOtJrheLbREj/4U358+NneFDHciirhlKfUAh9tSVnk6OmljWSq8NT/4nBETAz+6aKjgFQ5N/9I
Ln6Kp1tCxEi3TLX4AYRygN8uwggNaopYHUI1Wi0jQnBwH7kiUM/hU3TxUo3i1aNNEdeJGzRxk8IK
Cuad5QkxEoeTV5yn6EZT9Wwxsbb1BethmmqU0PknUM8kYRzdOlpPeRbO7biCH1X4xr7IVyne+Ujs
0hbteQMOVHreGPaz8TkgBcEtRbBj99m1U/egV4UB7M5DpJAZxX7+sx42rqIRr7aJ002A5Xa6OH+O
uCWO5sxOT7VeCaK6g0DYakullJqImm+KKUkAR4E5dUZ8OruOwC+6GKlhtI6/1n/rKxWddVNk8Iha
iowkEM7KTo0N2rhk6c47d0xeZQvIj59QQAIDUq9e8/893AZ6hCetk37LU7gaO9l6v3B+5J0BVDxD
FsJDX0nz/H5tL14qCQgxW/dcTLwgYHdDejGlOYcMQnRwRsusTElI93ZRbbsgTVEgXGQTF/9f1gpA
zonVMcJB/1ac3MUH8Q3I5xx2WeTd+aPiRVXhu/nfm+bfRdFArMoqEMhmtASmbRGmJGt/uuGXwOYY
SR3lkCmbMThRQrmwIpJ20HrSxCY3/X985CYc5JFyCYxuORNgkEIFTPMafuGp3aAmJ8HR3NGgz18y
nOKLkIaShXnJUzmjV9O+wPkCvk/ygoGWGmeFmV0FjJCf7/iS8/zhoXs3fScouagsj9w9YXWpxV1y
VFECDzNu1iqh1xAPnKUqXhwyvNFQ4zhSYDGJB5l95wyWAW44BaiTdUyzuPdua/rSSKetOnxfdaLN
ADNEzSFuQNppK5WXlePEdtTGxZzfdZLm2PgBv0PLzJIt/axFPoJR2tnHXw4f7ENoPGCtveg3N+KI
RKvz12PERvD1lACBgtqGQC/wAzcz+kl7mkr1RoF/gdXMwdX3pGxi2Hc+XXiWEKhxYUzptmw1YQso
ojXvmZGa1hNw7laUqWTE9aQdRqx8XWh3d+3vRPrNuycLZl/GeDQjEehhw+GLfaqWIWqqLXeM5389
zBDJS9vXY9+RpIBNJpCjZupREgYclenremhQCFjkL5jc8ifj0AbvsgRenKlIntKawsihS0roaN7N
OvIB6D5gOAURWdZ48I5ntBZB/9MTT58aRrvafKJPOw7sCF5QfLWPg4hgHELsqqwbL8jcaxoVWTsb
BmBy9dt74/5j0Ja/ZxVFHNSI2VEIbHkwVH/CFlIcF33FQ07BEPAuYkVZXkLYHLhCs2hAhC+wMQ6I
lK/s1lKXRqWH5PrBG/vxMYIqj2ottJr6v0IjsS7yue3YC48fEv90HoPNuZiMMeFdC2EYt1jkxSVC
L5tP9sUrYuWWNRsV2TSZYRfNVByblmRQCvixqgqYDekvD/cfN507N12JMgPeudqpczkOMuW+pqWT
Zafgvq75Ljnk+fkRaoHr8OInGnSTSNfrYjGlfpTbAnL3nHeaZWpVecHzAKCtnKAoq01n7Ei1cDx5
OSfYGr6Dx2TCCy7vpNVIIBPmDR9d+hq7Pcrf+ite/HCSgPWfLF8xY0BN7RrVQNdf2PehNCPjpxMW
DSmh+M9hTx67EeLNvZIzplcuEz8zQDbJt6sl5AK5eM/kOOtYDgIJaFR+LitG9lMleVV5vq1agt6J
L2Gd8ggXbPEvM8h76bJ4CNm0sEk8f6QMCNwwTLQSh+lHExhwqquP8O7xZQypLKKwprUlevbw76R1
alAqlEBMcb6aBbSemMD3igf+7NMYB+mNiPO7glMaFmAJiVE6TCXpDxcgCrKhUrbaDKfxz745adoE
KWPDMZSEuIq3S05wYFsggyRMoQ72R1oyb2B0L6GgO5CavWSyBig/vWTddYV3yWZdzW8Itt+AqBD5
Nh7du/UYzQbnUAPGQ2AH83I5xyMQjgsulic3yMuTL4R4rlzHcNeFm0fU3jaMoCCMx7pZ0x6icoee
2DgonikQTOPZwOEKHEQvcbMZMG38B5JhrxRCqDrLPbgr7lzrMJfyw/HRaOMxi5EuSp+f8H5qqwSY
UNf8c3Etp7ifktGFaQKTsXcmAhF3A3XOHRE5jQjaqREPasWGURUfVY8s8jmj6mbt3dGWsNMXc37y
bcYlSfNmrcNSrrgcD8kEZI5rBKrmYhnj0hwvq865Uyx9L13BTecyA4N+v3doEV6ZihpEhf+nL+9p
wcleL7gPX964pstTCNVyMGWED/90/QCbVfQ3N9ZL8fPxoRIwFvhcN2pxRKz9iXDewNEVkgYUPKSI
IO6R97vS5C9cwvSy+ItWdD4xgdgGimsUoNL4bhpKq2FZLZXI+CF+aZvpf7cQOuRuxRDYw131taYV
jBZrSG6S/J5zHS2iw6VcET62AVkQFVMZ7lMxFckN/gloaG3tf5by6dXEcPUoTBQDv0FBG9Mq9sjL
A34/a8FGw7g/dKKhutgFI7KzJ1T2T98kV8Sjem6wbZ36vK3uPxCLE3tmvYVCN3awR3ojCa5J16dF
HfCiJAy7nnMKmECrGjzGB53R08Ahi8cXny3CKuYldamTMyfxVvwxX4T4j9QJyr6lyHWNRPFHZDog
GAIw0SueDipeup+r/iBAE+wNRusne5rQTJxn51Vh3UBJ9Y6hH3HWMDTnEHMTWmLS7Jds9p99eFSR
P2Ak3tvvX4mrZdLJM0tbx2uFlN8DKgTXE1fR5PRwVbV12bvQq6ifoP86TPthP+1LpnfjM7esTdfN
7EajJ9h6XubC0PUEbViiVVm8VUsBzddrBsWjPFnqsF8MCbwZXQ9/XCd79pwryemAd9GIbPnBvliG
8fk6rJ9EKQZZSbftPdpXy2P5tnc0rDeDx142ovcJbfsgoGTm0pzX0lQN8N8GSxVMhg9SuDygi4h2
TLns6xWI96CuGQaYl6SUFF0Gf05QlQ7wiHrwi4HgFI6dvAEgbkjZ3GSxX6B3ZeTTt36O+bfU9bxa
jTiiyLvj0uBdrdyi9RKcoQlZ6iL90Odr6wB3SVcY+lJIeG7HLjNQrAlskVOpFdT3xx9L4BXKIkQ/
8+6USBiKST2yA+ozif5B4lA9XmVxP8OX43cttaBs9UvImzrnOlw2PLqeNGzJRdXNornOs9GxvUPY
L2xoG88V9KXmXJwhfIx225vHd+qyzsJ8NiTBqHEK4/nyfGQkGIUwi1WK3GzegnvryLGei5+Pimuk
qPRrMQS8fwG3a3abfYhuXBWCBR0TYwMUjfXzJH2smFMzWKI1B3lWJTYh/GalR+hn9+XpCXYjaJax
WoW1qkAjYQFT6wtNfITAyiaU/qkwQTasQTvJWuEFbKHzq7shNZin49ildBr7QQA2+YETDs7dOvIV
3wq9a76BYYCLRQAepeONx/v+oaN7jx6hI+nCXWlIaTcD8PLyiYH2knf+LgTz9t1y2k7UPOWMV2e2
BnCgQ19eq9ukrx4/r1lShZm5yf6fe4Fo5z5Ya2plXffRP75ZENr16RkRzjeCcju6O5vGKLmUZJRE
mhYPYg5ZACKzf8A2/bXRxQXTAqZ0OCoPGDzHsFqfvyfCLVv3H3i3mhwPUApjcqW03CzKtXijEr/p
7rCFQe69JxvJGkNaJtdUShe6uYh99dSvCDIVq5XuhF6nEDkUmK9oku8oon0TthNNIDBTYvVNYX2O
r/C3CNltdJh0Pk9dLhrKz9BT5vqV5xwomT1wfzdc/mOWYZVMI3aKEBj1Kef0+SggAekAd+6Js1kR
3rejuPhJL8vxdgk/b/MigwLm14G/63b8THz8hFGOWX58j2I+LkXxePFFeW98Oqoz1YsOTbBkY4YS
QXXn4baDzVfnh8cs5B43kI8h8JsM43LLDJ2a/ZolI6cpGrwBhOi8QkVcNi9DqNNXQcKSWZetGAhN
HgUMdhjSyKhQwJVzH0SV4IHpAoy8p917+iEABffldeoL0zHh0Lye5xIJT2vBAIYqq21SxNekRSwl
v8vf6sWw9Vq+ntJB9XVu2vpeU6PAmRUEiTzeDWswxVXDejRY/3aN6MmwXZVTWIxEadEyqpj2OAXU
uLMGVHLdr7+jYAokcova9jHf6k/844ZFOorMHZ+oKtIkio6mXVB7PlsRqUO3fh9ISmYVpCqaNqvn
5EaXNpYMeMuEqI1sCAhdZ/MtUdjbnkRRg1IQMBasDT5o+f7saVkYYXZtUhSNIz0ztv/g3G8xAhkC
FzyeFmUyQW1sSLYdTRnmcXTzy0OOlgy6QDT8xwWc18L5MOHdqGOnZ4F1AMIFHxz2a58GEtuhNQns
Fo2i3ObkTr44ZgZdoBR5COUu3yceEFktnP25jE0YPT4hxhFd9Ij85JtUXIRQPxZZKAefLSkKCzGo
gmflTRtL8iBm4tdKZlR8gJYjxo6Sys63ES8yzscxK4UBQIni5a/uAoXr/Vvr4PEcza00/KZa/sZL
qfs8POKT2yKWWEXbCo+KdQDN4q3g9tvKFKJfTRddX8r9Qkh2llFWYelfKLtuJVgWzTNmN1qWUHq5
C1y5wlKyDJaD1Sk7yG3L873HkTrDdncmq6x9cBCUBfqGUIJ5Ut0Zn7T99fAR3/TvcnZ5n8nhFoGD
RDUfvnpU+9J3wKBb42DfeTU/wEQmrkR5ZoM5RAFRQSm/ZM3ha42qWcdFxJZDmangACmvZ7/uAMMm
eypiQ6GOVicDx4lqA4g1vDch7ZIke/V5Q1pdanJPWxKD6jJHTyIxTgd8um0wckx/l04pN2ItX0oT
QrC2HCZdWn+ZXIoy6L3gzbyDhegKJTbhYdHM0n0BAqsfrldlZMoZY+ZdPVJeZy/q4cMClh618Raw
VDO5v3ma3KgN2kjRKW/Aw268mVLaLgd1v5SA2pTMIdG3qUb5lGfiqb/p0mqv1Ejj9+BjBYMDjWKk
uqCRDMeKzT271EvZkugqj627SWjtBLtgREr1v3vet2UObZmB/z+AW3X55acNqgwN5ICUeZ5N2cjP
maWAc/W4Muf71lUORJnCe4BDg5A4hkzzsOZK4Fp+VEa/8JMXXivSbYZ7IL3MuEZYSv6GTMphJOEz
/Z3TDZRF35xB7C9uxRGPnvJYaYZOEnFcFUiOPbZvXp8CcSsM3/FEuoSwvtQaWloGDIxlF+Uu5aTN
fm0JKEFPLLfvrcZx4jiAsLLZLCCUgLTblkF4tV64ydyV94qRR25FQk/8nvYkrbjTmBYAAQZHmym0
dkOTDXdI5PpzHCWtIJOWMgBe1VdRbOzui5eTngsHP+R0JL5spONbf628lUAdX0qMU0+qTULSHLcc
asGsReDetT4dm0wq/9N3v7x9u+5J3kw9nzknV5LV8HpgIby9qZhpMros0LvAx7T2rwia1AtSiIOa
iz4XPJty7ExVjrd6CV8rjXmUfkTkm83H72saNvatNXoE4GqCpI0w/Xasw4p+jJJYT342tQck4RdO
Sw0TqaZML0CN4J2p949lhRrC5AWnnjtcffX+/yCjThujrRCyjfNUzMoTyglQYUwOawuFMWRuE0O1
BPr9xx9hJx4OCC+/keg7QlJAy9BSfTAhVR15TZrJt9B5lLxznUsuR1kpiQqWqdKzh4YSMPE1L5fp
82uHL31joNnHYhre0zd/W63GR/3Lhbt2aR5z6C7HC+b9QwBKERpPEHIQNnz+7apznEkcQXGTLaqo
HCkN5CzI2GCZV0G3IpCk7NZ8TFTWOgiOKnx5UNlTpWt8lCpAlPgYdLI1VGqADa1npBRY6wLAKJjR
BhlMIKyet+lmjAqqhdV9L46Y1oP7UDU/d7QqPEWL0w2L9vv2XBLj99sw006AoX1LUAhOgip7NpM8
LhpEMRpWtXO//ZFsWX8x/UVqUduRDckrZDY8d9l3zF7ecZFtAJ0c0Gd2A+DbFuiHepc6t8XD1x+S
5GKdDqq5nbDxboW1VmP3dosGdncNwCjecU3teGAfKE3gyYzZgKol9tIrl3Qv+beD0teEUa9puNff
t+tn7d+4acYImEaapNvPsqDf3jNU58izp7P1cun/xm3IgLnSv7Rr39EPmWtz0vd1AqOO83lNykVH
kUeUYY5xf2+1ycboBITPX6ABh0esuwFhf01APL+NSHwPjVQd0VIl24ecTxXj8nJDbeB3Fr+VVR6V
1GoAMkJVXZoaQetfQhcID1yK+Q//J171Rm6SoFVZHxTJxdJRgG46r23Whk4lkNFc20KggxL55mnD
8XpO99kALKe00Z4L59+bUUs0mUlldDtiZ+nTNjSkn1gZJ2AlOPRCqInI+oU7T2GPmeSvsF5aRlPT
FouKywInQAbJwqv1hnrFGripD/bjds9W8qU/lFFQcjH7MlmUm8k1ldc713vbgO5sOGQVDA39QUrB
rlIp+K9tkbUa66+UN14F9UdLP6xhuFWyzB8a5/VYXjaBLFMOy73DCxjMzMAS86VNc4AWkuWyIG2r
soqE5C0w1a8iUfz4JMm7r5AInskP4BU9B45N1Lh47btZKBcZMnqESteXGJdmSYMPa59hf+9bsTVV
f8szL6IvzOXStGmgD9bhI7cnNowr7OkeOefL22y/vfD0Z8iN2qEj6TBVFLduwsNCeOTywOUKIfxJ
IKhlSO7X/rcoKIXSIUCmGzyGrOl1j+JR45xjkIDJY6TkL0Z/aO2/TWw9mVKSWKEd4D5RjuCmM1BZ
D0QTXPy2eENxDz4FZv+3NNyhz1Wwq35nw6YOZ38km5w/duuzX9fKTCMRyOx7I/fLFODr8KjTNtCi
Lh6T9sbstXIFklJ2hxDwzrMmpH0JWukOdDYEKzJswV5SGLMDVoO8FDLvgyGACLuCQErHEiaKyaQm
9yQFEgr8n7ArJj+KPu6DP+9gqI9jwllRiKQ9Qg0myMAJ0xw4W/HkU4igDgu+Zp6v7BM7lcAFiy4X
YjvwYqAerC35oDOfL0ZCzT9JsdNkELefHz/WiM+tGXS/wfVpiqhFaalQqRvwrJVofighnBr74/xF
+f3ISnKlRJ6/hXKEPYpuqdfDZdCT5KjT4N5pOYKL9JFoHG2Lc7g3X6s/SkuZDdoFIfRicSlQa30v
zpkpJfFQA0920nxZl/MgqLNw2jbpE1JviT5NAb8KFck5nDgRQJMr75Gy6QwbFMroRvD1VztU6q+/
z23Yfi78k6xXUDm4D6UI8uyGbI4pjRqILuZGGPqVRIYE05Umf0AvTJRcOjT6QhzaCRfq1o6YLLpI
QCfPD85PCNzD6uSxSoN3WTDpi5/nlEtESCg0SihE6CEjvBLtyz8afjYxIAhJQDezAPztwAcuZ7yL
dj9f5Tid23D4u3pr0yLSDNawxvs+0oMQQv0Dnq5bLVv0iGIbu12j0w6xlGlHASgjTRi4osdBGu0L
1NiwnIf9FGVebEOEHTgQZ7y+xjbNK7ZODRWXSXWIL/lD6qNGz6r0t0V1hu4Rpct6CyVqWbyv2SzJ
1s7NjDm6yF8UgCa74K58Wde7kiqLcjrsWXK+kxWy8kkwhuEbKpzvG8afhjKnggm/2BkvW6RcNG09
YipITNIgbSPvMqX9/apJU/qsOouKJv2ztcedtAmOi6nwniuy52+/JhLSO53HJUjf0yyRYe2LM2gT
r2wgHcq4pTAJIB8JoCu+YQs4TRtTl9xtaUmN/UnDJObFLhOGGioCDl4pkl3UifpaSu1LmEQPeEp6
6xk8QCsUwNc44OYGYuZ0a8YbBT0saCG85lDD0Lab6iQRJEM7jedCBUnOyODdUrluHs4PmAnLA9KY
ZLodvh0GqENyBjLSQ1eECQdl2vV6wyckb5G63SGcxalDsXCGLq2voEdmKyxeU+yeAC95wesom6Tw
vRxrgLPOvZDfXoHyHniM+wYCslUpnoZqEK7nCYm+tVylygsu/J1sTkyKRbhsr4niAi2SvMouGCz9
+pS7VAC9RqlG0BoHSbjEQ2vs2gwpKpJpV70xo/vS5g8E9mmGH3YP+SyvqRNv16eg3h1ClakK7eVd
lCsckVf2smy8gKfHmQUT8e+F1YswoAsGgN2PzrfGgHmLmY+50IDHDNB/3U/V2Jc7aaZso9tlBgeK
ppTApKqvmKg3DNRteW3I4bZOSXymKNa4tLrImn7AC6keSOpe4502V8dkAyuoi8fh3YUjNgavQxBw
rvi3e25504aZGc/6vjrStYd6l1/JaDPf0bQ0Qi/4i5HxROf7JEzZG5Y/TK5si8Z/ol21NDSA1aQc
YApVjB3F2eV5W/9RLJMBwX0o1QBPsifF69DJ3swjhpA4eaHnKT73V2s0fHNZd15tPFXDwKc3pvfk
rtbPX6YfhC+WnIG0Hu7yRuOHhBu7VpBzTfvCzsKYswqbMTZBVbmlPMqC+id45k7ZAXYxvmf6qXYm
HHfUp7fgg4rPCXkOZ4Vk49PepUzqTl6CqhwO0ve0UxpGguKrvNZCQ7ZqMlDc5E7rNsLwebTUGnwo
EuhsN41cF05ujWFqrmnu03cT9ekRylfG7mxB10JYLxa3n1EEBVRNboSl91m+Dj5nNN8bsfHRHTzu
Z7nSRCVBJCNDZ5JsttbjUNkSM8V4wNLps549D2gOxxYkfs8OjkCQOv14DaV6FmT18WMdfGK5smUD
AseFPlAW8rhE9N/IZ+fdnQwjPbAcwrBMcCfc3feRaRu3ljjmmyqdTwhPLXn4gECjqunOqVwfRuw5
S/XctxJAERreuAuWMZQgkvUI1regU38swFukx3r32JJKR3dHJ9Uh4uO9tAj46e+vTEeI29CmahFL
UHZWyHySUO7tpaUm9BTXhqYtkBxmDYLg4xEhatjVrl4Um6PkjSNGCwTKX9z6SIihrB4E67zyjifB
P8GLJZ9z1bMKz1B5HZ+625pA+MeQAHfJscF+hDWW8QuZq6l+e5cuyUBtDZu9dgzwXQBQoPXfomvH
4ckuH9wNHfvvpg9XwCy6W9gk59qGGvSrG0EMEXTfCmFI2W3jwSP/GZQDmxqNsbEG5o/KLLbFE8WK
5KVMQ3EKqCaOtY952mUWEgn4ataJpD6Y0xebYLc8z+uPHSuJ/WTZtrYW01GEOiQX2yxpjA/P/mEV
bzCbbvpcUAatRrL8z9jaAPgi2b39bOAtxIhdNDpJor3VpBJzPMLqyrh3Rj8DQZ6+EVx2e7kWGbIG
JRxu44GwZ0MwwN/dRnvLIUhp5HeUdK7LSv4U4le6i7/9NUJ7Wl7d+RIJuQnICFk3Ko3m1HAJE703
AZiWkAS9Qpm474xOk0KzxTbQ5JgBxyL5seDlW7WGWe8s1K59gQHwh4HzUDat+1yQ2VAjX1gVRJi3
lhrhVbVHdha4k7WvnsG9KVRkZusxWhJnZbItrOiY339g1PAICzqSH5YhhqvuuEtSN+ilZMRcQL0v
kyw+RvVw8lTz1p3s+EoH0Kgrmbv8/+p3w+xDHJ6eGePYqG31QIwB6vcortHp03QETmOPzcsjldGf
nJc5ONDhsvNWDiVT+hLi12qKcwd9BCMs7yuHAKsK8y+A7s5YqAz1wArbJsmMgu0flLwngsix8DWV
pokdzQMyUZqaolOsqsh7pS3AIG4TRVfYs8/npaYHyyP8HEAqdAa63F8PDRsO3C1YClLr0CvbzTRq
xx/aHjafaVUZ9KHzLqwAILjAx5uBoCvqHgbbErxJ8y+cd7u5tti8rhrmdArgOx/91BqvgFBs7JNw
AQH1oDITOVMvJLMtNIZ/vUh1LvhKzv++DY7vHZtDpxnXE30UxO8X2UbWSnEbSaC+npK7j2CCGA9d
O/EfFDwsQELy+rrbgomhULrnkSTl11BchSeBlOzaXBoFNrJepF8by9AVk2X3l9PpSXyC9K8r0wvz
adfjtXnnt068cxlDHEorUqo1KLcGCRPk+xKrdyT/RkmylVuJ/Zxc3z+URez4G8d0Nd0w67zHeDnh
lw3/lBZDnavZgROccx1B7e3QuYzn9yvGqYO+1299i9OA7tfrHrUPqrWUFaazQjFd99EB0fdlaBvS
c3HVKjcB76cccLZN0YUWMvUnT8siH7lep1+jv+Ar1QMzkQRo3HvoKZgTBIXjBsAVixyfr48v0s7l
J5t5pMT2F3PuqdueEXCR/nN9ND+scvnUnFSbZQuVGZevRKD4ty5Cp2oHc3GmWRSDaFd4szbU+wJk
x9uI/XSmsIlkSGDfj9kwUxS3KFTSnVX0N7OwS4CfvvJl0LAllX9Kqr4CmFn1lZnLhKB0DaPhhVGY
wegL8dIZSnyeO20YOEgjjdzxP1WWrtDl0IhzIGlYcmuKqrSod+T7JmwPdxKNK6Zigb/HGbdsarcx
ZMAd4hf0til3VTEQc7rv4Vy42VtHSy0DwA+OhYBFhqADUHkGzyKRY+uqExXyuAxhQ/Y4ivrTO/BX
edn/mFc1AmboulDAeaJEj0+ItF7deBGGj71LliWKj/PtN0mB8gju4AaLfbZCxv0pnyuuDSz/bGbx
Q4s1rdMxpheP4BR1pmtC97jcqYGHkZOG/1gcbN0SGM4TT5yabSwF5qcybn8v3ntTvEv94BRWOi/j
OS60iBga1xE6vzPCU9dLE+MIWSQxUzpJropi7DX2AyIW+bnjaEuXA+jzTXjBxSTaQFFvpv1w5ueA
Zwbw8eLiej8zfxFuL1iVqjrI4peMyYBKkhp03ufVa34wuXexj5wt6Kf02F83YCoNw6ZzOymSlzaU
uCLK8ElKmFOgZbwMZuTLdIWDxmiEB4z/crFaXbaLX+i/Kl4B/gaJs+fo1yGh1ZY3SrzAFAoMVHvJ
40CM+HqG0XqYUksFa9TyEyHesJB28MK5W6cG+tiFjW819jqshr6MW0tXXI/YvnZrVr69wHwU6sCz
P7hIUxI+oPiVVAHjwpyIlWQWiq0XXFxAYiiC5YcVFBaphC+hFBsfer1YfCSimIFkGrUKRzHa0Lpl
jNQYcX7f2ARQE6KYL7sNvhNiXQDn7DHrtLY8bMSkDi4A2dE3+qEm5KyKVUpFYZUXwWnlHfOswLc1
V7RidCT6k8fuapSa1vFZQYxekAHTmMDvSATJpBdEi52I0nIuW8ttxzaXxVPQRJMwbqhl7HEFfbXb
2VIzWMTthRRm0xuepwb/nE4yemT6geJbulkGrQJM3k3HIlAmkgJFk0UTkhiphPVchnXvrUdo3Eq+
MkkVq5U2d6NAN2B73EGF0CAoyw6pBoVDUiVU5qie0bzdNlzlPtcXeSIwl338L3LaYrE0sNBfHZVo
04Rm5huD8kHtxqihH6s2ougkfzeqGswh03PAXyGkuaXKircEVU7biHA2+W8HbxbZ2qfJs4SJtU5Y
MRnK5DoUt7Ywosfty9PPLwtWH8RJkoo4KjQErdi2YZ+NLXYwXe0o+3KV6Qf06ODWNrAcDQJMlKR1
MeYjv58onbZx2jpEzxCl1BMlox6mp0yWOsf84fdzz2hFKboFWF9oONI/3Yg04LKrnqbuNX0DjIQq
qK6EQXHhNgga7zIfhpwqYMUD9nrVfYgOR6VZxG/blBAnRf4BnGGJrpnamUWvten7vGG/5/CMUv5Z
Um2aGgyB3QgZAe3GKITqJKQIuYaO/wMiBiaXNstXJYnKTD1q+ok2CQG1/i2DkrJP0wz5qHz6JNCB
S30GTod1j+d2EchGt958ezIbPvY8v2pHIy7v0XI2igOQsmD9we5KlMWHDbfJ2iCsFJpASVs+hE3T
SC16/Do9cNjGGedBGOkB0uyqNZdkzbsrdySTEzbLhzC2cN+IXExeazdUdphB7cND6KECS4Q2rS01
/2l5YyjSyZ8Ko2HtDspiCXUpqlpKFeD/oA4j5mVI8qZ50rs0ZeECTZwHVvgNZ4DGDPzPWWdtgFyt
TgjW4iYbjtMD1vnaYBVxA++4hTpzuBEhPF2dcp70kVuSaqu/oKKrmOi8tKy8HedBhCCWF9rPeBck
eLumIlWLRQ/Ziigw3JSZ9Ijl+RIIcJMkCnmqMNAG4hPlygP5aNRtf6P6qfVwQ1jyxliSfjHYWaUs
otHXh/dg/VdpvLHw65v5Gl4IkTAlLiI9qO6sUh90BJCQvJvAtcKJi6fYinirDbMfNFAHa3GL13kP
R90EeG6eAi8QQ2dDO1ZX5QKRFBotNbU/OP9NnocJV9WOX24LKBgPM4+enaxReq8uFvDl5PkYWz4f
IzWUeCh9uhvmtpgRE2iGHRVhfVcco7xyBAYkHAsEn0/Y2jugUNUrTsAH9gIv+GKiOpQu5MF6at/j
Mpq+kxDLEy4lwpGUhQtL6VTBMGeXE3lr6blulGXXjQ4FfcaAX/pZc4hss89dGJ7vthyuR5QPNsY2
pGqhaaUCfwDXM6Duuh5KwvnjoQZuHJqjARs5w1PWZcMvKX5Biz73uX7bZZi2vbI3Ff/9L79cx5I7
TDwG3WX7huTc3+zzIYH1/EYLBejFdYYUsfmojankIc1NGXSCtIi9blCmAfd4IydSLE1Lcd3+Y6BP
npudCYGWOFOob6QtGVXzOPynVpCpA1E4Vj+Emo6T/DFQYYGP2blXUVkGaxZJdgf8WTE4BQ9wwWzt
ISQKnThf7K9qV3ndHckBSbdpLNQvH8wGGBl+XGuU4oin98fvOCzbMlfIn2zSonM0Y2Tc9yArUTQa
GTrZkMyHqoVCwHbam6nRcTRrdF3tWVk+yABLm4621YmMQhCFs2U72PJ/jy4wI9o1nVZs66mtNMFA
YAxkORzxDw4BzMRel/jeWY2c3woYJraM7d4QJSKA6vg3EhYhOkkcdIHY02E2CibDrCuHdG8eAiSd
TTI/NgYTfVzGUbGlVjyZuz5QUn5GBddpwvVa+PrH5MhzqTn0GXuDn2VpJJEy0aRwnebJw+UnsPuC
OEfJ+5KcWFnUDeP73gG6CxFR2iEESDvwIl9JW5hzocdWEWKn8veeI+NXDD4UirkXmOV/tRk7rFSG
HEMmTAwE6n+l4qY0qn0VCuStSa/8bEl9YqUZS016/DIpQv9iVNI/9iOtn9D70vO2HTkhqik2N7wY
1W1d6cJylZ9M1ENoq4zULtIi+CL52+W2ULCgW2x0mk4b/IhX6NG18Zc4YlihxfQsPuEa9zUW3SqN
AoSgfim8pyitqDR/NNuem9gLXxQ35wFpl/q90w+cJgGZrwIfPgYX+g6J8m8k8rgayLuqto3G6DOB
anfFY2hrvBPyzHSDpe2S6k6JZwpyR48MpdTmlgbJLwWvLaSAphUV7BcDqRUZqAes84kI9a6qHxb2
3k0ImsqshfsWPW8wqN7+cIYX9vy75CFiJbtA6ZgGd6dziDd98EmnIkLh/8Urp4Hn8osa8mNhNqGX
UnbdZmPu7HRaIwQ05FFx9MWmjCt0uD12LgM58nYew2LSp+rEjEqLbkApr9LcKutY0h1i5DEF2b2c
yD69MOo/noxVHrfUDqlaevkKPooEvgMy9QxtIOcscbWZi+qfrPfxee8PYIXJ/tKYcN4CkXl8y4i0
tdKpkNqwhD9lvPNRmzN27ZmKH22LQ8MikVPVM3mrY9JW0pErFcrqT/Ij6Z87ic4rdJkKSCVgjNHj
rCOQX3xIEyyMFTx9y1keB+7CBV4Rg4kb81coJnPcRyO2gZF5d0MTDDXoLiErupQvKqzaEqswwajX
QFDMnDW9NlsizlWRJqod6Om/LVD3hGi1OuYqv41M4Q/Eb6MIfu6rI2jmEyJz+F65MdSEeWwjVhgI
EuPE+PvXaPqyRzC/b20iphhicXGn/0XYNniXWSGyC0Y1JQnWZB5ZTMOyk+/SJ00Rp5dMx4LsCa58
9+oqqU21P4dSBhCeSzlYyy5wcurEUK79L7KJMgEsPCpEEF3c/MnPnhcjfLhHmIX4cmbRX7mYviwN
or95rYxgaAfaN85bNYHo0EmyXpxjSELRumvESs1ei2vZ4UhJB3w5zQBhTs4WkrKpgOowZsAzKjrw
gvmMKXXtmBB7Fr+T9o+eXUzTvp1GcfVDRacpIsD+tYB949D+UBZ7CGK6vQAK3xkUmxqD1qRj1uL/
yIawvqpteoWu5rRcfAwzPrHuEEtptstu34Qw1ixdkAWyP8HREIuOGAIS+D3OUVVgOSygxKDSdEzy
FsxsQJd+GqtASr4OIp0JvyPJr8Vj1q9jY+ENWtypyKuCFSxTgAJFXxzaA3bWJYekY6BgpYyVn3NN
cPRg8CYzjVkuNo4lgBCBDQmAbqsjHmQsQmw1x4Vd/dyXXQI8KD6FXqfFbArNs4gEVEDnQtfW/Z92
dqv+TrSEh0jgIMtNdNGFqZ5Zhdn1GiKZ5HNbJtJPvDFuqWpWcRsm6bDhKEaxgactd7M5OzipQtoM
3efG6IoJYyTeR1mV78PuQveFd3/u7NpXPLsFFDnBjXNK2D4e1jyc2qZnBWOk9nyLZDr7Vy6Aiqae
Mjvjz2zmlNhcigJQzMe9jwTByoiZJlXZ6xG74gWnOI9TKDcpVmWIgkjcHcplFGpVsq1S/kpL1t90
5Wi+8arOaRmi+EIQ1N6EwAqDpb3SyRMW/KO0FFy7w4KoajksqCXf3eXxhpfTU+k1AfddrbAHcOdL
m7qP8AeSOcryLrh7wxW9GJ4WIYFTX/SutHbVS5eN0ULHtIPn77PQ1JYxedNInmlrGVenh1aFIem7
XnT9PFQjvoapaZEUuB6b5K5qjWpY801oE7/CnaKW4uj7rN+rqVPfQdi4Zlq6ALYCg6sO5sh7iYz2
cvCE/YBo3kVVbt1j3nCsscNep8+2PnQ6cUeHKhkWdhaoLJYD9nphKkae0fgbo89DuZL4FmeTSa+d
lDZwAc0hyC2TpK0fI4r7wiH/LUTFxVdC2se1wD1cC/ujtze2grJTOVikxSKDqp+tqkbtSwMg+y1/
CGWng70FBfcNW23BNTsOEMngg2P2wRh33XqTVMCqj8xHKr0rPMNAC7nXSNYU6Vp6VzF9H0kLj2yx
UTyl/QuUrfVoInoCmpz9rXXD28VopQOGqCCC2CgbqhgLRrbnDEApi+k9dqX/J22DfqjFI5RtqDV5
ucRr3q0PL2hU6PNMO8ReIZVtR1zpt8qCtTKXUqgvN61Js9UfuapuatYvXM7GkFyrAfxNFXLxfsYY
20lLmyWg7IEw6APuXTP38GGTZjQuAR+H5hi777gRJKeGqnk2ZCtnmkexdudRKmtRivtaquIUUYIm
CCjei4CflIFthpCLCY9/HlcjepyPa/8tk4/bcGB2lJ0gjeJdPKhyCufC4GrDxxIK6/Oje03ztrKl
iwN3RmQlSov6hz2jpN36+uBgwBAfHVTjc5Sq2aFKpnEo/yjJQcagsw0vfHn1p9v6gQayMKn//CX1
ieElf0euRCRKBihk+4B7DAtgFSmnjCZx6b41arTDaUe7E6IWkC/IvnuyG7sGC0Y5rrlbwBbBVOzJ
3owmtDuaIBoGJmKPcNrm0NfjiRAOZIOA/bFz88kJHazAe6GsMhsN/076y18Lp41zyA/Rr8JFa0K2
3tegVKlXAI4kLMoH6YgT90ApdZceeBDpgO1uK2bVYkJ8oZoddklk8fuurDkCrQ2sQY9EMXEgfjHl
O+IYjeNs3jQcq2U5D0Um5iiMr11pmobR3WxCEdkH9JtR/OyUS8iFKns3p2H/JALm/u+uoiOB262u
peBDmoIWtFWqWeIBww5ZAxL69Ihhc64xNdQIOXlc3cUsAJBmej2ASOPlEa50+S41ubckjNtrbPmM
J5a0QDhj5Oz+Tj1Pm4iw6O9JnSIh7cCFzIacf2iWsluYYZgnpFmrRBh1oHrzswGpAm6cetKtw9/k
u7WszyH4c20JVc19LgxKLgy0X7byvzKDgYA8QCwte0eiVAWQUpz1TfAbJLWdcGilGcsQN5jJYVNO
fKK9oQInbLDHDoGuKYK1xUXgAbLpkN+1fzB9IgwuZfIk6gkPDdmxc8t83rl0VqtOrzkOp+KzfmIq
tGDeO3xX/LHb7bO421PgwuBpvRunYgjYoO4zwl2aHjKAUQMPd5QrFnvzlt34uWu7AU13zAOz/00b
/kOK91ztXhBRuJBtCOs7Rkpby4v1YH1GpUMOFPmqt7i0Sgfcmq0Ji8vtorNBfjajm+zREtdoXzqu
IrfzT6dm9LAEsRS6RDt3AhhXdZSXxDcX5XrH8KMJMOp8MdYkoCLtY2HffhJInQoGHZycgUQmtiqx
TEnt525sseKGE17KmYCM9lI8f8sLldgSfsLgtvQXiOXCknGKCX9kdF8iROPvnxo2BuIWslIgQyQ/
nvPi4zOSY/uvfvGf0bVm0SiLj3aZwR96GmoLk9Z2QfO/5CbIfahh/uSBdm98MKSbPy+LuOWrEAdh
fNqiiy6af3MVfNyupPwaBrE1AIXzwgOW6hyQUc5R7QXibA4LwknfAYKSfY/vgnkPFGKWZiBOitS5
WFELuqk8ZompVDVraFtcPBjEVhbxs1E9vLeZOYIgDxKc5Ra74Igt08NexMHKgo2W8xpqp77Qwzcg
ACq21GL18fqatrBg2FQgtgUrqPZgugJ1MUWJ9nLv+N+C3pKRFqpTq6N2tB4jFVuw+7IL4wTbSFuL
CG/nQ6yYdisPAaFUze9m6xFKxLaqd2eFI9aALrubAo8lMh6OyNGMPR1W3XRK2082AI4+vU44ORHb
ch1k2LhNvXhIcMnC424g5SXTr0KrjYqFHSkUmkz0yIfD5Q8SyT2PlqLNjDwJp3oOX1HWa4ekargW
tpV3quIK983TOSO84t7iTdTmyln1fAKgFm5jkArNo5BBr8kU7sjAC3nrxyuQTIvBBuBkIzu2FGOd
4UmwPhpgjvTic7A4zZ9O/XYln9qS300nRezrv8eqe1APzdAglvQkXJ2clO0i9nVROG8zsZ8enb4D
7Dcmy4mZAxrvqoNAP+TSZ3haFblTRhMq+c/zweU2wF4mq6veC98Q1QDzMXp8qbH5xd+uertGuv/x
PUlJpnOIykR6lB8S2mY4EvDDVBjB1znJlCX5PXB0tPtzmMo38mFn4t/Anu3Sf/kNtnopqWoUX7uK
yxhjMr5WhlrdUy+jzfHgL3/TVlJYbnqyLPT9KdJjh/Z6mCSXPIDCek8cPmH+8PIX0I01jiSZVwWu
cQoT7SjHbREWVGLaWWa9GWeefOtLXe7Ux4hGxMt7EX67iODyB+6kP+VubUdYVNqeISdHdak83OX5
uHqXKVilxvaEIZ7TA5WMF5rfU03ZUUl2ve6YTMD/VHT6qrRIKJ84b94iKXzgDSv+1MVPNiMfZpES
oVggcsv8KQvtH53aKQ7mVIRiW34o5hoFsP7oIUXT6jf6scmpTorRajtCa1t0Zm4e46RFaAC2fJ4c
E/f3+ztQapNLv9LeazK9xcs6Gb4uNYgiw7qKnI4sPEo2G8UFBQiOVbWdOuon5eSYYEp7yUNhD/lu
WbZdxVzwCGkq6XJ4W6UcmsDDHBYvQCOugO9BnHrOt0d+a4KRh+DVomRuy+Q7Wd/6ZKgYV5g4crTS
4Jy+2b7JHav5dBfSl4n9ECI/4HdbNo+3E1HGoWFC9qD8swhacTjcELiTu5zHYg6/ctamPgdj7ia8
Rq6y/spMAAKDw9+tMUo1v0lDFJksN71laoVykbye3o3sUVpAPmUIknd71wYhvjqj3LFv8Yg2NY3E
qeItnnt2nXcmo0UzckNFNW755B92D/jWSes0NVYJMxiOS160HBPils05DhKPBEkv1dtWD6GGmyaC
gFqHKwumsKJdEkc6BotM0eMGv8B1q/mEDhcR9NH4q7vIh0pZQoPALATw87y/+/eH6NL67lCDnM6X
nitb4apOm5grAO0jnfwwlOiP66VlVaUDWITEnLrKwD8kWRJUoM6RmOW35uU/vOKxlH+fDAmVGN2v
4rAICBBGrqZU7yp96IcppcPNhYA7yjahyUPie4fnhnL+KP3RG6Cl4bkZ7/uMPbB374VcDC2eNx9x
/tPLBhyqJMdjJrz6ZKR0RqQZ1Mj2vkTn9q0mMRtD6r934sMk52+3YIQ0Yi640j7tLHpJj2+E/JV5
njpX7YxRlgYoTI1b0ZYZwIQb1iigQ++Z0x20Pau64njpdmAccUN9kgL6Ywe+jeKM3htv+bLMzLIH
wc2y60IdgCSz++lu0++IK/ZLKkMmr/0pdxHnqEThP41xVt6RyC+KOj6p3OaoI5TlIQ4eYLtmwGe1
+9EmBLnGUkngky5/2z0u4DE27qJvBNH/INPUNVWmyvvn+5lvNl0abobtHs0wiVptUVtATFVuQJk4
d+iiAhQLmTarseuk1T2EiamKbnhKRt1YfLzZJ5Wx2l/IxHOZBXBXrcX7FP7qAe8i2PVT9CX8FsvY
lQHhorYWE8502bQqa6X48tNbLxdn4tgRg0gXt2nSl24jDAS9WsFmzJyueOx8zBu2mFIJfOszAJWv
pR1vZ8xp9vsod8VpG9UMdnvRvxKhBrRAaRIVAHG/DmaNvndzn5UNKcKUZla1eNsXLS7URxvIxRVY
ZLAxEr1zhjOjKvPmk6lrqB15duHaOd4JeSagy7IF74iRQ9kBBJ6g83T7nB7z58fvEbIkH2nR1jQN
zR3o4gKIu60C4m3P8gawaci/kRYGdlisvdFxZTwZBuMskFe83of6Hb6Py55vYOnBtDolrTapb7Kg
v6F5r9G4AyCyxzhgM5Cv3c6+/98FULNqQDnFZZsrGnBVdfsfnvRA3Yq6n9JsO7RqIdJOX6WtgpZ8
Rh7Ay+COq629vtuFuA/jjo8LhLqpZCjtEOCp06OXXOyFA23I10omlFT6L5fblYgtF6dObDaPT9FR
RaYggLAU6ZxlSrq8dcMfSkCPREMBbxq5wHEG1ANnJ9kntpHPVgCsrx8EsYQYVx2FvLv18zWLgrKb
uCHBNg4GVBJNSHUbUG+Stb92ZzF+6C3PCwUe6JvvfhJaCMFyL0/1UyhX493aLYT1YTuBHo03DwtQ
G7LWj4tZWsqZMnI8eBWIa+PnRXUsRLOwfsgMj5PsBJXu9f7KUJwe6bOGMmmImd3YwXwItLqZu7ZH
1FFZ7G7xbM5gdMZUV4u7I6Q6eTcNMsIR/6YFbIe5lIVYIp4eAf26eGouuYgqORB26fcs0CcyfJsK
tJfubVDbD2Wq+GcKbtYqxM1Wme1p40XgO2HU+1pB4yeJcxMezCFppJ2AiucOkiNhhV1Dgwlh4/xE
Z27Uz9x9jMZ8GqlD+SmIp3OwvEJuPaYPRha7mT27rRuCPYQsJL/96PNUyFLs1D2bl5R0opHQxQX9
NUJdQ++Q4P5f8df+9Fs8z9cL6g0xpkEuHbC03zqiRQUun8L9BJAz0iyxqWDKjeISxWep7wSpqu4O
onGia0xki/xl2dIkFY9czED15QLTZA95Ke20nUm2/8ea8amNAc2SPm2K6cJ8+IYMFWqz9duqUCvD
aCZ8dkqPBU9bs550vpiEc5vAIBlD7KI9qCxZJBqJF5ik8T5XKiYfQLGTwIIC9TWu9us44jSW2ZCw
elZ4zKL88iba54syVejaojFCwYWRgLjbJy9chU2lik80svp4Zsk6A7w7VaWaPMIbiEjKkrGdp6GU
3HiT1uKT//EtNOpOtjcTTHpxixQk0zFV4muwZClsrlYXIaS7/qkUuu8veKFbQBOce/iPik5MT+Zw
ctCLx0jxErd5EpLoEJ2JsMwIfzarTv2bipbU1aqEGE+ne7zGBxPhd6n+EfMoieORx3/jGTbdY/xD
gXIyZFUaAIrrx4AA5RUEL376VRaNMBKAp1S1Nh9cBP78gSN9+hWrLkLUW3RYYiyj+7LA9Egi6jMR
0P74hBu3nNfzoo5CpcIbUR1pvlU1/JS+s8nBGQ4dgV3WsYh2mu3IYeze5bPn+b7/I0HhQcM9b+jJ
lLjE5rIyDOCs9XGl9UsPvmuZe1UzLF+thfllBJocNK/p3NBK2iGkbayHbKRbRObKgVJGvdpfA7BH
vwnsJvSO6SyQ+YoezjfGoLZOqWHIYK6mD//j7Fc9x4Rwvykctd5it6J+pUPRMFHTVAmZ1NlTtJUJ
9YJujJ+QCEoDWmVH0bwBpD+ZX5/3DWqcMID3ngHFNCxn61uZ3aOXsNAorMC0kBdYmy0f3QP+f+sC
mg/84GkPf3Kj43/ie1y6qsV20fBJjbjVIKOrG8CWRxxsJD6Imtqjn1aJa3TvfyAWw29h2eKfzmMd
ybTv51MATSF+coZE7k1cV1qYTbxQ32hDOX8PkyO6en1006jYxH3JcxnAW3TY6Er4FnF4HJn3wxN6
fYCS5/kloMlFs4bOpk7TJXHnwSL3UsgjBESEsryQ2Xa1kLaJvhrgC77P9rfCAGbdkJiSe0B5ueZH
KmwVFDQ3ImITetBJ38qQAQjZBtZuJ5sPXc5D9bDtlAtyE8YF51fuojUWeRyC7GsvoBHYFC3Q+3Ij
cE92hpjml6k2xv0sNb2VcEDtCaielIRy1cWdru21b0zOZCA+0yEve9AotsRzxpaeWAJ7twD/hT3r
uJHPuGL0WyB0u52M41x4cpyGno95UATd2qOXMqAZAl5V+hrxUKSxDlQH1JKy0IFyPL4gei9/tbq+
w+LAeUVZt382nZEOOlCGXYaiEF8txqY8ftk37UB1iLDO5p18+ahsUHiy1CV1wOY8DiFL6TPJ8f7Y
OuSo40IL9UcgDUNj82kXWTnloa4g2/bBvY0Kt01Rn7dzu3i0TLO6Mni7zV+JzrtzzBEwSYj/5mRx
D592iqMykiqsxrrFeIk0EwuF4j35/7EJNpWe1mkztAnDiMBphRLa0JQ+uE8+DHXyZC/Sg6uvZWIj
4uz+JzIUS9XcF31lxAXjTADlWe3cnmhC1rt27q7fVlhMsmPoRWg+soWTJj/ZeD1W7+EJ4mdKsGFH
jPbX+nmkHo4Ejnz6g+kYEBGUhOU0RNRtY0V/Z6XGB95H8jedkIXAhd8qWv07qyipZFOtY2e5FDJh
p6guIRR9lIHghFQPNFyVetxSSDgZaI2C6n5zWJA0/gwdXkThSjrbxutCA/ujnY5apFo3r7K9gZeN
wtGFqFK0aPc/ANUVSbn766A4Qu6QTgcOs04kqsRpLUGyjuIJhhqKIJWKnZGKd9scy2NHY1gMjS06
27Yw29zTxrS+/wYrrHPrGiQK2/EhhX4cQLjOQCyf5jYxrZbNS+0S5uWkREdYcqP6OTnfgX7kAMfr
4KDjwtLGFjROm5x39xh24Ul3C7itHVHhS9VcovbhhrUB/1s/jKgC6aq5a1kVBCnJ5bwQdUFld6Rc
NKwjTbsMu0dQsWnY/Kz6asja+fPR3NFFLJ3O1U10apB4JwnXTkBz8X63TjkfJfSoIjc6UXwU+xIM
hhEF7kwcSyRxK5789llfMXqbEwQUW3NEm53uBNLHI+TBtb3/ooWMoSNjSZ8OCGZLPHL4cMLGX4dk
UxjQ+fpuS0kGj/ip5mAYtHRY79ikETiJ608qTtS62NqmoRyXPU2ylzq92pHehO6IhvK10BFwYpEe
oPpTveWyO5K5xxwUAJzmGJWEZbdOttJNE/3maxTjqInyI2SJG0u90ZK3pNHIBCVh4O+HNZ8K7+lM
sN+BvjabrCvy7UrQr/QrEitVc0Vb8l3mAnVQJlJa9htJ5sT5Hr2NCgdXfmW2OHVig0PxsJcTX2XC
4HHhRBNKgr49aD+4rMvtLeWAAbfFqprdw94Y9TjAAHu6cfrnIDDSmPa0IS4R6jtEQoHda5/eP+RH
TmCp87/taQD9zzGdYiY3ONzMKLAf7zKOgF6mfZSBACJMXFUjY+cKvtjjnhL3k2r/feFd9KMqf/8F
K3f94Chf5LB9LSRQZPZHRdPsFEPudjLMiaTbQtoRPH3L3qcxU5Asx9O3AXN1CTs2CgwC8aNyP8At
W3KBlpjwOR8ig3QurGN3Ejnbt0rGxwg+w8erNIH7bue5wxegtQCV0eYXkDCXE8gEsOatnHBol5em
+x/ay05dM7BsvBh7d5sOCG8FHT2y5aL7+gOA4EJl2fZuqfGJK5NojtrLWP/KPxlTWWz68tuUzid3
S33C6fPBYUuCAhNx9Cxvgl+GQKkQ7Y+hs54YZ7As4oBqOzLFtxUZnZBiU9yHd70br1ToYjglEYsn
wr/J6tYlxODaxi7iayTxp4pw0n8efL8vjcefHqVW3gQSJG66JhCUycN+m0W5u4UUHNebAC7Oa/9H
cZDFmOmZdtve31Quoas80he2g+fluVF/Lo7pvvDT0B4a5xdE/kJEeYFATvWOOLk97wH16+v5R9j2
S8Ak6aWFGvXYMJx030/sBSH8OKUC8wLoCqKyyKbpXPn+umohNPHy0Tr2RbOXr+4aOvk9UGucblHt
5wlb2YYKJ0QxKUW9/KtW+McMqYtNv+FOcGeyWtYOGEXl9mYOqukjomRtubjnqhOmWJskO6ry/wjk
jqJhQzL8OfqxGJgyfuyqxsUKSH4YktUeNj7IvGdzNBnoPR3Bo4+SI+t8c3GFr4GzJFrzOv1PZDw6
Se8yDWGKpaIt/spc13PsiIvT4j9EsT8XMIHldC79uQjfOrpECkcEnPlfjWGBEL6uUQa01oNWA7YH
NWED/TtB41qZ9V8WiIyf5ipsv70DgTb+wjtATpQuJkDLQGCv2KoiHxuuz3uKhGeQiBLnGpw5sxP7
8kJpIJ0qsTtgaXINx4f/PUat5Egli3CdPmWZ0xLrfB3JQvCf66naQ7KqTr6ZKgHpw5xlNXi9IXFl
fYIpfta0tito63XyDZQ4BcGptpL7FH1EZ6GHIZiKHEpwnFCtze9bwzw7udt1CkYTDu3MjAI1sCc7
sMMx5ZSYBRS/tGnOnczQhbUV8hAPSR9u/aVNy2feVZrNKV+gRd4mHhq30/R262+XlFFAw/fTLa8A
Phg/FmtW0+b5/qil8vi5Jv5sqUMnVvI+BAkuZcein/Ev4aBhYDQ32kBPgWjYc/PBJ7mBkMsqZjO3
bK3FgRLYLxpumzeBr9W568q0culRG95JVapyW5USxuHqmjgkAFjLbAuZP16juqCdVfFNvYXZgQcW
mc0jteCfzDKutm0DobcJd0v4GmD+q8W0C6G0IdMqXm5S0kW3hlFbq2Pb7l0NOwnY+zJs8EX5b0nS
KB1M+MnfwvLVPWyYBxD2HPubrRW4gDCC4X9+gFJO8pEVFNj4t5oanY+581IEQhiA9mWcqwGnJb5u
DtASgePBtbIWR1Z/RVZYQFsGmRTjqzIwqoO+Y9f7+Nxk9xnsgZmRlUCYYniYu4It7uoKe+mEvLRf
uWp8jpYMBmQSi+p2yiL7ApIA94WaIcv8s3azprxLxlkUgYve50cHEEaJWFa2yg5lnkLBjOreoDUe
gv+7ikGJgt0cEyNO48rvyIuaZaZ87KKrMuj3q4TkJpLi4btZ9OxwaQx9V374WsS1vcexOICkmyfo
iUlAs2X2kxQdDmlJ7a+U9BfC3Qn9N9F4yWEC3XozGtdRW1y5Kx/y87MKSL52/zd9826SFVrMC77B
+VwIS8VB+q7nK70Qi9vbrW41XDxtBU/j/SsI4XuXT/sOU5bGbnndT1lWq4VTZbsC6jy8J9J16OIk
HBO/88Agg8KraJ2z7LIbFWoRMsK/LHpmheJlqIn9rfRgGl3U1q/lEJRY6q8qURfPWdY5OmO3uNw3
cpAb8rG6/Nsn1lfMW013E+Tyyti3y+A5KRO9bo4v7Hzn3KMwJEOb9Iy9XuMEv3vMIK9zWyUxwBKm
XMV5d1s2c56gpaF3vjTmPMHKRUpVmhfpbTBuaWEiquSorSWzTRSOKSguzILZcuWtUgTTV1bqht7J
BHoQDmtZMKIwYo6vHiuTd55j4dQXOj4UH3tGFLrHBprT9pWsQ0MFqepOY10Gq/q8hb/ttHyja6ih
P4r310Ueyme/X/58kc+biM8dvoXy7z/XRQYwdhFohrolqWxyX8e/46CBPfkkmjOkXZd5wlwLhWF8
Nni7mQiyjF6iaGB8apBYqCOHhC49j9FcGL5PKehDNW/GaMRvNnVFbME+3kAtJaVmJnxOsdSZzWFT
OvQnheeGVylb7LUuvnymhJzs3mv8kIV3jrZ/oajCFyL/svmLzdNNSTc/USd2l2rdaSwmcA9gm/Lb
AqJk7gP6+4G30kFuKIYkFDk1LS0jYr1dff//+FzA1ULbJwGw0PFpVWRU5Rku7dotnz67lGofTlG4
Hpfmj3tKc3Kv4JFQ6pC0353ORRhKI/reZ/lWpdgKKag9USMz9Bstz8U+viX6c0zlLs7u4SCammJO
L8kJnaqA50mV6BgjwWhuKXaOUqTsT/QKtqFfUXRn3h0SfzAI5D0RbbQBpXtuvl8gjCTrY3wnZQbd
xQ8UudgHNZnmRFCN0UfMvns3ETW8pykirs3pbWhUA7m/+kuV+FFaZ6N7HtTjazVYeiUpr+Fk5Fpz
HRMe+RqovBw2wX/NJK5+qmew5/AaO4K1m+rrxitgBW44ehkFnVpIMOFYNFqpkkUe8eJfQVCs3VmC
MWzI883Sfwva/8zQJlAI2gsyN1LZJQYdEuln9N3SaKqv3P363lNlXNPQy9xBJxipzmRRCR3WXCI8
R/LaP33RhDjiQdFSwZdxthkczcio0oRqhcJwMsSrQeY8NNWF5Lzthi80W94GkFpLEmmsaVMkkGmR
YC3g4kLeDJPICSgZpFMBeJOc/amLMlKWlbNKc0OnsEkTU1wyrWg0ge8YBWtxBMKB6fM+HjweVxX9
wjo/gI9doH1A8oi7MO2Jw87uc8oh7W719fMlxSSdhnndOkRq56PetI65A1p4/hgMvd4gSrgO/bZ6
IqfFpqNjDNqMSSLNhsRH2AKPsl6bKuy0CUoCxDhjBXkuOeuyZ8M7KvTD1F2c+wZyni4qjFVsiFT9
iDJZtlrrxCUA+6AlOS7vZ1oLSWDtE2BnJiMnJ1h26YcqkUriFlFSpHvnEuEbid89ECakX8eKuSSo
48YtYw7PGHwOy/5Kcx+MFV7bedXFdBPMRvlwbbYyrBji4Uz36hA/AUS/dgNJ5oylzqShEy0c9EG+
R/EtvFYA+lIc4DQTbJmRQ0FB4j6+rkg+WUdvWQc5QauVD8YXJ6UA2iK/IZ2Vyt2vGjln6VJ1XL+K
CbsEV8DDKl9tbj3jEMUrR8w+9rYPwMIQYlPo2SkQO0KxFzwTzbZYl0sLVWyUq10EnbcO+dYEOegC
fbZTagPXuVVs9H287wyPc0npxX4wcqdlBuFlWWKOOqf5YuI9UfkzKdU7M1sYNBuNZHDLo92vQ2UV
nLi4kIg/3UxQ5chNwveuaY4UZ5BZ6RsyaTg/HMed1HiuEPeKF7iSspMQwckqe6UvSu5iuYOZF1l7
KKeeHzzkulwY+uvnl1vgHrUJg3qO/0GvvOhRlmZk4imT544ix4fg0KdyVAIm3P9guzIByjfnrygd
DuCynfL2g2IdzQzj+gIilVEEggCTuED4ACSq205iEqMY2ppvwtQk9MEW3R+JLA+JLr60migWwx9g
vzdNZYp1yVDv79jLblp6s3VMghZcWdp4H+iALDXUOb7OCqme/GwsG2x6zvxIIms2Efvdhp1gYRMf
2PSy0iZy/H05LdFjtbbVWGgYJsQntG7C9TQQ8XyzS1nteBkbQeXtkVf059HXLGFtBJ9+JGulihv6
+4zvn9GXu/fcu5S9aMxs/rcm7I0ZEtyIgnBeuyqazi8hZXWMaLb+LKwsg5hrzqNvDCDgvHNLwopo
U4tefjr68/RJDaKpiqdY3DjphBcSleHMFn59oFwMa83LAawP6nZoh5rXQKRHMTNA7UT9TcuJc/9q
v+SJkemf86zfn1twsenuNmSEAOtb0t1ZdrPPL/B2plWTpytNrkIx5IxBmtTrfprdHaComnXexr27
aJRiX+LNreJ7x4zclq6hWoQqg8m5sGOfhJ5JKAm1O1tMBJm8R0AjxSTeoCuMqdVfFdxt1i0+h8J/
rICa55tpVYRfx4TAiP7CJmW1NIaiuTL3T/t9FVhWPVfDQ6bgmhk3H6GtPtlDWwbLgTKlYkhv+WSY
hoAStd/wI4PZGnYQsOtsPfpeaXEfFClskrKdpy0B86X6BWBHpEcu9uK/DYc6jVIDPn2lUuaftfXV
LHIHX7jMNI2+eHR7B8QDnkPAf/VJJZvAtzUGFE8ZCMqOxADh7TXfuDeDmtKXQhafuxmDkQkValcp
SYzANjgqKf3JOZVGlQ+Nsjq1NA50XNTV/qJWPSmidf2ScnpD4HV7XDRxINUW9ZeCpuERywFaaaWj
N81oMMuL2eY/L+3jg/MBgc/m//TX4OhgYx1+lR9vSbvS+h1nNqKK8rat7fcku9/a3FarjYfS4XaV
QmLysOJuwx1FOdLU+XwYffyocjNHPwp70ocHgMTNgKe6P0cxWCPc2UXRyc3yEifeDvDNrH71OTlZ
6+X6YwmgClt920j4eg4GH4jx0YkjbrH9tZeyAJgSgYTnItbe+0wacQWX61NWWwCPkXtbJEMJyNER
hxfds0JE6nYojbiR09cMX0kg5gsUfTjqmFAeHnn54P6BkvW48bZCEgtdNDt/MRKqNqQ/dUPqjfLM
04IDw2o49Wg7dGqaKb2RHzYIhxrtDgWleFUQ+BcF0kgonKFCH2w9m9cTgjfS2B78XwPBkZC8Oy9+
0XDd8UwynFRZblJZS7GPxngPf3lErZww27R+V8BMTPTtP2FfcwyoEHKV6Z94muU4qSX6cwogeVZ+
MJkgww5cOA0p2jW7q5x5Q1et/zlVWcWwyyXhL5RuUOnNnVaw9KmCFlQHGUdxBkcE7qX0NEkhDaSv
eLpiaxgFGKHxNxAUvQ9nz03XyZpv6synx7LNljHf3c5815Adkf3UccU2v9wr4RqoAIUcxeVxh+Cj
d6oWmZk4Jypti+Ezeovy+PKmHALPsa2PBzYaaxkuNzLMzBWyW7pL3mhdO/sRoX9HwBbwHuxkhhrI
EaWnEKzbsFqsrzA8axj9jtAw7sGtBsRes0e/t3V34g1qBUA6gl6BEkEwpXBw/cz0HLhiMpJYtSxg
zeeZF57N09g/LmOTBOn8aoF0ptqjD8LJaTzA53cZL7FI6CU0wIPt/Von98KRXTyxUgNgRlzy3vAl
4CGLrJc3hbPT4uvi90vOzDiG+XUdWmlJ7N24Xi9YsZTsSfN5ytuWxroSPYiOyKcrmFoiu+AO2jn3
2G+JwEoBmwt8ZbW/PVtGT8dhO2VgLOPOXh851lR74tZkVlIX4QkUQ68w9VaFW/EUwHv4r818eQZA
ZZecS4R27rpNuqQ0uptl8n4faDLAa+V3PYfWSzzgreDYA3Vbn73fYACom1p8dGjxm6lbpXO2Ws2q
tM7SgOxRHs9iJpCmBNeVsuGqV/ruQ5cSpvfHEsbwUBtM8H4B5riWM5dfGikD4iI+A04xNEt66FzZ
AbNHktM8rSD0FP0u0079yVvw8pWs1WQ3MAMJAlgr5fJOCDxj6ZHvAbYstcLZ6b9dHP07lYcHyNOO
DtBME2ZXlhkxI4wr/UIkGlBsBV43bHwpHtfmmEU0HNo69/4zKG7QuN8Fzl1IqoUHCP4hc7eGMk3A
eWdcYYHDaTvvk7PM43CFYBUx7OUuABD8JutvVF9vRrRjZj2SGt4x6Kr9wublOzll2FtL32yRdT0J
o0kyyRFK4h7TrUMqrnBi21vDPralT8vrWf6Rh59lH5JvHmo3r7dAS5O6FPrDwTFQtlaSNXIwqzTw
c/HimYcDcLaVF46Aup97Bj7u2PjDy2e33uXlzEwlgovgo7slpyQ6Tfg4rkcFfo8xORuX+MSB4bv/
vv3AT00Ls6qqRnysuicS/KT+AzyX9BG4VnQwqtzaaBa763mJfpB0ud+Ofvv8QRMPKm6/UAnFsp2L
p0JnzxAP60ZwpfKH7U2QVoV0EmUAlFLnu8iUlJeIyj+sTXSzF+oa4AQQpP2am7Ji4KzoWuAFHCkc
rykaTo/GEI8DxHJpPkNzzXPcI0/QLt5ew03oOH/0Gw6BwXwgiHbBwPIOoSehGf54NZDG2XP+CL7K
CpyEEQeJEnh1sdJA3JkSAfCmchtJa0MTZgnWAUIORoGDGJoEMhcVhih4jTTZL5OSGp6LG8e4TWAU
tRzDQGjEgVJUgZdpE1BU1uUp4M0If2VDtHXhCmoeojFfR7QmX3uIMAWMWzgd00TTWV/n2l04lxje
C8EshbqhPECQjG0cICGX3W+s/o2Da6v6dGtJq3Qiub14UgBnJgbTtd1bcoE46rA+ZVkD+5PP5Ks1
nVXAcJJUxMGWjIkajpwZ8ZU7HTV0gza1BVeruTY8SU7l7Q9fT6D+nXgrX1DLGh5n72EK8vWzQc8v
UJVK4dI4xeKEO+HLDJm2ZRpeckgrDk9xXy2aTe+WysWNoO/jt4rTz4WSmTyTDnF7M0N/6q3BgKRn
xc4TV40pAXWAqB+Gt0LrsJ036IuoHWCp5gPNxukW66LB5GPs4TYMEyiDoCPwu4COo+w5IJIvzDm3
1A9t3NeZ2eGZnhsIxDjlNFDTYHJfTht+f9e8QQ7t6uM+Yk1MP8LL4fnOZE9dudGG2ab2jw8Qhr3x
Cp/GOz6oYfVPj12OwE+iwqzOhut+9Jf/JozgMvJdVXpz8OybEjb7bbFLzCqE1yAzMMfBrod9CbI4
rtUB5Oj3Jt1xUytN6fnWCEjUT11z0amQO95K8rJTo9kBLHRGBmIcBUsWFt1sr9TTuqgJlUL9IzrD
kQJ+qiMqxQTPySi8GqhQj/ysHsEI9S+nyc1cBUftuwBxOuny9+/KXMLidQ1IPOuClYylJW2832v6
AmWpe8dR7COSrwyDBo/FyPJD8jLIjzHLp9bMotIA4fu1NeHUKaLo5C4u7p21/iJLOHDg6z+zEzmD
WjbZr9h+2KGs/UfclSnKizFInq2ybHUkkSVj3Ye031SqdCGcjFVvRXuPiA7eKFZV4wPvIrTdImNr
f8dvQ1daGLffF7TOyHhHWCG3r+k0tUmFHnupCEdfGTP7/96w2m9oiRfKcS1M3LgDmPmE7MI/+i5Z
xn8vcMAUeyJcBPQKHs8+yMJRnLAKlbUO8QcbnPROmJ7DWouSylhbskNWADuNXgpfy7TCEcbD00+f
l+zmJyy5c6aUICETma6BONeBmrCu6INbFnkd2akjdiHpymwAhHtiOh5rGqjtAR7e3HIJxSri/00O
uCV5qKuqPlAu/O3Bw2kVSnKxDXNk1IOILuqaoabfAXAXpsZTyuYLDICKBbDB1izFhbeRNofUzNGf
R7y3qK6ZjrAYKByuZWqWQ/icW8+3rineAbr3FVw1lsBIQMNYyPMhg1nNOEWRXHkg/aXwMZ9OEmJg
pMlS6uidtoaZrVXYPQ9eMk57pi6MABGhdDR1p8FOd1pUWhTb5ZMeKm4EXsc4WoN5FdOMY0uUkvEL
bL5Yl2V9OkiXSXuWOKCnpTSo7R6F3YDjmd8UeRnteG3g7xLZC6p/Ly1LtbRgsvcGApSXjk+o9nl/
9r7MPj8BpPIDWB1Hmm3dCRuBjKoTf0Pm7DoCv5LKBtGff87YjeUIsCop/brqcjFBXKIpetgvtpni
UqTIVk8y3bGl1D2pubp9WEK1N9W5rDJ6gY6HbMN9gAgXc991hDjWyU0+JwUzAjlXwstc4G/RaR0p
W8/jPSGrw1ag7PeNkUMDeaC58jd3WwT8LkjwuBkwwUSKe7sbtKM/ZQdrpZBPhDSDMq2mDsHdwSYJ
joaLKIWeA0OChJAhY7o0GqM6jSh+nLSjwhf23k9JV1mvk4Ydfm+nYeSAUttkxrUR93vwJIdsCIp+
IuYUIQL6UlwlJMBjqkpDUek7zqq73Ae0wALGIZUnH00fBae+gHpo3A+44T6JjXQ9br6+UcBPKNXu
drhDs0Qsljxe3R02VVSaHNahz9OvJrM2sWCQdSDKwp43/YSgqbZaBbd+G+JTGR+nSM3tEx/Hrvu/
WtdpXwE561fDmMd9TT9pGwvNH3lDwtJrTkXwl1CykLfszfcTVy1VTHyqrCn34m2SiLE83vFBSbfu
f4j1Kfi2wN+VGT+E/4VO0/DbwdNZsvpoFcJ5P94GmnoxpZhFxwkvbOpfykwPTwN0yB6TGk4iiI9g
TK7RzY3p/v72S21fySZYl1abGoPbOWqc/AMUz+KsF+NWrpdIyzYZ/vVIMuAsWWc0a3at0TuheF4k
A/a+rIKjN1C4pdxsmAv465xR+T1IE1P2kOsfR2Su/usDVVyhWu5gY0lzWISlYsD9c0KSSmvIite8
ZoKo/XcsK/bl4LuEzw+Upqpk2/mDt4UnAGz/AWtBOz03UgHcQl73JnNHfbVMLP4R2UB07hLlFr8s
oyUTaC35ew55vBDX4pnm82dq6lgr7JAyRkZX5Brefcs69r+QKbElYnXQTqsI4uG19TGx2rOabFAl
AHXq91vQaI8zL+l1zEKmCzCSEdTVbLAg21PkAMg/dUbl0IUo3JLcHwdtGNLCLiSKh6cqRKO3MVig
iV41cMgXPrp4psJIKloREs3diu4WcedPUjEUHeLFPD3iGSJpfLFs3BqizwTBU/W0iitgOpJ9h1mh
DnnDnGrw1hBCawYS5NgiqW6CUBT/RqMyZan6l/L0WO4TYUfG5WKmIWVRIZ/gcuKEWASp4+6AaArz
2t+BxuR/xO9flL4310nJ1mYmnSy+WCDwh517HbMuH3U89+msk3Gs4cqXW4rUhFTPEXkh+XU5d57z
z8eRro8kwQuPxUGgEAJh+PL05f2eZecW418YD7kG0Y5OnDTOxQY2vufbZKIOfpgvE7My/seLKxMB
c7v8MFaYKwrHvlpIS8YMso+8mvS2PjQrmQN+gXUOrCFGsIy3nA9MN08rEwdRqpmVy2rg9rVpcgw6
hxSTzP9WQYo2AdwulmOIvjg4TuBv4du02DLW/6IteBj0wEGLm++uv37Ij1Fi5E7zq65FKn+TKnwf
oAPP/gu90ENLsCjcbPGghoOFQs76IZHDJa0Q9qmnmrgqlLZx38nZuqlM4JVLGeJxV3Ch6xvDZmzB
Nieqd5ma4k2q3zzZ4/r1j7ZqT9FkggDpPQeVFOx/Lpncsdf70+lDpDM368kv733uGHolfGR90xcq
JHAKCuI0bYEWYJDMy2vjJ3BOcxYjUEhKFqKYVxhUA9N8U2kRH4S8rwaI2qszR5GUSnaqGZ5QIijP
QnTwJ5lpjONXwCmnoOdrvBUIA3JRRB7vCWO2Mqx4GgjS4aG9U6h3I10MznphX9JXi3DSOMhXJxDs
sEa8b6/QzVt3RbE9eeRiz3bClcXHMCFXOCHRCLrmrQcLsD5HJyowLd45Hux1TeGjf4CtHHJvd9ln
CBhNq94dkehv9l+/bETkmaNjvpbcM2q9lYkd0HZdvP39kaaKipA1GOflKo6A4C9SbZJ10XCIk/1l
oqSd73UmFbRBFJkvxJy8CzlJIftdS+gsq/rWmgILDnsSP+fvYLfnH6achh/y0uKUfEFJjVBR3Mqv
VZCBW0uOXh0jp1UTMYVY1SJjh1bio+Qi5gJI1BH6T/rH5bL8vtBwDqCMCNxxfdM3ApMDwMFdsCKM
fs35KMkYXhucKKR8cdYdv+N+7Sebhh1P2xXvUfzggfPrBLRTMVoQFV/h/Andnz8eVPoiULpr8teE
HjYCo3ObJa/TRevpw9vamz3qGzpxspQaajGTywnQnSDBkZ4J85MNhcgO+8rod/8MJ4HmgdnY0H0j
AWvm1dVHC8x0P1go6iT310cbmc5ZQeX0jZ56cOowaT/o+wLWf7tJgDkJ+/T40HbifryGYxBAVlBl
XqgoXCTDVJEBKSN5XjnoUq/YUOAvm8QQb8M5VFXdf4afJ4oVhK/WPobOajDu2NGrgVe7vMAwdwAq
U0HRLD9gE/HyKU9ighiYhYFDWeL8E5UXpTlV6rDYUV3+0i3cfqGPK7IjJlC/I6HSEQr3lrIOxeAa
d1GnnLG8XqNmaC2JFCyzsSDNpeAAYjpDRplgnyGcrtPEI7uhhPHUpZSChGLrEg/rY0fLgfMx3pj5
xlWe4OYXobHh3LX/kWx2ykJSzAjiUtZjir6nXcGhI1eroyQv92g1tlqkor5Lr2RuPvTn1lfMrVHK
D4UwyqF4ykdOnoRBHxxLPr6LnTjfFKGKAY+WtAf4k40XJVN2QMNBjIAvbLp5wU9FeDOjc86E1BLb
01VklXdCf5nC+oFI+BV+9bQ44UxtgGnw+3poQSnF6ZY/DHIfdnNnRWolxfN4a3yDgHYWCNTHaY8v
eRma2GEncRjehWuLUhqWIftYl5fm+Dg0GcOXBMvGP8mEmcvYSqRPzSoHnvm9k6sOjLg/t04qo4i6
o16xIzo0nJbYkhVjCttiN82IzuxDljMoJ5CbbvR1FCuociVTarPxY5L2pGW6Trg7vjhPFpqfffEp
maTAqKhaWpKPq3g4qff9K9x0K2MaH+DUNpv8xmiZ2q4TntHsLva+ZnjWjuA8KlukGaJqSwD/cMVg
A1DJo1oUL+DRVIJPbisYzhGyo4n3OMEUYUGiA06tpQoQXeoqPcMNCoc6QrVDYL8y6NulX+bBHUoC
y088sLU1q4zfqiiuvkf19SPF3c0raISb4BObMUTpJsl+oAls3jM3WAZYeqsAzqUa6l6umBuc/1Zg
T5D2ctDGtIPzyC7iavowNK7+mUDEbRyFeUYH2Z121TKMQcY8AoGTVgWggxcda5R7iNPNaDunkAmk
x1uUGZkkgAVfOqrQa2vbYK7kiqybDkWLzk9LbbQWHqY1BRqFs7CQKwsa/++6BEomY7Qn89HU5VeQ
bSTgxzuUJTFEPDsPZUuGDmpATZUdMV61pN6J2eG9oNcOTEmZFtl4d6ArV1BuQSyZsHdco8u8C2vv
T52h1dxv5Fj57t36uC4PcAQ/PII+nwD/XpbjgimLHCmm++Fz3+OvqxRVtg75KQasC8ngyAcjK8J2
gKO77ZJqaidgNKHC2JpnBunqOoFm1axpgJ4cqu6maUxeZkd+e9sW9V/HBx/qVlzKeJ9wNXo1mYyX
N9G5kZaPLjAJU+xgnc4f74JaoTt7uaXyIo8gZIh1k15KWn7WjarWyT2s+j0dP//WYL3NqwkQzUW5
q1jvuQHiq8yEjiNOpvQJD4SZDLISl4XqKpwyEtyx5lqZS5/ZuLXK+an+pggCF3XDDXSUvlotEYQ8
0QeX6X+py+WM6dILLldGn7JHvcgXkQn/fBN4sD0poSN+fWR8idnmH6OiZ/V2ez6000EcbY/buheb
ZYFUb59pJrlF6j57jUyMWMlXOLjs9A5j2L334zvOKRIqzjG6VrsUp8JKdJhDxnaOFXckOLX+GPo7
AUhZ+A0fpniGbz7h3UPrXf44LA4q+8rTmH7boGh4WXZkuoHTQo4NdNUfKG79lFkY8pbCe43Rubgm
bjXkn7zcyszXCLImx1a8Db8nBmT/b8rIRVbovLGeT4bdKc1SOXJrjvNey+kJeJcgCilGwqrPO6KN
tGyBVagbUzBcIchGOFwvD/Rdqj2jZm5TNFglXQWdqWKL8HutvmaS57M2vOn+AnRVXbaYPgo4Fw1p
T+ls7YZawuoh3wr86GosTLgJKg7pAWO8PhklcSCcp7ApYyhS+8GaaAfIu7DEG0O1SZ+lFq/AScBb
x8jFbRcLUA4QJ19lILjpdGjFCyrN5+eB/6y/DI990CD3yqTeKFIo3uRVpRgQWgyFt1zK/piTclCu
TH//gx9HkCho1BWksIIcBMAHV+qL1LKi1kGUJvakmao7+pXq05j5oN6IETSDEmN57mp/282T0MG7
TYCsGC2LPuNIxrabf5YJXPMUS6vbFjf92IjXLTQ8cI839CfBjwZzEtFuQK8VznvdofJpJCcoYLIR
RVTd617xZHNOKuNSpK++bo+PxH+W+z/CTFKzs3oZYp/d548+AKSC7aNeUomM02YFtQ3zKUaoddqA
4mkNE4pLPvjhRgZRaufhCiv6YcPkdEkVSNfd6CY2+wcCAetHTE9VDQuLS2hfKOrU9uQe41Bu2EfD
x+wszeZ/Cy6FKrkHVizCQIF4r6xDe1xAKJEKhOGCEPsi6gBkqwLMCZ56h5n8thYMcZgq+uNejQw/
AKvlTsO0zn4D1gzPBlBxrpiYMi9XICiEKYgFIcRI4THjMFBiIxXUozZU61u8EdAGaSDz569T4l4h
X0odlUmF2YJEMtSVOfIv7odzEUXxsa6hKhFpSydSPbn1qSe30LcsKe3r8i9HOB66qQg4TjhvBwQt
Gd4dlqXFZ2jRzj/tQgoYBMymmYh1MMxSv9AX45nVqxDpGP5gNots2SklufBFleQwpka2ZzF+HZMy
QfmcKYxRgN8wwrFTs2YQ9azUDCbmwFj5bGCO67iGrGiVLR8i5XEu06PnWGib+TiQsT8LG6uAVnyq
JavN/6R09W6VwZtR5TlibbHvGmKWadMY59KkklV9UTv0R5hJCCB2rsBPbha1JqlMMpWVgGospwLg
H/vT3oKQIC/BkJI3sPXyncPBXHBi36U04OQAGsogkteIhcnz4WDah7fYex6B9iw4p+EG+piVlShI
7fCVvXLU9vqsnmPmUlAnHXAnvL/g5jNcrET8CLoFrLhwA76j2VLa9Rhc9ugnwDImQwLuDZE7fr54
qMBE8DhxbvVYP0JTHZhH3NpjXcm8pkjRtgz61NtEqNtl7WFeVz5cPR3GQGy1gx1SVRM6OFOUE/tY
twAs2g6VSzwqr0BvRJntvBmzs2DA9MbrxHQSzVDl+rYXkynaM+I6HHRrSCGMGUq/XUqpzUI1VVKt
jNTwEpkGI76bYQ1RDh9aZL/V2g51gTI9WzjbpwO7K75GbZQ1zfF+FQ8xZ3E4dCZLWelulJMg9ECP
LQ8W0Xz6yzKnidGCZTUBebKtNwimluo6dd7NfWycvxM1D0ZjHECEbUG/ixMXA0i9aMbJkYYBzgPy
LIZXq4dCZtzlm9o9rzKaU/juwUcOooVmpdDLpPsdQBQe5m8KnONAtcoXWkiSGPXXzLUZHIUFIJBx
aYV43FEsKQI5cM1H7cpJVg/cGghDo/+sXhj30U4WWbHMzFlB4Etd2Et7VB6AxxYsNMInrZCM++Y4
XLX4FqPRhvFK3LJ2o1pg45pXtzbIfSt6ic2pLhlGIADk1rJfvBPJqS3NQr4YhfG2dOTtbn9B+APR
sqpXl9qq2KTvX2h31Q/LxiCJRos99wyh4es22Pk/O6FE1f0yhi03O57GFaS46aIS5F4k90tQbVx3
ItD4q62kTZs0VWaBykPj+8zxVNRkUo23oYkyNt63ZH/9BnoixTynZCaXQ48t5uH2Z6jmx+JpML/M
QCiZvH3FF4gjXnYwqwaQ+iRWldxVKzCJNuih4j6Z1+0Eiji3FWd3AEwX0E4dU1mcTxTiakDiVNDn
j73biNPdkKGuX3a55YDq+6G50C0aaPzhj8spE2+dzZGVmM1CLEmeEEj7ffvvXcYrPUTWs9mNWY41
XrjwFtGlOzd5kZuN9YxblzkV2xYoRCG7i1WKYUUkAbWfGC5DqTXr2162XnqZupxHjvTQt+5ASnjv
FDfVh0Brp5zbo3INpUEhp+IYLGJfDWvpv+BH+zcO7D9B6WySx8pR6cgYcuBJmyuH5zIMCMLHU8mW
4fca2ta02uc95XrUtfGn968LvfOaACNUDmwB+sEeb6fmG6GJ/+jtkQT5J/ALxpbW9NYU95RQh6XF
BEf4cvvbnNPWXnNu6Q45BYY3iDgPg6+fC1iQRQ2a15w+lA3VVxm4DmiV3CNaCDoPoGSGKub/OWfA
NL41yybQgO6XjI1+f8e+iTfkeZuvRVA1BGyRc5pGU/85rFXFbI5t+68SrnFVfxM5MbSskyPnGtH+
/H5RN3aKQBVnNeW/7Dati48gO/AvG/bWtfn6g2gZ+nTQUcDivd0a6Aw4RDZKImEb/E3ZcV46KwqL
V/cwxwrVG0t3FqSPxTPuMy97qjqJISFuwwCIHiLZDRA6f+EKG8cLUGJzIoIOn5gieeGQcf/lEec9
DOKY/OMWAh9ce2XOr8bjdAZVygkgvnfMbePjBscy5DkmrkZ2qiV2QuNpmxkCc1q1N3qbfPf2FOiC
ZhiIipAf9Bc/tOFp/4aky8jezbtneTHP7sI9K1cvyO9titXHhFxtURRM61XF2yjQ4CPrXaSfPrtf
/DhkQThCnn7B7NdEE+AHhxa40z9Ux8RBhf95hnjES+zgpeOTU9H2DDdP6BFHKnYxuMzaLKNTxwMh
so4nftA3UPuBpVDHaGky9nIh0ZfEUL33Hd3HW0J3/17FQg5/xSI5rMAodu+Bmr6vIyD+Q/g4dh+v
J0vG3goK8jX1RICuXgTzgO0epo8R7PG2t6Y0uKSNdCp7aqNA28KHzBpYgYwzLV1cXFjQWxLn6SSU
N1W4CZdRh9ULekH6l2QW94bppuat+sxUtn7lkDOMwzm2s3q6NLNF4m2KxCYpwgjM4wuwtPUMRleC
WoNFujX2gB0mEM5g0sbTL6c6g3PYYyYLnaVzy4mwc9gUxrLODobkwOwFrP++6sM1rqmGss6KkahV
t9CA4hGu9V3+J0DhmldrU8Nux/GfkGhxx6ZJ7zXKTOprHvzuHyn7ctAU4rkN/bGShViosnfIoE4D
/cFL/gObLOK+AoUFkeV1/7/1Dvu5K04oeCAB1OffkS4CZVagXzFheTWsWfxv+dGiqeiLgefR2cGA
D8M2HgIp6Q/wzbgwSBXnZSAOUa+gKA0g6Xfj3DYNwsYqiUtiGrllmi70eFTauLoGNnXFGc4Ipklx
lzJXqRXDw2ObVCkQS3GsDdtVVdwYqNdHcJ1t9uMNvVyslM0rhKWVODYaqi7JPc6g4XPgd9QwbChQ
c18JqmKJM+SUKghs0X2qfmD6cx8RLLz02RB7aNTQxx/HQCVw60jan7p9rZNvdwepFPpv533TunzU
VrcQuU4L5cLRBmpYFI59GE/n7pcmFPYv5ge6k7wCdGDB1z5V401HM4jFQJ4qd/NwPIkG24r3U6cF
UY4x1cVjD5YLMAW1isZDT/lkKZjt31i+FcbIwrenOYR1r3WCQZmxP/keAvjoyJzcvnlf5naRjE+W
jfGKyZF0AqBiGI6+tlAXg2EwFfpAPuoWP9znrngFg0sYlggHYBpZsVW8tVsDfNx9A8QGJng5PdOV
AXdHnGXRYeZ4VYvGoF7+9RYlirTPtcitF2tNydu9IAj9DfR+hCPnF8f38g6elg9ZJfifiAMdsvJj
rxfnmPwlFrLaB0n4u7Hq75heNIgyzz4Q0daGy54LCMSfIULQGzXjowGwtk3gSVzkeokplpJCEL0g
ETfVmxf9Lld7hmoSXMXJb8QSyCSToqYq/fFwOOw3G71vf0fBvIICVQO9SW6sqGhpVTmI4MHlu2xF
03Udqgmr9aQr1uB3Fmp5c8A/+318PoGU8UyMcj2PXA2WZPjdFz3NwR2Wn3IUPr09kx5ONcZmirmx
Me8iEgD6kxgS5w3VxDIEotfXGR9TlJUnHAk/LRa+E1RkZzYeFQKQfQ5z8jMS89p6tbX6q11LLWfl
JvrQVzghYoGQ/gwDQwTQOhB33YQly50dl+QCPqGnH/tble0/XVbff2+BLcBrjeIQeFbpqnFQTE2e
wFk1bYpF0B8oXIXaB7qEb/XAIFcbaqTdjAcIuMDgDUYM1lnIqcWimb+G/1LRbWYaEh80wpWmLZYG
tZgzSm/HPVcfqW6bwnXCjX0VZ7Y64Yvho+Np0nYBMBlvNiI+DYIXg5CddXGmlFQyYPEb6tLlYSmv
eI5gfKURVWNrGiLm+0Z6wqmBTEsU2EcmH8xPvALxFPnzqKdEWoXD3+LgQItmDcnyzEMUvMgBf357
UtfgIp0wW3yMGC37YNoVBB+S9mvR81WeHx0qilFtzZBWWresLPAFhsIwGpY9EvZjrrVunrz7T9cQ
FMQO5H81g1g3z8c1VHv1253nYTPOPsdyWXIv5uLVcZxjLAfEBGo8oMp7g3VgPBLFMsnSHeaBQIK6
irZY/8Y+91CsTD8/QQYswEHlhAvGC5VeOrP8pv/MkGvF92KyYHeGbpiKsY3WMQfxROByMtPuGPIc
+I/4YYZip9VRIszimSUN9I79+hw+haQ7a7J8nAfRQRKbnxBQpM8pa92I4VwXmUjjLmA4pcxfQmE3
JNmU6MSRcs1C7HHhkKixVRsc2hthurd+1wvR+ULr7iaJrZosyl11VzL1a4VpW3BdI38elxmN/DIP
df4FahJvxCfFHdlPTtLzTT6LbN9XOin3TCXceRY4JGKfRizB+Z/D/3xXwISq42Swlon0d9mQ5kw0
xJ+VS+GqTjAJA12JdRToBc5+ncbTonjaiPm6RwyupREHH1SZSpROJ2uXa949lS8z9OaM0qg76kH3
wdV1NrvPWwNZeWGaL5UXTtFiBHJO665QcqEr19XupUXtxPw9BWLvpOhLU84usfz8DFxVxDAnKQuS
T7Kdg6Wsz0rZCDfIGMiqfILjTmnVb1YI9NcUmiZryRHAMtVUnPh8c/b8y3FxrVbqFULE1Qkx0ssb
cx7mbfT85kIj8NW9KAjjadTw8ZT/8KQOhD8FzSfgJ+neXo36kgam2OnaH4Vo+F3IecB3m6alzVA1
kpU/o3v4pIV1MMfHY2hAuOcU0orNcD+b5ewCTcsK5SJIE6/zMU6+aGxiw/lXQzWSpGv3TNZu+gSU
jhX1ilEj53sxpRasg5JuRjue7zn2nRrK12+nvx8w2ZKMJuQf18HdDlvKuT4nDxey3UhSZ2HDqw+g
LqEDZGdFitqtrFEjKaAGQFz1sm3P+CXbD9hGYDiBcuxadHvd21utlyzsqmu34zmdtqrMEH1FFKm4
RTEIscLzBbAQ3Wxx36tLI8kP7f3s1+noa4aSz4rDFpT8tsuvUMI/EoHmTjbd90wJQOJFputGZNs3
ZEX6FekG/S96MLmHKG4XHuWK2R/L9cJVIiktes6je0KzJ6ohVXq+7IkYuStrMAV2aVFdNCJzy8sr
Ed9y+tmCWlEQElo9KcbZbYH47DTTvmUF+y7JpOBBrq9iMzDFM4290Bnp0SXaWpiMLv2NmZgsE87n
qOvx9mEhq8vUG+B0+sjVPbwMUXJuvpXxJvwV4Hnoc/LKNThGf79NsF9dMGgY8ujuM7xbdLrhIJCX
48z7Dzpl8n4gymMDZegSmyeOjySgCRbheNCMEl2zJ8zH7verEdTADj97iL67sd3Q/CPujSsDO5cW
uyK+an85l9NXEjRa82BljmHiJClSyZcACJcVqBZay1R9FeAHIkjd7R2rTNrL4m0phyLJBCGA6SI5
aNbk7zDazG50r1+u5o/O1grNYm7DZeZAox5rdMO+VU1crpFAXfxzzmLvCzuBLSttm205I32Vor6Y
KVW4xO9HPrdw13pL/iN8DB5ZUH3KAAetAnUJdgauEnTYo8Ot2I4hZ2PMsnXKvB4anyX8oEsh4v1l
diyL5sQEzfabmtCMf27jUJE630yFgks1OYCRkG6f5QkE7FYkffddJUBCNpzycfICZ5oBHJzwkVk8
HEj/2VSpJyOT9YaCDNswFEeZTS49dDBqpZRQg41g4fcyJ/quPnlcTUPv01kvCIDY4j0HOV6iPvzo
FC8cd2hqB/4eAqU8VRqOB13T8AU1v7AJZpvGBIvcy8e/rg03kEjk4+AtAfFlIMFuc0PvhLCHM/CO
CFbH47XZCuX08hV6U+Ua1W1NmYm/5zST96bKhfL+k57p3gSCOjzryt4Q6CsPuDvxDByO09NHZXVc
aGs4bFgSLnuhxBZnSknwm4gvq36wex0e4szZZiHsbJeyj0eKtcpb2XJrkttaN7IhFirjcwDbKDqw
t2vR5kYhCzVmVnxbKNasP95HrpwQMf/RvC9oZL0apg3zyjKOu9HuE2hl6eZK0An2rgXeeHtEfp9K
2K22CAAchDZ8IBwTIRswEdrbyHLg51+pVqJVi7eRc1OF3QSJGG2Ek6WjeeAh+T6hBEK5s6Sl20RA
mX+/+IOgqTQHei09A8Vpw31eM87p8yvWl1vmelkQrgJrmroFR5KLQhURMPcR9Mm3KpEqwmUcYwhs
bukLI+c9YaOcnBLelcArFuuC2DIhZZIeTpNnIebW3ClqGHXDlx4OPgol5DETQyqLpMxK3s18pBwj
jFhBPzW6739E4uBlPPWEHN84L9+hnBrFxWGRmmsm+o5ELJCFsojFvJ9KnuzxJJIrhFcaYiK5BXdY
pq4yK6phH8j4esH2nxDceT3REMn1hJ1tisvRvve4Qpi6iFfP/+8hSne8caa08+gaerMXpCFcxK82
jpAuNr+eE00SR1wAFqw/H4lE+zC+TAvZMsKX8mfVPDzym0l3piSnH7UORs5NVLiMW+EEoBFdLV8K
/6x7PnVwRcumtj61LqDZf92TY7xA8mXX7BwWvPzx18nwRU01fRkVRQFDPlgBHFXGi4FhWf8BD4Ba
mU6eKcWaYC5500o9Ut3X2h1ZY5Bs3vFGMi4patqtKGNiUnwI46J5BHRNd3bB2l339D9Sn6eU4xTZ
fhTreFbCGOflitC4Vs4qJYU6edrF1rJHmaRzkL5jcKeJT/lW3Q5E2tpjKDI5DTFNYEeWDRvAdOpQ
aVQMYui60VmmO+EhU1lcyskNQpwMiYPakHwanctkPKvO48rK2E/s/0ZM51mffFks+/lC7obcSGU7
c73kfsoJrGND9FjX8eOHZZmH71gnTG+VzjccXm4Yx9C4E0V1mf7PH5EjnV5KwnNUdTUVwtcPmRap
+3BWyAnrQBNQsWIISiQHfhSAYwIfdkg4+KHdtL+DB79eDPH61FubfEE/SvSYKLPXTc1Yl0TDdcKN
65IsnXNRwOK1F6z+KPW1g+61z+Xl4Mp9Sxa+OryeR/puWD8Rx3ayVFPLDHa85iHr9J2kJL6qIuom
ZemJ5UHpIzrSEPgyD/88EqcHpdTR1bCQ1HoS/xa6Q1vQ4rVHvUyvRZ6yMQKg12z/FQohnVxBsm03
BiGvyKBJxlmhi8qNDlZ8D83D93jHR4b2PiClBQ9nlOiUQ2VngpfDGLAs1qHxajrAzcu8/+Z/Y/BR
B94R9fAmPkkSXZZhUdttGb1FjEOi3zF5KGnPiP0RZFQGI2GVWp5FWBPRoXLpRQPwdeuK08DkpruD
F5qvPM0+yHxstin6phYlSRVMB2MNHGFnApjocRoO7h7O0f2LFoW8y/Mxf37+8cflS7fL7pMx59m+
80akSXexf5tf95pCMQRTx23b74bsti5nUtpQDzg6YVn280fLNqvPojXPgih9FlLcDaLmWJ8FG5Fa
qrMhyvBKini9PAF3+2w83NSP+jb6HVrnmq8eUsjHxHSn5POIDo9EP1llEI/cEzW3V+OQumamVZ9N
1y5u99Ie6bRK1oPfCLxNEMH62fFnGKHENFtXRUmJqw7I6nEwkfernaJw1BxRQT520eb+7iM49fZ3
kQMrAhm1MlF6xT/TJao4TIYiNaEutg5obSh+WRfBgepA8LC4EzBkXLJ6Y0+XztaO3MHUSGLSvVH4
oICeeZAdYapO595MY+KVHax+PZvMY59TOeQrLgMbb0TCUIjwEq6gPUYMG/6npNrwJwfcIHPQslRb
Sc4Id+OCcn/UebNoRpqTlEYOjVuXA2Eiy6y2nyl5Ys9qV4mcketPQBoE3AHhgoNC6ZSJG0JvVyrF
yajx1WYC7Oc8/jbatENQBCtyk+pkvEgqLO0CrjNK35H7bTo56g75/GAN2omXUYxTr62O6HdwtK7D
XkXQ2NV0q057fh6DPJNkEGfe44t7U4SjZqBwpG8tGguAWHACRKSK4FLUfGAChyinIhlK0+9wzQU6
PPYF2wEwHhemFnRoH0N+QqTo9VyOD6LsTa2y64BUP9B5874WDIKDc/kkFMAK7fMxk1nndyQQUOCL
Q4Klm4/aydRv/6AQ4Fx/UajiZYY23CcIivStFEQP4pZTQPxyEIc3tqKLAYLvXwY7m9DwmIpwMpjh
k+DfB4I0o0d/BPxWxGQpPbwl6Ufgn+QIzxtp2izf6MYxpRC6kntn1ZFtZ+OLFBs8zQPVot18CyTf
H4ZLH5gUeqdhQhdqxPZDSFHi8SsoCkUM5Oi78bOE7zLtVZigTG2s+p/VdTOhmSt8p47/rGv6QQ94
yWczbr9WODQMH3m9eurr6ANgH24sCW279FVIkOJo3dRu+1VkszRcsQvUDPVBwikZvmt29aLMovDc
1qCs17vZORqZDWOG1A7URLD+mw1sRwtCaAlixSgA75Y5xp0D13XowVSDXwS/+KBt3QBaD4vbEPd+
uVl3UzVBbr3LhmEjpv7E58Jgz2B4qlBFLA8zFQZiF1jJqrMWEd6Ybsg9fkQg99KHcfOJQ9b1+3F9
miAYygUAGaGo1ZvQoFDqjycVDx9gtlgEfUbHYFw4A+zZgLfbC7kO+U590GYH5o8tYRRGr9Ttrzvh
J8lyPKS/tEUSWpVWPV5v9qCPsSFMtjNNDlzxG17FEMonTr4XqbGW8wweAroAshqNM7Y97G/M/t1M
xMVqrC0u1nw4nJxGgQeF2GX9U0Bd2oyvBYaS04G0zV8RkPdUXH2QNo5XH2XzQUxYSBdvs25JW2Ab
oI/HONiLZWxL+7V4xRVrIqIPNUT3P8LZ2j7FV7bM9UOhmpyOpetGOwq9M5ozqJ0KbjkjECIc9Vcf
Gxf4EwZntAkuLn7dsbk8161PHBkt62+RLcbo6VTCOjdvk54RWsDGjk+3FAYrTPugV91WtLsWMc+B
3Isut779CdBobhRlivRN1kq9oEs/1oaYo6nDkAKth4cNklqc9ZFaBoLnqZPql7UvvfPifaPOF28W
5qSpyHthl9uZ9wjwRHahkF2iwtwNxmHPlduaEfLj+JFSSpzVcmEaByonha7gqaQoBwne+xAf7bwr
ti6+atIBnDtwHMKsH/bkSli/meSFndw9AkjK+LWwO0+JonuhyT6lAHS3eWwfpltnRSot7UFjZDQI
IFJNEIAybh/mUdcAqI30ry3EQYHaa4OfkHXIZJitpuZBsoOKZwd+YsXQAamqwFN4Ke0PM3v79Yhu
i8ug0Hl8En1GMcRcSclxEWoNRqIVP/h6QK2wQIHnkihDx7pyyCm34hcwGxOK4V04n5x06aocbx6w
RRjMJDWRBDwYdzVHn3+iZAFcKkCVe7tMAQ6/8yMAoSEiKksfOsgXWWMgyxUbaaYfSq328vP7CQZU
Cvc/XplyhlKz0D9h+Az+0yLyurR91BgAIK7k5IYijPEyI+qOSuBv/vXs248vGB0v2k1fi9cJLPwF
CYt2vLbC7P/Sp+ObmSFVIUOM5VBkHu3YNrJA+z1CJqFb3ZltoMq1Lk0g2/BSALdr8TFa4iEnC6Yk
1Ujgo0B8QTcsai1RBbKkLHZHnrBvx0bqu2B+hmA86EEY576ZZeQHn/gK+sdoTvIqwqApVdBZgCD7
R6HFw5BrY2j7vLlXJeuyeuEhTL1luggWt/MmhPumYObEdSMpWxCEIxusWcx3IG8oxHDvJKE90UDx
9eeUae/kJQW5KJicKNZC7XIQ1mVo4Sy4QKu1hZpu4CgvVcyedTK2gqQwQw9TkztIqYqWGnGVanOk
7C4E3VjxjNSeiBXK8BLFK5e+MP9upiryPKKZDFvFnI9wSP4fO7gDY4KtPEiCHmw/wZCFI0j2wODB
U5aMfg7LkpMM7AnhhIZLbT3umkUukMxxFmXMkxl01eaMd+3p++b2Ne8jdW/Nj9jrw4e98GJt01Sg
5I+PlKiIDPF/tzslzS8lsEwPHK1gV6xKdqNT9LSLm/JgqduOUE4g+BAF43XYlApaw2eh78HSiGh1
HvaWLc1Q9F01r/K1xRoMijMMWK190+kiSJOX6CPU5tw8rDzz0uKdUr7lh8spx/Bv7mGDMZ7nsrKX
c7fhGKbjO1tS0JLEdro/2pTcEC7oeJ0/H1QDTcTgHSJHtYIXygQBw8y16yTt2yJD/oIi4X3v9UGP
1+zchEwVgvSgLCg8eRbksjk49e6Bm81cHyETMZSnAG12Cu6Mf3RW36NgPlCJ3DYH12g6gogObqIL
bUewLm2rG3Hecmw27VU5DLtTRu4MOSQXHpQA6VOhJiwcKyVpr+VGD0bdYD8eQ1sMxznwO5N/U9pv
+SOQ8w4QSCktkCvHnkpFzHazNDMuAUXBjET0HpQRJXKJP/CAVYSPhLNpDMdBgTk4x6zirnRDeztW
HM03GiGgNmwep3JRCzBGqPuWiNvCEeBMfNVAV6rTY0lz7DuBgWUoyxwTjK0rtsBbpdxey6u+d03G
74nD2WKpfkP9GmBi7VzBtO9TQeEHl0aYpvSmhI1UToRhEBlSrqGR1akO2ytpeMkDclS7+aq+vkQ0
DEjjzeDwyR3cwEp9pgohZavxsjlkn/z+qOZoi+eP7+tANhm5GNihEmLG4DNtPI0BXO7pqD+WYe0a
KTCi5tMItpigKIYtFhr4KdO5AJCxQIN90Xew+qEi8M1dP/tzYDD0NWYDR49EYS54lF8fXOFh06BY
RQ+e6s8sAr7kiUAHtf79kXLITcHrtl8lEJ0zje+Ig/7WWqwD9W1ZQFSs5jAYCeeVs5PRWSkjPbgb
IAdh1BMUwUdVEUjaLVCnTPKhEzemSj3E49cSfOM6sIiHIyknKzlJJobGn10Odj4RLgUvgmbZgZTY
eKRQbQteI9TXUJMoWGNQlInDyt9VLuJyhgyWbLfnL6R0PBJ9uQBBpbZEFkiTINOOHSISl/+VlxZE
gfXYKJdH0114kdtppgLH0lgZaev4jfxnlVe7g5yqzuZO0ZPIxGDO+RmCP92VKuYPORQ5ZlJdwdQH
wNAZuZ3ekHR/69nAONAyZtalAGE3Ups6udN7F9H9XjU8OQKdJPUm0G5jhYk55YxRyt1/jLyg5fom
zvaVd9lltaD4PcSIc2DHA8xf2yq7vt+KyacaVTqe7LSSTyPow8blRIld+CW4YFbz9XaaZCLFk4bT
t2LioNECYNtNqQpPeWDRkeiSH+AUQrMh7qOGY6i6p1REOihaBpyopf/CM4hYyOiJkcsQIjBFJGZD
HiXER49PesTQIo64ddFHD1WzGu4AaQFb284wkuNxFlmSGdWjV/wbyqUYXEsB8/yZeAZcIDT7l/PD
3BPQrvKg2ctd0UBM/9itV6bqwnaP86uA9NbdomstP00gCIQaYxpe5HXpupBad1EEpsfJP1Sq+R7z
k8OOOcJvoRu1tt8xEM+4wy7HaSqmZbRMJ91czHjMhxAhTYJntxCbZEOk/n0xj8bazTTmeuYxDzcj
1nL5dMt33biZ5IVev09WrqziIImCJnXNYZd7SdrLKiBLr+J+bVO4wGjW217wWew5E/uyoy2uqZgk
rRIFLKnnU9c7E2XSd09A8o9rr6Cn+L0pXLTb7KrT0uz1YytKy338QNv78CYLaR31qc3dnLoDPLKa
VOy7CmCw3ZdHy6VXTc0GA27y9sgZAjRIjQ+mi31NJzsKhR22FMeFmuqAXvo0eZm1Ca7TwcvGxZJr
44H74VFJfZKQY3x9zDgcKaY5v9GUyYZpqf88WBCemAocBSq1xe7G7CYv7vQs7aZfigP0MBVlqhrC
C9/Bd4Fpaz1AQF2XgZuU0xwbyiK0hhRdb/SOOk2gH6K3zO7/DtFMUTvxme4rqsXMItF4/JfAQIEC
S7+INvMcuL1takGxgZy8tcg6upfRjGA2UkO2Kj/72P761yYj4xy9CACsXxs4nNwPYf7R9CdqbU3a
NUxWaVJGnroX+Ak2cPYMtasgAkHzDlDd/HTQq8U4i5QyV5US7I6NMuPTYT3n3T24s9VJjhs3THl/
yvlX+EqI2QgyUc6/Q7NYN2ShBc48X9XMwP8YK7gvMP4abjNPz8+5oxrwG/cnTcxL5D/tf7cxVJBP
aykIteozMNzaEkbKsM4Qb3o8gQWDc+6piuc21xnKUoNr9BWpR6BRit3SvdJwqpqX7WAAP1/wBUsb
pxGjyYwP7GtajbIlIwXnFvk8fl3sqfxUlXhkoKNHd1gDC6ukrjzAZH2hLVaOqe4tzUZD48JZk4wI
9Fd1cVF2DqI7QID3inEphFOMQpDCkFsF6fD0nE3F4fz7+ZiF15bwz7ZQFdE0MwSKcYxidfxGaxXb
W1jcqp931qVSu+zI9kPNYGu3h/elnKV7PYgNmCxFLx9AX+9chJ9Ak/fv/PXlFMBJtKCTEukk7tXp
U0RNNGTv5ZxUIpV+KHuGAcO7V/aiadHv4tcO0xKV2AZHydtXun0KJvkLVVPoGCMUSWQJduxwh+op
btNsH8U2pvNEBdrOWk+Ig72DTQC4Bf639SF93eJfwhK9QuNP+h2N4ZFhFPiVsVbJVNHH1rOM+4KY
dgZHJ2+Gd2o4duEZUD6KVM7bVb8DHS4lGFjUX/4j7FadyeIB5Mhrsm8rppuG3UTNiIowTv9Fgm0/
1XxQ7GTNVNpex0lvc8HsX63iq5TeFxte5D8H8Jmh/uZq+RrintbLX+2F+dxA97s6IHKC2uwLZgvN
vL9aer9T0wtd6KBfGWDR2dQU5ERxuEEjIeUxSHB2Pu245Azjw0dKzUf3s/u85ZPmj4EHxgznuBVB
jLIkB6RZLlgnC73Ib9ibV+8pdwtmfV8cTsHH7e/7D152iydiSIbYw4siTCpCQte6/o2/lH5FPCll
CZv7rIAlKsiwwbQxf4BuGi8SiYSUIwCRzvItRbb5WFtKdjj36PMWvt1sUpsKgQtBTDJISS2zQH36
3PgorM1jqfq4jdLtL+Y3AHOZWtMx0hb3ozEUEU24s+7Zz4FuxE4/oxkv4ydp/OcC6pGZww3nqEgf
DoKcMQdiN757eLdiZij13u89jTI+txnEhHhST/WgTtkZIzffL2zW1QBBc83QLczC/ubb6dOz9VGv
Y8MPQp+2ENQvCo/JTg84APXWUyh1BjdUm8NGDrI0+SDBn72wwg8/vzUk8mof76yYPc6tmLCjoszw
X1yIlDAMqyDcqydZnr2PC3xslPZo2nYbay24L5Tfu3yQHgVNk7hn7RT8DeVDi5sCnjxPit5nNMtH
iS3U/2I/X3qVBuLo5CwpAjTznSx23qWEzMgVOmNPaufKzldHLngt/imM3TOKZOkvvF4Qy1+ndNd6
qmWXxjnf9i/Dv9IpcfHErWaEG3EqGVxp/6tM9u0uuY14HLau90WbpQzFisNjQcngRsTxMuM6VWOD
CEZH8Nn301nb4zyQMNOXC05J5yATx544AbIVrw6WUIbfiHW8uI+o1E46NYtvye/AzKG5Xee2iuCI
VyNgM3YE7bWYPq7PR9KxJHGIlhWiy6x+OsO/mDncM0kCqH7twD7LoBVOYwrAxYMZ9aOr5JpX1uI2
FgrXRDDP6rblTi6CroaO36tG3bkRMm2e3vY8GvEMqXuWEOng/jBDci6l3ZpmBHTKyRzIQ5Nt7JMC
z7aKHbzYzd4+XoscuuIBzPo2E/hSrFs44sxdjTH+qO797eLg+D0bV/ei9Zjqd/Xujh1d9bx69Shi
38mPb2FwsFZZ848Vi+dt7WXMRKzoE2g1256xOPCeRH69GW15XbPtt4WVG2yAPQ4zUoGO0WslgF8v
1WybX6kRt6KjbV7ZpoEwz3yG5oOmQ/zwICuWWlqYix77Wx54rYaNBHxj9/fU4Z+LomyrVLV5sZ8N
Ro8xlTmHuJFHAZ3c/ihA8vlQ9qyMIsSO+jtJSfM3kpbmUZ0OK94HJ2JNoRV0LcJ6yJOR5VU5Ropk
Mjme9FH6WTLoNugE1TU0uI0D8a4qIXEbtF5ouiDR5Suw083Aop5bguBv69H8ouy2vFKnwi1RY+s+
BYpJGcQ5i6FY+2+1IINnPKqBPrAB1VjO946QbRSj//AiO8zKUWATRjCr5EFr5DaDEhs4VnsdnU0a
uLGd7g0cL8zj3nrvgCq/5VDP8sNGiRgdwU0JJ/rJYfzI90J1EBCwVQo7CCGYFIdMIuFkgOCMDYVN
DmxsQAUeAhLMglmAA7p93PB+AhV86sI40VnJjFmc9Lnj4GTYM4d3h/97kafVTnLA/tz4Oy4t5Z3n
2Ofa19S/rcGsBlk1FfefVllYHZtPj5lLtStv23r4ahGCOxlZGHJcXw3yRPOvyjOzHWCcRwXSqk3F
27Ch7gUE2FjdBfltlGd7P4lVS4YV1WDCNKishDGAyT1M8TXaiu3LWobSU3TPdOPYq6s2kjVPYG7K
n9sYibX9M9AZyOTwhlAmazm9UuALqnI7gyO07T5Z1M3/rza9u+8H3N0K1/LqeJ0wJflfjtcDyAHQ
QAvElpfXPyjBqC6yAJyQ7GNwWzFAlyzxACH/CcQGirCy+lJnTDWH7WRBty2n3G5rWR/4AOw0bL3+
yqrEElrtdmBMv+lSbEbQaCIPd9Jq5hD8V1BBZiDOU3tkCcUt3U1bNBeHxdnXcjPVldHKXWKvkGfm
7Xwa8Xg6AMGdH0UJt3KPWdN3iUJQXEfmn+adh75MkjLLASFHrZMBUw6QQ+NwRl1o07ERQFesh5vT
Ct0Aqwk74BTGXcCjg3DH8Kj8UhQRr0DmQaVkiPEqBqJAIJzPrYqJJs+e+5Ic7J7ZnFpK2cFtGeJZ
BYc65OgLlhE4QF81H4OdcpmSaAiSvESWoii/Y+sPmGVkBIJA5Vnf+0s7nqLsBMg8BgBeVqMuKftp
ENk49zv2cwS7QYdmz5VK/acib9YTC9gb3A0qbCxrAh7EIXp46eoyyBV6Lv7eyCrQ524FZK8T3mQX
wolP3cvSg2r6a6NCXed6Pch5iZbwwNts5cqedZERpjJNTwnwXvjodW+8y/emneRdqfKWPyjl81f5
pekJX740Xaol2AEJ0vhfkzYqvXa9cOdzTMynvW3dNE5lITD7bw94vNKr6d0zlfVlIThC0k0vjHOc
5m4fRm1hUtT9NXfkgN5uqgfSRQuvPVOORpQlGfhIDst9oQsY9kB4IelKPDX3qGEKUQRgEnETm2Ot
KZfTZJdL9GtmCo/SnSl/dwzpcCXGlOMGRwu39+3GeuLiPTjO1kLIm7/OdNqzgH1mfECqMeIP9qEG
dDfn9PRaUDPqNy6GsZY2iGPyX1axuepQ57PBtrOyLzMagHZsl1UUr7y4usoJwzfeBts9KpKSHNWR
sqxqMoAEXUX7CZ911e1ZokSq8OJBW0Sz2HEqJucEgV4V8EW0eMUqc5vNgrt+NDFAlHG2uWbsexz2
A+U1vrgpuFb/aA9xAk4efJoT1/h061jAZmWGUh93l6p0mc0wyhQH2zNxqbIamkWhl0Y5C2/Zs2yV
2/igY9um2odE2NQ+K38w8RbVdVVG1cHQGz+lOC2PsO/hZFx5SBg1UVxEKkhzrQkG7o/CbSaPMJ57
O+ywel/RiVbL3S/nE7H7SQKIjuHtv3Rtd0LXdHhPKoAfirr8mfpnAhfzKrYVVTW1QHSVxYwv/XOM
Vhh431dM8C0Dt1cFzqYms7wO8r3cxBKdtxqmSXURUw4eZhrJ4S9aNL66MJwoy9AfzbDxwYGgKUa9
AzzvioOx7fYDNMVThs97FethHY0JEFFlclSJ299rXa4yUFQ1/7Z+ycfiGyENzErIhJpTpBf3Ntcc
IKYDXZzwyW4upBSmJVc4FdHMqT85DTZKGE5IMWnyVmZNjEYUrrergR7dsGzCW6kGfnJfE7t3sJ/t
s0XtvrQufz9A7ODZCRSdz4H8AMl5Mv+yMYmKvY70E9QzcxXUlTahAQzLQNO3R3rLHtt8fFSyOcoc
x//Og2rkZcqec71MpT7FSoMfutKdjIW/7HZhDIN8pxvTY/VDMWPmfFyw9304t0rEqwdbge4RfqT5
6jlsZhwAvxP7Gfq83t5bzRkRW+wjB40eoFq/hbaFWg+kQo4l+tOsjUxnik5gjF5IlDtQ0wKSaVB5
8d27lQpTY62mtCrnyC1c//74fu02DcE8mD2ugLsdnmVokmYRu5Gg59x1S+WxPNl0ZHENlo1v1ZGM
ZwAAHnBDgHupoy0CuwyZjZUa4i4xSfeyZUlUbAHv1qaemfwiC5WO64sJgqXHmdD2FGJBieukGX96
gqICS1CZNj7IroVNIyq37vNsXQVb/68eiPcRpBW0UDS2za8Yz+CfszTiRZRdhIYHbBan9WQIElaM
qDTen2gwBFHSQOuWgbG1cNusM83NKx67ZS40AXU1m7x51xAM1GSrGR5hSVyxokH7RV8onK85TquG
fBJctqw98TbDrcrL06arhQXqFLCq2zDoXP5d57k19R86G/AJEMsZwgwmoZpEb0GFyKaOaCeUM3iu
QF8rXUlbI6uDURITilhyKrh1N+qABR+w5WYD5d0+X1EBuk3UG8uo5Uhuky5dDALbkaAsTjYNa5jc
IbxYnwfp8rb+9gRxcbxLl1G1gZE3AYBLwkV7OwFHwBWZQSZfku5IKqkLXCKQI+wm5Lh8G+2Mo5/d
7w6NM5cSn8JzdztcRPbhXCmDzlab8mCHUlnu8Mx1mBbfpQO9h0h5hT1IkLDQVYDJzKxJpYHFJVkb
qVs//IFYU8ykuROz35ICsKn14foNZ2Qw5VYaQifhfs72U0RbeljYIZm6mg0btKi1CtTGL8Y86ZLY
dEZ50dwyjZbj071A7t+EbfrEMZE65x0ghVFq3Cmkf6jV7Ip8LaSt4TK0BLZSemzCzrdAOocMm2Eb
MZRb+6zL0E7ZNsHzqCo21La1Kvoby+zrnwr6AqngR5Rt5ziGfpoaTGH4xb/y+NhWES0N/CNS6ZOy
+NmV9kRXm1a9MOGMYk9efMBy0p23R8ci5Ub9b6GxSVeqczjAKeNfP3E+TPCjCqMCVbv77PD1Brr3
H4Gd5VJ5a62LozsJjMFSsgXfQ/jW0zSaiu6ld31nLD8fjVZH4DJM9EAdwsghv8tSNTnStMgL/8bk
7JCuzcLx+kMkoAQzpctqlWWLAvMM71Q1m2QQtEHhpyTFMTgBZ2cAZUdijlkC0T4Wg7UFQ3U/26K1
0+IUJbiYxI9ZcN+N+4ii9Tzk96KW+FclG4vDEOO4GmIGYG9MmOelrzX4Dk5BXYKd6gsI7sNm09xu
v36vSwr0YaLdjzwBboX18jzgFl3++huQ91GUIa9PjBKZfYuNi4MrX41dzL7CxrBpr2Csszth9HnZ
X2Bc2kVfuHBQhNRyLiYEEeEzDx1usIfptIkl6SKF2Bdm9aUTdkmdbJFRsKGRBla2m4oPxvh0Sk+i
GD95Mg1S/+PEFIFGzhjIJoE47eWgurV9Qh17RZe0Z5CmyDpC6hf2mqWuoSPudiOorJUiIITHueI0
vnKynkJpawfObC9hft9s+e4AjPTknmg2XPzGqWPtiK8GuWuRgSTf6KCDi4MSnxNBG536DvCad+Ot
A4ulnu27DIJXs3DMJ4Db0wJ1dUlIQ6mDglUk7oKSAYLiAVlPe07VYnBDHZvB37QCK3PKYqZIOV82
sL29olsUSYRN9TJ5F6zxpwEwfoEoHmMWTeMNcQXalHc7NNtV7s+1PH6zNP6LtDg34VVVLzGUDD3d
Kr6EDxiQlFAgq0OEHW3y3C7wqBRXh7rsuoqHD7PpD7Gdi/L0OuqPY+LeGTHTWvWqPUBCktnliaxa
p47m4ChxSr6E57l7glqCEVlRbLC+fzUHzQCCaqOwy98DRBaVcMHHSi7IaEiRn4jdnOnHmLi1s+Wd
KVSE6jRN1pJhIDmKUAoIGjh8mn7z5eRJNQQUU9bj5J8OPvEKmXDxWy9DTRMXGZT1YIWYJhPE/NBK
c+1GoqEVh9O9P+c/7BajVmblq0BZEVFVPAPHu3HDppCeCHCAmNB8EfFGxCT2RiZRr3VYCZRHd++6
uex+ziPAAbkv9qUjkQA+nfx4gNeWhyjEwl6s28+yWgZVzhis3ADd0PWR20Z1Ili7EJZd6e2mGsCT
wpMQ76rXHmUoPrz/nVcCsg8ilisA/PKPG32SeFzcO/wl3YiiGBkpim0wA2H5p9KohlMTCFulz4FP
I+vbZPW22NMaP+8UsIwXFcpoA9wFn69zQ1yKFwDhuL4FrVjdzzgRf+JjVpAlfTUAcZSOJuEOK+ft
Jr7oPDn4RafDxvjfkvExjGXfjT39XaXbpQ5UYorYtxZ+PoR+TfAYrW4+XLvKKIBz0JwHnEraNIzf
DBCRkYNMQXPX1QuH6elUdekKmov4wnFVuPXKIih2duqmXZK6sL5NQSJKSobqdZWFI9LLca713HNp
v9bFbo1b0A/GH/plTS8V/7FJNNP1JelqDCVDXLRfWpmBy4jKGTWRo7i+OOx1/88WiOX1szVR1m07
jO5goNTWyly7F18YG1qeKY+GefxlhkEBSwz6Y/hMbEHaQaruQXSe52C7a1QiiHx70j3D3UI570IW
ail/KRQyiDrX3z3fRDG9m718J74OUHxJzYnWmUr0/8dCpayDfupw5ejgMt2bWsbbJrIxgcP4HqFB
QKqvi6sW4v+OjSFDm3HD6nZ2+2f8AHQbMqFsVRwunMxK8vdQ7+6cutm74uCbOylq0VJ7zP90xVNv
xwjQCdM2YbgL8jNrmceBYt/7q9v2RPMi5OKH/6SFzofdTGEXsBgGn7gAZ+FzxRpSr8MSyXq6dcTi
xjtkF8oPxJFpfefBHpoTYRJVi3jclasEvPmR/+IJ31I4Qu0y5icSqDN/jFYgNoG6IqJfLC3uAgzP
MqQ0OPWcJiG9dqItqaNMtuhv4AxZqr60Hx1exgr97PwBFQteCqp35fevoURN0Ia3mF5uq/6sdSF9
m70pBdws1qMjKWk1bkKE5YI5/4ZXLFG5dwfPOyhp4LmqRVzi7Osq5N7kcPZqA3XGyV75OUuN6UEO
fYYEbk5MvlMQ+HRjljPiHtJp+ci9+ndvcAq9HG9ZyYtxBR/KIgwXwKtu/PNhvar1USxv1L9TmBcx
holNsV03O+qY+nODUXoi9vBFZih5jL+UnkFAb4UzeHYgwNdVCacuD+0mcNZomGH0CGKeamIb3lDR
qgyUORoTiu8Gk05u2oQL9rIExGsm3l+vSw8FjdwRoAbQczeGxs4uPjP+PZz5SOeg36sUwyxGDFUA
OY2q0Z0+ZE86iY+ijkub7idpr7X+ETMGMvtfZdwciwZlNlNVdO3++I1V9C7Ex2zjYsMsUZdBAG2F
zmzTy7wdD7D4URwZhO+wXm/cV/+Atr6U6/u79hEUxXbRuLK33GfEK1OmIF0xQ8I7Bbo+pnvcrRf+
miGHAxKcgUWSMrUsJbK4EuBqVA8q1mXu2SZwwpg6rOLxerIUt/TJ12SgNpvk1HrGd762Yu+3q3OJ
+XTFJ1vZ4BXs40+rcrXKitw2oZpGVSaGZYSb6W3GCFpryiwjpzNFaOFGatDF1H/qLKZh4tiSMHhI
SaNMw0fP670EmecBTc3ntyfGXDbV0lQ3/PQfz2Q4AiH+in4SO54KRREzD6ezp6mS5bbUYqLF5Rsq
T0e4ODSipbfkkKMe1amOr2FSZRl8p9A9NoO8ikXWNsFsBiCZZlOSP3bPe/seqbi7XXK5QRGFmriI
/YZF5aK3YsDupV+EL/uXElWkzAvQEWzm7pi6V6BMQM3L60TRNO+CVUcs+dJZMwENkT5dgjByeA9d
U3WvHNm7+5ol/9TVZWieIyfGoFCTd9AU04fysiyb3fmpz0hQpWoAGcicIZ5Kk9XMMFCyFdLnMCee
G85QIrFVsMkfCLq6ZUiW+ZErUG7mDqdJ5Krvt6asWZzcNRVsaZ+yDHMc9N6h5ro8G0xoxKtPlhKU
4daidYjfRHgKlwfhqo2FNDSLLxi+FWTUZWCgFjeqNIFXB7C9dm7szZbG8QL6kOZ4AjU1On1xIkdL
DOaH6jX+NvE99/yhIuoDmGbJOjJnJe8oChXyV5l01gmd/BvAo0awqiMlSsXDdH4SfoeoA3E1/4kG
xJ4Ocl9IYZlKAV59to3474tAHELw4XFTGT2+ZtvxQRDtGyBdzqVRaXIWxxM5ktZFfPHWGtv4TNrs
w3SGIM4FM5EcFT7KssDH7D9YdPlMbwHDlKRvi/Mf7dZZaElE1LJBib2RrrRE8iME/jhX+N7mBCUO
4nyZN5ZzHs8/lT6IyJLVBEeb/CdT2IN/bMrl0TmdmzsuH9nWhkT1uD/8AzRKOdJ10pLiZngIc/fU
yn4242DBjF82UN33PnKFjZzyzLWTq6c/gpodkWGZeXaRj9ycUl4RAYJYaOgHWfQhBc/j9wfbbPj5
9sZ876EQbihnS5dKYo/Frtli+DzOjwoGWhWPZAjWuSnS399wdAdWwhNOk4ym7FowoItg3EinCv0G
zYoME9DirNqXP2BCoZY62VHYaEY6aox+jLGZJTG3EboqKnooSX5cntWshKA/9T7kHlc1fYPNhaC0
MDmhist77EfcC9jH1thR1q+ckbyTaEaIsluIbwEB6Bhu0yJtCXX2qQByjTTS4KrDQDZJsxkC1c40
113nGJhiV88hcye2IHkn5Ob6sLgYiNpEWrg5tm7SCd+07x9YNI8UtF8IcioZrkU+pHSpVRCLtbQY
o0GMER9L9EcEwy9CNYd350rNwIMnSVtdpWt9QnIrieb4Ay0thIDyXyNmBxT96bBduSdwP9HVYuGq
cerrkG9d8w3K9O9gYVlaiVHML8eG1GL7WEZ7dxRLsA0irjkUl7b+AhOVvYFKCa+tfYG0tFsd/rod
8sWq2xAiX7YqnX3oW2j4+aF/Ji65Snvh+IUsNAe651taTCX+FEfHas+fbNrzZIjrKraEMDVhymgI
pL90I5MRqiNIDhGy02QX9aTAGkAMCrEb0b/j/ReX4ydeJr7RygAJB2LnQMNAe71DX6NFo13vHgAh
hW4nX+PO0+AXlnv93/hQCpOvrb+FIVihqPmkdMvMp+3ZUTkEiB0+bxZXFHw64l+GT4N+V+gtkHmw
IAtS48QtZxquM0vfRrcV6PjM04zSIK9Rry0XVNR1WjWqdwGgdmTPcsmGQZVQv1ofiBG0J+Hv3gn1
b8UqtLoOdRz1J6YbH+fmrZUj7p9WRBUcvI3bD5OWphcDKmH7WyAd9Ezg/n7aoA2EyjnGjPQYiUdU
sLbG5IzX8d4AGVxTjKGMKfmTioCMDaWq/09VUeIy+ApVxZU7KUT634bsrNif5iwB9rU+OrMrKrP+
rTlq9JZ+p2UB1BznWnyDSr3Q+A2LIJhiZzZn/PbZw/DBiUH3tnYq/AKsxGnQSQt29ebZtgFp6AsC
1ZeBC3lEQa6ZHAfnoiZeZJylykXjbPJhBYNKlScfPBl+jbGYJArFNcyNNvbkHqJ1VpfrMY/9LFvb
dlbWG5rMmUbwwdq2TP1UU6aK04cfaJ8AAStIkAJX4zDZda6LDh0CodaITp1mrZ4Fmwm47uHvizmR
jswkxTkRZN61STZXCDsqVRWBIvXyvoqkRwK3SFkyFn8cP2WRpHlEFIrNqSck4NN892rzUOGLS3kP
FQG8Ah0KOnPLo80tan2VHXB40SgZnJ7rgPrAAfae4fgvioUU19WPwhEjnLskcZcLTgKTjVc943AE
oz5BaW+dmZm4/rArWjnQTh7rqfb6jDPR6lUfZQRJ1ggFTQ3VPdc6c+NI/B/569nRab+qTcvOmbTY
ZrBvS0KGUc6I2IHVGNpXrCuPt7erGbeds0Mh3nfYwAKDY413k3pX+Vq6osBygDSCnheBhjgdXY/C
zLhz1Pl5vJgc0VjLFU7MoZgLavUumkxp9GESQYl9mKxWa0N5sbkDnOKcCXqLV9alwLQTJxURVBiG
1NIEsUJoKhfDLUwGX2VQrFP6+Vosb/4cAoSC8H0Oc5CQqkdQtwP6cBt+pgGj5bKncXxWsMpvrn8J
Xp0m4srD0kS+pEdHF7m5nZGJZOLpektImKA+Axl9YFetDxT76TOwWwJmuTW6nKnN/ImF9ulxpWaL
EmcJ8HFYsjbQs2a4ZeCvbODcgeI/xmstZH6o4suA7SKhopEb3hMUT4tmgvqFEsa8mdyjOzNff9TL
GtERioyNmrcFASK1pqv1Gz24HDo0EZLAVpMGVW1lXyFRzgAPrZ1MKalEdoYkSF1liH09yYkn1H3V
8yLzxmOXvuGGGdn3CCHhuV4PYHPceRGBLjJgvzSPnXP76Nmmyz0kN9sx4rk8h/IKbH8XlnF55NyO
NQlAy2tGACeb/uwY3egCm5s/0QpgKUuAm1/DZVsAQ6YLyN8fB7qnuE4WV/iHGtFN+H/2rXf7q+UU
gFt8IAxWAKvQd0938K9Wo65V9p3ssi7+8XWTXCKn34oP+eBBJ8z401KxJ745IsSl6aYbBXAbcvCt
kDq+f45l7Jx9dghEILtFh4fsJHBa+TeXsMeWIumpuFJWR6GPUeyjCOOYnzQk4Hzy4VMtUj0uTFM0
dYCjnkVHY4LCZHp7S5aAyeRguYQGRH3bvt7Ihbqd2fci9xbDlk13tsZZIvuhk6SBLMSTCAG2GMzT
ipHUkvUJ5yz1Sj6Caq9ZoM3my8YsIyisZP5wYH3TqFxDq9vs21cbJtLFG1urB0qJTkcS7AS3l7WV
Ns34UeheFLyicdujw3H2usd2z5BG/n6TOVeYDt7BNtKGUIjAzxJVwoe+ikUKpS0hu1vuZRFwPSdp
422bsYCi6BVqQkWPWGAzly1IdggYco4P5efW1uJfk3SGZ0uDc49ts8GXd/RqHWHQYVYg2YIbrKc5
SvyqrJT18QBJ19AjWeJzxKaVTGOOTCeBtHPYywrgebT9GwwSqQmcHjtDGo33WWAKUZaCsJqSjRZv
lnqWgDbImHlcpzk7n0HQXpTmJIyPSlpz4sCgbYr/iSoxVw0pmInMiYEP8phi0id1AVSr2pL4+9ju
v1zuHQ4TQbKBJpwaCsaa/bRtxwCnI2pHjKFRu1j8Ry/gtL4CEhCMCtwhxyESqQSjyshNUo+CYT0h
aa8BdXQBmYod8T7bKhRhcH6+nuQ5Z7siRiWr3JAVj6Ibbe4znZBeQbWQ+QadZj9hl007mDj+8hhk
NugpflejMOOjtMKIzasxf65K9LwgpXTbAeXo2xyVGygpzQuRzeLN9KbdoOE3OWGXe2xtBpGDpT3M
RSOjmy25zC1hwVvsGC1Q/I+f7uao5U9lq32cASF3+ED/r9DnrUUReDuUhjyqnXhYwsCw0ZK+NaD2
Pho+oNnCWpkb35IrmFSHdQXbO5RpuFnIK5rUOBIKPlA2Q+GoBew+3HbUIiuBBpNXVQrfcyzkQHpE
/gyeHa7gzNYt/D/sFBmJ0QEXot7fbfVtSFkaijt+tyKmM5AaHX4SWO0pz1uxwap44ZIexvvWCjS1
xR0wBs97NJc5oMqV/hgPGky8dX1YsF6LG/3cf2D3GFvcF5gGXm6KlKeg6C/fLHr1L3IAmbzupm7w
zG+1P1177WoUPrYN3Ra3zjDp/qRmHzguUk9IH2Oi25yrMpz3UdpV3RbYV7ge6DX7uI12K1qUVvE5
1XexipK7Rkq/F7yLM+MklQrhCDIiKHzUZtT15ooRBKQfP1Vac1EIr8iFISOZrjPLIrXzJ3yrg+q8
cqm7AYdkwFCz1qYfOzhVf0rH0mPJMubCeMJ4e/beGaN/gpRWttZe2UxNiXNtW34/o6tKOpt1sbms
pDsewzhBnUw1IDiiGYF6X2xBT3nkP6+CF9JAef7/q3yNt5yiE9kO8Nytw9H4rMxFa02ID0cGcVCI
Zj2Z9DPgM99FVUfVOu9rqIEp1Fx2roJ20rLa2WkdF+6Rq/AtQg4kFZYTzGuV5BIF92Lcl05APDKc
++FCW+08IKVpJGItWLtvQiq5/YuTDj1eQEmx8KMginW3+Y+Zb1GzEgGWXTwD4SVyD2ETMlPWPQdL
uH4wIl3NMwUwRYVpEsuGmw6WMfzt7lOUg6PqmYtmAkzz9UmNb6WCiTpKzd7j8I7M4yYZO++tjbJn
MlhbY9s+o8Es3Td1LEBJXrJgS0bce8USYvBASPCN3+4ItVC1f/DtzycU7HWymrfrX5Na9MXVTTqr
S/X8UG1BIzPAno+Bx6l5xXOOQEE518YO1uoaueSPZa+KIgo7zTPNSmt0orBbJx0Qvedz77pPSO55
BMS3AWd8y6VPbWXDlWI+sOmAMifsq9lMO5ltQaBgPhGVVvnWWZD2msoJRRBQTTn18ZO7O1kFhOdO
c5AbwP9pyLxs8+kEztra06ToWEIV4TZlvQ5R4xXly9uMWy/aV1azMu/0FJSNcib/xV9VP6k3gQuf
x1R1U8v8xsRZa9KA1WRh7nc50E7CSQgbjV1MibzWt14cThgwEmYyo3dPmstsnouJEIY+xd2sQ9MJ
UmsHm2C2GQVe5647D15UP4lBSxkXP47gQjeOPAJxyo44NhiXNSs+BYBnOxg6SbCYsIHyrkHinAf0
+CGpgCmVWs2mpYiESNzVsFwXbWUHLYMbGbpFsoOXTAsuIEzuGR1TeQVbdpKzs+lskJOHUSnUoQIi
rX811Kc/UQNorj0yj9TDISbafQZpz47qhhY18vr67fj0XE2vor7OScI0FekwEfh6G2pN/24Yo919
DLzhISkfAtjy8yi5zGS4i9q2qyDbpiKYskNnr8bh7hhS2bT0mYvyUlLXNp5hKxQYB47q3Cw8B+p/
RCy06s0sdFRTXBx+OiDsGx9guY9TfPV/xWPQvxXkIy0UCKklfK36/BuhijOVTG4HfJTCWse9HIp+
pMwCmh7nC5Id/xR02O0iG9wqtcxuSC4VXz1SoKGI8Xco4IMHDAKyyUczpPpQTD6mXqh/2w2GCWQS
3s1G9cZZj1aLvhlYG/EEnHmatIVYX2alMsdhvNHGhcT9GFebkhbOrBpYsyjmVLCP5ODcMY5uNQ3T
h9szujIWmcyjhqE5tZoU19LY3vPcf/4cPLn6iN4SeQZqduaBGteEBnGmaUnJi9oc+8++X5l6uWJo
to0F6633TwpMEaJG17/NenfVWGSYMfvEYMkXfhcOxhfQNC7HLRBI1/bV5ca5AIjLK+Lm5s5Q4tv8
HJJU831tMeXtZMfI5NTwR9BUFaa12Qkr8bybSvJxap+UGB6aAErf2mRjwJo7dOQ5eDkRZelURR7W
B5y1VZ2GrS9X15+1GBwVdrRE0yTpElQqpmBWobXdXj4G1Yd4r7/fqnsHjpUZNqrvpmAC8oiK8eGk
V1yhaxzHLfMMf6vvkXL1fJOrHt2ydFZS9C5Jcb97lMIbA1d+CEzYgRmv5Bn3W3bmX7zCP98lr0Sg
QrHmIAacoz7+fhuYFTmjNnLVZdpzDNdTOsU8Q4kcR2qdQ9y17vOqwXfCQGmOHvFh2g2H7IQYeIcU
Z9mAj5ddoFyBtkiLtcB987HFLpcBJ3MlOHZffckunwseWRr80rUWNEEP3JB+Hu+LCajRQIF74pGa
9rF/HsgpmzcKi+6UsEMhDsaAMXUt6fEcgvSIeoBXwps2SvQ9V2BjW5EHcrFMvHU+6E8tRIfU1t2f
K0JxNIEcmZLTOBEIaVqzKhGDTGDTcY13T3TAzM/egJNzoY3WcH7KpO2puXp4cYbOIBTx4PM5LmiV
FbZD4bhAofINokJyJRQCv471ZVpu3RVR80F6Gz8nRf6DVOqrvH1fepIAlvUs4jFQFVpLSgjLlSRl
hh2heW2YX/EW2iW5cbOR63dgS8s08KryChXMXQeI+XlDN6kxtPEe+yvjaJrK4XVDXlbnsXjyI9SY
f6hXakzry5zHRC/qON+t1YHvp+HOp/AqPit6YwlXiOvtzU8LG50ptOF8reJyQ4FPV5YACndnECfG
Xdehp2eg/kV/ntkzGNKQyJ8JQK1L+Ukd/E17aoULI+mS5fWc+XKr4PH8CRp8Az/8LPZE63ay2p89
nOwuE0ayoE84rvVO819Xv6XNfzfr7DIVw8eJ2I5v3GDqHre2WoXY+Ep40cdHrWYMhChVAzRR0yBi
D5NVFGvTomNViccM1EySksLpuhsj2noDlZA5IEPYLducMFis5aRB8UIg+1fq9MBmUPIurGxB26BF
OjKBdW58lQgNJtyr0Y2CDaCOieVhzDIVTfAbKX6r43XJ8o2QqaRy4VnE0Mx2pCzf9haeo96Vpz8k
3wKhkh7ZcPNJIv3sJ4WNNyJbb1IuUh3b/dOGSR28qwfj1eR2AnNA0st75HcWQW1RmjmkXczfv3wv
mdZdN5a4LXsWZCCPQ//beWEoSJWPqX0niIcIi6YSYp2rChJAuUagxJvoWoAVMY+GMyGZu0BZl7sJ
nV95IybO5qzsfsoxhAe1LQYZlVjLT0mRrLlLWm80PhNgYUc7tDYoaC3KNAOXYystImQWV5CIQQkP
rE3YEBlbgyiKkVwuvdDO+uv2tEkWEFxqqoPpqeQ3edJkTlu+/WZfRlyTwD6iWmzC4eizOKVmH5KK
3mMIzUaz/wQXyQELQhfgVS2yJOfpWH0SnRIVyoR1vm8pCWn/3xr8LdnZfjvAgByVmGGMYXh5CTRU
pOW6Frd6dNdq8aiOmYwx4ghI2qojYC1SK2KLco0Fz3twBn/Mb/eQlrmRniciVbThA1UwL4q2EYTb
WDwbwU4atJB6PuyTxV5ualUGgd05qDcTrI18etft/NCWf+N5R15jvjmmhujSIN5PcgKiob9RuMkc
bmdK4iKMKCNq97KKBh9mp8ac6ZK8vh5m3Galv1HNczMobrexXDfl1oLhN6YzU8a2TbKYLUPjs+T5
F7aLIsgBc9aJcI8ga4h7lHM6++IC2NkgZ2EUXvDgbZ1DOEWT8WhdTj2MI1m+0j/bIqZ/0T0fzS+F
D/sJbsIMM+4ylWLxWAYW0e4Usx8Dl0JCMLDoWrQSchUL+XGSmLeTwI8IqK2Eto8Byuq0MUz4E75l
9klByhEZigx5ddqut6y24zsrX71dMCCH93EfToX6zScZUynRTegLzNSvJNOGiKsKA5lajRuBTyR+
/bdveOIpUXgfXpDR22nLrb/C8gr2J+WfO+BL5w9XecNi4bVSrE8zmvxW42WQJDLQTT0ppkF+XUJo
4xbnhrXGfAmXKOwIFv5P52LanMTjK4/sw1irfbkaArH/rMCOZZz6NHoPBdzIk7ku205mZMvS2inM
Ql/H32yQzmiXVcH8fnH7Bggnbm4UY8asHG/rPCcuym4WYnWQqPmcHYO4CDnezfkgUomH5eFBdPCg
ivp+19/unagAK5i4MpjldOJt6q30BKlJN9JlbuyuDdtdaqjQn59Pentgtc5Jx1aNI11atL4haizC
P5WE8jiCFjTAOTbiaJqCFAbBh9JOhDOOATZq1WpTaxVfxEeIjbMcA3gkvslhsfvaq++fo/zIXKT1
3XurOWxy9g3C8+Kgl/xSGNuOu9ayDIzPsH5CmCiL7P8bDG2c9fgYzIkjAqfBjG+1cMF1h5OD4X1S
r/O+FT3v6aGRlsLENgj0hoByqVfBVEv4SA2nHEH4iThm92VUWzibeEnNPIPwjUQlNZO+H9E36hqg
EaolZKsQFvQlhX+oulTnUgvZLEoT2IVtZXGLy6PC0ibL+I2pzWemLdDdy7omTdhLn+kQjc0C0Bwe
tnrxNrW4oCwvzOwnzMElVYATwmS7A85c0uVHLDQ24yHZwIi7eOtUG5wJT+Os217LKU0aRHdCSl3N
Mev8eIdSPWkpCJV2/nyxNlAjrr+RIs5IrW0nwphQERIxFznns5y3vvYRaoSTVB3unmZM5/9BiaTK
i03AJ5ytNuTq8YtmOqkH7r9LLjpchz9wbgy5WsjAO4tsysBpy125SzPrkpI0tmt2cBbk4q4t8aiR
wPASRAftL3RsTjM44Z7c0mrs/XbhhEWjrFxTQ7dl+V1jvqjCFtRxuZ+mFPB4vmy/f/grE5PdA/Rn
RhZfHWmJKhDFV9Mi4Y4fA9P88BiSuYjMxVANuhR5yTqYrtEwsyQum1k/8sDDccuMQTAdeYFuKp/c
V/MV7WK0cOimr7o/L8xpVrPMZJAMwANktzbQrVEBDsdCCElHtTFMcVdIcaVgrWexfCfZuMX5nu+W
wcaBS75Rqc7BtxwQIZ64n7LqdxeheD+Lk4UBrAc6TQu+4+ttbY5I0wk/MWX+e35joWfV2YgTjAV8
RRo6BuhOoyogrojQEJ78QXKLhQBnhmZhl+LxY9mCc3AqYb7Dav1Lb3Z1ISf1LYBx3kqxabwFswpb
1gyc8dsp9CBY2LReU1Qur0gpe8E6MY7+nY6m+Ddq4pvsuSs/xWYKGaVSVTkqGaBx4HIF+2miGlPp
8U4TrM//LxY3RfItua5woE1nbgps329pakIkmx+vJJ6V56aGJg4ozq5f/jpko5dl1NSbk+q7mggz
MsBPvBMq9qOEkfSr3m/0lWM1etwoZ27ifFUmo4oRxlach8o6pDwZXgYul9HYG9skRF2uoxABHX7v
hRpwyUNx185Gv4dmHTBKsU71WAVgc4H1th0UQMFGl8NvzAhI3uFJxfbRW21w3PE0IHEGzcRybLcN
rVhcDZJPtPrKkv82Bf+QmhSKfGHOaV/KOsrJ0Qz676mwoT264iAL8yqcnSPuJsZ5BpkWAXV/pL9R
C2efXvR/4TbOp93cFZuNl/lq7Xhy2HttLNeTSYu8/oP7YCpw0WRbKzHMtNtKPeLWGja8l1Jbalpt
cq4WV8oEJFRJvdCRbatMkoIJTrj55oYFF5aL8AaXEbf2GEqU3aEIjZGNaXY32IakiTszMlJmi6W7
v0YW3oOb6brWcQq/XU6EIXVNM8DZFc6SvG2ZGGFNVhQidMT/QzO73oUtl/9i/tqslx1kFruGFa5c
upbo3HUmBkhULeZwHb38fbItI4eqBBptNFl4Kvc+0Tt4VcEUEC8iBMgsACcy57VXNPc3tzei+6eL
ZePNYojr9vPTcDbcvvl71A054UzoxGHz+74Zw7U+YhBzDx/AaOrx7mrGsXh4Q56qfS+rAY34Pxf4
pacaw+N7I8W9H+G7DbSF5CHA9143T6AhdjQY9OmDn5l0v9kyH8nVRQcHqBCasvHO5MYomH5VBq52
Z0DG/PE0F5Xm0nkE9weeIK4KCePB5iCyJtj7DzMr6PoxPlDJ0gzGov9IEmB9cCwzcXbQ/2cVHwWi
Aio/I/d4u88DHidWNV8IblgsLL8XkXkALhT345RbrJvbYia/AhKIUlGXKWaaNvDdgdw8XE1KPKU3
hTpVgTI4tOY/h2H6DdoaVdSZ7OnjDXKAXIFC6vY5mOfyKa9bqTbOM7X/ILfNyDt7gX5AE+vgdWAj
wSg9g0P4L6gGIXVrL/Gegaa8DE4TpR9BMBcG2jhIEzSsp7BvBuEp6w6yGXKSIHxZxe6CDG4M5NKb
F5pmLEnHNaIUE0yW/E/vAqLbTx8wCXGWxvPgIhXZ+mTgKRedCWTXnM4Xw40yf8hP14idecDvqiEe
TKTjmqeLGZxaogoLWmPzOmXz6pIpxL8mEuQZo0W3OHN92CUq658aN+hoTN/yHkZIRxTDKHqDQd3T
MOrC9QM3N4qSPn9oTQEsgr+DnLgv3/fMsJa4dLZmtVEsh1ZfM8yKzPVxMIRPtia/+IBmpRItvaF3
49eAoEqk/emLc3R3BDYiM9j0kr/jOEi/77cfpkfIrkK0oWoQYJE3wkCKc0n2Vn8XUUaZLzKkO14+
C0y3hwXOmErIpBvavBKhA9qHtPHHHZle+Dki7ppktvMZ1XRb2332geQaE6V5k+Qk9xsUoH1y/h4R
XBLSGLDao1aCjqhBjn47AtjcHpxUhsJi3tdmm60UyWmSs6qBC/TaugHxP9XbXyEHOtxW7RaNJnOQ
RwgE4NMyjkdDNf+eVxxC8AwE8x62cI7ro7zJeuwX6ltTT0W8iespPlGPsGpPfP2GWIK70kAOryvM
/z4OpNFAQ62XXL6pOA8sUzKKTG+vd7yljsMNUpTrWaPyYDV+CvmntYSkGqQl4hm08y4f6n8ooqob
+0No36u4ictAYm0tu780yiNuUP0aZm4Vz9fT1hcAAleEC4pME/pRriANAti7Ps9Bd632sZOaiWcr
d8v+rljf72ZKZRzFsMU11Ibmk2W3XDa+dt0IAmZTVGovYEy6RbUH/6Xq/DVQIU7oLlQCTExKX0tY
HbWOjFeCqickm5UwMQww2PIL+WNAsvd4XmZmdi/RPAvJclcpkpQJAXT/bQ32c5LtyPtx2GPruD1E
zjal6PofH+QiLUlovg3+EDuJCnSQ86R9y6RqPso9z3j5YX9hV40Va6Bni4efhVtSlsrSzqikBESU
X7G3ibRPsDQ/LJoJe9d1SYVDfH42JGv7eAnSFiI94NsiZTCL+M4AHfrCaH21ZvqLdkYM2NYHx9E3
RygzPsi3H9D3qt+aq4vQSvyWshkqfirwH0zdSIRWF1Ygr3R9oBcWieJN/pAJtAnTF0sVQIiDLE6j
aCezv+oZ1WOPQsrcG791Jtg4f1Xc1mEL20H803xow+4JM5UcJVom3O3Hgf+ELojFvgpoFR9KvcBu
lnmcJ8RbeAmNaex2avwu+AtXOrod4vWpDVc12IGpRdSaxfJBDSAa48IbhcXKSFcDe/5Jfal65zx9
91/pOC2wAcRoSo7FZA2UgES+jObFaTS4Vqb4ecAxmGoV9UmCTUezi1PbqEhBhJBlCoUAGxOz7Qvn
qi/slA6fT3bV+pDeI/MyxXPYmVg4hG1AxqA+aqN993ftBcAFHxZt6lNqpqV23RAbEY30iWjk+mj2
Newd3HhDI9uTysvx3uogq6eoVm6Cwci/11I2GabtRF5RjxaDXcFEKFTxHQiGyeFtKz4dQDBwXhUb
gmo3/0651RXFICFpT5XBz4D6/YkGngkqHBPxAwOw4tMac1asJyCdhXW0nR8h3y6MGZj6uR1+b2IP
OccR0FmpArEA6IPmB7YOq7r6sjjMpGywes+0xLlyABq8tn75Ahp751ruy6RkWpd/Ar5VGNqLZlVh
MWj0G+9SxJKEIHri7Fi9qYOav61jIoCcaEkNmGTsjrpfpm6VrVsOdncNIXK4y76U2/ceXboqQMZb
F2V25i3emVB9OwQZ3zbPadQPu8eBAX/Ta77XgOGIo+BBo/Us1erGkJ+am8YAOQ/5K76SFLLyQGx/
X+GSUAoU6EVvB0XZuzWjTrEwMd5sZEhNrl36RGpsqyZBeN5/DOmty4PkV2fnnX5VkkF7SMYYJHoN
+rqpH9TUEQTiF/xtOer+3jsZPufs8Zuj1i/nFDCrIQtFxRdr+poQAWxV6+JDsuaaQwlSb90M+d8e
eR14SmPCBcYjAEjPCqe5RFGaFJ4IZGleYAlzBmi81/3/Vz2rJUve4RefPKte3/RX6uz0QuBJw10r
JYipziXp1lZ2D0VDJmQixENvZ8yXa9ynZZr7ZMgoJKtzVME0eM9kQiYibaL8XdLXiI8GaiIiZM7h
SsNTKE2DQaFTG6WwtM3pwAvOknG3B7OmA0C75eoO3UxDZK1vgWclWkUuPpidGI8Jysi0jb44JlpB
1Dko9kNlM7VXRHC2Sf2VJGTJ9XzzXAbXxQ22PBRjn9zftzilD6c5Et4cUv0NrXt1oMRgdyKmaGgx
byy7b8pKY1Kxqpprk5n2oIsXFMpsIWJ+SFkd7T00fvq134HsykaSd8JBS05vqGWAxHJbl6bisJPS
fO+hYLJtkLxV1S2OWr5+fHWxcR3cONZMj/PVfAa+7EHeoLYXrETUmvDNxT/43pM7Zp7eNJU9jl/W
Va8aWXl7q1t2RW7nRnKPI0szjWk5QTivRVvHjF/Kuh2OhrKdN+xlerOzhCMV9mdRB0+oOnfT1p12
j7/eqk8D0CEiB8D1LurIm0S+cq4r+HIOw71u7/7QxecTu5Ho/X+kJGoIA1i+8xLlCLlJlrqvEC+Q
pJ15Xfp50WnTxvgaDq7X3ezqvDS14WgD/v4nVpg0wIdm/3wKfo1x43NpWHAFyE4QYPace8JWtuG1
RRL+NAMxuZLqBmnqJPiw8Ah9FRF9RibkyHpAo/mwW8lLcITY9aHuw3IZjB+Uf3Xnxqoft22Y+gje
WBIXmzGndQEW7H1bx8ta7GuQUkmNB1g0+gf79ARv/bn3RJrC5ZJuekVATmD4s1CN/XRVz1chrMvu
9ZRnjRYZ1jPrfcuf3kS2Wn/MkpIANaAuimcB0V5F5GUcg/CXYfNY8boF8DrgjggRSLJykk5l5a9y
5K7maArlEVWzDFFacddySJy0KcBZkLghePqqjHC1NuQ/s7PeS23xaQLaSBn4sajWpF5in/OOgoqz
vmXskyzpXsQzY69CFe1NFnIvWp66sbdkHZ5OSWtp8PCHuY+sSyw4AngZw68w63Bd8MPXjMdcDVQI
3unw1wQoWy+Fo1apI0L6h9Y0md00Bq/UBrZbhXI26IRiMoJmRuEwjs8gCjq14BFZ/SEPdPd/CTiu
e0jqMATTOQgENZ20hS9YVlRO4529svV6vxY+cKyFQN0X3QFHbczblinRF5XLBBbklOp+6fn1BX0J
OqMpP4bYX9BVo7/84zFKuWoSiS51+BZ1MMk5EXv3y0WvmfKi/AXoIS47NoGXyv4aFTRC/9mqcf7R
mso7gWsLK8vzdLV25oJbVbngPER5SKzHD8t81VpXduVAUSYJFRRrvfXh8mULuUGrfTEfJIcGDS6j
gQT2GiDHmX094D7NWfEVdxGutEafBneDGZSK4AsNqjbHsQDM88ytlkg27dgnXJFDAckI7OTZUTuw
fw/IhdWTIDsXqoliUJI4lWp5gmkuzefRwUEgYrVhJMFPd6zT1ZthwqwCm+GL0JA6pNh7iCODziCv
MjpzoaGKYdgibCRB8gNiwFrdwSFVUQCGUJWwriDvWPudJFdxUMoz6fYje+HC2wQ29yt64nl4fqGE
9a06fjJWubrgLGSO9xpspCROpaYhtYAYg1c286IAROTIWeqUAQRXNn4daG8jH9/H0G2JHU2i/nuc
GgTmrNcaj0deljQKlDDIuj2FTGCq62DrgTjpLloiG5iopuv6F3bG1cWepLO25whCV2XeidGzObLU
v0MYcqFnp/PByjtKYBky57RoTYhzTM/tYxvnfMfqzrWwWgjF0EIiTaI6qS52LGFS9jVkpSRpS0Od
6b9X3EzMiwTpk6mpYzuk9q1dGvVc4/lSSPtXyAszLAoOz8TVc7ZURPBI2o4DzU8BlAcZ0s1FYG6y
R0qOHsNYwu1SGltm6ShU8hjaRc0wYKWtuE4h8UDdXTDx/7Yy/Ybk8Jfv7D23+sevvlluSadnXPlu
FPQh6509DHlW3u2lfvR1VntR0MDdAOrY7EZOSuo+AqQTvojcg4Mh6kkMNv6yjjnM+eROC+JhU72B
5GuFBkNWaIMh+j01u+OefVtTyze86WQ4JBF8KDA6LSQ8lqd0MV0GdbavLXKPTDu/21bN8VbX2KO6
88IPqFumN2R7e6fp6phFKuOiHTzcWyY5jsYs2LTT62+/uAh4AcuLe3338JOcMBq+05cVBTfLk+KS
BEPGHOOeEmMdn69TL5hx6sXnEhhQ89qvycSd9yvrNlJe6TQPCiQ/rYDQtCNlsxxTiEM3E3/6spiG
nxdqYp6+FCzuwqYii5y4bRaPG7a8RFS83D1s1XiK4n5LpNi0qbnEBDJhYO7y6hclsdXwQZLjmVi+
zMY7UothuWQ0g2tSNaKYNICkw+PjSApmu+04VLy1quCJmlYg9Zpbvl5FHunjO+4R/oxxcI+thom/
UZeZLvSilV+1GzZD2KCA1ax3FiBm6r5Gb9U2TyRUzqq0eVzilb4+17K/jJwiepxJMZqE/UdxAYG2
iLCZPJSxFKX2UoLs5M+e0QefIp9T2YKns+AtrOFDjUpVOZJpSRpvx+iw+aacYUTo1Ufe6eS8nRUy
QOpj+BhU74ze41JHJrNgakihwr+oZSAoXx6ecJEOc4f6BdN/sS3MbyD5X2Rex2RW9/YJPCYUVv7e
E4dpcijCjWsw59DEqMg5sRcmVy3VhSlsHq21ViKQO265ACImSkJ2j8x3U4JWI7wpnHHsiiWIeGEb
qLwa9EhCsrUyEdPN5dff1yIBGxNMESzt3dSIMrChTFZ52aerfHDitkVu+o7wg7h4312lBPIJTfBM
z+0bGTgxUouoajdS39N9e78QvGFBNe28RgHyO+rhfC1Q9efTX6gSGjuZ5flT68HUH5SwKnYwLRmH
D/s2ZpNukFllZeByyEDHwC3eoxCO2U8lwutkdHAGKsM7KOaM9dGIv8LOCz8SOq2DXgBMfzoXVZjm
C64rZLojCi71TCpdDTfgmlyI4yXJ0nrmXFXe+YbdNnS9Lr/Gy/XdvPsaI2DvoCpz7w0mdn0t6xC7
K87SnrnMEWxnSRZapKFSpk9WrLRwmqEzZDTGEiUqEWpFAC2w+QvygGix9DOFRfm9fJ4TP9XZkbpL
5WPPLDteRKqPvUfF3F7OaxagRGsZPxlAdM/JR2x3sja5Nj8Zdq9JuiDtRsNdttJKp2F1LILKWYcv
VuaES50MpNuwjLM5yENraeLUx2G/Y5Ce/OA9JXnz3Ip2WNwBEJsPH5/FlbDPDM1AvSv67y8zRG6v
CXrE/iHfKifWdD0TztnRrZDKHl/GMc1hdRHghjkYmw2ppGB1PONScv/wSCPQjfHEbD0Agb3cKtdf
8Q3QjKRQJmOLsw8cgQmbV6X4oKSKNVekmcSzW3waFppwaBcSRXTwV8QIVQWtdriHeNj2CKMf/z/9
YgWGRs9MltYfRxof4bg3p9dJC5VyIw0kxiyPXKqQTExh0U00joWM7V0x0abE1/Yn7/SfkXU9TEmK
OyRnN3kTd8Ie6Q/eY37dFSjq6z3QVW0voaKzElJKKIDN0CGb4zrzqAx/hV5zoszK7VI+WsP3Ye9I
tCJzuVju3Uy+IeUmkAgrC1avfZ0FfsmjEL2h/v98eXeOiEaRkNVhv/A/BT+USUmepWruy3ULfLxZ
9I6NwRHzv9I+Qet5C9G7OLdXg5HhZxdKjRVwDuaumWJu0jfe0vW5/ESnHYB0FaBtdbO/g7oXMBHJ
shSek5AYrxh1X0jAmbG+J0e/VCpKX9JZkaWtU8iY6witN4fxGpAqLZ+SogbfWnO0Ey66XlpKgnWv
lR2ReKH2+JxFSUghduiT2V9fDvzz72kAjx7CTXFsRHJnufu79X2oVYGkUG3anlox2MehBuRGce1G
eRhcQish1PxOtX3YLgCz0GhPpxgSLf0Yv+Epypuyd2bQs2ochsuc6ncqj+Kttj5JP1jyGvZjUMG4
ZYoy+7SkLbmNqxXI8dqgcSj7Y0gB2IbDEBms+59yrLmX+23ZL0MlMX6oXQXikE02E0wr62hDbsu4
68gPNE45XXaoMQmAaSJPW0tx7dw+Li6ABH/VD8fFo80jnFA4JHqOUrT/aZqV4UIpLVxmMgmYz4Sb
KLt/0vE/3SiuqGE7eLAeVaF01EdT3z+l8A9T6JN+wm2hb8MsxTHDHSNaGvT0YYTS6AYXaP+2aO+O
1i43NUATfIBvZ2iCZK08Zr5Hyo4wo0MV1/u+I4HZU86dVP3JkB/M6OTok6CrP75sINEkrgNlzX2t
V3SH9SWB9Rv4h6Qaz8KP3To8gFaoSo9hNv5ICk3fMFZzb4RQ/omjO2yl8/bsOXeuE/8tHMeVpEM6
5LjT3QkrNGJe7KJXQ/eDVycE8pfT00ja4Di2KoMXqJhibo3lgbFCg9rb+aYYzput6NeCjmRM+AM3
VoVARrthGdBAGHmRy0IQglqGst0C2iKqAHByFOECDWP8P5fWuhNKZfCQO9RPiEBqdPK6Z972uUfJ
2f4WHbpL5C8QygHAP4n+PEmnDOd6zDvKw+CHC8M2eAf25AHPfBNcSQr77W2yNOdxz55JxXl7nLZM
N5HQnLO5jcVZSTTpjw+zO9xXqeCenFpakky0bJgZcI/Zk6f9NfIstMu3eEoRzGAhIr56AJEjOfPy
OnULakte0UhoCSXBJm8LuOd/IWY4kDyXNTDUZSJSOnDdDpPKQjBqlf5ADVKRGpPZ87ds4TiHOdst
FSUKDJdDmIC9QcCeXmtAfgocXk+mR+zidNUsgPBtfygmV4ZBDB33bA2S8yhlKAkxcQJOZSdjfcwI
eJEhTupqmmDhErYml4oHAGa8F7YsksBVGXy9pLjRh+0F/hPqIxVDbRpB+qCVtP9fqZZBQVOR0QgD
26DTPNY1zpv9+K0FHbOjJ0+wnVL/EbjbcX3kImi1BRD7A9K7+7p4aBwx1Agj8Xome/i8DmLxvsMk
I5amRb4RWRLrdjjz5D2k7xUzp43c3FIoFqZ7bbICpOe32pD+TwhEhPqhcmZsa9O0++Tp2x6p5z/5
HNmF9gF0T8196Ekw2Kmlc1fQYxBK4wJzN0hzqK5QHjBsP+70X7N4umo/IDmzDVJIure3gRUKbLnL
mRaZ2kZMgb9EKo/F496GsM2ZA0st3deTtRKt9m4AENJRKgPm8WiJ1hgT+bzwLhbHwUp/kYTRsMP9
xQGBckAZnHpJMD54hBXbgUmiwyxRDw15rh/T4CIx4xXTEIAmlxdQAIpczqFXFKFTM+13YrJAXK5B
7ip11cPbsvujgh+DAV9zeLbDw8edDTLDnbAPiOu4rSoWV+qbZeg2fHV1dYhVDyaqVMv6dslLoA0i
Q2/la0QHGo9vm3HRTMog8GtfhbDoXf+wreISLlDy7RwKb44u8Vq1FFzZ12sTYLt5SVKhvXxC10EM
xJ35c90z8egRuIYXyUT4XYxv1hmBysx5j/ERa7V+SQTBF1eZoLCxgvV/bzwffKqGCP3Gb0CDG5qm
PRIzp3NrzULK2sH+CsRh67XbLD45UzjOjt4di/88sqz4rVRL6axqJ5vmGic2kRYr0RmrZ+71t1TY
JpKPThsxHMzUEaS9a/dzPgt38/GxU8Zrq4CIeuh5gGeM5dyo+KG2bqzQQBfJOSILgIT8oGeXkr5B
bLW+Vqu/5doWyAdDCpqN07g76hhSQT1b4jxxySSCLJA/qgc0CL0Yazu2ujBjqR8Zpk6kvwOuFP0g
zhdeVSIWANY5PNTAoK7sgUUjZ6ta2qZKspY9HHefkAdnqR5BmVAaXG5+6R/6y0t9KWJvbs16DAWn
+TjHVevleMKmTJENFCDLOFsGYi6OPG2/bsUGtM5qLG3cWNLI2ceduKK8s0Iv5PzTVrzVCMlOgvnn
YzKECdfhi6LmjxDykmj5LxT40nbtIr17fbtC9T++JxxmxII/m/wv6E2J/g98UyosgMJxRtBnDFt4
n2LMAQ552Ti1AiOuBLO2Xpg1cs40kYBcLYWs367a0/g5YbN4Y5a/kbbZqDtIkwqiKd4enwYocctt
pWaVK0/CqKACumGKVhehQGjpiK1amgHffmmosmdfR4iZXx4OqToWG96mmLsQNl2nlcmhLyLzEAgN
N1QQgIiB8sJ2U5Xl2zxpQFHDMIM+kSThOxukl4UveJJJHjNWnmCVVbaa5AqCLI0EmZuuxjrQWPJd
BeFlGnxhnX1h4+OsInuq/MNbacnIs+CM3APoWoPqafGnMjBDqPdEyPUaaU30UO4s8cxPwdyWQYN3
HWTTShvc7GlabVSVw1hSMA9h5+7xrTlV2AWivE3TQL1UDBxST8zCGyrB10jc9WvGYweGUowjoTBu
VVlx0lkMQPx5IsG14qM03clcft4pERRrB8zdH2gzbh4gzz+cZtbAx6/uJjz/jmGD9MfyEC+Z6HE7
YR+ODJhbdETlIGH6HPJHaX8gw/ZgRIDJqL5BGhwKATkEh15iTY4AQDjCXwulMV1FHSYANH1eHdVa
DwfgbtVk3cp1vonnYKeLcwN76J+8yXpTztbcUX0L+jmfcE2fYAeet5MMCINkybt4klaQO5WZRjU4
CBFr4dcf76+mXxgKA5OF1tn0tPqeEu+KL721AhWASLae87koVTGmbTXWJlJse9bMlQbUGJrWtGxc
gbJDbMi2J/LHcOZl1QXT+Lrsh5VHU0QEaN+Cklf9IYsii9LetnEsSYQQJIAQ3XPZqgiZKpnp+b6D
mYPHeNsYOAlUH+IsMHBPWmhCazClp4Q96NAQS9m8dGHBiL73z4lrTYcBRgTw4pIc0OW8ZQqG7e6h
LGEu7YuiL14cEDlgZb76DGv6do2eslxHcgdZOKXJC+FRxQJTleVQqixvjNthsjTS0biZLrKPmhq/
bT/W5qsTZWem5cyGDqSgm8CpFBgkWHMcIkakhyX1TT+9ZmWifPnnWAGc/aO3Zf1pItAIeGmJTjoo
UQC6fAj9TDeFPGd+ezv6ZwEvhPLU20xi1aPyJf5q/neIVfMhCbc3xIGkPfIdFxoI6IEXKOninc02
wRDo4NC02O8JEjUiWOhsuWFE329pYYjKRePXr5ASBkR1b/nHPpp2+QqXXwnv0q3LuHd+4T2lJzWb
ZVYDI853qPqzoB1UnA/2et05ST/zv34/ZoJ08mepbcaFvDQQoDc8S6Oq5+Mr5pA6n0VOe7/0xuFP
/AwZExKdevbsDc0i1RjOnje/fHWWkqYjRzJOGaTVmsu8x1DV36aeAwHK4QidM3UC3BXjU113AJRb
P/YugmHfq8rGh9fIVsBUZPv74Ul6ngyo+vuEfATInRA1DoiC1EW6YTIb/Y459ldwX1HrBCegBlPS
hRdwd79KMMsotYwarKb0mJYz1OZc5HYaK6QPVx9a5sK0/HLqZ+5AwTny7JbFuwzT1Wt+jQYUCWtq
dLSxfd6EsDha3zvjS35enhn9CxF1IofZEEVeHhmCJVu67e+TMSkdPh1yUdWfIx5EOKU7cL8L/3w+
CzOChB9h37yt6QbGI0Sugqd/Fgx9vomZfiN56tM2j1WPyYR+elqKYvmpqJPQ8Vx6Hiaar+pMgFgP
71jAoI9OUg8Ug66h8+oVjT6AmZSvMJlrC7voCuCp8Gi4pOGTHLzquzywax8DMPbk5MfleDUX/6ac
eKIg3Y0YlHaZuTCnzb32XHnyMuzeKH3bJITATLyX57alBmRjE2T49EzAg1J42b43suVQZ7ytmE1D
6O+mgSiA3SeswQyHfydOXMeCZh81UAlv6NxqCRUQ3WgdFgTgG7d6co+ZRkT8BVxDs0eXwz2BeiII
M4QcMwktPxYlt7Oc/9nFcO6LFoxP3FulWrkgaj2RPi/473CcvlsqDH3/Pqk6IRPinv+VNbqDMQpR
hoHnDk0WGqvquICuQ650IbWqEfDiu1zKuBzHuI1iCLg9ExInjB/yk2pCatAHXD0oufBSVtjOEPXr
dc4Qso4tBh+fv9nM0nV9BJPWqFLN/WD9iEmsQfNfyMiMKZATIJdO9zO81CJcTLgSPsFso1ffOIOF
jeloXRamkK/w1pi7qdd8TD10cNNXeVuFi00xmkNyHrvQtS4JhLqR4LZJNI3NIThcIxXcEk9htpd6
X311Mo0uIjRguClPV1Ie35ez0hbIli/jihdvERcZsa0IjXEZAcnrC9Tbc4TDCQCUUUV6f+yUw5VX
O194fPD9n9zE6PZ1X+OPMQD5+FWtT/NSy607v+TuSvYTSKZX0RtDO02gC4ACTu+337jzspkiTpr6
D6GX/5Ea2MRlAiA/GxbRX+OfrK7ixjwxivwKSNbvQ15Q/Wx1PNVM6/bsyYUpbym4e9ml9DkqJPs/
NvT1feeV1GMSpysUTPR7or1WcUVGIZMY65Gjy5Dmmur5fAgDC/+MMExL6sphZgxUXLC7eAYXqWYM
OL4lRa3sK3qhniaNKck4kIi58m/osThnxvTIDa0Fa9xcNAc7Vucp2sobrQ2Fb62R7L/vxemUdJP/
C4eFgPy209inWG8DLeY7my+mVmyzdfDb8QQScjSBLANyrZzXf+27+QHC1jy4H9wREYnp4gjZzXDn
/KNgwpAXC82ijWtT6Idy7Y1HHEqHGZD4Cwh2uT25ZOIenyxLXZFOMDKsIAojrohX9BCLYS5d39u4
gvxf30GLfVmqJV96hD0vgbdbCHvZ9kqJ3WP2F+TGiuUQhgPlIvdgk02JUdjLdhCKIhW87lpMDYne
3KAsZybOYgn6yJKU+SKW5s4mXDB+rnv2vf3ER+gNqF6dEdjU/i8XW75a4hJwVE0HEjhFAmwZl05n
p9q+JCcg18tC45rLYyCrEfN792yXxN1EH3c7J4/4TBi7F046Vnvg3GG9HM+dsyO+C8m5s5eTcDDf
qIw7ABXO0ZBNfLoLLhn7Qo2V77coBGT4LpwhUxpB144wVmOGUx1n8N/4VYm77FvjnFSZz1lk7NGg
KX2TYuUWf//nrL5SjRDOCUjjBXSNr3YOGgPGkvbTf1aU1gCjwz/LEK4218/LcJB0Typ+v/3mBcrQ
x4P7aL4W1iJJNNAHnvgZBrsCbhpEWpWrOOB4CMWz6UfmAHqc7e0/8jytiXsQP6MYDiJE/VTjVGux
/ZPkS7qUC7toux4T/XFG3B/BQME/z3t7rE4bQGQvKW5Je9Cxp3NeQ+OlgwCr9Ceg9xzASm8uDvF6
r1ruVe8qEIMBDfbQPjHi67TrWB+BCvyzL6mJul2EZqhWRFfoB4fG0uv5m4n/Pz+49NvmWiHR5o55
cfzvPnFyj4mV8+WZ2m5azpVbDUtjqGcqfzhDVaP9awzZ4XoBlFYp952XWDiragnw/QaRJPymtMRL
qxFyPPM+Ov4iLdMZmNRghBQHV0iVqfPFYJe7koRbFrV6EnZ5zsjlk9qO65IREaHI4H/H93fDCwdi
NxsDn5U4KySZ9/GIe3nZFDo6td6d10Kq0ugSNVCzwqQ23TsdcnkDDFAJM76ejIkHComJheOKdN6I
cRdJ7wFIlbZ6SPVPPdeB2/nLYIjHL4ugVqMWnaf+cXi+sS4TuU4voH2RUIuZd4IqKfygN2xI8ZW8
mZh0z3OwB3W7dbpo3AUZspTgROkOwWok5fNvJtI1sRgngzSrNz6oRcsX0S2kHOibyrKQhcLvuHa4
zZ3NZc2k2UlaRuK7u/sgIEdrR1BKnAHOdeCyhPMcEekfjI9XvVJBsoJuF5MveY5cr6CIsTnBW1+t
0F8uoFHou4lvG/QpHm9QTKiDSAcwRinQGeT4R9Q4mEKeDse+XOIOcg2h73waz1E9N2wOzKp1V0Xh
PcLmf8Z/blwwa3qT2eTW95FRpTG0i98JoR9WiuxpD0IGsRONocgBOXV1AJaWQSke9tTX7ekNbFhi
P5C6zTXPWU1eHgH339bxJgWvfohPC9NVHHYlMZYwhlDRQt9PtX/GdBMoucqQ+981epz/vmaUmZIe
MJ3sNu7X6zeOiYkaRDLa1WbYM26H6FV4GMM5t8GYnfxjs14ynCh7TTTbsa8k2M7qWYDMRcDS1SEY
cKLJyz4zZMfYk+IMXMXY6jF5X7X43aiYkdMEv6X7dWO9NsWqsyDzrCvR32DS9XcDVo6HBrSZ02EL
z2OkM6pyFttdCL2r83XFD2nRRVRugmEZsqkeLYfNo2VuQufCnjs53ENF+WjOytdeHD0D5yOE5LOU
8Dh9tt8oEnQywklDyqfLPxquUNbQhv2gMNWUv/xkAQvzw/i6u9ETbkJcqrYZHsioa95oA8saZpXN
s9EMsu9cGju+pLKdMqMV8EGHFB+JFleaJ5yunop+aTFtZiGYDtvoDF7ZO1w9H6lYJidqYckLxFJY
zzUPAxGcd85/IdEr2/k3KKWWxCG35KVAkFl9vxx07FDrCvU9YaW7hCC10bPO7c+w+55fCrO1Ms6q
ab9mWSfuB1HM8qz4XoPOrVwjql+rA/hPX2BhNTjGibG7uZiCcvskj7WUb2L7DS42pNk6iewSp0OW
fGHFNDJVu/ZzvgkQBMouMGwfVok1csrOOIyhLr4ukI5kRZpYLlRrX3WvMFhVflBi0AWAghF0npOk
6HyCKuJpACqmkGUOOlZew/by96VELK7p+5gTcSc8IrJPxRCEgr8H+1azVnerWIBAhHoWfZUBkKiw
HqsGoIJCoGVJMYz6HHhtDBVsUFLIelt09FcfPyXsgSuE3MqFMbs9ojxYxiOn24toOn16p/aVmS9U
P3Pv12ZWkBzaxuSfzOFDpF7ZUO/NJ9DC8vVdA4sNa6QT2s6zxHVTmh6dOVut+TZNcNxE5O+xbYIj
Sxc8H2GHip7xse6P5VjMdXIEvt5z9luXvkqmHO/FD5UK8YzY4Eaz1LnmEQZVWPQTCFnQ8y/XAOVB
32XGrUr0GO8ekjQndTmqcAmKCXOle1hUphHVHK0Oy9C3pIOLTEBbMSEZfdxy4cdDQh61nypywOSX
NwYpWbhN+HJoboK4B6C/cI/+dGTMXk6hH/poyOeF2Cd4bWGicXqpYobiIyYGxaQvfKkO2oLy2omt
IPFwrMQzs17smU0GdCjQRMlSbpK5u2hMNZr5ECeyeHRPv7dnS+10OCHZC6Za/hs27dFQvUO+uwJe
Hb8SHWjU8tg6Z0QDXRtLaeu5Y6+YHt6G/5kgpeWjA9DLxXKw/6hnM4YURdGSb6tZepvHmujZtbMN
Py3Dt0obNtfEPYLVPWHBBTrQr1Fo4huJmb6Imw6tsOTpbtyKZNsIXKVish8TvZLhsPFCMwwOPUIh
ume9dH0Y4csgjoR18cQVJMO8x5rlu/DIw9I6dFJcZrJ8eTUvB+WNM8BRTO+qCS9u0kolba39YC/Q
ySe9g3IrtEqVoF3E2BeiJ0ou8s5zv+qWylXlsYEwisyRDgO2R3Z5OCOpdwcpHWSNuN9oEcSe06vW
H7q35dAM3UDjMzEDmyCCDBW3O1Qm861InoSKEz9wz6mh19WzMWJ+MSaZ/ALtaGCZ27uHobsH18Os
TOedskAJXlbSvRYw//3GAfuUB4PKpFUDJSAGKPcIPGaMBXUgPscvY4Ip8qKL901CcswW2oEX6wpk
Ev9OGqw/zifYUcv9eBKWIQGHijGX2PoQTyX0pyY6mH+b0Dbuba9LQ677mTzCg/S20bhWHcCE3tnD
J/phyTqsHeBS8XmwjdNyqgqQJRrFWJkSahavmAF7CZjA9lm27PfjkafjPQSeICvnfijGBZ0gm4Nx
8rxpEjFGjKEflhYiPOImAvqhtJ0UZ1JecHCZ0TG8l2RzLBr/YEwKmPyyhxKFlB222gUw6V2zk86r
f0lUQqgkT9dOTYqyQBTm7EZhZhziK35733g/032EomhLrMXJuBao8BAwWzeNUC+olAlyxbPNo15o
uWfZer6KOvUkuGT4nf51LYWCDw4Jqs3gXFcMKXPD8M6Q7TQKIVMUln57y82sI6O/eXdYNhJh1rMu
ZdcCF5RUcjtbX15ewK10Ha0+XVCP1ABiM2sh4E/3B6aj5e7XUGpmM7qGXdhZP/VHA74bvlpWW7vi
gItRFgcNHXejnUQufeZx0qNwV61wUjAs40aUanHPOB8eVed7zETmJBTcmFFKVPjQCbhycUSPguEx
dz7VsMUdtp+7QD7RXmY+lcvxDHfnrjRa4//da3db3q0Jvv0BXHc8Qslyac0llMgFiACC2UFS3oYv
8beOriNvvkjufpDGjrCI88HpK1vfKcz/6nCrqvoheze+taun7aCHYrXKpY/dTKC2Ow+EZ8wQDnyy
aQ04PEO318ZNAe3zwSsfeaklzAJuLrx73zbBA1C94hdiUss8NjB0b5fPmUxcgRoNNDelFniqK8fJ
if19qR4Fi7lEyeMqVHOiZhhiAx3Tcn9ULQVBfQZ132awypCJtYbNIPOCDQtxYsBHtUu7pH69XOPW
JlNDl3spfZ4tevnXWC67evYmDNoCyCJL/3bx8q9XAQkMdiOfhwCKEkSThaqiAF3rlXLZdKwkdVsQ
wyUV5OEjej/+47rhGGH93OAzGCDO3sYhI4aXZg0P1mqQf/zntGbODnneFSfMXKTwSQtoSO1X3w2M
kwPf8Z7bTbhA258QB6YnlfwYy4pvRCpzCkpDkUdfh3v/6dRE38cEh4TgUAenMbaHQmHezFfDdvmv
+b8dNWq0bceKGlPOaRF/VkkbLZRGWxnMpNL97sD5B2pULd2ZTVdP4G6UlfHTqzJsMj97g83bN8H2
cXqEMhB9y96wjl1gK7mTFlOfs806/AJGsM7A7jCC6gEaH4GG1GWhhtoRn2YIB7bkgdfUtQ7tIAw8
BTPglM/WSOUzA4QA8wV+pOC1V24uqsw00V+FKRq3VhYMo2Ly5tUu2gzwFcIm7lMJsjzUMa4Ml7zJ
t0AjjVGeYA+kjWyGdf+Hw8hMNnnYtD99iMpeSwDBTNjPO1pF8gv1YLXuTuVygXjaiCY01INycm19
eI3a+DoR0z7XZP+c3h5DwoirXAUSWjQHhF3wp8SqQGQaEBRO6Dp5gp3pkqFE2mcnKD7l7M5OvWkh
HBqvRKM1QDC0ab7HWivxcYA1slbnfOAOGjlvg2Xnao1EibPFmIYqnaVvvN+vWQt1Z1nc1ZeWX+bp
LVYectKVD+L9AQNqTg0lDGyugEZ5GpX9jYbGhVkgJCaNVAkZ+iHOZUA9x5ut2szOQl2bOpaSB9M+
dcfBSAbxVROmnAJZuNDVOWlPfFabGUdPp0EpyRiRziJUWcwV6EZfT/zO+jJGRQGd0U8S7n5HGQUR
rgn3B6PCyls6+im/1GLmyp3HomcnVt6+iyJjBbAh8+7QlUINHS3qnx0rGSoi7BynWNJX2xJXXivP
GsoBfJe0Ko+q+HQTTiuPxBaf00XKlsH0qO0yW595eS8NXjLV/FRd6U5i6aw1Xkaczekp8CQSD8Q7
xdKxEZSS8lfnhDoaKUd/LR55DQNGgfzPPjij7GKuCGo6jUhl00HSMfuEXmfQfjmQCaWa72Plk+A1
rg9PIF8kXpZZBbqUU8xiSCHQajw+traKNuj8TnH1n9sWhpjvGdhucm8XRNokBxD/MUOS+L1QwTUy
evY8+fBhY7pBE5h7RFVLY1K6dMIaeSBA9LbWvWYZt0+Fwd82xg7rsBUGfEvOJtoqQplpYI/rJ9bs
1LEtjlB7hnRfU3gOdINoG4Ol8nnsGG3MnbDX3aESJ76wDwCOOroA2RsrhBX/V/nlpxWiZifevtkj
sWnclAG/lQ2qwJRHVVlApMXjtCCCoKGRr5htf+2+UgLZjcqxSADWVS63v6DL/ndvB5/LuC1/Tcmd
SeLZnxLGtF5uyrDUel1vpa2Es3l1ns/CkSOqjNF2aInE1NwBUXJHrb/aA14VTEgkgtBw72xYZFiO
9nBUqpCMBr7bsDtwmd+UHJJBgognvAYaK+93gFtEd6umRDkPKVwGxdlys2bhRcNlMAX11GXysEn7
QkU8tJ55wqvQwrXu/jEKzEnCXUY8FdNuQ3Td36l8iXS1S1hh4apIwpFigtaXEZeNhwHSYugwGib+
uDLQyDJV7MT3U0hp2On6Yz88i/aP5e+C51lqkdg8R88+6DUBtWnHdKY1RRfxqKcWQMgvEe09pUMg
D0XpMfkK3IcihLul4Y8x4QoKTiEMzbQW1DONGD0Eb0I1X2rDkeJMzVIk3D2Elq/m8piCecmuCJoh
X4BVlb6wHF17x8rkF8G1l/2ZuXCpy6OxoZV8LFsqz+mZFkZp3EWm01vI/kp6RJ4OjQ8RHIQ/+NlO
5Ymm7Zu98HsOqmH92WxVXzhfSZP8jJd1l99AsSTh8TAt78lxDEHHGUkAXOGz3FWA5FsJzZ9WDOM1
aOuhhkq0Lpxi1HvUfJ5ZPEhCcaHs1Bz12yZuIfHdMVFz6ByXwXqTpZYCCgTOv9NoM2BvE1eMoSXp
0lI8lP1Zf47TNIBJPn7IRGgfZSaXQ6tWpacDyapbcpAIAyVLllbHXwnYFVzF2my2shvJ8Gwy5lRG
SDjbsHGr20/duyT16i+YPdsYA1wmRw1TKMlwVXwHMqWl2bUwi5bDn5aeTUi1j+MkIVFe3+Q/tXHg
DvUkfQJj4QWVVDpGYIKsTsh0BhyzD6zEdRyDHhCSilUr83fCjqE+jIfPxmM0MTpBIbuANu9tA3ZE
Ia/I0LcYlZ0E8QscuCWXEbyHmgDG/rphZCTvjh95vI6xUt2noqKnAempekoLkMyfAmfZp7BtI8RQ
KR+IojXr6yx0cC91H4/VkLJMCF3HMcXfM0080SxFvuGlOReasVnZSmVb88tNZ+WCsBNbK17EWCGa
0/BeWMuKpAxm3Dnv0fxYc14BFC/ouoKuKAZCc3VO+EtYTEIUGeD6We+VZNwO47izPNOe3eruaVnC
kXqgVlBTLt+HDyjn7x6JQNdUA6AvhTHDNM9WFqjUVQMNpgMlgisl7YYz0ktXazwoN27Z6SDQsuva
C09KO4P7jLDYSRsP1bgPTCRFlcH9FqMDHNsFbDGnJvd3Xd5/C9B4F9xTwOpUl1XCZnWfVU7tVPJy
F+TLqb7wD+vDWatq1R1zZQx8VZVnWyQZ3RsbFHTc47S0qZfc/F2CTRfNY4+bdLo+UQz76Ico3/Wy
WctMXQgOgoLj3jtgUzpl3KFTzqeu+z3STPCUJqJYyc46g6viDD/FBtJJZf3q8S957uINN4BVD5i7
t4IrtejKJR/XGJqyoeVA1r/4y65r20SFJAhumsk7p/B73cYKAmdGXD5gAyISqStmtQc/8sQlQ3ZV
TbLRMaU8cvOMVtIsvtwHQJJ7U9x4U2im5AYj6BPmL//MD0Zhc/yRfgW26ReR0K/+flKUQ/CMzo4f
YvGnYClkXl4MX1KKAIMnK6WkWjUuwRieVSTp4AIV9JpIFS+N5mKBE1PEtdd8+6fDfM56zf6WUZSw
2bM4dzEiMvgRLIx/3B0x4FRgBB1oUH7U3Wuw6it3Amq1s4x+Sy7CSEzJY/tEisP9FRoFFMY/0I/J
79+4JLRPiMbm6r1+wv5jAikvJZtIGCCd0Sh+7PVGtsx1fWwvEd7zTCUIiyjE3C6khwE+ElfZqZ7y
RZARxNvOT3tcVhzpOot/TWLFo2bBBV1e2rV5+aAIWp6PY2Jo1qG+XprG9JA+BqqDYhea7er46bGU
d7rTgeFSYg85MA4Drrbs6IkVWFYDCCQIqQaa6rRdh/UwDqAh/5tChw9gitaKQTPlSUnrwzn1XwKc
KgRCP7aDiZdsa7498IYLrWZLbuQmKZPqplK4nbJHJz63d0olKsEHxn87+vKEkjC0dGrNI1C1ETcg
TEJB0/g3EQ5CgWSZLf2FHO40Imqe+5HTlNRpeLGe7tmdiv+OLVVgxWmrXRHieRWm0iqHqTc/1m3b
hvaxAFI3wOoKGhQ1V+qH62LDfWFWbZMUx3VQQXUdRFwSUO4AG+hd1sc7NXL3suC6Yx170dv5ZlKh
d44E1WniSwTS3RsHl+61oCHB4HcCoRnqY6XLYGWMA97Jw4Q8Q9jf6XhpOAShJ8UZOXzvmM5DthIZ
Wjg9JoF0yquFeTjWQkeRukWNUUkv4HUzBvcntHoY+Q9kh/8rFnuQqE3ozt2TdiK6heXj+4CunEBU
UD818fFdf0cvQIVuNjGGc6QKop3gUwmJHAFAufwLHjT+jEj6wUyBVb0sDnjIgrTG96x3bGvN/iW1
7AmkrdWFZ3ToIBXKkKW6tc/T/hHxV74MOgLwSXSaMrajd5tWu6VwrX599obeC4oXRLuU8xhUHdGb
mTFQBLjBUxtkcXXhREraq//64KrQgLbWz8iBN9rUZcLwAuvnK5ZIwsN/j3/17gVRwjommPA+jD6N
m2aPRH3H5XnUN6tzfH+FrPeiYuqD/pn48eB/TZaoNKU9+eh6KtasIBDnEPGgeGri54u36JGavyyB
qtFKWTYpUdrTviDaucViZ2wMZMKNAmUy0lmkw3ng0c1t8CYAjsnm5HE68QOF/HOiyI3dGi0uwec2
EqsYR/dnEczDjX9/4XvYIfKK2JF14E74r+38vARK3bPOUFJeusAO0+8JXSlMKTu96qpDLpTXQr2Q
dAq91aiWZ28BEwk/hmnNeD+ysMjkiIOafb2NrkqUHbytLs6/ZSWJMloTQbaVjGPF9bvUd/Bhi8si
x9OBGrk1dbXuwgroLzYDlnK2Hu5ZZeD0u4YveV78P1YQJysjt1Aizqd54MfG03K8yTyNDLIUSgG2
vQd3F5ZzAOigmDKgIwnq8gnDDeciGsCqqVw5zsbNzHZQlmpxtxQ/HvNKO4qLBvqdH7W/DSHARtib
OP/7s0qLOo93CBlNtzwDlPwlvqjuCCz446s9hcRK/SmqiSdXxtWM0uqikyM10qr+Ni5JobOU456C
Wm/uCfRIGOE6D17qGExNdN7TcKi9u1I5YW4/IaMIzRAa1MppHA5JhNTNyeIkL9EY1L4r2r/+ETiu
mvSFwMFvKAVoGWvb+pAgONet43uS4d9OuPbwUGilpHPhNRlwb/Za0rWot6yLezzzUrSIT0p/V9dr
vPAlBl7zMu/MWVHNnC2Sgbxjy4SzA8TQmH+TL6bWT7En9bUKC/fjPvYPx69Gp70KqGPz9MMMDFbl
uzTqaRM3EXDYZOctDXXKVOH3JxMrhdoHUQaWE1vZtq3/Sapa9735YXxV0Y0BddkIfnsjBc8D8DW3
lmlPidrPKsf3Vw29wwUw3u2rSzmKGG4YYbucMn0H10EqHSRULKV6ek1vEzIbLPvfXElt3KoVmdFf
6s5AsExef7UsHPA/1yA7BQmh0BtW9cHRas3YKaTSartNRTjzEMh5MNtBDkc0LaFGzqblC5ARyzZQ
xUdJ0RQkQmOO8RSATl0sUy2kjH3x0QsKgbDD7B3Ilcdel5pot4XBGI5VLY7WMzJ8a7fEFQxN/biF
w8TqPb7zbkeLeWIgQDavh9/u+2v4P0W5uuqRFegNAVfqqCR6KAF/W/+4ul7/It4hNFS6CjMfOxjJ
ci7MTuTW8ItmHb2K7pse3Y+q5VlVZzDlVsHyywCmclaqwuSAv/5XsA19oNizgWQjVG59LUwZA121
c1puFmDaoSP35HnN+i10uczK/haT9XWR06Lb+V45pMfmkIxpilBcRi7T1sTPETzBvVetU5OWxj7e
Sr0SqTl8x5bPdKKSE1KpNh8JdzmjhiyVFrmtzb1qaUT/ilS6a+Mr0oalZhAoYkadMYMwtp+iCC/1
XliIsF5BUn94c444zX7+fqUcmM8iVBwmLfP5IpXpgT4LzdgdrmEuqNvWVq4gXD2ICA2brRbr57Ho
JAVT4awh7AdBNcrHxCVyVD6GixU33ml3eKh8n4EQY0wQ12BSzMbsDYGCM8F3+yYbheZrsB61WE4Z
t44GWg5h9eQ2yjdsuoa3SVrT/9tEq5vQLxgmR5ibU/Q68e0T7orjdCUy0lJwxCMkLxpAurfOB4V/
MkmnUBTnh4Y+2f//WSubSSrG2NVtCyIU+8GgXcjgPgB6VGNyiz5CMl4WDX84/8cwiJD0h+L2SYCR
ahsUnqybNgNaZz9YefmeJ5hG1id+T9WFhuH4wYFcnVrc6odu01I1v2eBG75vGSz997kvBkgIcDp6
Oh1z2ZaNbwUIOfUmzCs7/6QSJmZmwPoLwe6U7gBtuJc3SnaypzQKoNusZ/0H9oroUBKh9pLXGTGX
8kFCjfFDd30WErtciQDkPFnruoa8DhtJujQC9PpgqdqlbnOzczcQmzECa75GBd7va3gZ+t5mWH8C
BZ4GJcmSk8T6lbL6ZDjLtaHBhog6SRQpHuDlVLIAJXSv2AgYXeVxwTqpTdXDmaZqlqU8aLW/oIPD
F+bMCOocmxTIogR19wyoWz+83MNnW2WOW0xHqRK9T62D1yml+8uYWKbPpEVLlZFhgaI+jLQbO0s8
ybmsVTGCkr1mEultfjiArRnPnIglm4WmGyymSchzHKm4/wQUFupdaWtfqo3YSwMW515Zeu6gTGmA
1op55uo7Cb1lMjYQQDBzGLNxRMgTk0EZHix5qmMZ3Ns2a2wlFBX7p8UCbMbhKkIXy4MkPUy9jxGS
i4rZXnPKzSrFSmGgeqiiAG12rdPf6DisU5RJ2KPAZUCtvN1IzRX2jZSJk7NAtrfQRhm5bM2HyfwN
UNgGB15Js1Oufmwcfyg0iAS829UV5B8co3KQHTkBHRderociWfzF/1CTIeb0MYorVMRMKECnLnbs
l/rL6x+VWTRbD0NOovxc88NLorO3niYyqr6MSwLpIO9tAmtGMXBHxgViekedgTEKONWZwE56GaO6
pbiAmPhd5Co6/M29CR07H7crbGT3H+rBaoWhRwNUPpsqtqF7HlN4ADxAispC2JvvNDeR7aeudTAe
Y2xKw+lwRr1rxqoDdRn+tG58HxS8orRZ++i3ocyOTAQTnjB5bbMlscihD/m9FkuspzNlyXtUVy6b
NDC9AxalKdWJYCBjRvfIVw4s/CAUrui9dHec2m9Do5t34/eiXODJ4/8gaDNGkFU35OgDejiug34G
GxieRLyUvQ0Ax0UaxE2VmibQnCdUr0FZ2AAzbOs27aFbm+XIwCj2NI0Aycxquk6gPkkQi9tKOwsy
WjWKIi1YQWp2V7Utp9tkzbvpiSyvTvRFBYHUQkOPHIrsvbQMBX/RvEW98nionLhhb4NGaxNtMmkE
s/sEvIzr8vc0X+kvK0ugS22OPnk27sxti9QR1CkpjmD7504KmtZaNZ9cBqL/t1xtP01UnbnlRe0L
cAPRI+Ugdfj8jgd3PygxrHf8VHcwREmCIbuIlWaQ4BgXJZV2nJyISRq8yv+2C6pMfkb+3XdOx66S
sE+hNA9Dlg71j98fAs5wxC/miwK1txzj0x60TDJQCus3bKP/7Derahl4y8JN3aplWH3wlBE+IP4L
jIJSw5zSTZp9D4xlfTBaPQ8ab8/XUSuIZPSb+UsW1RmTLU0kjT/FZjvyeHqYdUnYCD0x9G0FRre/
hm3+SYLc0OUh5DVByxhDnpmNw7oq2E5vVSah1pv78dmJ4vib5YfjJCPR9kPXDE0NoEV7Ve2SXi13
TeFG1peA4I0B64GUwwyVIqGsVQ1HTk1Dz92lPP2yfVrYCdSanfzdUlc1aO29MwNWiBGpAxU+/igm
EvI/Aqe9vDPMtM9TSjkv/jnaGAtmusqftIUVEWzs6ZkAbqi+XG24j9bp0GJcd/tiqge8QTgF6sxA
McPZv52Eqkmm7lWUX9HDzy+NNAE3TjeFrx7H5f7WPzgnBGF5TWet3nmyqy0wY40hKNIsvF+Ph9Ga
kI3bz6JJFNoxsq7EYSGh+fv0aSxKpTAb/PPc9iXbV5a17KaStBA9rMPJhfQ6geulkAXWPtDcTKhe
x0eHTNk0977tfxDDv6tAYlcQIrUYBT6fmHc+DvzuJKMrCG7rjf3Mw48LaMu5U7rTnaiRZBertbo9
RDLfc9sd/XB6qE8j9POYLZy9s2ubBpbQRO6dLM1NBw9YuoBpx+BpQ9WYP0qpMmB2IRzQrOZMGXA8
qPd45whB20x8dk6tTt0UzQPAd3B3Z4t2D20Y5rCnMCZmvjQGCt0d1XjjrcvwruStIG0ibEiOrfIO
GY/soTNqmnr4cuPFQ0RNSS/1fA1NMAyaY4zNPDTwzPF1rB6qM6zaBNXgL/XI5lYRhqoBRjgCLs5L
BIvIg9FFlkeGQyE2RGchVr9r5EPLUOK1p9/PhGDJasGIzrYRue7MofinfX7lMaFbXAgIoJwXE7mP
yH6lXIH7l3yN+Jj0bXNlAWiCJdNtRaSpnzDTCj+8J3rCHfkFeDj4REGYXFzGYrYAxAaYQ4jMd9Y+
In9eiTdBd5Sd2gr4+zquFp288Gsc/eDPzZXlZKV7XzH3lIMDStgcsZLXGdBY8zPf4an97O3C69r8
PXaYCzLIsUhGeK+gr4C2jW3PI+twVSEx3mXLpPiJMOzM3LrugqaN5nTX8kYssT2fGZ8KhTUiWPLi
xYc+AYQ5HJbWNcnvgdc9JYricQ7Dt6LrcwDpnaW/bxu5xTE2e9h4gd1aVIl6QIwjquFVhlt+IJzQ
E7RKSvU31mSFn4UE5pbCOM55s+kMSZdx/hgFFacj8Q6HNImUd6HODHn5G8jjwkIhdtQCemxy5YYK
lOyNmbIMG4tLLSRIjGpn1+iay36fFfIN3jvrO30StXDSFWg2OismUV/lLQkFfX79ZOveR0qRGoog
SsV+95RZU0QPwr3/b6jkaLStAUSZC0RU0YP0r1jkOFae4PP9/dlkOG2UKKQbgk654Bsow9wE3rxh
OoG8PPAlZkZWiDFeFhaF/UZQi3Wq0k+foVR3LfcdaZt0YVXIe8xmBV1cdgdY514jSwWfIirIMEtu
puRzYG8ZpXpxVC1JmYH1WnVisQCs34fPrRZI2YGDml5J0nvvq2NKfwGaEaQSD4kTEvcZIAhX5q5t
m8avm8dj16RTlL1Q1DSQggUkkCTeMbtamabyAs3vzKlg+QGRDaaNqcBhjXINp2Wo0E+npCGEjT19
VS1U8LluOHiMrQ5KNnUY8uD24ltIi5HlttE/ww32R364hJROaVTyO+Fi9nAyfIpU8aVhsMraSjHc
r5KJlcLRUISJzW4foaaaPSAQTTVF0G/mcR+/JDhdmhgsjasufSiB2UOK1CgAIdCVEVv3Tx7PM1TB
neA53TQ9Nq4NSF0mAahGAVame1N++7uQgbYLO6HnY/B+/mBKAKjuU9Ylrh0rdaxJTJOO+NjAcVm0
THxrAJFpj2hg7VwPASkbNY83EQ5iZODDvQGKi5QHoMSNwgu8gMt5yMFlmXRPFGvuKAE3WHzFAL2o
UntbDnCXrnlISC1gNXVm6/7RzkIEmWuu4GPpCUZhRwtUMVFrm5ikt+IuzZjSSrpgEdU/WfWcCtds
Lp3CPPzzi+TCVQ74BXhL4auwK09YklAonKVOErVqUJR66rr891uyVpnx2q4FDRVPcVSzvoBeqnAz
mWabppsUnFQYvo2t8VsZrZCe6M9azBuih00j4MUxZ8bm6JImcwF4QNtBoN0oxp84z75x/M/+G2zG
J5Hj0LOtudYfB0EhNPjLooaweDEBvPJDjT8cNO8wxItbqdPmAFNp/frwQTr5e89+Uv1YwSvMULrE
1Bnlxhx3oQ1JvLpHZgbhLAysHFS7wR2Jgv9UzSbJbwh/Efgug0CVAAPGxRAhW9bHIrukysJC9NgU
XUBbgbuqXOXi7ZLzQg1T+Tkc571NQcSgPUbOaFjXe3E1exTa4pfWLVO1w0276yQJ7UuG7wHWQ0hw
LDo16H4fovKkdDRcxlcRUh4jQL3kIAFsIolpdiay5xd/gMgvM5EduAHSjhPMBAojGdZ95Dbl2fNV
XTA4JzZGaVpJgKzYcpN9XSA62lNBvEPuqJGvcOjuq2UWDiD7fQ7MdiU+TtPebBuiUFvLjIukF+AV
/+nEec3OzN0RU4SfdPcaj+DO0edf7f41PMcKzKT2hMDgDFPpjzFGnH0h70ZATGtL257K4X9MHNpt
MfAXZ2ttbjx4s7PhIVdjV8sDyvtZdjFVf8fyatK3upxH9EcRRYpYyI/slL4ulbHycHL0DUkLDg5g
Xt1fRM5V8858l65ULO3qlvUod5PEJExuO2eyH8LA/IDnV9RWNXdtTsd9zwcTYD7vDWV9/Z7XFB+4
EFmmOv8rUdUwfoVV4DBl8h/9lNVC9xo1qmsP3npSIlm2t5B3SVr4uLeB3i4VdEHjlIyS+60RpLkE
tTKnmlvu60bCCWp2tCyz/Zzuvl9GhSqoVwHrgVWesIYWkARK12iNftbLUfkGrzcExKrCsTj4TBsC
3XEQiG6k393ygldI66070OOOgjtglHsSyhgzrFyKERaxuNUU9PQFa1RhXClet/Uv+YAsepMaMDGm
iD7/6yK8KI4YYc8hqrBJrRzMqGld5WSWSjwMgcXLXrLCd3zAPeTTDx4kQnHvozVXSm8GQBlAT5qg
A2BKixIl/H3FFJf/nb1fV9wE3SCu3YNw7ffNxVdXG9IXv1jMYtV231d4eR284yuR8zo89bkylxrr
JrgqQPHMz3fEtq86E+i2Z8VtZA71A/qvfRKhbhRv50EWrscIGbLgYCKEnN7aZw7+pzNXV6KFkGxz
uSvAHUk4lY5Mxx3YuxlxCSID+8OuZkfRT+Y7+94Xb1/hCLm30KpMe2/pl8MrZPfGZhxtzRQ9HF51
BxbOiGAlZts4SNAuV+Izs03cZV6Zm3LEjw/oVFKpQtLU+/hSpn2nPyN4ebQRtkwZ/3PcgZ/klpeF
pgQF8E0wQOm5+EYDC/wPo4m+3H0CF6eCqy350FqT2K8MAebgZgoahDZuCTBUH70P8Q8knFVMBlAQ
6bnEbuIXU2l+/lhrjPGYUBtQAzo5bwZLoC8r56DaH+9ewIMcyKddZM2yKXlfdA7tQRjOyYjtP4eo
VFJRIx1zkXT2X0LTOJQ1ZpbfrxPVcvuLOOmiyxvkYTTwNxawPeM5koWHBn/RYN506lh01GGU23mj
vm5Sw2onNzt9AO8a8uMGWScyMJGBTR0IiNoH8MBN7ECEsDzpl+JmYXU0EoF87usP7FQjpA4A6ciP
QspturYmrVw9pPR2RrEKCPZAQyQfiVbNY2m2FBYgW0eDDWmlkPYObFDqzly4QMx/jpSnqtIYkUD/
5If0deKp9FSB+vXJ/oEp43k06+Yg6Qf7IAoW1/NaX1dIWzY7JCljm2TRtzQ8ccV0IzfZXZmJNrTv
1cgsOrR7d0/MmK9YJbhFiz8Mb/fty7Xriy2N/ZgUCPJLHtS+HpNqIr9XXj2a7m2EwDUpKIhPbXM1
8yNw6FFN3yhekLlAx3Y7ibbx6EZKb+ZzUge7IYjD4OjX3iqvng/Zdd4pp7z+78eDoBpr/Ohzv+1Y
KAzqzo0XT2DXUM8x4q/3/AOKHr59S3Y6eqElaHTfPHPao3nuwOJbiZeIKnV2l12mDkK+vQWvzBzW
9yn7nbj/91ft4fIP3SC8G3EYEynf0BwVmU8Uqfq0I6crHoz+0QkatG7VOGmJtznPLyPxKMPTAsl6
p6FLNzFzoGgp/wpuxsZURXngj8LOoUFUPvDIRzudCz667vIfek92eYiVMdL8f7PeXJlZPD/mG/TR
md+/Klz2H1d6cZrfEGhBl1QPWJfSvW5T9cVwKBh508RNKVsmMAOjZ538Dp9tAKxYAQZQXqJrA94r
jw6sQVRbbZG53woF3pfScuL3DumWiwluxENf1rGDob7ZA1+RkkI/sIe+qztBiG6rRd/6UTnktfvh
Wccgb/k1kwEphS37l0HWyJcZ5EWxluujAQYUL5kN0BW/5Ocg28onFwVIeWObwXj4PCxElKW/qI7q
UvsnMBvcuv+NAv2LAVX3p3oWUhfCyss9019Se5Ou9kUbNdI1ewHWWdh+64vM4FksdlDpnZ2LYFcu
pD4E1St6o2GSzOKhRUbrad9SWWLveiZY/aCMoPY9VOujMnkfzElwCpxKW8/hmeyBv3eVx4WEIPbz
gdN0Gl8SIzfFcqksyJomerCe0epEtCA8RsIPLrmpclTJOnvj0zY5w+SWrKUBQcZUCTpWs0VclIcK
s9O8qO9QI1qoWbvrSCOv5JzN9qwbAn3+JCPe0qe5sqYJ4kbz+dqQnaGAsEW5Rn7q23iFsMSHRbvo
ZPh3GrGxpLhVs96RRUF+bh63E51gC98vwaOKnyCQS2ydUta2f8c39MS0WRx9d6+eHBZjP/gfCX8i
LGt9Kc1nvyWDqwfDdTgUtq0HutL6dyfrc3g9UpZ5nwzWJQef4fS4KIgt1TJ6NLArldjsuUNatMU5
VU7g7HccBiVBjRzLI5GxNrLUb8Wiqj3lmRmN1vI+kIDY7zNY8ENhFnP8jCe3k6y3++D71fJfn5Hp
4Trdh8aRxmtIpCe8dHrDhu40DsVwTkKVggu78e2YVPKwmIyQLcsx5xYmj/E10f9SI3g0Wf7mWe2G
DvZlb1tQ7NzU1Vt5DsKmvu1P+V4VO6oGjx2/3gYLVdntRztNutYhg+zu/5Q4sCLuPW5mp4Yy12nm
bipf8dtEOMzlu9ffPA+bIEiC61rnXCdasj8/CVvpM1A0RecDQSh8Gpy2/7ojx7BqRC5TPwO0lnnK
0a16hFBK4B41fODKYU5V4UTUDLHe9KnTAJj09GL7xk8a0az6No0cYOYxugD0sfT0k5YJq9BEIrDZ
p9axEPp56KbnD/RiDoeMQdtrBw0CkaaDvpHJpI6zJyQqtVsFCbHS/icVEjUujD4rINHcvDZ4St/K
BWC8xQvH5wmdxihlr90BxMMEVvrwdfRV72roPG7kHPLZ/hdSCo5dLAvw4cCGnvYZEYRl8p54CqT5
ZCFhMp3RvN88OyPy+zTH+z8BOGFx8Z+n4YfmVPJo3xh9C6ozl30rvcuSb+mRXnsaxq9IjMnoI5rr
e0MW2f96GHcrC6rckVaWt341rdQccMgFSZUDeBF4IqyAvn1vjFJRl9awPKncTUozujhHodNrBTTa
4RCeN2SjSgZjCwVC5Q7Wpl4U/Uyj+ByAvPwkv3ob1v2YvoMWCFPCynY0h2+RAr0VDz+/MTmvJLwJ
bPXXA6xzVQHAL6IOGZSny3/L1L9ztCe9200D1uHsWdPeAVb1EZ7Ygjp3g8C7iGGaqJohUCf1gGFz
C0sNH3xcxWyMm49sGvovN7BRWYrfwxe6WlKgbugP3s7t/fmY53Er7AGjJISElMTTWoG5tCtHmXc+
HgPCH1pqYMf97zmfvf71e2QCknoSQ9uvpWh6bHX4x6UWaO6jc3HNKTd15lmJE5g7t8zALkWXDQN4
CoWy65v0Xo3bhsZ2OKn7vwcePCdNViPy9jr9V+IJTGnCN3VAa/N8iOIPx3+lyimziL7teflqGqKw
b/pmqMTyaV9OPL7GUvRa8skcEG0wt1GDRiErjn4GzCe9N67QEaGnplv5UARCRKItKPUys8qN4M9j
lS0M6TtYPdqAO4/ZIWFFKpRz58n7/On6rOU0Ea5WcUDABe7wMamtkEqhfVwAhD6mMoULYu9TmG2P
LxEq0XlOJTH6e/4fPm5GPEGdrxaKGhA+EW7RmLq5CyneJ/VDNfLGzJMVrundp1nk0/XTnx/mq9GR
GhQMwPZ8CjB/y5AszIGuEiKV3BCQOlrBtQqtw9mZrR5SanTtuf6ZAqaG1ouRMXOKteFSa2LMOXVC
77e72crEMKpyzjWhN1ubgrsImmAJ+tHycr+y/YAPpB2yoTlSJKqxeMi81+nzljIZExi6+PJ6uoUV
vBDMACoDydrfoyVXKHIum64ZnEig2le6N3gnYo6jfoXueKl2C0HScRI/lIROGD+FkAVKhRRvenDT
WmgqhVS/9DDjSHxm6PLRea0cWibVuDFoir18Znew7t0yL+IBcKW6cbIstDhJE3yAMQp3TFm3D6tI
qpS2Rqsbxry8gcTvRfVZduKi9B+8C7ShYsfd/fY92jAEwjhoFyXdldJdQE3PWjZOvNMom+G+LHdu
4/FqJIQJK5OyN0/U4DOQe4n8xVDjQkr4UTFsLX4uEmR0tGK2/9mfX0pSwktr38gNGAZFJ9Bz7PYj
E8wK6BrJCc5UJbTevL74K0hfhIaumTYFFWJRmmkdCGcD802/uew3oyTpiqMCDmwbkFhXRm9Qp3z1
uhUMHpmW3asAD+R/8XLhRdguZjsS3LYn0TuKn4BBM8zxsEC6yyya9a31SdsUXLuvhwSdky5GXPRS
7yGjNVcHztzS0+z2i7eKbdo0C0FBjFFvMRm1xsBbSSEQQOF3sHk3lUUm9YbZf8BVy4J/gN+9bI/k
/pHbi9mIAtjWAuhMzbEGL/mbSlqzsJCSmE35uyA0gAWiR+p8blry+frzB+GcHYISjIFxZKtii3l1
nN4yPKpVzRJ4gMae5aYIceDvLWvisNDyAQKrbKttWC0VWrINLTTtTbALr2exXbicvPk40AL8NlE/
3PNhXpjWX5gnSu4S/FOs3zWT00WKV9F4PSMPag99j1WIZpqr4gmtycN1DmAvowNfCfxcXwkyCj9I
O6ljkJm3/lxj92cr5P3roJhyZ/djIuEJhjlw2K4y5MyskZ8w2+jLxS6U+tAU4hfutAZglziOpM1n
EWkK8DY+0ziaiZ9m3QkoQw3qL96Ivfr+7k1RcTpr73dXC7f4RiXZ2G0/rclIBtKhIvtJsFpBslcj
dX1c5Rp41cL6WePM543EfUt9KdLAPrxQR05aaaCw90dkQpRutim2CMSZfNeJx3VEc1sXyXA865dI
ULlvf0bboWU9sITvFVGVfUFGslwfzUW/Puy1J7g6QYidNQ6on52KKG1mVdQ/Cz92MU+PyyCt4qvk
J2nFPw5v3YiiliVnHO+v5EAztE0NVCTYY5+aShQqwElO4cyB61qbkqfCKLH/i8gXONyE/5E1UQlS
JvCtPz3yGlttIyWVvhxPVtlCMPR6sd8X/Iyhp6GgGzPJY2hCOIr1TKsTBarXxKo5RKhlczVLaV0m
Q9oj053WdlM4kmfL72hTVpqmw/eDyDjw3l0cDlWYetsAnNwrrwwuUKrP6liryy6wx+HNHn02WyzW
NSMo72sl9+CIDfSEcH5xP/qjM6V8Oz5dM0+UcUOQM0/ZdfHMKBCGPrsEByKdrUF+ugBUx1HHjJKO
tnsZLOyxqj+FlN8S7dMvbA2iLUzhU89skUWgi6x8EDkAQVqWgO7GN/4owROf2TS9vDsGYFVV/VJl
zUT+vlyDl1wU1ICmOyRk9X2drVT0eUr1Tp+yqClcLWJXMrUwJ8OkHEJIIgkRmc5zTGpfT4GWvKXd
fgUO08ZFcTv4hYVeqEQSlEoAG19OxHiQ3j7DYQHXZEE9G4hgnyWYSPmMlgH9W5FI7SWxCXJiU+w5
q7Y4DUa16l3FECsF1HXAQtUg/hH3CTzEIy0gwAdU2XdZB/kMuzoUpuUOq6U0W1vdZ02muBVOKBa3
cfTWW+bmiut+LGG+XN6s3AfsgAj4w1BLb2b+DVuzOTnr7sf77ROLBm+TYqW4IYYK12BwVWMfrArV
mrswlHNxbFAOG7Sbw+5ynDjWK4zE2Gol4O3jENWrrxPu4ZZKP/w7KXFEHp0hBbWS3y01hsT46p2w
5rcsyK4X/JTLKbUaYCGmf9a7CFGXlw6uBW94PeAtSaPMiUSuRhX3GBdFwn2gVUxaVI3DEsqA/gM9
7ivppg+OYL7EI5nk8fWuHZKZzQlDe/snaPn2xHCxiXLoL0G5ohnm4r+hb+NDQvHWsh8EJB/aNgNL
rnFRsgWzWlMtU5y8JeNe/L8chNaCPK4rEK6pN3DHAkNuJu1rfjQt1a9sRUkSz+dCb31lziXCvKYA
mKNMmqM8cGAJKimVBPEoHaIPgqf1vXefVcMAXXpGv8Jz31qNzQrsz6dXTPo4MQwyryid2h0DaZl0
YK+dTYHztca6+cYuJZNjftg6fHRIouSJl8krdqZMzbbEbOG520TSxKNt/PSWzXRgRzE/7z35sDuD
Aq25DEkYO8+yBNL72/xV/HtjIi9CuwB4l7ErR68w8G1HHEkclNdBewYU/cKUg8Bs0PikgE1ZHhvD
J9Dvh45tXheAfIyzHXgucbY1Cg9yeCCy3ZIwGsv2xemEcqQjYaPSHwJlKcanwDYcZlsAwaSAo1Df
OFMH+djkqvz9dVNEBVD+I6BKp9mhbedkN3LkIsawr2rvVilX/qd7QTXIW3ygKXj5GoU3W4MHycc9
BjO7ZDBK96utj0O3Eq7KeiKOXFMhbf8nPfkVUscIA/9XvlSEXguiobLXHoFjrOQN8ibcRKV1LCCH
hV3SUOjGAnzCYBhQi5y17RdctNZ2y7UAupKGUpjIgPo1pKSh/dfsm+0ar/JQIrg9O5qxsH+tWYXQ
ZhRGlHzSLZn3+kc6x1c3CXzAoindkMtk44p6mX/eDWa4/IzJr1bv91npZx/Uj0yMz42u4Tg8Mpn5
UA+EdnfeRMJmkRv9XL7MaTsnb3OcC/hUCybRPT0+Hq6a+bZYU3BT/YsE5ImqpbXEAUx6RvapeWjD
Fdn3oqb0uF17kOCQyBK9WCZqkuJLoDvh++ScU03EWVmBTSzg8RUxV1hydLQ/9Ve0RzB4vKvI50WI
ea5hAJSV48GqOhgSyMySxOw4+YoJgD7lrIz0SJa/lkilf8FDHBucglnRO7VhApRr9wk3HtB6fW2F
uamGqznwzFjCEQU8Ijt8gDW7e3sMuhX0bCllh5yUFbAHUDfhIOgFjJY3aXWTed3aQVNmLj0BRWqv
etHJtx/7kSGg39cp6M8JgvuU6BiVC0ToC2bpyMUfIuu0oe7LoSHSZTS3dR70Nsc6tvsZkpw3X/iQ
BnqAfT4q8XQi+b2gHeOzg61F8nigdornEhQZkHK8VxEd04xdoOHJpcehq7JMTJjlQbml21g68zQD
0X5KYj2hPA6tDJrX5dX2862NtIimxPNoGVZGHmpYaBffRdznzHMlPD+P0468vRyC16188sfavP4X
n8LjD5GaBgLopLQ2CO+v6g6rQOSgMp8MJ1ky62Vk+qguhMFwLWmgBiRLVkG73dZwN6PFduKefwr1
nJ8hYPUeD2/bx8q8BR7kOhhNE9e6USRV7pjy5wK/X/ehR3hiT7h0hN4qs1EgvFxO5P7/xUfgjgBk
+IIQWf778v+phSh0rGJ0+LTInbcQuvH93elP3REKW3wVU2UnJbbgDD7rUcPf03vInnqaE3LrETpN
8mNY6LbPf6HXGzISmzwu/uyOYbWZiy8NG3cPYhJsBxzlodlHo8xGV5HvVXayFbPsMpMsJbR92Zsb
bq/3s8hmY8Tl44Sw4cF5SBYRfgZSXWe0KQwQlqiTSJ7uCrW6it7Lz828HzjBnCTbaiidByuwvYqr
xcgE1aLAmg5s/h0L8/8Yflkhn5mjmq83zvdZbKGCDhr8T5LwFG9pgHMkP1qvrHazvJy2EC3USNhs
6nKN0/sIOEWCNBygvhQvC6aLOSBYoRSiji5KxGx1ae5c7r1QvDo+b904k3528r3UtMrziB7kym0l
jRxpgkF1bz/5r0nBopgvkuMEluy7w75/e2okWxu3xJbkRxR3OAzURotYfcQSMVi6AvOFWmnlEMh3
9oxBgsHkZEr8NxPPVxc3ga313Rw5Mg9En7SCqFCNATSPqjeSusADTQkqXe4FCq+2lV6WXlLoDfVB
6mEbbQzjb/dcbai9vqupKawenTsLIw/SCcOES/EjrAVWMmDLBZBfk/Fo6mEJ54m+m4pk9PyJr6EH
hczL/Vpviol3lcFPwLwLKU40dGmKAEhAhwKYF4iC4uUUK37I/025xxLaLAgZpuOhjdCEnWQ64/jO
SZ+dnpDk3jUZVsupp4rb5ClGND8y5U5Tdu+BEgGfdUmDwHFVd9vfHIQWtCIJk3JgQ3D4OwsB/sOv
h9VcDV6S47yfXGlEHrfo+0qwWP96Czs0XhvSn43Bt/x62nv+nUoTHh8H4FURThm3tOzmI+iRzVWD
HrruG9XxDnEv3R52VONTSrfwGU5WzQZnii4h9kUSj+wXVv7ian+H+5Jp1A7wqVhk872jnumcg8Sb
IyBtEyzRvOEF1t5d9La96/nTbvWGXsB2SXD2+nq/t/SvCkL9xQgAvOohZoYtymGEDvg8ecm2/oVy
lhIujiUWDj6KzO13jXmeIwmMZ75jR7nWKrE48KI3CWziDofesIRRD542hf+c5ICSJbWdkIWexeH4
PZie7bHYkXdQxMGj1NoRqO4IaVAKumC6CIYR5wU6wdZGOlJou+ciRupQjIw2M2NRVRoNEmKBRBrz
9w6BupPuD7NUd9CRA7+43tOYkasU1VraDUXp+Zp/c4mvrrMNFtQhg8PNaCdfD6H6EA8g3oQCwkkx
aEFtbx/w7Iennc6tRFuiQcRHbpXvM27a03v+3xaPcmOxQUvBgXX0YTySMQ+H2xtWRfxTiaWW152w
62hia328mwyhjxUfv788nm9YT1gBXWcjShhtomfU551msvMXeX5uH+VgZGvA7HlhNmYsI1A0M5GV
mm2LNlDJpH36alK9WcH8n22Ve08F/HjOpKXeLvRiFXnprz3YnD/1H9qEaE7Emsd31av4/Mb+8o6W
0IphVilFXu+ds02uj8XrP++h0qtxgUmLgUQz0brZo0EwyhRu1DeJawyfptLRMbLdynaAJwShNmJB
kV25H5Ks5sBcaV+oqgP5xaTPI5vV2YYcEgDliK+ehXwR/hgMCuBij7NWP/Jasiz98bMqFIpbz7xr
rD0k6BWdF2PgYxv2mhCUzEs/Ft0QYfYjU7/vRxDoj4sZ0ofOjBsdpDdtbidtlg+q6Npob4jmekH/
AuiW7a9UbU4T3NUcRYdqGDwnFw769WDSTiwcq5SqNI4ZzIKoxxI8q6eiq+VB+hHpluq0nZ5gEDSw
H68paNN37WoOeLKQBYLtOWnjKHj8D3HKHcUkmXWBWhVZL7mclFsfaTe2B5o3cdtVGbnIqOyB74+F
QcdaciH0+bwrM8YnEF25I+2JI4ybSho3LViWO1ONe3/P+djinLVpqUzumaFBNJPVg5NiDuLnntNM
bnsizq87xNbW977DvpJL8VOlmr2G8ayiVBl9xmklOqqMQfb4sVmFLkxAXO5xXoSoOCSdKyUaSKsK
5pGcJqRu22I9Glp597R6+2nMQ/xD6cdbVPRGanyk/d07rHdxOfbD6dNWXgOp4vBjTc30jeooj0LE
0LQV39w0IZfWZyKsxIvlZorchKYUpgJlObYkfh8xH1FMdDXEZ6IizR3AG1no6rQMQVl6IwUK+0gs
K5dfhzL90vrJLvyhifLBao+j4v62czci2C5vAzfQF4wOWFeo+MpxEONHl62jJP86Jn3rmm+v4SeI
/OMUhUIjfZTWYPYmuFzKJ8VwtPUbuYbj/Vk8bmL8Is31kSR/gvK5DD8eAqpDhVgVNnXb9NbH9sWW
7PBN3VEQc6NaAvg9QJ5KeABIRZpHhFAbPe5+L0tptvoBw8DvBSEEbK14wdxCQtSzFanSSrWQR0p6
2xtF/PtYPFh3XKE6zKJhJMaW3OXBut4EO1eH/RBQOJeDJTihSAKFiyd+v5mQ44qv6WiqgijR6AY9
5nUAF1c4J7NbHEovgYdE7XwjCmVMV/6qbYYSQ8SPiv1Lkh4gbjE+NJudQcgOfOatyWO037zx2qvo
v8R+4WY/MtqKTdCLGlWogRMAE+Ps2TzRhg/nXj8kGbE4e2pXBKeQ1gcP6AIflFCXq3AF0kRNw1GO
qZE9rWQbGWRQvV9IXRiIKLkNsph1MvEj4oFjKg/t+cnUR62omjD24leosma1yK4L41psJN+v5a1d
T6NDApoFoySOgP9l+m5xPbnpZQwih+by8Msc0uC/LEeQ2jP8lo03EvLhcfeD8FsvkxdiLWbU8eVu
Oaz5Cl/gYTczacjtsF9HrYjVRn/VcR0JDwNL6V7jyme+rey0cgcS7VuQx0ojdOaoG03VcFQ2s+Cq
CefWqtA9aU70gj9jT1Pv0nIFKL/U52d5v2RMZ8fsvgS6M5m8wpcPn1G2F2tLoofE7dE6vV5mIHCa
qp8YtOYdZXbWRXMgYxaZIDloE4KjVsHiAQcz/VWmSBK3AE4rVVDfRnuWPQTAV9WXBj9YYWVnok6e
n31pQ1wkocuxRrbyr9gdjmROcvbWZVQsbdKs2rYzXZ0vc75O/aqGixtKMtD25SeTnOAyzv2P92Tl
m+4O7GoVuZVhupeIKhr74AcksVmvvL/9wR3lxJP7RQQQG/xbvjDsIAF5SLJmdQK/PSwB1YyI//yo
u33xxoIRb/yu5lh9d8tVZbgIiLaPa1UV4NxFjONt3GXZrUSbHLYd1PnuwuLxxtbP6s45+xOnSvnG
hxN/dAZymSQEGiMlqT5ucKiELq6YULrWQMur38QGZDdGaL3XYF1FOqjzfk6kWDAvTtr3U7ZG7Zyr
4X0UbJGb2aZBTFG65RT6hQgJVo7HDKyGYNmTTRjSXWCzfCEWsfqR3U0mDYoZg2Gg0b3R0jf9Vkll
EFHZHkpBiGCjxdHzloNfAev8ESx5Q9sonp/0Nt7gjUD+0Hy6ZMGWKy+vHgHYWWbSrKpoKIt52NXL
QA0tC9j88CSy3HezI6WRoK1cjyPbkRHwlHZkUI0X1b7VLC70GBwkb11mgUbwWhTt6NX86nVUMUqM
9mddpYgKOLI59Gui5fBeBPPDZyXo3Vwgx+EfQKqha8fvGHctOY7YQ1CM0L7b5NMQcPK3RgQ4p6R7
pCwtmmXOqHu/NocPPKJ8xlDjMxPsRCWWJqaYXR9TiywzWrqeK1sLyJW1yDA0SkAHd7IINl4PStKA
u29BJe76VxeNEIS/OIz9EG5Swd6AVXMYczFOt+Q1JIUpsppnLXMXgmS4wEmQe4dDb6UT44LLv/Sk
djZhC13mdqfPi5FhxDXKwaFi+KmfUA/LJrIF/NQmMW9UqLQgQxRpcvg5LgE6A3J40DH3j6IxiyAj
RBzvCFa3Gz7l9WkMB4Ff8a53EdcImtclRFAy//t7MYbc98g3UByfYYRMj7TLIIbxnT9CbsQaSr38
qJ7wCE+XrC7rlAMBVIl6WWI60GkHS33/FuyR81Fi/mUTAdR0hJpky0aIPcMSbMMXwqlXkg1/4uxG
UgObapH97NfKiM7F6Ub8F8rU/Jar2EemFr2NxBoa3qC8Dc/vpMPv8+EtWclqnRzAYLOPLO0F5gQF
4QTDb/8hOflo6NMBs8Aga8MkUzkaK06dWtwFqU/i63pvC2FjzFrS/mDXlAA8RBei/zXbez1Ympva
OslKMOdHO3k+6v46lQ1Sb041f82C+dyAGUYu3YecRK28u0kNQXsta5qcW4ox1abH6VRSQ7shrtQz
8iHqbQUfpYMXvgT6Qdu1LwnCD96NyLFDG5ov2Nxc2fg1vB0tXyMpexVwPgySwKj8r1+Pdk/WGPpW
CBty16UJp9UHiuakJHDxquPugXGVsRgdwQmQQ/ebusMu4f144pB9kF1Hz+GBwEewK/gQ5Xs1N9JP
8mI6/iGwduAC6REAZTA7fuOhBTFELi0LVlFR1xGGXx7MFfWJB4fDLK2mA+n8pqaf3qaYnFoceCky
DM/iLiyalQ6NydcZEGp13yZp+3kMVLgync37hJoN0RmorkfnaWIIg84bBgXY6Zwy++QrOo6M8wwH
Nky6jXjx0K6u+Y4hR4WHm5H1kPDNX5P6rzd35YjSgSg0xehhkFb1xtXqCfw1Qr5ABf1o1ZtZRhpv
adBRYTKWSpa+OA8Kaz9/9bWJ5rgoLOV2uCJEEwHCXrfk42i0zpcjIRMFHehqQyiRnYMM+la70PhY
M3KtLwlXiHfTngoMHYXxkNqlk8Ku4tbeYpyZIQiILuslY8lNCEL05mAjxcxJKTDU5pZJ5H8SLKGG
eot2hDPSDCrKjmHe9TVkMQW6aiS+RjRMTQZeN+8g4YE3KwtV1+Y7SknFKUwbNiRxTGd4mEXjJBUI
1sQQj+PCdaCzrd9TXY2n9Isk2hvPtMQ+sEV1XOiO51J/bwiXHQsI785ugvnrxWPI6+570eMcS91k
QM7ZDZNizXcKPB6yXUL1ixMtPE2rocts1x7mal3UxxQ/fPS4xrj2BhI1hf60XkVnFvl1h1jwKcao
iAO703NZYTl5LMNBnpX2QomipeQIEDCFiv2tBUerRX6BaE/4G66tLMrg7/nCEU58FzfKpVRrUkuw
s3rqQY4ybntARJs4pa3bqol7/65n4ibPKPnVEKy3pZd3d7KYveb8ADNiFA8Ym5mq6Ey5Ips7gpEB
nAjk3me7Emt13jKaA6VD9cgs8AeHhaAMeACqVJW34mzyZJUBe8dJZ58ZAqYlx3KviJy7vfM1eFog
+mnqwFVNQ8noZGIoE7YtpzfP8wIGOlzAVjw9HLpzlC3xmSsuCMLYsrJAedrqVB5/y9PI8IpNFVZb
8UeZQ/R6CfsK4m+lCFm5ehAzsOZ4Zwdi78xJAdllwFXl0YqqhL9Nx2LsmfpqycKt/PqMxyFhLZKG
MEbOOa8LOa5MULO2Hq65t1f6rKDi4GC1FiIO33fwOGTXTP9bT+635qglrW7EEmj0hFQgFo6iUE4O
dWm821OjoMBpEhRcrBLCrei5JiXFkroCLLH6c9DJfeyL1be8R6VLURJKt14RMDabF6g+hNozNbqk
2K/NquQOVUwKIvC8G3r2hEdIOt0dJltWOaXW66SDU0yaVPAG7LWIJSWRe9o3a1ZTanLsGsJxlZM7
3WH5gIzi7MVc8FrPy7erplJA/lZPTT+GXLiwaDVKeTG2oIx84cyABCmU+mOuUGRS0gFOT9re4cFX
cJajZ3txEgpD48PRY2fmsKbgY4WQo8gXwzqsxphFKXBpQKL4KNkIIzjLHdPoB94TsC3TqQoVeymc
qqWKV4O45Z2EiFDOlYRjmr6PcC6juiE5P9zrTDchwYxjFGbLHI5n1DXsM/oTjWtpccIfF7K28YZP
ZCC+QWtYDgfAJwxPS9oJHI4t2tR+f9IA21nTy+U9et2wTEHczkvQwGLNy/yqeuft3Nl4NKQe1jrh
FYoa3Aye7RXxit7zbn8HtuAz7qE5zhRDo/8UO5kBC8huJlut1/0dQAFE4tAg1UhlyRK2d5J54cVU
iE/X7Y/wM3gTa7ltupQQvjOhDso2ZFvzExciBG2Fih22+HMNDG23A7GO6H/fiOTGrx3G1n6uQ2jY
8xOzk/M/sf+3TK1PR2EbKBFSfG/qRvj/eaUgcVDRmULbGigggHzOWbBqJpgQ21BwyIML2oWRYuT5
NamLzhyeDBNtgms9W1GSiQyB5qqsGTBz+1ja/ad+Kpt7lx+hH7YTYqqbDBZAmvhnfA9bOl/q51zV
P1iqnA5LdR8Jeq+sdsU2PM31Hhlwf82ehGGfcU4N1kWt+rUQ3NQ+WfaHt/gcYzx7kl47/BzPFWLH
f7xHw3tIH60yOMD8WVp5MkuJCYQK9B/OSHBG4h1g4qan64kLhXhJER31IUDToJOUG974/V1t1vLL
vlhxRdKYVLKfSRgm/qfK3lmJ3mJAWerJWR40eQCW2uMRDJhCbLYSlHdR8IBzSgBbIVEzkvhM7L4W
S1mRST5oH3j7ir8YyUj40z2EazU0L3B9o9getDL6rYpb/9oPBkbdBCFt2YU9athHwe1AlBFjas0Y
KeXDKzewIXDG1oLGLfzfqNfE9NokVwQWH2+4NXyYRVAz07o/554JTL0K8qSTunYyQt513zdlqFD5
cTDqpEJpOd4kxjeTZeRvD1VpoGC5q7YvrCfX95LlNHBZHcGsjvPTfHG2omxmtM42KgQDRTsqq+Eg
qd176PALUkUwVA9RDoOFqBy2jWwB3r3o113rwZH4CcmJsUcNsqpAvgat6H2HAI8EBMfQxR7wc3Fv
XKHgFnnIqerqS+BMBvhiyLeAwMD84b2cBs1galJ5At0do1p0FvzIubEYP4R9p17X9wnT84yJqrcZ
+xsum790zQJ3mZ9d4uJksqhW6tVIMU6MP7GXzzrWRDmJ/ALCpA88skIZ4f16AgCs1b5hSAkzKLl1
odC3HgWxhi24O3bboWF0YPyhgHvgK1jUba8/suG3hyaBvh4LWlgQm8kzIMqapBaCZ8CtohRW8PVS
F6D/CEIOL/krB5Yer3ONcHAAoyHYTt5OjgYBLJONfKaLPXSgxttEmHk4v06ff4/JAB0PiLk3HDnT
CCFNKpwvwtGowKchMgZAOxAQkmJOCaRrQoIsS+7YlTrcM0l5hs39EDUABP6Pgz/3IdFGQkQqkY8K
es9rohlg9tLi8jIMxfd2BD8FHyXapY45XkTFX0IDXWsT7UxfVxjxlTnOLGD2FWC88VHFhuF/kPiq
wzkSbDNEPvQ9VzwFMDnRuCrqB5cIyab6ZbF14CHUk/8f1BDHR4xvajMnQuAZsaiNY3ylKCruwePX
bduganputVsDQ/puW3C5GB4M/Nxtkf8HIwxQIYX4JLMlnZpxIb4cc7hxSI4WEsvytgtLwRh6xbI0
T5ohCUvoiNQcW2JwkP0ZcarJsFcG1EjbJr1Gep4wlP97yPXvebVguW0TWyiW4X8Tb1uhF1z/7NU6
reN8QxOraieHkrM6sBZqGPLwcib9R9WgDWAcUgXmhfDjum7NOTya0gEKzmlIJk3C7ZhA3GmSgHE2
1Md+18/FXJGFutKUwhOsJyNpJ449ePvd2V1FuqPHT2/fmyabCJt83KvA22pVRWdYYXSgRj6wqOxh
gOZfeDoGvbe97iRMxXv7uhrAWk5zknIcOaAlZV38hmm8yDPj9HG4P9qjcol9nrcK3iClt56GUDs+
I2WRi8IA0mIKM3FLdVGleoju7dy1shMyVLKVsqmMEhW/r+FHlQizl3Dx+UeEC+uv76bWQSquU474
ZSD+XqyAyZWmlrEBIP1wPRn0U9wD9fmW7TStJ+m1bXBSsbou5Lx1/nif/aTRwYq8fTQBuqZgza6Z
+vEP+ipiT+j76e7z2SIAbIrT1bdfktIVLos5/n0w9tUfhTAnLunP25SB8OFovR+a/VZAa7Ppv9AK
5o8/b0UBDYaugCx+tYUWZKsFiG4EWedQ19DIdVOyfMy0ByeAshZeztcbz/yNX3HZD3BIEjAdSa/b
IxnnLzj02bbVVCo7Ws9vh0FlsaH+LjhBbhCFkLHMHNG++8bvjcXmHwwzGV6P2/FU4Wos+krSfZeC
p8qWsYnVTNaAEZ4YeAiekPjLlNVwi10Cp50L6Oaqx+hJJ7KmlGUXVEO44HB6VCnJ+YrrzxNN21b3
oERPfBEPuiWAbmLKD4uOF/o5KdHiI3ivmGwWRumSeOYLNM4d6p4dJSYgYezcBL1r3UfQws0VcpNu
7dXM5mzTzT/9qroLLRiF62lk4EWUudF/OOEO51cjZMHZ/EP/6Jf7qd/FqQ4iWWxWC88N2YUW21Ht
Cn7aiGvDdEYQge76Bah3Xy5yd2OI0/ukkZys2kUqLoUe24eGvHiLHrSvjfPIopomwrOlwH0i7ARR
pXedd6ZHXkogNnRwsr5xQnNO6sDa0X37TIDdlKdyy7MuTaBGkJGIB33wDoPMZtcfA+1oER5A78PS
VtvhsYYGSGYobBaXU3rDTERSCYcy2GraMYvAcvcX3gkefsOxO0cGyuaYoVVaIHGpM6+HlXIW08C6
hDRcC+sqHn7YcMwmtyDYmACql8CFXdnsQ39M9wPTbtbGNYgfRQSQQeR29GwNjZTiI0vps/oZNZpo
qIrpFfLzaZLZTkQPS2W+PKXbWzrQQ3YaQPhxbjzkOQrU/rSVhKRMaLc7ovBzD38ULdnDm/tkAJlN
vbbsxx65XQXAkPb9L7cp6dTXWmvE3ZVKceXIyxDwXK4zbADp/rAi86gGVQCTDmEKiHgJBpG3WL+9
FoRw0UVXw0VZ9XOEWJw9H9uNHL3p20YwxIVf+0V2qsh+aOqH0/wXNT3OrCZRDoUKBfxvn3OCM+aY
tfRpf12jsytnsVzW+dmAEMfGU0S4YsTJQkh6lisILBKXfzO+xf933x1MOv5foJYdDl+NfoqQGrtW
ama0QQbWg5NQYYixRLkyHC1ljLHoA46RAG+H1D1WNzGnWvsDsQeDyD+Kyd7Km6DVtFDpkK++mApN
Lohas0PpAleHN96lVemEjCDWWN8ml1eAy/PvutNrUU6nLQ4PYumk3r8E6/xqgOrIPWmriCB2/zWq
pOq2/pCXKmUqrd/TBNePRF/b7CrhUCcYeFkLT0Mm9uX0SydQYWpZzCwZwI3pJAkR1a52YbdHR2vd
pD6G3c1N1n8KNeBiq/ssU22p/gVTzQfoVyQHPyd84eMNwo8S/5JLLGxW37ldfW+Cx7RgSWiNhUAl
HomkmorU2CkDbbqs2Lf5iHnpLFV5pSQ4zDXn9HOqtGLB4av00qgRkt5cjWcamzDcuBW++APOll6/
kuscQ96ZGFgCdx0409/4t2pK59LMiLLDX6EJSHHkxGOHGxMB12acjdKFtaH4tBeBkCc0mCGOJs0X
E9ZFfpvvh9U7aFuSUmkM5B5FZBJy/XSrI4TMN6ZCzjjhL5igTEspjHkmfxnkjsJ3zyHV4oTsRYXj
PBlmskvqz6CWg25iCPKx8GDBb1wM2/0z8ecgA4WHn2xeLn3g9OkHvyc72FiKr08cAD+u6fJXzNX/
2575o+fnPMYCLzhxoWSbcx9YjFiwWEpmGN59AjOUA7nxSYDyNnmIZxYw/T/M/s8VdlE1R8WQe150
ypYsrjJ3hUHX9lAVbhdOvDO/y6QMl2bjRAuLicco8y9002eQumFEqeXUu3h2T0md/JcPN03doz2g
RG8wmMzUftz+1HiwpjTQ6D6hy78gsm72NQhUgbkYDMP9fcR7pAouq4lzCT0BFI/P1ZgFCaX1hCPI
Y58orQmUoZidsG/pYxjmY1PV3KJ2Im9a6zCqWWxWho5ZuUfYefEn8deEBa1MdRnHlA6wousrTdue
4tUU2bLkopqGPFU/tRaH55y0ttH5K5FIUE7PR/cxwzftqplCP7s1Lik2xfXcivrB84jlt7khPy/s
t+/h0+hAoWE2rzereWMCNpU43c/MdJO+9BMdECbI/zeIq/zKPUFAhTgA8hexBuxX95p8UP81YQ5r
+RGFKWa+Dew+jEQG6OSv8irluh6vI73M8muHUeIaJEV8b5Ft9N/Fj/Zf2zq7SOJOU9Mmy0OB0gW0
sOX254jGZRX92d8T+28cYovXKHqE19ueknFN9Pr3diocCS8vnbN1EuN3uyCA7NLQ1OtbaN0pdVFw
MPkWzbjZ7r611lYgQMNrnUWjukcN1LeVsu82UnG7AHotXZlvMRs1+G7DIew7D9BIa0C2RTnm5dtt
eeEaK8wMax5YpbDu44QrkwyKYITglGDATjA9wPMrd4897wbftoKY8wxKEMpP962NeRB2e/BjbvrI
8tzeqO06Zw71zp7Fkc9mWclMiYy2ShxQHKb177LZ3kk7utVT548llaSCmYUjrnZFz0QOhRhDeY8b
VKNUXY9M0PaQU/wYkQhb0LSAnehHrmRzcHUlRQy+WjMRiTBg8BUmNyFqreRwD8Pknbz3Ld86Nqoc
ZKGCWA86e7MDkJy52HhdgU9MQYuSHN4LD1M5k6f5DmkfpVZiIKOOjNVN+nlO0YRSNzVK9u6EjzqD
eSejORK5YaTNLyOxSUdiDLgWg9/A1/TorpGJFr5JmYyfgsqqXnfnzwKQeEkvu3RRPSsWS02wX7NR
viXmFL5ZqgeiMF00o181QWuxqkk9fRqY7gaCCk/5kyN+gEOUGy5s5B8eY/6jhm14CHoK2+lSgWb3
I18SronSZ7F2OHUZCcA0SuNHeT4TKvb+Wl1aUSP/UAMhCipn4VAJQ714kSP3iIGgOFkfIsH5B0Qg
yY+J5zCgRUgXbBxnacNQSRZnHbaVpbLtGCrbwZHyJLwHlqt3oQwnZ9t5SjHG4bjBFyY2fvor8gNw
SrbExUAMMmu5EhfXVOiICo/ck8S9Hp034sUApmev11rOqm3UAI7SP4d2B46aZOZdtPggoMLCyBNJ
f4oomGonIloGZVoKjDoB7PZK/2Nqg9nUqwnVxkj8n0ECsVC1VhseTQI0ZuhpwC4HLEXembsaGEE8
v/NgSMDAwhb26waQkAwgvolkfJZCPTFwF2exYHpZVKRfWwQ/KDii5OxSpr15CujTLp8AKqNwzszW
QarPmbn2lkcYB+dxxGLz2ECRnUIm8fI0H8gIKtUmiIdRSElmwjNch9bQQYPXbhJYFodaQxN2h2CG
CmxDr9NEzAvMO05yv6V5huRR0LWS3sL20Q96L5nYuxoWO2X/1jgxnbw/mS4XsAk602NyUSABnvZS
5f8erNa8t/sOlGveYAa+iPpSnfLjm6BGiIKA7cYz9GimxghNKPW4Gk0akcifjSJX7xUn02c5/Jtr
eY5PkE4UgY6P/tCgR/SrzCwtYwOdc8uqfADpj8mCaKCIc+BUFe1Ct4jGAprGNUfLYHNTkgNV6SGH
9uAR83TAn189+KG2LdqbAHi5Bel5iF+a9vSFbbIgrXJwnWjzwhkv2hwXmY6+hMxVaxOG59UJpLHl
8LhRZH5F43F+Ax28/f5dDwuWryn2xx4AXtbSADMZuAj6LWYe0eT0Hs+/OeU6O1xtC2x4gUbTvbCT
a9LFz1g3ZlePrldwXknhDAJmM04iIpPpwG1mCwzgbCDvJc/h34J0hXVGf0hBIbZN1ZPINHEiWGdG
q6wCqr4hgpW4JaK3uth9/jGMYSDIcsKN7J6bPI+8j1oYho2Bg6kkLBgD0NAwqfLQE5xjmt8UoQ6b
BQL9IHVWJXgBNSQQTKKOt4CaHlXQMTmu5NTEC2kDB8FBbbUTUJxLVO46vA8Cq06FerAf3k040sfc
IU04oPd368yndOLTAKcFs++PVBoCdmavcdb8CLsF42Vic/V5MbbRzSDcJ2/g3M9e10Hm1V4Up4UU
XabczDYVx/kUEWktVwt2RXCtK9PHhbrvmiEjfMrRi5Z/IjTdkuOG2cIF2X0tEUtSUSAZFmfJfc0y
yJ0THHBHW0WLzjSu7F+td/WE49GHwkUCZCO8nqQYOcynSWbwfjhB8dzfT0nXXJVdpI3FaP/5Eae2
5kOw9wKN/Vxwk1HFAQpIpj4u9k4qrkbpFOxnTwO0WUaSGPGuHFRzD09cORDyQ4DNmhYTihptL6eF
YxtYKCLKCEp2JUpTy9J3PSa+ftLuyLHNHgFoSiL204BrCGP/L8upy13AtW2lowYT0mJ7N9Z4gKp/
R2EIalWsh2tbHGGg3xaXrYrYxIvNacRfjN5xAVKQ5yyPlKFKyhxeb5LeaJC3C6hcnSaV+2qiZycj
gVoxMsGQR/nJVSLoliyq11KJuDuCG+wCVul7o/f5bVqouhebLCjqSnXLBuh3klObXU6BzeZ6h3Zp
Vro75vpDR9IUWdvE6do9csRKJUxyEoUW2QaOjfmfHPu5w9W2g3rzIKwWcaT80ayXC3pz55u4eQO0
80qZV6t5Bb/iVRH1fwjMQUKDwPx0WlCtNZgpBLsrdm4S+ojOMgkcvmPm9ZOJChwfUB6lBVzmJyuX
E7hzJ2PZtq4Xbwxy1vOgul339qIjd5sit/TcoMwTVfF0z0tj3A2v+CMNMuOtg5Scaui7/sGEYVYk
rh0jWkcl30eOen2yx+JQaL45P4edzvJS7f9IBlcuphy4QdAX18XANb+7eom0PWYODzbswxsbK7ue
XuKQuRUFn+CgCu7ht+sZLVqC1wQfgZrKoJdE8K9bfMDcixDvUFu9SGyvCjO8Gb1eiINYyP5zOVb8
jIIcKiVTfuK2IOwFmXyJVAY9iNU6nUGOmKec/v0KmZNZfw/R43IFmrWZC+3NH3Z2+izt8JY1vVZe
8TraSNCGs/JtQFqBBy8ipjcnR3T+oA1qrMA2w6z6nnPIUEr/Rr1GZm5uRsA595YE5zHBKLTbqgrK
6AWrwe/vz/2D9pY6f62vhjdCrOoWrCAz7YayS2ehC73vwrGzDIJISR7PDOD0pw0wMq9DsDsCUCsq
qDnMhKFo+tXL/w01rkqE4hqk9kfjp6v4LgJIg95eF5F0hxZIBt6bcknfmIWFex8WRpitMN3oIP0u
kwcuk1I9oMZCbCZ1ByywuoZpB1mxVe+TJk9TacSLT2Lq2K1zrYV5M8a90SnJs532xapAK06d8oSs
yOdQBXMPeA/Hy6wIbpayn+OFKBTGxZ9yk3ceqxLVsZMSCf4uUZLV29SbGjaRu0yIv7RwPZczDSL2
G45AxA/g1AZHG0kEWvZbK1olijrKIODeuAlrl1avGx2o+BTcfD2LuRrLfTGzTTctc8/L37QxV/G7
KH2Uh3uNa56U8dhRqz0tAlkXeGzMXlV5nVLYAqBcKNA37TzkffQ7m5g9LsZuiXYJ/wWlBS7IGPJN
CUdAD3vWJF1NT11QTDBbQnljZ+MIpE97Ig922u+9r6wQHR9k3Y453YJfE1j2NvA4YtLkdYF5l0dD
4XK46VnAVQE07wH/7kB8nSgoKCrhV2zCB/QLJPflztCUcdM4hxO/rL0da7kUN1w7DMH6r15DeoOo
i6hOme+8yt839h7wJM264YjIOnHaEBDcbEZ7IFnZUnwtoufZTcAGhhAFppnibOKAN188bvTaHH63
QJfiA6QDIaxw4FvTsQ4fRq44z2gPWL46lkzgFTlkW831lLT8jMH3BcAc9KtioS7D3EdfNM6sUzYV
c1baZB6ogK9eaVD7nHd2bUjDATbUEiF3gN2WESNswdiH8UuiNnVORvEbqK7Ja+pwYvLrv9fz6WuA
7yQWsRw2Dk3lyrTLTXcEr5S6gl/kSDZ3Ww2Ot9JMFelrZs5Ex95wYe2+MgvbnFygYW/oAfN5zloU
1Xllfgy6qGBJbeU7OIH3qpmAChofW5YveI5OjPbVE0O8boN3T3Dtj6DKFZGDnHm/G8+VIGqW6C3H
aa1j0/2cA/JxVB2FAhTkWeXtR5FB2I1AlcSzWd2EcZ//WvCfzQwkE7xctD3m48CF3ykbjuQhGQUi
PqoAqp948HLNfALNDmID3PdlyJsQVRYaJ1xtRKbTg8MtZAhEMt7SJfOvRVf5XWbt3bnvCz1u0/qb
mGCKONCxIfgTe4e5hbzoLjiAKr9Es7Ont8/ecIMA7+/LrTBxnoBocIhR7DtyYAE73VQE1FdxT/6M
2VN5EKhcE+JDsoKp/cPxPXw2nTuNy5sm/Xi9Vw55FCYwuhlVLM2BmPz36bO8hePZI6g1pVSL7taR
b7KJZvMhxfVS/mFtIc7fGWoCuPZS5nH9Af2mc9oeKmyntaBVybHEQe52OS6YO8qevONAQ2YivqMM
qupQ0AJ7n8XaIovnWrq70AOdDzRChAM9fN1b8Gbk4io+MGVury2udsAFNvzVnvJut89/BZ589Vb8
si9zxt27jCFgaP8Zx+lMf3eGhPNPD3FRv54YIvJls25nY48MZ+FHgk7HKSQozM5Qq6i2wg/vb9QR
KznTr5ErHve5c2KTdxtZLLit3+G9W/UcD3zgeChbJDPaW2AXAT6RSAMcHxsXmR4FTKukk4WEKLH5
rtdasrImDmXyJzs8ibI5eODKpkONqvWL6B0yZ4PRytRXSynka1gqL2eJwLfvDwHpb16l0dsVGV7V
1SDSt/zrfy6UT6jJTfDFMpXhAE40l32p4wtkut9xI+2TCHODyBaZkf6Q8zzIl5dBp/PB3rDfJGoM
UzEJ7HuPU6FENoXPXWwcZDXDT9jIfyszGIdc5AKUQnWW3MuJYGKvUkKcAnfNDAU3pqQ632o/kxqa
a9kDTlfOkZDMhv/Nw+h5eobwnRm05DW+MtkUw2KN2xi9adj7txB/yklxzTNrvimfNlJOPp5UgVfq
rNOd/CjF/4Br9s6HD+YAbm3q3clhC/ZC3Q15+Nxl/FTdEXtwspzh+1uH8Q1bZPhrp0tZYR9vuFSq
5pTYL0aMm41xOAMzJLU0ppVbcj4Vk6vNsijP6iWgPBEuGTxoe3zuOSSdpHE92FNo8ABwqnSIifQR
wC+ALolo7MThNnnfRncNradijs7Jd1qAW40VY24sYA3GpvMaKslVMV92M3+HpxXMSK3lvEfDm56E
DjQJCtlz6M+U4fjyWqWIUk0O3IHXYYe5jTgu0pcolFqON+xp3JH52s/RrqF82l73ruI8+Zn/8Bm2
8ZDENCudopVcO+uANaXn2MAsK8sD4tSgiQdNP7UT6FI4JqzUAGstexfwqhNhAVemjkmLKWPlhIoQ
lHdcHANGUWA5P6kP8mFj12LVeOFvtR27Um2lxyfaY9YR+tcgPZxiCXGdgZa4xJ9NwyoUoQ7rtJAo
3ILNRkZcP1Y9EpKDo8NP25QM4ZNYJxFE6jWxxxsNZkPe97wbQdVM4hrFiHweg/xxsdqLCK8pMaBC
DLVoriFCosDPIfeP/+qmVRiCCJUEbSLkS0CGU1qlCf+IGuBd580fYatzjJS9CWsNKavjpRHI0g2u
h+XVEM+Pu1oPLCiJSKU2bR0rrhLgwPvmBoOMbGHGYkoyJS11hRM/dY1dOgYpUcHsfCcPmlJ4Zk0E
issvPN4zfnZNW4Gs45ZeqUBHHk0FF2wB7ITSCfiOjmNIKzfYoMT16aGPZjoY+3/3AHgxIer1x5Dc
gE8uvN5hV4D8rpTYQIZlHBTqwrLWI9zBLR1si2EbliwDMPx2sYbPHexnaRFniYg1j9kf9TL3gkPg
+PQJnUBQMOWS3joh+xZ4xf6ws7jj60RMl2PW7v5Xts3xSMVXt1p2gArVXTGlJN3f9fIInRtXq++5
qEA2H2ikfeXkQ1+7lKedAdVjsXUV6or+0OirkcingE2WvYucg8uzx6j4VlR2LJ2w5nHCazyXh2RJ
vI792AaNieGO5aLHNCDvPO8vxcAZuEO9y+Mbco+ov/lokfnypzjL4v5Gu8GZqdy9youe5VjjLYz+
BeRO3yVDj+3qpmkmJQMqeKfh0C+cB7Jw3UJT8pvlUVtJKoQYD8hKZCmi4NVH/37sTM1JKZCqcO4Y
mdZL9n/cYUnNliElvikeVycBkwGiZwNDTu8Gc75kUzs8QEQ6PqoB2dfDjkty7PBXqObvqRm9nGSZ
T6zISTk2lEqt8eporJgXQ3VYi0UzWri7B6HcMiTaHKHud07ec0ucyPg0xyqm9CjrV35SxiQhuEpF
gRwcKWIDida+MBAezlsHqqehUydpb1rftDI73+loW677vZxQ2kl4bJeiLwnhLHGvQ01Qlzv9XwmB
YkjuqJIKxR4J+r8JmoZtqXulnA45qTTH8qcTKOaF6zIANyz+XJttYz+IrY3Sn2cmHC49OIp2nzXP
ueGGBhRJzNB+3UYs8i+fXbmrFpvoBvzq6xkudAj8LnhHHdpf9/LGbncL71GIqwF6JUShHbHxHf4m
H6WMUCYx/fwCD6mHMKGX3E6+f5o5q6CeilcA9SbQnI8kbbTItz6zAVyIdDMJqzL/NVIIIzyhNigK
jYoclkrNPag4Ae8E4ZOyE5+LbuZdWPL2LV2Vtq/IxA6U2Co3xZndQfM42AaAbHyHpVAdjrdo3PK1
K55olD81qO0I/k2S3Bh6zEUwpGuqwO9/Z8jnyyMkEV8x4VOOFZSdCHb2no3I0biZx0S5ayF8lKvV
V8SORPBdOPQnkmxqmMwFwyJVx0dmSjq8oTYN76rFEo4c5rtxjm/dIJUgHD2zxYXUPxNLgDOKXQv0
nXDQAPjZ0S303/MYKMw3mxupXZvfmLXeSLZcgbZuMlH9SglNaXBm/9z9NS6o588BTTWd4WfmdS6K
vn5mhjZbRvhedxJxeoQsXbelMPJq5CP77TdXsQb4NnoSAEdXbSlAdxOgK8NSd9JQpvolG1bNk+9c
JL71LldEgRB/AHO0TKWqQKPCXh8UmS82UFlDqKb/NcDkIzZHyL1+ht61DG9OrP9NPG7JGLCgYQqp
DT/274o8tnltJDeVrIMbOJ9lLWZz1A+F01cW9Wyu/R4lyEOEzzDCwHUekE8hI9ipkelRGHGzAjIi
gZX+FQPaPlsT76zwV/tAkWCTFJLLO19QpjVBwH6Vu7xEFqdSo2zCMtjj/h4/af++ULOTb+u/XZf7
dtUi+WjusUwbu3NwClhziKBFUmqYhif3/pha7kub8Yyfzonraez4XElPRChKha7Z2yDgEgNogbXw
v39WwkRcYzAtyobAEWnW7d0KzljKQn3hcDp6dNVXJmxKSlN4sdCLO7KO2vPbzVxEQ2ImZWEZwGgO
6iKWl59d/7C3Eqbmh8e3IxA8oC1PO0pmpUOv2VS8ZUNvvR2UFva16aM4Ju4wyVAP5utB3qFvpZCZ
NjmMZlXy5XoTmOgCjw9flJsWGIzZ0ZmuGLzGvpy1ix9SRyQ8dN5Chv/0xCM8jF1tLY5KevIxTHDR
6ztHuP2T+CcSJlgk2MOhsVp4rtvtc50kf83DMCV6dsczvnt+LxxZ88gzbHfkm5BEMgrE4tR0HOwn
9RDyw/UcGfoOar7OzfYTz/8Jyw1i6VmqACcKUrJzlgP9Qaz7f/5Te5enqZ08UGUEiX0YImkIMACN
3na9UxIttGTrD92StQTUL3pOvd7zOQJs3yA3jYw+zmGFV27nWURr9npyGLbRFV0mUL5OnPzX0Wzu
VOgAvppUaaMtdb3bKWZ3sjmIC7eDUgfbIBf9T+Czfbokchh0JASrGSQWRJtcoBe19RvNGXUQCYZv
gdKpYiu8iN2TDgU4TD3NwQzvRLNZgr7oNf+rSJHJSNwOqSUXCgGEqhYjxYRd48TEjbDenrpGEGmK
yCuixwWKYhU3wytaIy7l3R/maGpdmUDo31r0t9wf6xvuea49eIgdV5nbnlz/SPOMPSxYDcos43MM
DXsixhZuEDFtRlmI9zuqzlOy02EkhtY4Y9uEZGaoTt77Ch2TI2piH0+X9SYk2slSbEuSImiBU5H+
eEgTQfpqFQ6NsdHsLL5k1xp09gv189kNgQe+CjgmZyadYlKaDUfRpLjY64abUVo+4EthMsIhBU/e
mEbeFwWjhPBe2+UqmjkIeNqviSqefxH07vmGwF3Z07+KtMJUXVbqVXVw7VwNGV2waXCHIBSbgE+v
/A00+7Ze+VIOQw0TkohkHI49XRpNV53n4XeKYUIB52LRVwOQIa7g+p4GSFc4QvODCABukVt0AKkE
aPsKP79MMPjvJJTCrxD+K3k1Q9mpaclyfzYGw0sEXjUnI0PNfkHjBFiRCHQ/NWQI7hrPSDTFZvpN
E2RkUadsjx2lERfGX02kbproVZp05s2hUWng18USY0hZVxPzPEIj9yXFR3WfCaKA/TLBRclAhWS9
fXZulFqyFkNAJnkvQSLr90lpYVzd7FHW/8DuBrJ/i24ZcjEnomNQbKgVOdiImL37oE78Cy+kR3Zi
LgNjMe/y/vQmsZFQgRiusFAQRaIJTpVg8ZR1pbVRPpmu/naORng/4b5m/H5O1fH/6Le8EJXrX3MH
AQBmLGNp6jKCdFrPechOlfuvKxLKhwvzeeYImXoEq2gdVkir+gyNL3W+XieJmClRcAmf6mpYZWrr
UeO0Gj5f8M4lWkoAws36PuswB8OtLIg6PAGgcuW4W6u3s/BNhCaNOT3zpMIZjooR7M+mdk7NAkMr
lDmcx3keClb+uC5Eg5Sr8uGBY+v8DVdP31Dpzf2bnbiZ55ePeh2g0ZqQ07cNju0ZyV/YDhBzeDQP
EjiriKdXT7JHR8Nm4A5SQi4aZBDj4kCmFnND8qB619SPOl/kBf/AGFElLXGOba7q0JGPilRmecML
aJoCwwWrdE/P9fohPE3CjNs9YOI2tDbfp6+Ft2UqSvnJ7rALkLsJ7i2+FpbRdGcWDjxL8ktUUCxV
a/1D8KNY0w/QDC8/4UEXEf0hk5PZVKoe8hpmtog08yIEWSixX/BSqqgpiq/BVphhXxMTvjDtxP6J
Nd7HfNMhGkgFghh5HYo98mJiqrMcmYs+oF+XgBvFUQZcXNxFmBRnoSlYzSpy3xTXvOeJ0irM25zv
mrE1HesYNDOgMU2C7oWL79lqtrpEll91uX5BlqFlDWYYEfYvyUKA6byRIDMZHiQZEfPy3o/5/DFF
XY1xU94lxHBUTt5MsiBW7JyoNDwhu/sPdL4ZpSTwS1DIjKrXRgQpEH/Jrlr2bEALSLzRAY494BsS
OJ+VESyt+oJq8OJ8rZAPRju+hNmrZUE4UGYrzGTDXY0eY469TZENlwETUyo5bTtF5OjGkASW2AGw
Rv6XNQqYGGqvIHry1K0C2CM0TiTFabEBXT4ftFr2pSnk6HBjtajZh24xIBZ/fkW/5cAeV2qkqlAg
6oU29zNV1h9ue9+PDyCg3nmUIYLiByHwRlz+6IKms3E9z+sSTR+0caVJ3hune+LMVr4avsdxBVUl
olayqW655NuyvtDLzkeHnoWPFGdx4A2ZuWy35dL/yjkuALNrbc4Rbnu7aGpGg7UhmOj4ZdPn5Doi
skzWmWSgx12i6x75vnx/OrXYKrZfzP01qJSwMx8nn4SNBQTpSyC3NnuXceYuj4S0gnezfaq0Inph
n6pkIxAASRR/huRgoPaOJQE6d4l0Iwgw9fzwXRlqfCIJZ3CENy264Bak+zm6a68jwGwYUi7FSffT
5dzYnb0ynXqgMB1QYtz1db5hpo/4pL7rmQ+/AnaQaAXGSHm+5If4XXHLWfhOvz/HFOSOoz0YA0Zx
Dg2Ls9xOGotbZITItBTU+9MMAftvcldIRz4HjH0aE7bQQWJMeBNLVr+3NzO4bjBS4UVzJ/9FD8+Q
XdH62iuzdywQ34f+ydp6KeEen0kW+39C78GdXrwbn2FbAaymxt+QkH7diSccvQ7YfSSn6GbmSCoY
uyWoFskXVOxjzHjpG7YCSvADCX4+xKa9rstAZq78F8HUlhEeLaFwD7t8S3+kGjB+QRR3hs5adDV7
XjBDJtdc3VAWyAYsLV934eTOGWvVO6e1QO/WKZibP+qNp+7MdlJjI0L+dKWIY9GHmP0E2zIVNQM4
q5nH5L7iw7k5RiAgic/q2mAe5iOek3oqP08poLqsR0KyvB43bk14n7LpDweXOtqOYYFI/yZ3liuN
po7au6GHDOXCnUnPIE+NAVLdQJbvk31wZrbcBniCKo/w7bCQduuWD6en9oJVfh/K7OF4HrtxYK5p
JBziXFtOsaKysi3n71kpPoGtx9Er76FE5PFDHAPYrXOx3nMimZ89iA2Hw2MAC7wyNLVTWNYYfdV7
GoV4yIQXzzY8STXDXgOy5Bt+F2g7xV+/XZGzNtYKjskVHt9QYg9zQmEyCJ+d0MMg/2sn8ZMIvsnG
jfBjjPGmgcAIlADNFF9iyDRtWpYyaCSbWtFXTqGQjBDAa+vtRuc2YWwyeZ40c91GDoz/XoO1QMqo
+dVQwdBVx18XVC1pOEVnXewHfPfllKXAanxycsI56/GSEbAdzx7oz05on5tcikvYFY+AqpCPXIRl
64PJqJO1AND90qR/ASi58ZpB+BRImQHJoFalzUN4WfXvEjAzLDLp0YQU1MwnY6DIyi5vb9adxS2Y
k54J3+THWz/02GvoxRvgIElIbuqjUmNjC2SoCu+cZNoaF3mo2Nl1Jef0WH/lSqwhtpf4JBVrQ/rf
VmO+/AWosmNNknNZHvMFld6QYa5e08CJDNWyKAF2tONd1/ZsCLgxnetqcgZlpCxuMNH1DbjlNIag
dBg5i7ZQkPtV1cSEfIb8xQlN0UIH5jlNMSH5Mi0IDCpNGtuHzli/zLBQQ972KB10bn0ujHMuT7na
5kNZ4n0DPrjPVvQmW4s3zEHD6PkCoDpemElQX3EmfTTJO++vxS1S9/QaKYEzT+uCbP0Yr2fe3StO
e4XNagIPnuz7NdrpwwziC0y4c2jt1wKDK9kOhKih8mZMNEBmn1i030eWoBPLwXWs7Ws8p5w+0p+/
L3cwXjPjnzISiBsv5gId7lwGyC5S7jXaMpNFMfLcGo6RjXEfKLMBHS+oOuwk9cue7230S7FPSkRV
0DdzYyWIZyffiwnV+Ey56zyFoJbOqkZKlsC5i5l8uiermToOKEBjNbOZrFTUKtiqTv6nNjlqxDrd
qiF7FAzcl1W0hCrLnzFnJpfmDxpWd8J0Wen3owu8gVAa4sc9dNoOEe+IRUDRGOoLPXI5RcApKl6e
X4//LO+EZK3a9+Iz0souh0jdCbew7HMewbT0bns4XaRXUZe0BeQLQCWBzZy5vBsvWEDe7LOL2Bf6
jbxnsat6j8NfOxw4EfOESR17f2kZ9EB7wjfCivjv+joro5mA2Ea+w7TJ88I009LD5OxBwbvrGeFC
f5yRW4kiugqv2qoVB9K5xDfN5L4aKpAYvzd5LL4GMrLD/W5tjFC/Kulcj2O7Ds4Fjj+9KPK/Kbp9
ldP4cNDMY8l9VaaRKc0WEOGK6ktHK5rWrrEtG/ITLQV/nXmNGAfdYTJnVY0lJxbi30RxwgOumheZ
YX88c0eiZpcw9F712rFjwnC4pd7rzZnp+ugzp6SoArVx7arJJ5ukKwmNopQTyMlI7n6zLLl0iID3
aqDtNAcB3axYjUYL8PLWgANN8Q7ua1r08MOukfuUb5KXpCyMwYP/bXCEesGH7qjXpXk18fBxnlm9
sfQUTeLZ3G3MmsH7sNaxQbTa+3Y7IiSlTPMksx4bh+GkKAYvrHjEnijxs5vl28jP3fnVDMEpaEIj
qdI04aRl05y5wow25L8arBmws8W0UxsSqIyEy34kAib3lgX7j1tj4GTRTjVBydeVD89CVwwVsaT6
yVnMEuw8C+dlhvIS2PRC7CHnUWpPP0Yu+bhxbEHjfUiMx5OUYOGblVnzJ2FerdeGioMqaSW72pyb
OG0nFxzF8+XivftpT2+hkSoUjpbuH9kNfPe931cRZ1k+qleXxiIgxjU66WV5w4rUw7TV4feRsE9Y
2+nUX8mKUJCJ8bmNwweA05uzvJUCXrMMTegi9Ls/7x39CIk4Mn/G/tA+m08+wlyPZPolLUTS4GFL
ekLjvwrjNTuxQgtLGJRBc0fWw4+uxtzl2qPVuoV3CN4/3h0wymKPzKy8ztCSPz6rQcsT/uRuxvNi
B11sEqgEOE4U0BtaOs7kdLA7IwPHq/TVDjPrNuSE/5inwkX61SbdGJJjN/ysVUHtmcs1DXnFwb1T
l2zbaA1eolt9hJIrcEJCUMHwqY+PX4kq28yNru2TB/KjiaOvuWrO3YlBG0wspXHvCkstS67GROfz
V7Y/huu19AoJ3tQkWrZKyHaIyQ0oZyK7ZWxNP9sXi0ADLAG4KTauLtv5xJhe86yuJIlZjXxvX2my
LY/uauK6fOgCOgbwLb6Noe5RtQMVDvGoAPnp5ugdGXnfsODSntXq4FIqckHETaNQe/H3CLCYSHly
57UlkHlWB8/Ubng+AQ+ICtSpnycTO5RJ/9LUOAD+AR7XfvpjvDvV625Qvqci3H0WfxGZTcpD6Du0
R632ruILt9k5b+Q3HfiYdsycHFVvyKGs5NFkGgGuc+TTsK7JgAa+AEXXi8Uk/v6t11uv9u9mnV+o
b6R0yGRcwNX+tu+8KSSg9QZGhmRFk2lXRflPEW4N/+1sBo9mSF66oV1qOvUiopSuq3lHIWAZgqPH
Hd95ZS3C+0nZmfOvOD7HeeXRU5PqSHA1m8AWHCda+s0aJQwix33Ds5/W00g0Ibm2e0ZzbgSnMe46
P/Fa45Tr2acOHFC5e8BJ5S4Sd+IIKXG3HnK9z68hYSJAuFyk5GCBI4lAZSUNboASzutgPikgS8l+
AUoVDVWUfOAyK138bSSGnz9nS1jXwvR3YQrn99fmUa/we8YjKTN021xez5Qq1iw3d00FnWm6gCFZ
15xqYztzpfss809AAJJVfqkKal6EGxWxax1TlZbhxYQZAUlH/qajn2xWNT7rBtQ7EKdWPuv7/I07
mkVPSqWkOo02anTJp+XfnVKA00h5SRMMQxnTfeqBBA9BjFp4TLgAlIL24K8/MPD+gVftRnrV1VG+
fmMm1gVLzgiGowDRAuygNGWL2K//Z4u9HRfGvyq48hqRMXe3+viG9DMknZcgpJzoX8oCM0TzX0hM
p3NHRi3jbZChk7FMH/wwLOIzAHYtvTRXM0yUIgHfRUu/6G9dg6XOtywjAZEijqj6b+DGOTXKTGMf
h6if/YS8UvvCWWaDoQmtZsROSh1HMizNp2TUuDR7H92fM3KSIymu8S97LMLHNd6D3c2Jr6JItt2d
LuYzaB8HfpYTSG+sOm7l+9lYP35/ba2rQyoWQYL7y617kEV+1Ij9eGxn8WhS2tu9L8zKKaeuLYQz
DooPY/HQKiKQxE/qFu06KC66R5Z/UjOW2TIWnicL0XsTqXyD+c+Pa9NQ0aexP9uRldLft32Q88m/
94Ugx7MMRpV6LKqQ5P+nfZDJe5DEK9FY0ZxUz+X0s892ZTrXB5sdu96uZrVCbYuympurWIikcWxd
LxfM2o667YC/EyjcGjjSx5ULs/o9cRk9fRMSPPHcjv/q/ssjFUJu3vZfRUfzJX8X5dRQS27Jsf58
EUKVjM6Ytbj8iDGccyBSD4kQsVc74ZxTgJpMeBtwcHQwcjouI129YlYjSLy1SktKs032sCx9Taek
vte/+mGDkfzAsr1TUK/rgtrUaJGK38jk/tPVbNW/RiYFSV5+8Ysl5CRSlXqHMjBHYJATEnfX+lSE
1drIOiFr1UoV7mH2US1TfVbmKnOfb8mueMcmlJTsNEnmWSTwbtEHeKsE6Qh8v62KRg9tjYvxN6PX
N5jkfuTJ1Ifv6mEoIKpnVRjEUckSKBTQhuH4+zLG0NG8dq+9qUQ8PnOep/jogWa+b2lMLC0312vp
6lO8jZUFWSvwY2PPAPrLuk/4XO2f4tOV81PCB84WUkrI/MAQhCICn16UOJp4/FcidzAyH33uQv+E
U3IGSpfWqQn6NE36ub0cfrBy0MBBA7Gn6ADzRl6dFFpCkUOL2VkAN0eWadjGKEv42L6LJlszdBPC
LfRr4rDK0UX1IQNEDyV8OGVqqc7mmVKTO3I+aBqfxQ1kZDdD4g744B8ETUYr29fT7Mtvuc5j6mrm
LfL8Es+HKiTa/mV+as3yw67pFqKk24T/BPhVAQlkg5dWTKYcUBZ2UyBYTa/Wlcc54TwU3/tAVhCZ
E/UtfIVTWq6t/yjkCVxi60vHL741rVwIL/E0+fZO+RabsakuGa/AEaNoTztPBeTIJYt8whrn15mU
h6306kmfNxlv0ZxWrobYAJ+dBB4OqO3qMWq4eH4IUF16OkVJP/AO36ubgIj8kyuSn0Wpguz5qc14
KxWFpcQOEqTE96QVkiBQMBiVFmCoRnmFxQ5PuKxNVIGoB0AyxWOEvK0JRqq30Tk8/q19gWX0anBq
hYLQnW6w5XMU0dY4QIs1YyApKBPAsDQsF5GQYR99V0I6YOA+Xlp6DiZKr/aIe6c2n8R4+GT6moTc
luAR0zaq3Xoh5+cYjQjcA0Th+Id7RbZKTSEp+1UXEGKB3zhhkfJ4DQ3t/39n5Qp3CoGVbq5dFNDo
eOYkpxsPuHRMWuTpw7TtN30hnEVHLDlXRnmWlxz0aO23YOECYZRbYRJ8mq5TMCYzhMn1XmruFQtA
2u9NFrUOVsJPHw40iv5KNLJ6K9920fETEc6c0bh7dZU46FncC7T6pj6f+eaSOD2DZOPXtOtnRzKO
ZKgeeAslXdrYgNvzqARwFS2DhSWN+vcjku+Fc/7AfGHqwBPZ+dXUnXStmrVyX3gWDoi96ZDzzcSL
aLeKhBOcipiGL9PZOX0FhUeTHXSDWZSooNMeWbH9Z2DVNbb4at32UOif8ze7l9eQub7nIyIEPkpf
wG3pPZoxvap4qE+VPnMu9rAhZEwClBMjK17SBX+5Z2geNgZnMMd0LFw4BAgbz09j3QV5CfgfVdRa
9+0C/Jav+z+5yZRtCbbsmSvjJuSfzZOyWlx0Vy8mczIi1b+n5w3MZxJCRQpuKT2oYM1NnjaheyuP
S39h326p1lJqQSgOlxskz0fgDHQGvacsh8pZzXJ0JwU8zU82ydxXVIgxrew+DaQk7PxKMhbk56ni
EaU3qF+s/J+ds3cC2jMxz38KPLwDynRGQssCb/R0vc5Bm/TzjTbeDl5TussqlEZiE7xlecAP2t13
qmqh/gMde9VtqUsP18gRRzqHzTNhRrrggKuDl8LycyqisY/mjyG+SMYrJQAKdxJGLUNE9oNn5P0K
pAs2c+tAqSItFDirYbig92P2+A0mAfp1Vnaezwwg/gWEj5xr3zb/kuPPYBEUE5KfIRRiEQd2pobS
LNs9Y+Ez/j8lEzGi1oZJJgIIIPPZHe/cXANfBnmJR0wzohu8Z3/N1NqcrFvQWv+u34ep/6p06d+f
hQlhlE3bCXZe4ajBlaisMs1dcmq+c2zEHxoBH7KgnI19c5ObL1W8K70ectWLV2wgUaaoFBNaBSOc
no0/GWRbBfgU2hb0TWWkDPCU2cP1AU3eS1lWlvKx3SJMzf0igw/0pts0njiYCq88ABVIXY8ymv5U
L1cghbJUvjeaDvmZ44a4zZyNMtfmjbETpEBg71riKlhZKUmEnp9zjkweOU8KpNahHRYS8FVOJue8
9enXTAOA1rFJ1OP1urIkPQzULhF0auCSpYtgTblaRwThfIkI4Ebqt9yobaXH+K4KjW5ir1VhLf15
UHeF7yTKy3PcrHBBnhItMUoFSG/W0VV3dBvoMIYNiAOEJERfkXt5+t5gTreq8c3S4Q+fns6wm1+w
EBfqtq0w0mLsDkQc/93PVNmWKUePGOp6dFHtnxb8RigfGK6muPrINXG3uL02f/Y0H3LpQm6Huxl0
UCvBo+kUyZ6UeaDM47XpXift5mB6U7yEWpKxAChi+0ZTbB62S3KA9GRRuNxBe2HCmVQOtystD3Tl
2u0+cBWnDR+45kg5PHhcdV+ITcxWNazAp8Rv/+YuLv2cAJA3gdPGrBSeoj7ojKibeKg42eQs9qXc
mxi9H+cbSdKe4VRWx04yLJKvAFD00T5gSySeRsrpiZcZPieYP5nXX6cuFGcInRhbS5iw/nZedriR
NWlWeWF6zRp8f821dLeF0u13UrgKQwD+sWzdQZOEUC9aUtfwcwTaJzhQVMptE+Emn5Iv9EOsS52T
M4zaQdvdL+GiyYPzrjzd98STNY2VMgaDyp31qqtdzUmNbH0AYG52BjTuqDnXlz2L05ALxF7schQ6
MFRlCGlSL806exvX8ZiDQUrVV47Bg0ltHifYUxP6o5pl3pHLBOwLdP4fCO/uCeNxV4hThrzJCi9b
D1ZwMtBFRq4ivBtyjNHiYFd5QJX/hpVS2QdOv8lCVm7nLSiAVMWmATfhgUS8VvHx3gs/J7zfHuvO
wb4CpEFG/gaHKoHEnZA9yH1nEaGzARqW2HyaphTnpiR2LTDTOc/tbM9NlxXjAaR4Gdnw0q29g9f0
RJ0j8Dzpa6gcY8V/5p7kgXxvNO8KUcaZejoChaoq3qPNCZNFwGfA6EfRftYbcxFqSdJYt/+vEFga
6OzfyXVtRhRX+kv4WZndm4BjuRoSCGkOuTQZu6LNyud1V5IwBnrLsLbkBllW+aY70Jgck5Y/P405
5nI0Bgfg88uOx+b2sxewgATcPK9M0zo4v9VJ6d716biRQxV5aQEBFJXEzZ/zXNuOcPX4swxxSW9n
pKFnDt/rWLt914h2cGTKY1mThGSQHUG2OUScTgawFjTlTPQIuL0jjs1aFIpmblG2PCMIZRD9Rp82
mG2WHKchnW2ElUHdybr0vpiEIxt4jafMkbsJ6RBu5XCZvowJb1eWoymCqcdriHtHnm8LGYXIXTih
67r6lrXTOCFW6JCiFHGfxtJjwIgnTGhdCD/KIAHyO/Lb6v5Z6VjHRRWOYlmsnJ/QlkMjN6AD/EkK
7ehWEEH1VPRE2Hdw6yV/OvdvYoBHnUnFXUL1u5iYJR/sUOSQBtg+hygJMF8rYu7mCPBdQRDog1lS
3111voj0Kj3HhQIV+BRCpXfm9WtEa+JdeeELPPX9WmBMN5WqAQFy8nBEym5JyVpO0DDSTxdY/HFC
c1BIWmymfsmt2sXQBcSv9FlfwhEI1Fdsmxp6rjYcBhB41fSdt50/Af1yFTfsEf4BFbJz/3u6I21w
pPnFWKtJ1cBXOxcNqCu7//KV3zRhILDhuQ5VE6s8po0fnnvtP1v4Rv3jBQOwMI0js/xfknbBMEJR
wnK+KFIbAh+h+wp8pHIRuP7eGBOclDHWMaAoHhKAifhzWNGpA9vsx5CB0iB35xA2SDGQ9EBStOdm
YokIPExFDG67kUxVc6j1Z49GiYmYKL0Q/OfPrphkPYUZU6q0htiokSFqnLykEmRBhkYhUgRakWuS
U3jQKCiPIMKxqclqXrhu6liXXGCc02KgKt0p+/HEO2IWNU3m0ynftGkkCpnapLO0gG4ZwG1zp0PJ
6Ir8dnNpMUPVfNSfgg5804k3Xk/mL9F5v4HELAx+nOTWgBa3shB9ApysCYOClEucg8kK6dmFtLYR
Mf9K83XJvEyQ/G4IwRYFBq+R0Ddas5v2hE7tuDz7okKpQnslvYmbIxEBgPuRR3aPn3qGw2GreWPR
qRIaCs+8koqcAZuQtLqDeL+wbCf13KlpeI/d2DE+faZIUupzBaluxZNSCycShfKWCEiMziBzbVQw
mMogmaDhaFn6gkebIEX4BJc1aB3ezcyiY3h/sJsEHxzTqFbrJMrGjCqmgMjZQThQ54GUI/h35Fzr
xlssznc+ghOfnJeJQB4LqwYEHH+tQI/rYFeVAC/RojdZAb08KMqeDsrfroMaK4WWUH6vWCvVFUKE
3WU4nvTDtH5RthqxeL9Nm2KCcvgHXkJRvcwZ0mAgm4jvqCW1x1Pu6hQ46ZDqkICOYibx2PqL+CHl
Gj6lO4ew+HJFPOpg243imngMTr50uwz/lRzOwOnfPR1wD8+Q//YB371HmFHghIQm0mRlAAk28WJi
6XOa8XUYesVqoGCxJr/wSPGwYi1NcuYXcLuGfFD3vI8QDoNqUZ+/IDVCRPte2D1x6Xhc9vjj0ngL
y7ptd4IxzQImV2E+UcEnytSNNy8unJJxFj81RPvNtC322rBJbfq3S+YLX0mZZD0bysoyOsAv6wV3
Ooi8CZMGYir118ctujXQHNBNm4HYSgyr8OaBRvYwQB19f5eV+QA+WUNQ7psQe8qqVwk+OkdNRA65
WPBTIgBJhxA/fZsucK6CpU0aLPy4uQ5wWwJyfrVlGxAiMR/XwDtuvYPbbdV27p4OXipCB0rTnnQw
nd7q+SThLZvwZfbQe2SBa61kpbUBrR7PgZ6Vh0sTOl4qLHKxoaPM89gisJxhlErz8ajdictALC6H
2KYIO4qYwVL+Hboe/SG4Ol49irJXOjpnNwbGN4SxnXuiitAUmXmmh6h72sJv1KqWg7aXtGkHB6ht
Cxnawuct9MowXLlIyz0/RvfOKu+8Vwyxr2b/Dj3vTJTXlQhQpc8YalMiGoUEs0ulHaanlm4tzW44
JhW00ppKjp+N9+SeNd2MXEdNIuQTNqefaGf2ezEL+lOKfTEs6tpzEn94wWI8rRFiDG6LZU0sahys
5GmlYAi2DxKH3gk76ig6lSizXIc8NuINnUkLFaPUZqJfetvSlBJa1WugS09XJdkKoYlYpKNtW8xt
mDKwmd8A+c3FgJGaxr9hmno+eKDUxq5V9jygnLdYw2ijNe63Uf184fpnGg0dcJ1SUCZvwxZEmdjk
xL16aRqhP0ZcjnjFC4yR/RNGzPOr5NRIvWJFL6F06CAL39qcltDZ2r5nS+K/zXFGjC+HyxK9sq+C
LkMH5T0aEpDHS30WyCIBA2orHTNEFb+hsfDvE/78YxEWjMfs4+0JsOq1wB0cXEPTfSt7SRM1vWdY
oSpropBfjq2DBOd7AmwyzPlF+x+aWqZtxZgN73lEsf1FSSdDYO2Fq4kn54EQ33k6/nxTG1xIlKHP
m6JddBTYCqLmJTIpNkEjD46nXoEyzrjPOk81/7zeRcD6GhEVv9mxRO3hJLoK3RgyqggJQ8ngqCrA
2+wz5kw2EpF2GlKcPvHv/Up7uL0ruFNkeDVc82sS+q2MKHs05YZ2BBe9aW7hcrfRAkJwKJgXCeFt
Q8gzme5Kc2PNxCFF17GnH4Xa2terGzhUCl3V1fxeLDuWGKfA62Nkaavp+MSaiFJG1FZF4hWzAVAp
yZkc3c1dWDKkHc9YbXoOM3agoEeNZw+vJkcvAtAeRiFKMJ6cUEbbFfOQM/GS9yy7uKg3Sbh36jtX
DoqSyRPxP2M3gZlRCtLcuW5kRLCYDKkKZLFk1EichCWiR9+/ObchM/XvKZkkxLDZbeZW06sCkfrl
c1VIzNi4vhws3jh37Kai7m360rTHe8H0CCCigEmBDqadpc+HOwbhD1TXrFJCcBiokYc4emrcBkUz
y8Ae0HTDR5KlZh02tHL70gy+JFF64OWoCgY7lXAeFvl0E0LNKS/mpiJ6qIQ2AzrzXonAmh4UPjnS
kE7fsBtVqhRCWeDAdESVsJkECJQTjqWAELvtedc0d4PBLbxRFkLhEQpPpcU6nzx5Dt7OZDB4bYlP
gMEhY71BZNI8yEWaUdSzhHTK+CYKthOiiLvSwIBgBD+lyAx5d0rtfLwboKG5ytopOtQuIyJs3EUo
kaxtUQ0JaxAEdiKpQTuhJOIdx74EQXhNG6M94UG1mn3fVphLhGJRgcepho6sZcm1Kk7fO6/OKBMz
yhzOt07iDxr3xZSLieUVb0J8pHEFsPI3oJ9DTHWOjtI9fibgfQpToe63A8Zb36afn7woF5M5mH3d
OPrqb3eSeMZBEn1YKRsnM7bammr9h2E2Xqou8JRdW0klyyw6ttK/FHfguRtYmXahRoI0vfm/VJP4
pC4fwow/xzaK4fbUoVdlU8NABhDCJ6usX8QvadAVisVp32HFZD/3VXq7TLvo+lVWpDxiY28hE7tp
1dVyY7zsBeK/0OhTj2b0c2N+6lIm20eRnqZDe5SpQpUFkSygBcT3/hF+r/vLXL+qFmvjxfOuurg1
nG7ZYprRXzefNKsciKk9UU9FfgwR4A3dPHBel2DTPDVV3NhjGt0uVkilaQFD2pki0Ar8dyVPxdq5
2GHRAQzTaUXv9OBi32Yu361xph35i0JrB+QuLa4CnO6PcAqcep1jBl6vzX08+rNx3MCcQsIK8qN4
re9CLcYHvlTxxHouGePG+rYzpRNJ+BUJ5kuqjdybRLgqT+rF2PGabv84GKdOuGpjNSknHoIKIBkL
UYkZKHhr0A9fccVhlnrN9QSYhfqgOh7Ai4Yxm8FT7oMdUk19f0WWlgADShlZkk9HvAczbq1p0T99
BhTeQPHfcMrW54Q1t2tAvL114FrzKf7U6oz2rh4EpEDsCCQiqaG9thPDxn3wMHKGlhfNTieMdUBE
hgj21y/c2/EuuLS6GQuSeCyhwSczLmZdI45vTG6EwMkf5SmXxtUV/yrXdeplrKN9S5YjsBEbtwpq
h488mXHS33C1uPG3Ff6Nv60sY2azxFBGE7aFqlOIyTuUd9k4/Tm/j0XXCyqsrWe0TTeQjKosrVE7
OAKf2SytL4Yh+wfH7zUbXpTR6eBM86/jKHsMwDZRBzBkdZm91s8JvybfxTGiwJ7kj5Ek5gfoPEsv
XqOb+PZQ/ItirOzCOJ5ywzaY4FLIwaBouzA4VhPLYYZp9C4NSAGYyER9ArveQXlhw5eLwQCYlbMt
Hi1z3MaMaulbd0RyOuiSq/dK1HhSwWiraJOlOvb+wOKbSKaCpWgdU0RdQgp4uzvZINRT4mJ3Ez/d
pkNYgRV9gyQt5CIVPwJCv3v6AV63tpxbWfG7ndlMVU6UVMMHLGIu5kEu6fRCiJWUnJkh6IGfA9PP
j8FFX3Pt1KeYZPvcN4nYdQdtKMp+5BKiqtDZkfVm7Awc95klknmz66L5+Skawqaa9cl3+W+gigxN
CeMDMT4Bw3UG7gmysZRlXXJZ1AaaCOBg34HVnsrwXY2Mlbe6JgkS2jXN8vUgrfdvflN21aLxbjgt
BW6LzvpD+VksxWpH8AY7F25dFr8/m7K/tIM5IDF9sUNMYT1StfIoS5u5xKnV7M7GYvlIH3K6kCV+
5qYJu+Nef8ojqunqi1D90azkiAOB67C9qIv1hvAMqmEIcByv6Wml9908heSDWlWYiQhDA7wUGoo/
9dT++LXHEun/68RX2VJpwVLDagorvGndwFUQcpuppYpRryv4IGAYIu5RiIBTvvdEYuYKxZIignea
sbP6XvtSed/koLyK8BNEU3A9JXqRWPfW4aSg30YiKBNEb3gDJPo8CGS0GPU/3A+x6R8xAQEDZN1J
JJrH55v+ZV32leBMwN9kfLhTjQhtrxgWwEOuM9kOfeTvhpByhD7nmRJD+N5ezZrnWE0Id1f7wQWP
Dl3x27ozS7JkrQw1KwTxVrwwRw+DG+gdo4nwxmBSG8n1hDK9VF91XrFZ00dw2mTPEkOxsPlGpF/U
k3DBGIe6lduhQCa2qV5t9j2ZE1iJDkBkOb4dM4bqAzCI2HUsKEyEQGFwdn1cxBo+gqhmV4WOBkP6
5KKFvuXj6HdPsSMCzj16xuZG46PjvnjT3c2Y+JbVXOY5lEJje3Iv90lG8Oay43OlGV9LQvMl9uvu
i96NTNW1Xrr73Q1rFxGfhhxhNVuyCO19VQzCZ9eP4etatX/FW2eQZH6XK5avVMzu6vJ4BFJLi1h4
slLMLmgW7yjVWyg5wLmNGgyf1U4x/sLK5yAuXIvge7tbeBo59R26P8Zu8hB9dRgrcdYhqpNxcEnX
/IOlgmwtM5ZXa8+bQFHs1s9vZV1VDCq1B2/Ha3b54l7N/yo9X0ADrDXU0QWeLhAxq2qX9uLuWCG3
nZb3unChfxiyoYNgEp77+LigZ4SM1kdUPF0rVDHm0Id+rhTzasA5Ov6gq/wzt0hXkh/8NKR2M/ie
UVurcDJGM1zWj0Mc4SkeuPpVl7QBveYfuSMMoDayfCTkEs6mZmEDhF93o0bp8TxoAJo2CP7PoR/3
FpyWrHqaENDC6cbZmAl2XDQQDylLNc5l1uzIwd2W0FuZ3AsLQWZyb7/Vi1eOFAvex4ScH/g9hTXu
fFjbQLDq+bTlKma1DlKEMRbfWcFJGYSqrwlJ+kMjTkgilhjmp6lb8Wd1YmY7zkNOIFAyYPINz6ST
f5tavVxim6RVAmeGGw5I25fkVd5BkxhJjmyy5SVq3MfVLrDYi4Wnb1nLK3kueu9VqLMNSWmUN6at
eZfgMHwEhtx5GHlfHDE+SEAGnPnXTFHXoAdyCyBywmwwj2nriVzM/MgIYXTk9FhF4Jckq8nys3nm
Ro3NEP02JvPk/0ZF8UN2JdxSKanSHLbnNKIP3s+z5iP3/FgOhHhQuw8vU8FebmEg7Si0HfhyDV2b
N2lndKKLmPyvaQmOfDHqr5XWy80eZH9qWxHfagrNJSL8/rM9lMTwJBzG27GgFU1s5HQT1C2KWV1y
Z04peQe7OoE952P91FSUSXnLU/xmd4INIIsmuyz7isUa2v3yCT8MNrsfv3c8tIi3nn7rKPiT8D9I
eS0M+bP9GkAxRwgrVkJlbosKp3B5gXBHQOsrNfLg1aZX+ABJl3F6pSWdVNetm2YeKkPrlpvS0kfT
BbkcHQwck/QTG78jnLEPL5I++iKzqLlvtAu3k2CzN/ZymsaQt1Mwe3YJYxXbN8mnKjB0PRWQ3WH0
gzkyKQRanGtWIfaecCOLLToIlx5bqwMjj+3on4zBO4kxRJa8zg3f73O4zBIl/k3Pt6WYHgG8TyXu
D/SIsaWhvuSJh5ctdxyxnKjqVa6AezUXMBPtFXAHka5piArLb/YFodWhmqNOCLzv9jHTzCtS9hT0
6D54gMENEmawT4sv1IfH9owUjk1NpEIO9CGnrooJiF7YaqP70DR2GSR5n3YbdiLuA7u5cpo3vR2v
VgWUKC9q21rSRJyy/6JruSH6lO+pJI4EU5WNudlNZX2Y1ya0rrvD/ryIEfTqy79zHzs9rEZrx1DR
l2HiL4YT/+N3SrCyqYHew8TTyhlpuBtdTwRwyR99yAt9qVcutmzcUhIEP8B2DoUOnByjLjo/LWf5
sxTsAD7Qe9SqNi1Kc36bWDcjPk3gQehKvsifszEt77Sdq6qh/rxCpWa93YqfriCrMQrmd0Sj17nk
9dtI48PBxN/P4Xzo0HvZ+ei0zXAjL+JqDfqFXijc9Msn30UwvVSHNr3zRkP2Egef8x9L/z5viqIu
XjdwXmJHh4Rf5eEf6rWMn5AXf9vaQOApYQ34Hp3O7vaqr3PsigjvVEt8ozAZykCDNrTgEaVJ09Sk
CUuy5A7LXJ+xxRfoTYkEa3yp5APsRnC3icLfQjDjMm1AfCody3JkOJvKUxFZYylYfNwmMsuZnSFR
LUGvU6hMGbjP/8lA5xlkvDE5h4V7Ur80H2+j2iyJVQRSscXfu7e1fGmEQngvpcbI24OJ1oueX3kU
RZ8+gk/DSnHPHwPTyEt05cJD/Vq0L3xqj+tqso/UrMfwpykNgyro/02c8bfEHdCOSQgTnStPqagh
kW1ogQAe3rGbPRtJVmyMArwIdt1zc91PX2zNlD7ev1hbAh9qlcsj4OiuAelluG3evle5qvpO+9uD
2p/4vvVcN29carSN59FpX/lep6976SXBmYq32B4xNe0bwu2BCm9xhbdD4tFmlAYnAqABuuhPQQ4m
+6potCQ1hEwBeotBAd0FrEERSTlQOl+LTfoeNoRIXKQ1KgI/CQ6RzC7pvTo1ernuPya5clPJkSMf
cFr/yPdh25T3V5k9t75MaJg+9lrrch30oxzQ7FrUbDNVc0hon2lFxvF1rXOPwVRK4RNyQehCSnyI
gvYquWB8gUKmuUjb40DnFdKET+2qN/D1aRyXNZxJZl2qY6+/OPZupo+xWxoeqx8ztBJguCkeCUsv
pmaQVE3IJlj+zet6pCxvmgHxAWIchkXiA8VGdOL/PaTMpehBMENkU0v/0d9fHlBrqdU1ZoXWS4Ew
t84xRiBSKGPc9fPRi4hLBYMgdji6o7gfAFEGvo6pii+q3gyg7Okg+I6Tu2fUB6ZrA8DPBcyjXsrl
cL4T6o+GVCwADB8nRTu5EboN+ciP5GTTd+wAeAyfpuSrO5Q3+G4if6NJmtcv5pR86zGCn3UEbEzQ
6wuOAExInpsn4lXoAJuIC8YCKwnFijsdWgvpI50o5l1NOxPfVvGd1lBdkUFhOWxHhwg6by7+Jwjv
YQkQlQyrh3O1YAAUw6FiP2hcjtAmB9Y02xMAuPVQ9RZ+9aYnEHGP4lOCaawsbcOKPvF+lCQ1NWf6
i9HEJttLU+462VdN+nTtk5deBkHVPj5E5PpgX9PT4SSe1PpkKSquQwRyhiW517PmDkQlPX0TJHFh
ZGPxt1YhtcRu6gMrwfv/XbUP9gUTS3akLplsqoxka8NlACtjqbPe8KrVnGfhMTFOWHNcep+VwRHG
0YH9/VtlnQcRZ4Rmx/YFeBX/0vT19Dhtm8teFV43JVzPpileakPTZzYRWj1ZKgECsKtyUtkLj8Cb
/QgC9ZcQUfI2fCP/kNl6mu6PwOCM8MO6XfygDIZtZsUNoMSBTe2h+3A4LzbcNixFot1ubfK/1llW
+5aXNS/ahDJk2kiLGAO3FiRWLyliIuqjP1JB8efdm1JEkYuw6Kr+hu4wMlopMpk7PipvaR6u+nl+
5o64a95sgL0J3PpOugpJxJAC25WGSQkzOXvydLGtgeCSs5BRvLMnmdL4i0T00k98N2jOnNYHiFgj
LulKd0f3F6A5oOEdwcBKe8ibj7gkVHghCn7mZbriHoQrkbjxaZ42EMT/p9hKb5mMjruPTvF+Sm72
SQLZoUcMTOcbJrNK82Z2xAbJHRDvxj4hSW0IIljRtJ97lHtMXecg2GMWTdsj30jkjyoCcNpRqO/j
tbCU5KHxHhQp+ONscJv18Rc0o/QFG+cxX2cxFQ+O6EokA8SOr6R9oBPfHHk/PkHGt9guNlK+Jz7V
5NK1dpd6OYtZJosTlvxOiWkq9CWK5bOt9I4XIc1ZA2BRNcrpbb2BUIpMahgXP4x1yiST2I9KZcxI
yATztvSzDtMWnLde997eOM+CAIYcxkHVWNpPeSY7KsrmH6V9cAG+P8IoI9hTpqgIrkiAs0KLDIdL
andxe7/AwAXq4gC6qOluctnni5FIMzKTT7sTYkGDbw0dnNQoLOlxdlMbjbvyZrv4JxqDWdZ4vLPD
repSkTaugp/SpB1Z8ulHFsDT69W8iGmOs8UZD2v6MXbVfOwbZGi2UKet6J/odpLiDtlrK28vUVb8
4H1dlQnsT70THGq+k2DQ4wPgMLxpxPBa+04tclXlYCt4BC5CNnJ6c3TvgB/cfzLBmc3lLvgvhI1J
LHC1lMshwoPWiLnOaFoDcls4OrHkjUWo/In8a+2g8EBeh+n7kotj922m5x1KMd6FQcZoDm3D58bF
p8q0XXwq38psgw7rEm6BBwbb4nmp3flduKJq+rchyo421UrB/XY1xofeAOOflocxp/6te2x/Kacl
qmljdBtwIhsvG7lHr7R8GuOkZaCRzZrFdj6xHMdVRbn991tcutaPlUprVWioS8obUjVQ9odu/dYS
dnAvJWfqTgLgvI6kDWBsSrz9ynqUJY05jwf/TKvL7GKZW6fl2ytetbxFpMymWPr6/7e4zW/20T+K
AMHJb/ZekM+p72su2pZkJ63FEXLyo6BMqaIRzwT+TefnkE+wHmULWc/ztaQ4aLebgvabvme5Kzrx
E56YSAb/ABvcpoxdLy2xTOPvAwourA6XNeEqc+SalI/knpWpeXh2Q7eUomhMbDQ7EX1tIdoni6LP
vPQ85uHPnXdlPoiTTzGDelxOL4KaMKxv5X1USVLikfbKr8pfmLaDJhvpR6UWwYd7g4KKmj8Bm9yA
c4XkkYNspnzHeNtlqooYwEtBNlCG9JMY6IDBTnsqUB4WsNo5zxA/IMavDJ8l7GFKyDtBWvgbRRrB
NeGzsTwP7DPDWBLwvZ4vHPhabb79fRp9Af+E2uPD2hchld2w8Xqjm1o52Tts1/qZFyvwz8CqJuAe
IVro+JfjDQZTebgTeSshBFKVwuCPmoA9kbwTxso19xGpjeJNvhcNkJVZqN1y398iaZROeiiWFBm4
gH9psVPl9mxNTFZ7zIt3H32y/piyl7ohyuNzzhY+b4D94QoidBIBVsFPvhsHRb0rZpdLUEOCauls
8ShGBTxyusigLk65CiOdYNSyjFlG6DJiF41wb1dR6EdhjMPfXl7E6x10PXc2+vuLJ4N7UN92MiMR
KIACCVUyg+7jJi4sUgmoBd1aP5wFIAtgsiI7pm4VwaYmtatpZjjbQbViBP99nbJPlylCtGxxOZzg
tBBJpyn0O0csURRWuwiHnv1UCsY9d/dfQFOaA6uyJWnz2Ls3afERlN2CsXQmJXZUhGFJZ7KLHTn7
Zjj2fhUYCbLQFnLA/wdVXDpCTpZrtOwKkNG/3epOKp/8sKtH63CRHfEHktmYdp3Av1mmmokp+b9D
Rf7LfnbzKF5kzAeJpGJkGdajfKbMpLRvcTwgWwoMamBw1t0mqyt3rlcmSjbv+jZUiKsDXYC3HDKf
GCk4dELxVvm4v/EUzeMdsr54DTjgdkLETP909PfC6ppujSKQRlyjyx/6hFDgjegfedljIvBlvJBW
0jP0JkD96BV5Bf6Q9M0WFI/STVFJ3bl/OBh97e1VwDHYZ48uod5U9lI16xcasgXfmAerf1GiINC9
if04syeQMA7jsjj/2x/2YGHjlwapF7Q8IxZ0vMFAlg2ye4A5oPrjlQ40xRLq7fAvPPhP9JqJ+mdR
/MOkMUleL4DyhN+rNtSv6qPt8V8NUxZIv+Llzbe2iiE78/JFTQhzDCdGKa2WB6E45eKP+TMwUATb
jZoK3V3CfQWChBEmiupUqGVmnSZGTk7Hf2jz1Mcy3QbiUgf10sa8QtqVE8nyVJ6XgG4xPPzyljHN
Vr4kV55olF5sZhirAdqLUhVnbbfIKR/x1UnMNCJ9adYxWHsUJu2DLqZszCBb2BavIzvWCB2xMQD0
W1IIm0v/PnYxY5BOGQs6HKOdal45iaNkbMq5LzF2gs2VlsaWqqy6WYeFdL0dHyqXHwLQQGElIFop
rOkJAzgTDwvq5c5TIDFfNb9zt0Pvrm4zjEHjnjZnY96nsUm3UB3Dy4WQds6VOFxWuiF00OgtH0RS
Y1DLe1GpTvrWuh36HxI6ltGSwcjv66YLQ6dIFk5UGBBF3eLGisJCQ5MYcVTzeCgGec2yQHnRLIdo
b5tA1Gr7hfTjKBekD9EOQr0ltDjxHGtO5AjrJMD80pCVazfFRvJdjeQCkmMCr4+nt0Ki5VlvLrQM
hU/sf8FTbWqlXDLtDC0gjqH+QdP/peuKcDSDgioR9EGFXFVW/yci8PAEHJ0pbUG2Os+UWhzp3K+I
/mSlwDFsIEQvPppHaRIYBYk5wijhr4eojbsA+pe4TNmqZ/brqPPLLSai49icrXpDu4wBJEciiFT4
I+L9rOpB5heww0lgUjrc0a9+kik/oS6TrSwSN5mkr4A4yf292+NMZbcNmJAOi+c8nbgWF9QFu+iC
Q9F9blB0vI5C9f9M5StbzYupM25xP+0lpDLPYWwoYmCr/jpoo/PcXT6Z2eDgMsFIS0wUnmjUuci5
/4GiZCjOPyY1MfSivNgt9+G8oBOZ1aIw967f7kYqxMH5OmUx5JUUTNOkOYR+VaSsYjNWFrTFMFnT
AQWyUiqpvPCWHqfhaphcqklP+1t+vJqnynLu1WtsmdqdrDi4HaHJX+mZzXK8dHg33P4MtSZAJfQu
0emaYjnNSCjJkV9YIky51VkRGOONqTgGofVoIfNVZVAlS81YT31x0/ZAdh4u8uLpzjDrGJPt+5rE
xEKw7HdOc81P8490vLBoqIuuH5jR22iLsoiFeJpjy1yS2P9ZAOiECScaTT9x0s0+prdGzpcQXJ1B
8mQi5Z93ZRmdjPP6GKb94zoGrHh2MU9qdXPCxI9wMwk7oXnGmNZajJ1qQYzrcLGLvi1xcl4bDH4B
r77REf4/d2kRAnGUPb4Sy06HpRk3WzafWm/KvoADGAzWplTkj6TENSfXifFuvUafE6OoRwCRMWOv
TUCBtKdt8X1TnMekzWzUOI2bp+MUUBTe9YIaAZpxQmDfYja9dfWTJrCOsY67gSWsb7EeZFmmv/3X
rho+HLVJPzNv9hDNvzolDLTepeQgjnXU0QebQc5QCcs/KCWdxd2O7CatGXA9kjJi9BRydhDKo9uK
c3fxyDX6q87HJKmMdL3AdSuheH8LTUPz30MFxqPxjBv5jz9/qiQ0w1X1JTpV90kJvVGrHKDgKYbq
qupN2oUsGIFJ4nwzG0Zy/a2WQIcaiHrbnt5hH573Q7Mg1elH3syBeLDsiUZ4VjacIko3ObfE/rk+
eJuT7bWC6GkMpJ969EyM6UAxUx8txcrF9TAUOxA98zIbskB33MwQ1svlqHOPPXXSrD4l1xoEl27g
WuMUpt5DM370zy3m1bYy7sKvcxgXzILumiSn5x0CmdI7gJ+bb0eHfPu2Ec1i1DVtUf6TBZhKNz61
YsdLlaXeBmIEXtEtzktyP4Kz7U64I2g2LDV9zFSDoMzDD8MbpiVtRzrPWiXr/sWsYAyIZ/Z1Rm9D
ASgRqpMN7QZvcMtsImj6+5+2tGO/G8KN8fdfLbxpaDcKkajw84bNXMaTvpJT2rhJxqKC4hp2LyOH
Mt7NimR6z0K8xjzqVHyw1XmCdvygtMjSYuG+J8bwS/TzNX25uhOMzUmCPkzvD2ZE983PotCUlRkI
/MCunURQntm0kXgLBRhFZmKKsXf6n19dEuxFdSIkmv6U6D5GlFxBCI6NrjGa8WH0hIwB6prn8oSF
dAYd4nS0PVt7nZlDGZCGw+AcfCgeG/TWsAHKL4D0KNEZr8J9qnhPOzopmIoKq5ZwmMTLWARmaIRz
vXOe2zJtQrDD5bL6ndJBmIFV5j3BJp7NXhbHknE/aVQOHluapV6uIyN2rhWBcYSctHPpRIb/VodK
NpJ54b5d1Vqbcju13cLjOEKIyNZLtW6i9cz5nh+N3ZK7QEWiGqFEZr3OdQEaWW86bVLUGfmak/+o
3F9tUbBRc7G92OZ5YnqK8wzXIsp9myoxSbUEYXeC04J7uTd67IeIBd4cHlQBqSiA6q8h6P+mK0Au
fBd755wgXTAyt2bccI+KuNoQBJa6j4S1UhK/WXpVoCBU3TRu+8bzhFPeohQ2nkfu8tH06Lxaz7IH
/N5S9MrIv0vQIzYH2cHG32QHnibicAJ3gM2Lc68CQPrrRxRA31gRy8OZRJq83h2PDUsaMsQNaehh
ftDtSm4bqenKWXjDBSxv4OVc2MY/GlrrmNSfWr6WuVPRX3itqLq860SeQJBy2Z9njWqBqAR6by5O
YCsUCfBB80TFKewUHlHRiMcswEwjFfvwjHiv16jQwzaKbs98NvVmz4Jyvlx2lBfjXhfeFywI4FSB
WOQEJ35zoDljxJaO5gLY4iLDq/xb7OfcWnqz5gc1ll7OMYs0TjkBC1Kw5d1SC4oFVeq40eqBALsi
GAvq64zhmztz1OhpPz5fLVsbVcT6CWRoAPiJEczulhEe67kGInyJWeNw3suV9J1NsN25gLyqek0w
SyHZ/vqNZH0V/GMPrp6pQ6M75z3sy9cIO7sUDexL+O4xJG35Aki8vT/j/nQgYW1h1yQRPS/pXGXJ
tCQJv7vakN3HHrcDXbQPoBpuq9H4YHoQKJH5YQUdy65MWWzpnIaz5mga8c+Q95n79ycwM2vBaOKn
vsRiZMgRz46kcXZNq/ofNBBPSv9xnxhrxB90BaCaXD5ZxBrmwu38GbXhk5/Tl7Q10TP9pckKQbZo
BJeJf4GoW2HwUi8ycDyudmYccuo1rPSARUdRAPrkyncDsMSowD+r0aTrG58X0hwJOaJOpFZ+BHpH
5S7cHNlQQWXwlqIG5daHzDIClnC2yIM8KKP72voHXQ009vY32xnrOkLWF1S489bRU1Ai6oReA7Ji
bUa8dOt6FUCWi7n48edxWI40QVcFxNxkK8dxVjHUgAgybdJHtyg7ND7UitbvOsrGnUCLVSCNxx/a
P/ZfyALdHFiflxbRoHKUYnOlv/9inXdzX18zHQMG63HROaquxyjxpvdgHCwJvVoVlCVwfWPkkcRj
h9+TBzBb95zSRi3UaT//Z2tDMxYgIhOwkM6rdYsbNo1y3gM7HWGTvwGxrhRa1OzxHdUKqFbX6Epp
4+9iaJt/GfGa/jFonUEWOMmgq7bMf/ImO9Jn6r2rU+xauibfD+nL/KoiQNhGRd+kjDmMkVjILdNi
QbmcbQbR5X8P8Toc2BVfga9sR3iqFzW858hYCOJA55rCCGxqfegLbssENb+DLkRT4I2LEbsAOViC
dzbRE1lOVOryi8d+GNUUkphboT0BB+IeH97YBVZqJh60Bu3UWPP+2yW2lwsyHQefo7hFVHJQczUg
A+HJ2bxjDDNHUnKeOML/bk6cDu9+jp37AfbdMu8QQyzv5PzyV6RJ7jqput0WHwTXLLsb/cx4o3Bp
SLGEMX0UNnb1N2QDuQADwXugIKj5eA8bkpWdfGHoCeDUKHC0RairRKriSyFSNv1oF+njp40B8NDP
OuW2GKMi41ufeU+F9keUMMTHPenMb7Y+izw22Sv0FpBZCmtrlinvJrLekAUkwmjAdvCog3XSC2ki
ZqDK9Yu+CXin308I1lopsMSHpdGETMDI8ilVzxifsYMMFCqTJvTxBPYKcqKmzY088NIxb8oUufIC
/bwaVgOamlPTD0rAdKjuD4u3MUIR3HsSx5OdsB0gq0pbb+v6tR9nQaYHdITlcDb1G6Wgm9w5LwzL
TGy+AjDGFD09zyiLH/dsO2yqOelAb7JqAoomHlnAbEv4ZfbIGUmeBO0JM7Qmw8oP93TvVyuJs+Uq
eartwD4zAI13EQhckZpl3aGI4eI3owMxc8/0lvcb16tFS9+SwW96oPW34/+Z3ZB1IlsjtIKNnaRs
lCg0MyJOOYXz1y0B2KhYtsXlXrDHTGkCxAyVxc/V6VIJCNLt0UIuwaVuXkLLIjsH6yGtsY065b+7
NWUTmmIzgv8b1FlVkh2EPZeHZG1oHnxL2SvZrTKm0j8TANGKL+SGSd3UbTok7/LMyp8qoZXyZGI1
ErtI3eKgJMo78a7hFCcv3CrtMA46pTo4HTYI9eWTgWiWW85qiGudgzCbBB8TKYYnxoOAu+qeAlIh
cwY1mnIiz4LrdVpsDQRo8v8L4S7+zhuQRk2tqF/mrb/jz5UWDonJJARVhH+CZG6hQPK9QH9grkTX
JQDS6Ls3Jt70O7hfXSGYSUsdgCnjmw5Zf4xFWnxl++LTZNWbzT0EPMjUSr/rYCYB9rX9ul9JpLcK
1Y+upny5ri2yuARuBIJpjg+5onqfoL/OC0cJKgztT31hX/zS1N+PuvvsAtEka+IJPk0w6NZffT4l
x+FU4Gt/rkJ+xGZdgjL6tTr5bLi8GMxIA32VwMA1HLj4umCHyvkQw/KNxQ8+eznhgvPSUfpdeMMW
cF4730g23VS/3aVlJtTsRB22sbdPqNL9qLGO66XRH5Z4vtPCjPzj26ZWjrNgVrJTMzYpvXLGIMY4
tHeDgXTFjqtrwYuZ7GV64SWjeuch1peqV3mVxpW1nc85ZmMQVCM2gaoMpA+FwjKwqjd3SlTt4GDi
nmrYiHJsjjpUsBGarJgtT0DTy5Ie6017lYKPcNvI7LW8M7h5lC2XG0Ei/dRhw5pffmnie66TbuXv
xtLQ0SjyffGtxle+MsqahH7jURcEri8hfs+WS5AWdCZZcIZaJjl8rrj+PFCIQ6RUIRgAzO0odYnI
rAg1XDhZDD7vq9dcp1Ix7RDcCPQsAMPRvoZkkvaHqR6NhYhzAsfOfVAD3aOrGp20dCBV5bRJ5hJZ
SWnMcNnAteG9tp4mme5KdR9yjo42pd9sdFCF0rrGthv8D1GoOkkAtGLD+HG9QZXzCaHouGYTdze8
pTs3bLdVXDVuddLKkjmHtAvJbd4AVKcQLmtWFQOzlzAWDPyv652UWkpuWJryy3sPuTsNSg82GdGE
XHI8LbBPUt8yVb4NsEBhA1pB0esuTl6tZqrKKueYTa+z1ewU3p8YnMHixQrb3TSQncCVLEKgofyQ
EHijArTOz8W0p2ivFpUaP2VUcjCAqB6Pwfy1FGZo1P9XnGfP8bKTQa6s7cmdJA9NL4FzawEmiyAS
2jABnJJ6RUb6prBofLOOYjiDVN0PnpYLyXgZ/tUQuOpHP1tQQSXmQjyl5+jzHoAG3KAMPJ6MxKnM
NTTfIOAh/+5YWy32fD5jE4g/Szw+OskeaFJuLsIOZzN1dT4NL/hN620X/SqWl/k2MJ82njcVHjSt
Dwj9aMO4zcJLS4JamWnFFYuQaJg+DneK9Z+bE4WnpRTKG1rLbnoFvaQes2CXHRWEkpqWC6WEYNY2
Z16BWFQyZhCo+dT5RvSAFOxCZ9sbMiuwuevdGopbIlipk3UdRBn4GQ02AIhqJIMWKgURFyDXxw0P
49ZdjAnQLOv6HEwaTOvdX0lqmwhWoVnEkiUSqdD81MngYuSlsA/J/tjLWMbHA39Prq5x/KHOXKd3
0WDwsnrdsu3pbDzMp3/xzso/tNgVgog8ek/7Te7Qje6vvVwaFWL2akckLuGVE/uVHe638gxURYec
FUVJz9iXVLjtPMTuzI85N20MCS4CUTepLX/Q23REOLJdehBJDTosssMbWuu+ZEYqX0NXmzjmVK/R
UmHLL70aM6AMIxyyja+rSSk69Ptn/l+Rpn8t0Zg15XYFa2Rfhm48kIB2YZKLVSTLs/BqJ49WrH9U
o4DmN2Mc4qZEO6VVZ0c7NuOc1/IlTgqKr24OQIt4TzPwhKCwryxQP/qv/eBCop+ZmqCkREGFTC1o
HMpmYh2SGjLAqr2L2+y1dT2cV469Afz2DBlWUj1aeV1zzd8Jy7sw5pfFulh8oyj/E4yS3MOVRQGY
+g1lFxpczUL4SKCvTKhcMEVh6GbnuR8qFRTt8sEl/g0pYou9xNKVnT4wMRGzF0hh6Si+trjKhwzY
ImKIObRwXbi/6HpC8AwddgDmh1I5v3hssvxJWvFLzTJNcBhJnakYeMk1syx56jqGJPPuiRVj6cy3
laUskIBmI23iDNY5iKbqG/W3NGkVEry2z6oHHdIMiiqYnRQsCQaNs5Xj13kSQ6cKHEUmb0moVcJq
XRhJC65KLkDB665aC2UEyAuXuC79Ak7OLqrJsK3uEPDO3dMbCfs/AgnDrc7YeKlbduO0ex7/oFF2
GpZ6n/KJPIdwJuXdWAohQmk284wVlGvVUthQGGNrVfClhrtSHnS8aR8S9DqQ4MX3FSdhLfYmYgeu
UwXVi2xC9B8XGAo4jTlT+ABnC6hwlZJ6R6JCwmEjiO+u2k4aT142a4bi9naI69H3ms2dwieR9xXr
/CfSmnZUy1k9QtsjQuyjAHoDOAsZaic1OQiXpVGNsm40fbFE9SI84+j8tsb7LMwOw7wXtXs2sQQQ
ELGbnpWgZFpbudONUYy0jnUPacivq3NQqJPeaZ7ML7JAtHNzeZg9StHek5OWn/A7eu46gJ4RSFq0
/XbQr8PaH66EmE7oOMFfYCx+DltlrvrUwTK1WY5NcbR/o+FZwJvI/EyausOFeAE+8y5EA9T1cx1g
d0/eyvzUOK9G/wnWJQtHR1NIXm9Qch/h7L7a188J90SvQ/6GPUTLe428PRYyZE4Lr5TedYqdaEEJ
nugr4nwfVerqwgjy7re2muMs6Jzp2BdEGW5EyUQWPLQMzEc4VkYAzC6vcUjwIB2Q6AaAUtgJL3Qn
vOQV1qA8tPk9lD70/k88A8CPDi4EKr5zEUB2bK4fdvQ2rXPL6m6KC+lbnaejRaUmG9+u191VzphW
/67fYirmPLd31BTFZHBE6Vc2NG70efV28bpCAHOg/G5Fh7//T30uho5h+rX9FcPI87/1hb46v3R8
xEL6AadAXIMAKl2vKkv8SbqBP1iIKJ7wgW+ciEuIkAxFKIj2EqNrlbp/z9SFKxygkf2QF3jjOsdC
Kinie1TWhSER31zuHXWcNz74vG2Ke0eRs39MDFyQXoP2MvlYlIiSiQ1THul+iEckx1hIIjdJMVej
SOwJEcXaPseyt7LiiVL3rR7csBy5PzJmcFmSmGU3KByF/kaiQGceaDMI6xGen5JpL2dQ0kCzvfA/
nnWqVTC5Y4qdE1Rf1Az7y0VyQk/+HuttLaaQugNSCMNqAwW5jmT3yWbUkRuw0thO8YyXPuvpoAip
PkMSacvrkSyDI8D0brTF767uQOvxmTL9n427r7ziFVhRIEAp+XLNw73PjXsqQIN4xiyb/Xp3eRoA
sfBB51BlCl7POoQa1pv+ugX/WrzMVVCAFd1Hrz5GF4wN6dWzfZlCADkStud1G5uGFbVuONUc0s5D
5NYoQZ2aJtSXn9Rpafm041C78XTLhPFLWhJS3ZQFINzZp9j/XNjiZ80t5hEN9gldeKz6p+DPTBtt
mHXWLX0XnRHPBbuahNlpUImKMR3Udh3b/5YvdpJ7MKd8Lc9RwFpYGkRHKAB1M/ILiAxlrkK4Wkkw
IawrKQ4k4MIlareqEYdqWH9yz34RpNX7h2LSsr6tqPaTkLy5v33Uhm72c/2bKzKx67bU9L8O8pSt
tOhsvCwrxroc/cbeoXgBsMhFyf+UREBm/7gnMux2PY4Wv4og0CSnOB2hRxYf9kDAPIL/HmpM5afA
LYaDgVyXTr6aJNDRjSTfhMI57AyFrSp2xLXF4CQfG/qNY+c5oLQq1a3/bjCx1ufiJlnHfKRVlALp
mgPAAmxbrs8SsIx0JmKJb3brwiyGERlXUsk6xjttxPGEofUyMNef3M5UpJNZKRaXJWOuwhAghEQ+
AZGCe0DoZZB53L4HkHV1zXfraHQFo1OXyYhZ0Tpb0HHWiFjA39DnADpKRqqNm4zvzzauzl2yPetf
gooY8Y4PrNKdAAmvKnfW4YXpMbYxHAq5SV3Vv+df/QQsrPZf6WcWFxe6j0Bq4xAnD76Lvo4E48jB
5mN/GaXkhs3x8cRIimR64S13gbJHVg9ae7vCaJXPEvlDt0AnX4dhhL8DUr0Bir7cSQ9/J+Iur6zE
Vpkp9YL5ng9V8jIwBNWyS+16D1zJsQJ7WXIduX8jH5eb2R/vMPhVF5eLMQMJDUnQGkNP1iETj7Fi
qldibPYBX+8lLf4eY6ap02mwSexUPoUfliEfexYIempodKICEwdyjnVckYFUSaxb3yErN31HD1OI
0WyUbNAFmIwssYE7Vscfh8PJ0w5dTOsyE5FMMsfw7AiqBr9rBWWq4sJV7Vsf2jOGNlhR09ysLKaf
vQ5vZuRC2jKj0NEDeCbF5PpzwFS7Da+vp7FflkvAKVr3EO53V6JY3Dx96b0A47j/9lGPjkjhW/KG
IrQggLoUZ/SKsr4YmxfvsdWMzkyVMASuz51pi03nrdEQCOOQgMf56jdbdy0NTPojgJ7NINeneMR9
UEx/3qJ4oBUyTnTmagcIJSsuQLjea7MDP2OSb3WjrDMiKYU+36/50VtoF6Dr4Ux4hiuFnk9FjzPU
EldLyY2xCB+a1FWphWt+DQq1O9I/yjhPlaLBF3qKFTG3CumtYjELaAiwYN6Nx6Dtqis+wvZn/RI8
nFfbyH1xtTYzKt3zFuqNbDba7vsz/4Y1m6kR5/wHcghx96ErHzJCSehKSjZiDT3/51ukIBrR+hQd
Fx3ylyu4tF9bY0dXQCVzyzKESqznEaR+0Qkhjv96n+ppvDCjJBWSrUHgZ7V5jwkMsR5fSd2LmnSP
nFqfIgZlEDX8De48+rr48iR3RUbDNQirF8khS5oaa5qkwNfyeeF+6TcDOsj32Ow04zzH5Hsq94A6
cJw/yZybodE263+amcDfiQeLJTP/dcL1vqu598rakb4FYHDjoqLXU7dfOSGF6LEFRz5Hib3J+wXf
wk8t1CqrGWa/IZBIennqXDNmFlWOTiGPKzZrI0dUN6W28lQm3lMJEO5I+sxkVYh3TJCSTXL+5PjG
XSLEDSmzMVFnlZlBJNmEqAID1qorxYJjYj8m8MCLcBX8rqSPcdyIhk/yKpZ+IxNU9Qc4SxjSTT4D
VbqiDFv+xrNH/ruzelpMXAAV1JOylk3Z5/jJCwzz+6ZKnvpKNSwemf4oZR4DTLSvt5sbRi8ZEu2x
h4Ymlcl9iVlrxuN18fVGdTNYzkV6JAeNunTLV8O7tIx8iCOhicOx/vcAa6bsjcxPl4ZC622kcvlu
vJdpx0xDQ01K5kQTz6SsB+A3ZgIvmlbXrKElL9cNI+I5wrXlk1h6gN8XaOPW5H0j+kiHQu73D+TQ
75oA3bnbfNNn/Tw4fGJfesW6MOnzzVm8ESKwpVEkpfmqfe4Kv1KysrN7uVei9mf6ujyzN2XhBHpT
aMGw5byYXcnZaMIPHIRdurV9rDtheV7vZMrGcqCpUWd6s1X/bJOUUnRxZM3nAItmJCRbFBLdt+63
tYSrgfuU6q7owHOlda/C48AMFcuorpSx8fL//SVKQKiCDf1uVypNg0RI6o4ulXdyG0G+TQ6iKM7b
t3f5l9KxKKy4IPQAvrIeNGObeWArV3lm3SomukVCqoHqhzKJrZpGfZ19Pxk96SkqpsdpUUKoQN70
Sth6PVe8ITqMK0wV0uZmvdOqYR14kGvYzM6VCGBwDYC5vDPQFLaqCo6hLffFC19OkjOtpJp6+Z6O
HRXU2qfVWo4nJbpyQ7ub80RHh3S3zExaEmUV8OB7MorgtD/pxuSwUpNxgmVjwwHnnUM3smgw8ch1
ZltujKN85z2RJKrGIwea2lr50+5EVOWqcMEDcaGez3WIDB6XaQDdDNl24INm/OQQw7fCTRWpOHTE
QfevVt+ToF7ABfHU1UlBEcH5TIPC6cZgnwGQIVEPW52cww0g+EtVSVwO0QO2MFrQvhbihpoQhW6r
9Jui6uvif3C2nHShUhKGtuUAlnnyFIh4OfFm+f0u8mNcA8Co00kleclguBFDuwI964Zu3xwhlmDG
qQ2Mpkx936NAqyye5SDDgmpKiOu4BMd74+OjlEwOpZVreStjR05gpmvK67X3gbF0HaGXWFFuxfSl
ykuTaNW+wgPjGcrhmrJFx+qLW088DpZHiQSg8p6RNIcjmVGr3Tq77p4WcXfRSPVVb+AnsV8l8Bqa
AktwCn2hUpHQGDBOVRhuU4jtaycG2BeTJdGh4RU+bTt6b1lOfx21UrZTs28Fx6XK9+FuiebW7eYe
Go6ktiXIJqODkQx7nvAonITRsZ6xNZXLLEsv9UkFS4u33Y462aSiabohASGI/BHzZQRIaWYvvJVw
9Vvw29rGlAvc/AWp/iqVR4FQHa9fWtNwZbBu+YN+Lw3VlYjGVqm/3gkMQheoFI4ZqQnJ6NTajHAO
eqWaoqBCXzMZZh8BD+2bvBa0b+tw1QL6PS50CpK7G9u0AOhXkirMg5PF3UAxaWlXBDQZp6JyJVaR
Eu1Vh403GfN7/1LnAe5hIgfCoZUzOqyNyGotOCCeRLo1zcud8EiELRGlCBMm+HNpa1NLAkmHmPSa
Bv4V+IhqDaUMoSQO/bjZJjB5qswQC2hLYb0Xsn+0ASQC1e59M86Qvx+gMjZtUfY4Qh5Yt0iAvsR1
Cyow5ZrXeF7A7N5ksZNRhd2wZfAJypaYU4oZzmvBozz1vTTvCwx+tU7j+34tUXqeoOpyvU9pc9UE
jUaFW2qrg+uIwCxulSKQfS3huudfxxLWrYvmUD+yXkLGu0iRA8aIQjD53wx439S94aXchy7Roy8H
L623Dq0bATdbTUxU+50+U+FEoq6dov8oA02Cr/0Xcqkwg5zIzdbpBcHsTyL/btFDFuQe2+VUkQG0
jkqOfEXxDhCZ/bC1rPvVUO63xnJ3yWXyvwZu8RaZv1CUOUxsuFG+JK9NotKdzRZxp4W2bEMko3v8
j8A0NDaIqeIPmN7KqgfQgTmRh3A5POfA9SgTVqYo84JXCxYJZlMnX77xzPLJdMYwhPGDW4rd0rRj
/gtqtVLby4uUCiUtAIO/KSL/bFuUjix/sRBTYEvGkDHP45/Uauk9+Nc5jdOFHG33qTEUxqeAJAg8
JSYlCwT2yTNsq81IdJvSJyQFQG870fMrf7+hBmhSdhM5Gk4hkKyGAvBemFY2griGgcOoyjy1u5EM
9JuAUPmt87fIG9Nq4MwyuwailQHWRwZJ4PmwnYL7UNZUlfykSLmlKEFxiVQU/R6slLrPR7vbjV7X
I2G9pVO54uUy+twNSB/+tgsPGZqXHskXhxIHh4uCN09flN5YiKphaoH7EjmAi3pLytsfD1FoAkvv
/3+grx+IKwgD6FIhx3k/AVJAm30dpWmsl6RHzytSFp8C0Iuo8qAGqoVJbv9Gze3eMJx6KrB5VEfZ
P57excky1oi5WyQ3LJEF76+grsLoVhvJGlAkJ23UbNkU0tNb9OOfUNZjNSrWgjKfsLOPHSlo5e6N
qNf2gjXkdRR5lb/3mfIFr9V0ycHcRQhf8hvRG5Voh7FPolf46H+lgNJ2RzjomeHmALozIYysv0o7
uuyRAIa68v32i3d/nSh9B3XjUG17waFNblOI+MQaoNWC0tqWidg7hDudLicOv8kJE8br09OctTgA
YRHIrn9jWjBEvLmQJP6/3R3F7N/z6MCo6/Vjcxl81tIfTFtsaaltlnYLemXSS0blxQbc8pbbTV7c
yEX4apswIRUTCWK2BdCVpTwM0cYSbNll/wXVr66tby5tMEvhJuypYmhn0RIuDtPAyX1T3hRaiBO8
TPkhV3JZ0L7MQi4aMkzWGkXoJmAXWqGkbR92jIJQS6sMiSzCkIM02gRDNZyDEE/ti9gkiaCwfHUt
6aPLMQa1N7iXcZ23RqgQzv810T/GufQtZGjPwEwGb0aYuna/fXPZxEwAy1yoMPrqoLsq4FN+mi8X
4BfV0PrZ/oUy6g0Vhlem+bEadfzuJPgizGlbKu0zWz5cqreHtpB481YYhFMFmR0tO+Ff8+wsP+KS
lcuE6oTpyggHuvWkN8OmiqzcAXuemhG++nhOMUNLh/mDTtiGbJrORiU5GKXyj0IAYA05UK4F4tdP
2W17x9PyzSt3gzshS/HfPLroG5ABAuyaZXRX4VFb+Gp3ckdhNCmyUxzVUBPbq0QF8XEbP/1f4npI
14NQL3nIeCW/fpuWRWenRvo7LqtLck/VCIsdnO5nca9iKl1dlRn9eEkxqcvx1cRHNq+9Q79gJm1U
8vz9sc02E6xFwVDUsSCW68Gc0fMuYL3U+FkIc3qKiJZtl2Jm8rW6S+qgmt/SVq3C7UUNqa9sImTr
/hDs171QF1KqGNLIvk+nkcI35h4NZTTk6CmLpQ0zssY6koVTb8tgsrYr2qLYYw4xXpHVMtkjxfHM
Fvs/zBIYD/LN0BhezMsExudK+fqXV8zOxLufljrM9FQjTx198cjsQW1PiCNHA7FiFgu8BpB1cEH8
2dpBr0zAG6N1ODHzLZ0EnXG7DUV+2wte54C0SRK0gDUjZHwnB6W0DDmbzckdEDE4mUJsGTQFwUjt
o6fXAl1o4t1YgiyZSgQd3GL7Sd14UUAv0p2372Ll21hPnUSPfx46N/o+JUNeoAtdno0o4OpoCG+v
rS3JS82AzhQqJVD9Wb12B8NImRze1uzroaJyRcCSgjglBNMsoFUAtvXlXbuhxSTjb4DQ7mn8qWRc
vj36EXdjgbFzEF1tDJ05jhOt5vuwukCQiMlwjplaW6uiJLxjID+r1vTY4s6hGL98Cwzd6+XCPEiT
3KcH6BxCMRwq6Y9CzV2C1lgyYwoAWs69nSW0LbCz4r+41Y3m4mHsJG1QhOA6XWqzWDX58ikAdxsi
qmWwZPkI5mcgF1bVqGXjUZjvnKSc3/M/ySHjMoEtaRGHU0a2VDGMViXRVCKMH1hHlNDWoQbgeVeW
XrkHYH+SrM22JMOz5yamoMqfWZtgwStXrxVvnrxx9br9B2TTEHHYoeNb7aq61t7MlnptBAIu7kK5
XCtZ7drKqn7K39rs55vTZ/TQSHLMlwfxrzuEybWYllZ42ubbsMEHLyaiaUVLOaqhyM2+Sq7Spw8M
635Kyw+cx0ACq1a7JwXDPO3RY11d5XD88ppiHNP1sLg5BCwUJ/twl/t8RaZNAzGl/LrXcV3aoD5Z
dogsL5YBpyIGfZV3NTS8wGqGB0TpzkqGpmgfN4NkRPSBaS6uWrYviodd6HDY0pvfols1atIHlZbJ
cBY8qbkakJT13aXulcLR/kKpLIh+HD1IkVb/12/LS+IS4NpvrhaYRWLrhkvAMfvlxfyfWUnPWDgn
/k1gYHk3H1YprQXwzYKyoYl73ui+FiIivgLJAeHYvaDYH1JMkZu81MwmYCSrRvaWMhh8ipL3q3mk
JjywPioBcLEZZONunKUA4mEhxojPq2R0w/k6/bP9lA9oi2mhSUFHoSgRU0kwcqdb6nvnkZW3ebsp
gkzUXIawgtHGNkRrQz9R4FVVDdSjWJGRika6YY/+0EORToRIUKev3+HIQ/3bc2klzaRGp4rxJBIn
8PQIGgCTHnKgeWaZBBBnyBnwmXBWMuFPRdLu3txFmeIENFFxENkD3L0KNgRzOHWxPO3i2YNRiH50
/5DOhpwsY45N/KjMsFOtzbXwyLadWY3DlthOwQmhRmlq7qW7OHjbngfhwhXgaMdDqmWbCpBNHl4p
gQvoKUwd/mvl+yWRQWJxOPi7V0usAkkxWuWCgjRAPjwobGAVfL9I98jX7XG0KnPf4pCKcJgPdj5W
T3evhW3S0xIx/i5OaqgTqbD1bnjjR3eMWPsJuv+IPAcEpx09Dw1y5mUVcbXZXJM5hW9RsUDlbQ1t
TS2IlcUKghRuQQWkmzXfJcictA1mTnsJ2lZCL2aWftSGna5RTFkTGTQ2GWtt0TsmY0sHdluhiuKN
lVFkQpizGfzHs6cACYCnEG9MpAwBAkqsEJpO6cWTQ0Z/M/henqXiSmVhDWtS/zh6wnf0hD2C6y4N
XRE+BGTJhFWnTb053qOyuPUV+pOy3tqETrOCwA8oSLkPeFOwnE/EBbg00Q8ajhyLTS+fWZkI6o0r
NuANpWJSiAp1ZRqoLPBwF+RhT4qoAoLnOua41ZjkHBr/gyIXTanNlEIVHVOsIjuUDQhQyrv3PuYn
3peWieMcPweg9hXH9rz6RSJoZqcUPNv9OmAEcexxq1FnnFzoX/+RRTuRuWftfba6WcT8PO0WJBbA
1vU5uwQlEmlo7PajjHsjp60igN6j5zki9m+UjJeMg9GEdfXDTB+J1DTNbGdzhVXW4mU+Iz3GZXgV
SZ3LTHJY6RR4CiZjnfV4T48kLysfmtLP4aYOQ52jgsbzDD9dn1cte+WQUsYgl3h8otp7H4EX+EM8
slEiuh5FU3wcdyAqWkC8xaf68JhcfPpnB3Xemu4Er84InhwlDDQU4t5h3xVbiGmLKOrsW5mB6o6G
DXT2BD+EolEyIdSaK6V8SZjGTcVoHFDPZBB0p2DGNa4N7hfKnb1CV/mQHPgBUuMR6vQH3ukdwa9U
pgGG91VGHHIf90WxEQnt4a2fFrS8Cq4odH/VPKsshT68sUh7R+802omAFxi2Uz0LGy/4zlUZsZ19
FfgrPleXXJRh09lPOVbfijENGmSG1HMN6J3YjzhtiOvGWhuzHppmKaSBQmd+wsmGPNPX/K77JPbt
x3b9NP35oZ1dKP2QeEu0jYQKP0WwFp1dvBX6yR2Lc1wfQgJOeFju2x1jEl6P7lXWVB+jDmlgKIk7
fZ9jqW7D9GamxaRm1Gau+v/Ej+VvhEPBVO9VhXd3uGmRPbdYARkc3JxvqGTL2tnFFQoKwF0rnHaB
ofqPuRQnZKCEBO4DAg5UAu59kn4jXnNxCcrktoEWT0x+pLCIghfmuyzR2o4ju2/5Wkw/cC7hccCl
G3tt6I37hKIWeDrTETzdQGnQcpMZbqnr34AvuUR/pt60gGhNltrNuZKYIKpfua/Pv8X/WIITcaBk
oqDF5+yfFhScJEKEU883kwi5IuHaODpznDZpE5bST6k9GnZXBLUO0+V8zm0tvUinEnkj295nEoDd
51R/LhSakObeCDPEdu8wNw/8/E0icTMNF47as8CadO0Fco7xH9NNyutYnGHrLtm3tjRGacyTAmGo
ovB8aG0dO5BLx3sMmZBf99UIq2vUdrupWoyowin+2JlL31vAhD/RuftqO40KfnfrNh+pX3nGNNeR
0Xx8iKf5BOCmSYmJCLRCP+bPYAsIxNh+L64q3ZN8gS+IZHwNKq7eKBnGOKKtcZWqfdLquq/XmhPs
nyhTClnpQLzDZmtf4xPLGebd+6l0rixc4P5wF66618nxiY/7c9GejN134eQra9fca7xy2RTOARyZ
nqjoLqruFeWi/M8x2myP82A2vNgLFJsbdFj/AanDhwqMSpTqR2gV0RRSGFHdvyaJVIjWoMLbzqDU
DGK6FIuSG+lIw7tMV2UOKbVYkx0Kk4XWy0lRJnJgbaxWUw07vMKw0iYqEBJtwoXrNB6NYVXu5FBP
B8/YLNKMyhvMzo9sur+WT2gBm6tqRxGj08CN82GgtsesLUaT8cTXb3xVJ1/C6gbiVOZq/pm6gjgn
b2F5lYu9yXvlshRHAs1YZhJS3BXdxxhsBGB7UnaNHSS6nQfmL3CbQBvYkZcsHgQ61dngzfNm986P
ywqApU2utjSox2Hh2koC39+RtM6rmSQDbh9dElcaHb6atALWLkWCblA2LBG3E7eUindBXD5uoHV9
0aoD9L0yVNJ3eq6hpflYyak0OtuGNv39OUICB4+XQVm0xPgHG523NAQuNpDv5od6HpotlyBdFeG3
leauh4Rm6agABtrqE3OoyTJ4MZvbANQGZBOGRe+VwdCDHwkKQGqwKfAeO1axV25O4O6ZezqpWjFf
lrOQ++6tHcpWKNZX/n2wxgX1nfETNzx9qKY2tJIYdb5/x6Iw2xN96dkrLIjf+koi66pyyQByoWpF
iAG2BjFxYpXL3cewb/B7or8WnEOf4PH3r/TSlcxpuHvAwS6u2qAJTaiHK0DvKytJ5CcdlDKUO7yg
Zw077vVvq/+/Vw8p8DS9A1LFnBICY/BLfe6WlS6aKdHCS/hPviBKBMOvMlE+AmJ5n3Y++0XZTa/h
FVtKsYy3Z6GXIEzI2WbiRzNL1hk4CVYE45A+Xl5qCNVL2Q4/b7ibrGY96HyvJoyaV7S0zUA/sMMl
xoXMZFTJLuqK54MUICblMTfyziAt84zpy0dWboSUQkDzcwf2pA+ycyL3o4OrbnyvnuCRZoMuAznW
Zei0kbGFqioaXbIKRL31gGLtv5mVHJfWfzaMq+6JFhMGkpUfrLvzuw8Rc0wdBJLcmMapgwNL/ZrC
v+5rqdoebTDd2PlPsdiOI28W/RCo/BAvvgnMIiPafMUueeh4Giy/Dl1065DhNJ5ZihWCIzMVioqA
tQZxdmyeVT3v2RO5Q3ICJ8Z3CTGAyO0hEph4a2MfzaXZ0MtoaOP1i4crxV5x8IHY2Mlv5LwZusDY
VCCHbexSV/aJGDtrLhSpQQAdX+n+DFj+ZA3DuOoT5QQdQLJRSp2iTMOBVkK+VItH6s9D6tLkDOR8
tVfixGCsQM/SbsDuUI3kSnV8DjsqlVMdQkCfg5kHUJKJMRkf77wmm+76Z3IPMjEaXQvU13+ciO5e
Q66MTtwc3aS6a7RsyKgPS8mGUd1vnwDFPjuDaXLFbylRtVlN5Ui1YrRkfXNsfqF6DnXqjr9fQGYB
JtVy4+jmpJ69JU0UzEwWnVdpS7s0NsDyVq+lhDsmdJAcQ6hEP3kJiHqRUkfCjmS6fCu9vjsFr6WL
nh+K2BHdFeRxW24E/Sus/ABVMBBH31nxS2YPfWI0QzildVKVC95hlS8gzl7XCj+doTnG0XwrKnFJ
HrXx9YsxMegA+5Rfkxg5mp8h9p+Dmc2DTBUOYIzgKytKFwH173NbjvsTnsjGddiG9M8VeSgZXQkc
NwYc2jxtO0t/AWbLdZK8TMZWsF5P1GhFTKbLiffMvL4khqnwhTrtsddjQsVY2DofeGB6oxGSIJ1f
kGh//W0BLydHJJatVBH/urufz7Owh/spmnJtcWxtejuCealxB7CJyuLtxJx2/UruooQu9gjrWWLV
h5oxl8O7UFmTageTgIofYe0VJsE05XQ0C4qH2FZoSOMeVP8OMoS6oBoWYQQaAL+QatYrupetnyLI
tkGUBRqkICcE9J4R48w9OpIPLm+jvASW6knoeXzGScfvchluideictJIgqvcXazsCwh905cjGglv
ujzHkoGFpaUJMgXJQuSO7tVclk3vf/Ryp9COjDZ4XMskeXZGNjKVfqBPzawPqyz+PcFrE6B50gxC
5NM1mORbDNy/rJMgxFwdpH99ZXi5qMcwd/t7EDNJM+Hv4SIWdKSwjxMfzc8Mik4NIlsi1K0p7MSU
bp90GyFwKen9YNpuAa3UlW4L/fJJF9SJZxMG+CDeWOde6sjsq3y7ntnQId8y0KuTEihlwVeiSzBY
q/hi+bShjc1FsAO4PZlmrDBPtFe9y1yisiZRMV35+a2cdWje7oJWbvNdf/KcO8ltwmKWHdZ5JzoU
T8O7U7fG5Q1f4m0L9IlRF2HaljnmJ53eICSQrLGvrq3QsWGZ+metaA73rdDIZ+dSc8pf3OOF/yzs
ro4p2VfOkMoauyTp4UvYWy+e20qPjdX8j+o/hmrG12MoJqmtXW+Vpb4DEXQhBtycVaooVl0AX8gC
K+u71vcNr2AhFWmd43YqNgZVHyG2/2wjiZ65Smqf5lslvYqUkxhp/9GjWGffqWLn3ot1UnIQOmSk
nxgtULvk7bfCoylawx1ZU1L0Cu0jED6DnJ6j7IxSd/frKaRCceoy0CnBfagJTlRRbRBmAZHsmZPg
2fRPiQGFSJY061vxcC5TKsZQLUNgCek1oEf+dT6UQtS9SARF2+AUWBYnIC7WzJ7xhU0/w1HrKgYH
5LhxB48WDf1TRoz95/iRk8Akgv4B89YSfGAi6X4eF1aOXEZXk8QG9dch2v076Cw9XxoOjKTG/WkX
IlHoQifu/RXSNpURyMVq919ClTTgNWLfG63BQBKd2l094Ovf8N6foql+TU8GCf2OInhM0MYdqtKz
0gBV+oKk8Nsw5s2rxPaanabmu6u7M6AksH0J3SsyZtOpmJ/MpJnzEPH1gO1iie0i+PXq/qJhp98g
9EInMfO6MTwe9AKyQIWQgS4bHCnaEZeywJtFMzdYqYVLlB1UZdfJKO59vxB0vM3YbOXDzUcZNCjo
ZilPqwEzwyiuhU9AKPnYmZRdwf4plt//ReBemaV7f1JAxhoqJYvo72qc52F9rqOTvZfgFlUNySqy
3b2KbZDSp/g1+vOgrStSdssam8bGpnkHna7oQXNZhWEHqMq2uF8Sl6uvVVD8+bzJBOlFmsbAEUVG
pJhpA8/VkFpy1ivdmAfKkFiqjGBEqj86Zu+SbyW465VjtU1dZEoI+Tik6cTXGMbLbwCWuvH1nyYv
vyzqvfVbeGAVkkHPbpQCRnxAjwl6tb96rtHSqGuKJ9A1eJr5P2LBrZw7MnWvVCRfFu3ckFa/cQ46
rLMpkE9k9vbWG7KmQzK+wQohAm6sEhn6AP3yHq4j4+MUiJLggThwdRsvBZ/eQBGbKyub6MPH6F6I
21pqV7kMJ1JswzJF7D+KRPQmRKSc+M2rIvg3VW6XeT62h1PCv5LJd2a7LjVbD4F7mD0TMj4WkcMb
NT9U9csHgGt1vMfLGp6DPqMSK3cMTHEEovJCMqZBoTY/44/aZzITGEXM1nNPoqa3qEcqft1EIHFX
51+Stnz7+nn63KMqQ9+dnJ2UpQ6UmyRUq3SPnMmV0yM2UphlkixQi2P8Kq3LOT9czA5EK1ypMUMG
/wxvVDMQ/rd4IKs7Iw4G9ZId280O+7Z35wqgd2dDyjTsml8+0WGuuKHh0miNqSnXRpX9s4/R8J2F
Y8YT8DK8teOqAOTJydiCxexar92fE+/lSu2RIUUmFewBRq4Wtifct83cF1pyzi4fJdKKbV7djOyL
S7oWy+rwlR1y+Ijwnu00tQF0dj3tbkxB3Y1bfLRcnJuh46hwZ2KdM0SotyP2VMU0A9Vzw8H+E9XS
ty+xOZSbDo6FdLsPc7v/y+g/yghg54je2gRkPN6PwY5Tum7QkE3Cu6RrT2lMZT3aFkvBgZWSQ1qf
BLtuNn4bXf4FaKhfsli3XD9Tad2qcNUu3jtf00fPLnksgTYf5fVc54SgK9NZhAPdK7X3fN6DStOY
V1jKZuIWcQ6Mp+MqB0ELm6CQj91M3qUjv4Cam2tOmyvyeT3qjaSlfqHKm9TEM4iU1A5osa83C+lw
2PyX2KiVCCItOJHYoQ6WFvmBq2R+igjhjutiyaLzb6st1h6N0An7E8jdXzyoZZ+VDqnJtj6sGJ4r
9K1nRUBUrUs68u3ENCH+f+lsCm+EBPnmUPwcnswxJzDuNeNd+fziaG25xyaEtXQvE2To+tBUCeKC
OVFbos0+xhRJIuPnP5xLZo37eTWHTKIlzYSRaMsLW/7S2Kwu/JM+nNIVT6FyjH7ObZlKfKzHzS4y
/UZsQrgLonui8qjCcDd0a8Y+gtBRFkIaum5VlBR/6JjiKKLxx0VHkHLHnM5NrBHxVHcEA8Ao/yGa
//5xYILGQj/GOk7co6ueZUdZgFynoYHcBRSV+e6vISwzcFpjvg5UgO8kYGd9wevVHTrVN1e+jjt9
raXj2+IeLyCcU5dKAVDR8WdwFEuRQYWlzq9aaa4wdteZRkmj83Kfm3JQ0LmyVqu6ro27P5Ira/5w
djU5xL9MZ5d84xJt274iHnSGdMMZklYmdXX5b/JMpqMwUUV5YCQ3UQLfIwLVIwAZDcWwZW3r1JTZ
GU+JSTZFtl+vYxSAzJoko1dQe3d0xzfUE13JadoLeFUF3fyOKcLb7E83GyZfSTpzWKMwJnHpwKEU
tBCYv39YE27eF17zH0I79kwrJod4emdoNPQd5qsm4BBvtKDv3rK0vSTCuTrns4xlgQVtZJ/F/O3L
qpm42YRaBKrpxtdqtRSQyb+Pjgi1i0oLsNxGlLatTHtDQ6vsRu30dcPl9NwwZKbnecgaGTlr/h/Q
CMJtRly5/MrU2wwnA88b3dAYjgSnWddDxHjx0+hN1prtHLqUIptMO95HvpmQboR9qPS8Ov32KPjv
CoV6WWU0Bs3pSEf7X4O6mmZbbZUTzHZ9wslo658AFYzIg6ha/7e0F7SIaUmW1UVU/49egCtf6NCd
eFcuhNPyTBVVg8oE00EleLqDt6rTv3PpYhRfpevUUjamXuIpvMR5m2taFAAaAbA30TortFOKyGPx
Ws4ndSPmu15mWj66mvPgoO+K13OUrjWqor6qiCrStK6F+IT0xdFXQtZSwvHdsb2pAvyoxAj+FKnS
bTaGElsia+IeUcj6ylGSybigyKv8oIIKqaekrwni7ttgF6J+2E7tkbwvJToFV09+7AdLO2++VBIS
C1Okv0ICDlkikm6qdb02Lzv2RPHAVfe2eTNg5xxzciR8wYRg4xwF504HeSQ1G5Io97nsiRrMNmVX
Nt9jx5iDxvHSgbwNnpsaEwmnpiZkvKdpEaNEjXVgWFoL2LqEjbmPQOTqb0XUfABzFGfFn56DAOj5
06VXXuCzCx/5ohQQZipWwGw8lbz6fM+NwmatnXgIRk2iHbjRN4I4iUIciCkDQjXBTfGlJDDg68ag
hMHNMfOfNqpu5kgp7iQJ8a6WgD+JXY5iYRgaDrYfdUoJ5R3nmhFIycVASW9hIznC1K86IWRchUtQ
cr/PBD8rmx0kMj82XaG+tOl5APkkISLvp9XPUFbEirpBQTpTL/hRdOnVp1+Lb8oMmm7EsqAeu5Qv
QkByJdEauVTqo8Z4NuD2SfW2lLZvt43btUfTG/V8k1ZC/mNSn7PeD/vR7osA8BAFuiIVBm/inAC1
tCMrfH0qG+6eQg8v6hYiBvr+8VLdnn4tH18wZ8f6JJcyW2tJxVcdQIzVnO05t6R9PjK47P1C2an0
MgUJ96lJK9iApTMSu+h6nsDVzFF2r0w6CE9jqZ/MlfShFlkFzq6CcHJr3LFwajTIuaT3sXZBZ1eS
iX8Satoh0uP5aC4IeZaSnMcp1BnmiPpMXNPxNyQbjTxbpUYJtcO8LRYvwxnbNaZYF5Jp/P6ti99x
RkrSnzTbXsHMWuoAJu+FY2h542scAfINHyv7sr3e8EbVOSloCzW4nJzngjouvoz4c6el3/5MFDCK
8pYSP5tEHDauahk0aURWnBFOIy0CLSCLPkfY2xhbx5vPa7tNteS+QrDeMCcbEFMMGLie+w/q2iDW
lmYbBHnJS6sUATKeD60TmBMaj6xOlZH0gq9S5j7Ti/M5P7VCyBJ/nZFzT2zN4Naoiro0YrPiWLi2
+VmYtmpwrnZH5ArSm7cv0rHiqjmd3FUkpdCwPqdqQJPsI4lt32i+7vtMK6IcECwe4X0Huy7ZXOeu
Nx58vTEJLOaFvfzj/s5XSh0RigenibGfTCl7vhBuGCMBDia1PQsgqCwzriEs4NyjjqappwiPzgPg
emIW4aVm/YxBPTkTOq+MkJmWCdOoMeZrUFLmVgaR1Z4WpCJ8nfwsd5UJ8oCdmXiYH/BMOB/TYMzo
yoMgRW2WufQ8M6FTV9L7XMxtvzcZcPQGFuzSkseMVM5iXPlTC1XGHQ2I+qOhgG5oxcJo6hLhwcYd
q9xOgOaXIc/7zpb8cFuyN+hA6agRH7YWtdvDIgxQRi1zANagjrfkln56mBC+PuqM5gP8XE/tSD3k
Ijo2iCEsCB7E2nbOMUa/UM+2NlfD6+V8Mk8gflL7o/4Hi6QyeohvRkifbPRukQE2u3H+BS3okuk5
Wnv0GBXXeW9Osut0INHEiAb6gJtJ6hype7Sff3j/RjYINc8Mvl0bKrmyf7YTdMqfyJNh7CGFlsV4
/UiwMcyfaNKCJfF39LYgw7AEf8AOI632NE5jy6pt7xu3N9x7/bkLpr62vdoP4P9aGePSyZfCAqCT
fcJB2sSFHTK77qhM9+CCblDFHQKDRFK6S1AKPHWtguWTImeWPRDQNncXSSQ8CWsYbZ8LQ6jvxCKc
5fzn9f0uaDvx/Xp6S6H2YP/w4R+2WZVI9drM+e+4r2PKE9T9RaVDUZs0WFuqy/A3FFA2qaQs9jex
DDYQD+4mzmoYx9WKa4UGMe1PnPS6oCEGDog+PwyOHDj7DmE05TKF47bPvlO0T5bZ2u3cm6rktSnS
GmY0CrSMgN2Rvr4F3yE5YzYVCW0ZhRrJXr2VoYa7BtfIgNc64ih3rDKZ23AH7tMyRaW3r2yUMoCu
PytFuXXDAVtF3Dbp/2jA+VOPvDfVWH5wO7hafKXIjhpC9r8Xzn8DSQii3kXgKoFhU8/ja0uex6xM
wPgHqlR//rGJ0al0WYDaOIQTDHbIrHv7Mu434FACinjUV9GdmWpRQSL8oxQ8U4rpf/o+GQyAil0p
a/CBytWov+GKkDLi5jiIM3jJI2iZvDHIATcpGOierIkGGmQzKvVUf5TGdh8k2s6LNwROMIuW2NZb
piulmT6Ll6A8zalKQeySp8MAQxuEJ3XUld6FY3NfwNetK9l7TYnmtnmwsE5AsZ94KSRVnz8mTkq+
Fceib7W1U2QHVjACdu11hejCecdgI5JVdQoI2VIvZ+2vlR95e5KbdtgfzZ3ZxaZewhb2xUW2vcSn
RuKpn9wVMvA8vZ6urzlzN+YSaQu+giCxnViojF/SmYcMD9E444mhYBFk27q4PA9o8jtkUsi/NZBk
rK1l1wB9igh539ijUoGkN4iCM3o7X0VWmGFfkHWX/tTz5CqTiEoiOkSDDl1Q4XeV/7qKOnHUOg2y
elFClAu7FapJW2eRjhdu7GO2GxQoVmAH4F6jQENAwB5/CrHN/0Fvx3Gms2aXXONwEJsi1uXsFJe4
oblw6QvH07VU+wut7BoTdqNwkm65L4EJ4Co1P1hjxrIwJfZTASvOUWOgFMpMwVVT8Ir2sO39tczy
TvCZj95w1rth2ltzhHFpd9FUnfyMwqAmm+akq2gzoAdE86p1qBnqYGshpIiUOdCpTZuoC/478Ujy
HoEUdXKheIalnB3Bs+L+P/6CxzPQY1ORI+0CAEZkxQuIhKWDA39+zaOqDj1IOPd8ODiWBlI521on
ELy5hH+kQvwBEQ+3GRdBaWIYbR24JsDrjgVNnckRN+aUNF2HrseLSWgHdtspM5hqMOHBd5N3QjyZ
TfRj5mukXWw/E2ICm6+cT+z0+/2EqmxNWQwj1BOLzmg9V6qCAjqaIU9hGkOJMSSTL/smaXlTGyaZ
d2qkDYQGuhV4+o63/oRP6+gHt/VpWmu0Rws+VKcjZ5Bgiqo+lb6+YNwUOMg1YZlUPtIANpRlgVLJ
gpjr3VtRtQ7fFUKAumOGiMAGvrxWAf2rts5xNIMtSihwOl3TKJes3N3tD/NVaB+1yIYqVKdqrjZ+
Z9/uGh9IupwXnnxTTvhGOmpbbEp7eeE0joLOa9WxAAbLsXmsSKPDWh4es87Gs3rhOCVBKkpz+v+o
7tssGTBtbCJSfN5ShO66zGTYSv7KR9lO4DOsAYdkPlv7plDSko0yldy+/IX1RCwuYTQpCuTYxeTT
g2323YGGZFchX3O6GEY6cqyS7oobl4Z+tCvpLmIRRK5+5xHSn2f5rda4FN8aW0dsqtDAT9l3BM2V
SpLsdO8nvrqzK7UYz1f2QJsmxBgbSpAwc/XqOoyMvK45vj6P96TpQshQAXdtGupKrm8PbWPXs20w
yHPokX4UxGyNWihfm8DFGdfS9MDh3eI9x3W59ecoIABF8tmEeBUiy5bo4mV91T3Cf4xOkNtJVWAe
8k7rOD7z+83izOsOogflWvPLS5LAfhsQmuqZc3TxS4+NAy+DA3kfuxmA49PmL3R2K/5rJ+L0URoC
Il94ExQnei3+apGLTYdXmeSoIQP8egu40EtTrUEv7CPoKQHR6ZDG3J7NpeszEFDv8l11QO7WdGFx
5zIXShFZtVhR+GcowReQ8yY9tCm+KqKtIqBRD4c1PNSgUe3xQh0ozzPWwfP5ACxQ8vY0PO/rkesT
L9JSMe0+9sWrelMbEC1PUIAPZlA+RaZZb6tN0ijXBDRPcHxIakjwcKtN/830Wexdqc6Fhqr6j9Bc
g87Uzulgff5jnwFtx8HZfg2+BrZFykR+5HKEwzc1bD3amE/ypAvjNN4EjNABEDzB5nOv7exVsUit
wttd3y2xS1uFXplcrWO6UB8BgO0z/N7DLB0/6pLFOACNuAf3RUWbRNMjwEKIsCaxtmrGlowFb0zn
KenwdCEZJTA+O0SWdULKtd9twu8q3RsM1ZZuTIqYiKKa9otbfVuQqOhZ9vjumad5JRxUBP4gjDjL
aBUA8Umx93DDqtoXc8fYPIFREL2hcI+suJSIS6fJe/Cku7tc5Ni3J7PZyvEDEKkWXmpG6e6M1aH8
CFQ6N0DVLXRujrdCUYdL3sR6QQwp1SChJeviQQZrnedH1XvIgRDx5lcrj7zb5cHeLDCcXsmp7CGp
4A6RBR3k4by120N38LdXVcD3qalEjUFXF3wv+32GnYN5q/23eG00i5xG+V6ray4kh6+kUNUaej3R
Ki9O2jaSl3yBK3l9GT+YfBn/MTK32sg3bSkBCFpnT+yVZTxR3QPoUFrZg9/9MmUso7ui1iIs/pmR
JzW8GRmcVU5C0B6k7/lAl2lc6BFG6SYNAzGEN5Tkj+xNhsVV6FCd0927TiII9Ea8SyjhxtJvbq3g
5AGqUjWyyGBi+nUH9bz9z1Iq07xxsMJXwQj3+F+2N7mm1FmyRKlIzni7fIrnf6cRsD/l8OqpzmpB
9SeS/jTIZU1ZIDjEGopQay17BrnmGR3408jYFvXO8wC6ewXnQuMRBcUoYhsTUHGxYkWzGxRBRkCI
ATkL8sQGldW3ze/Ec8O9LfM96kpDvFhsKcFnK0yhcM6Ax2xjH6+bPN6j2Qj2bxb+3BjiLf6C0ZKn
SiMc8EPf5SSnwlzNDo1S5ZLQkcYhMkLh5l7sayEtRWi6TE6blOzy+fsRX2CLJhHju9bTvmYRHLG9
RwCqy16mRZ1ySgk5fadRPOfzh52TFke4H+lq8P8PzqnkJt5TpbXee++VolJrdbjT5E7EIuCVPJ3K
sfKIcecQGDfwIKpOhDRvmz4dPvJ6IIWWocwEWNZ5qTlKyTGfhyvnwmUtRjA4C42B81j9A9t5VFeD
WFnc0eSi66mxzrfVU3uFa9t6vt5Pm/ifoCDIR1CnIP0HcmIJplJdYZMf8LIN28sOlOy6oHs/TLxg
X6C3V5mLDVq4o+XtDFhRiNiOAB7FtLvIjoaHBtvrZ7ThCMhtTUEvI2NTEKYOQxG5dzxjHVI4TWeJ
0OhObU6e54Zl5LTewF8nMXr7eOlWB/Hltb7XCUhxipTUsNtYI1WgGZUR2/tcEZEDPYMa4Ccrzg4S
SS9fBhtC2aTPFPgeEbKoX20N7tQX2nWZJZgxbI/LKoY/JPh/rFjaWBGYxhPl33uTIq3Cpv8Ecws/
bUaxqgTsap4FaPbDHwWTeiATTFw/FeN/N1s27rrV1CBbfBMbH3iPO12Z8pB9wB029AsEm8HAQiEc
qmo+dcvEYBtQRfgI6SmjAjVda5zmo1DWJsblalGaruP5A/7MffhYQMW4aT4pKwyZiacbNazXjDB3
nM8XAenbZ1Fg3yuOFZTIjbwAhO1rpp2JkYKn8McnpNRi1AxehVF4cOpIxeubzBEMklMVMB6+9mIh
EiPqWDADYXudP7QZfnOt/zmK0pnpNLX5BtnbT0ptGJOv5qEikTGhYeINIAvt+gxntAvC819zGFPN
VTLhztc+AeeaX4MoGUgwyNxVRfPhsnY/llyr4kMmT1zd0eBr1zmVnvmcI0wAD7Ne7Kt8XkVqFNQk
MdzEfPOzoL/LAR6SWGwKK97noAjG3dQirjj3mydpO268wvyDIizSgmIlBB7+hCArzKmElwtJRzjG
WfSwgtNANt+po80KM+fMGMj6netg5WuYSXjD2xiPRTs6V+vBVeaIycVcVwwvbDHHcWlgWpS3imNr
wrtwRXkYUOGRMAaWslCVR1dfwTXQXpQUzw+6XpcdwZix8rw+8L6j98wEiyPGkSC4CstJlIdo+An/
FTbip/hDR3RD6M8NTno3N855hJyMnrspgpmzOTn/Nwkswb1AsYj6X4ceJIp+kO/MJw1uFc5T4dNt
52aErk8CVXyyOPzYPbPyBe+y7AW8JFn6/FSPH3vO6fmr/QNXSpWPXR6KoGFjomhBZltoTt7EfHcw
thGLkYqin+r31NEtbl5gvq8EnE5vK4zb0ZmouFOxMkaYGuXYXEVNx6pC/2S9qzkBocJj+87Qssnk
gwPu1mUJT0eMQUioib27eZdHSmuNdmPJm8nrsFb/2Ug5fV0grdTm+riD+gleXWafM91L5CoHam7l
TJDLuace6Zi9s9ObCRW5jJ9omPIrXCI/tJ5CvA6R3YtHYaV1jGriKkaktzAoDpt3WIXdNJfcuiJb
wSrLl1FPZsZlNnF5Fwc00JAqAKf7n0qOFqFKLFLxT2IS2+FT3iQqIFsAvY6BBtsDsH5b6a9Bq1BZ
5UF/ir0B4b7LuX8P6i1xXSDAvBZxjvBbSTwppUVVfFU+QFhpUroVT8l2Ne9m4T4SV6AIzAMp6iLF
AHOBOR6L0o5cwfKnGBv6MtHwCNL8E85TnX7e5xwtUTp7m3thdVZhClHJT7mK7aXi5opwS21rmCb6
TT8y6cfU22ZYe6R9Q4U7ZK8bImc1SAxSe7DXvCX+dNey50dtpy7y++FslJXaked5EG3fJ6KQTMl5
Py6zY+wYI2bdPzE7IyzN+zu6qzbrxNz2+QyyX6wiKBrC9BpT0m24rYZif64/Si9ETNNscUPOQc0Y
RcQbd4SPaBOWy5/nqw7oDHvcVtmdTR2oNEuYFnMlBj4DtCCp6u+rDIpwSBRudvBfzGY/RVX61lR0
tFE0cb+ns1J0iNkjpU4kiTm9oU+BiSHTWFuQOTEuR+9zulx20xyj8J4Ie1oxWEQJjddp9A0ZoIjD
aIcKcb5+KSXMsIdKZwtHi0ADDF3yyU/1KojgtljDopgWfm+pqr1e1GE0u363mYCvUh9DBg4aSiql
8S3obspW/VWF+HZdZb1/aJeKw7l+6+xEUqc6egIEnSh028fMe7oZ7e/xE+XfYjKoLEZ9ll2MNW2F
pMeIMZU3nTsZ+BR6xrPkoELw0R5hVre1qcx/N4M2nEC/E4db8km/jv5Mz0ymuy5/BJgr/Axza5UX
dEswZ7oJNHQjUv+fBChpqu1xXHDWJiPL51sWxvKNBUmT0wyRGMGnPjPOt5e8d+rDd1QxZkBLv2+0
iBogY9Zf+JlVI6Rx/NAlOIGumlD/wqcy4J8T4LtFXSo8z3XlfnbplHRjfnUKztSbqABOaMw/peDN
oI1smzdcQQskvAn+5nbu1kzRwmH9RdqtT62ngXlJx4lpNFidT8+Uf8BhQbEggHIprzWIAXf4VsKD
JVmDvO4/1PD70TKq3Ovtb9f9l1Kvn1grngS6oh0qChIsPvOu0QM4CaKHOEqKK0nGiAJnMbnAd5J5
WCwczFFjlgTvTKDO2CWhD/bf2LM6N7ZdZkIM4CgIqv1Z5VuDIqnRQaXhpIR2TiMX9Twc8A87+6Yq
GRGqBHkFPFWnMyfDxFXBdCV9ARmlyd8xgYFiIXNF3vrBSErorhn2lLQCsldqOBp6h9Yy4S6n6DFQ
t5VvV+WcR1LsIyJiS/MD6GeoclEG+SjDAmzyPgw30D432fkogUCqryw82T0QzMY5jjtEcOowu1i7
2abANsowbI5lfWoXw7tFo0u0lGEO9dkybe4lx4pEE97fYJPAOb4Mv2UNRpv43sSfygIBqkkR959I
r33slcWUDEyp0Ro3Oqaac/NKlIXWs5S+cjqCZ5Inevn+4De65wNIg2WmeRd1cOrOtRM+sIyQwB6R
1uoDkSLcjPpZImCTLSYV5FmLekdMZRHxpg2Y5nVokVOwjwR3xtHz1+C89vdQDjiK7sXfOL7O2PRU
P0pF0vpcHfPcAXDwCO7yzSRcarfsBl+Y2IpU6LSqIlLewTA5i1I5BZ57jD/PJ3WqY9BDDjsRzbBM
+6kYJ1ilQOpY0izPmzLAv7swz1TIW7xsnT8FshIyqx0Wa6ACFWhhgqA8ohTXARCbfGWMkDuMOALg
YTar2NzfgPhw9XcAYw4dHinxU2fOegtbsNi15GTRCOQ7sGPyW8gTsYqXEX+5CI/9/HxFymzoRAV0
X9t1WuYeROljtHrzwd4OnBdxOG4M2ynsxnbEOETq7xgNBfOK3JhjBvpcyb/hU6nIdHX6F5UsVMB6
BYfOOQVQJ20Fshx2hurFYf6wvrfemEgXs+vvixSZarrAA0G+E9Ql0VDunsttWIrgB3y3GgDpSAol
X/SnEAijMSVsEWnf3L6ofVwKVz61mNBbF5WUuaROcNuBr1qxadzC7iFYSQBw0FejcvimVgDATi3j
ru+r4RsMhGyhQtUqqvR1skVojp7nZLPrVuj2FxNMY1QQuFaIgcrWpoW00Oege95LidL/By0Kz+Ds
GANiFYndSNxt4WKweC9aGoOKueemX8yjBv09Ta7ELBpUmccBPdp58o/uIwm8ruL32mf/67iaeSak
OC3zro0Mba1JWdMsl/JnrvIJItuAHnu8d+PJykFvCXEhVcWKrGm4f+UabBTPRWC4NV//o7DjI4yH
oWNQn2er+mKfDieJihN6Td6rCypDLnGC0dJgBMLTiVZ+0aNznnWCoJWWcSv65NjFV8M5tC1QK24x
8+b3i6WzbjeUNM22sSs6yjY/11nbw8/hhxytWZmcDvhLng1OHp0CYZjaphULF3/y3Ve+nPhM+tPw
UyJ5ppt+OmZyDj71tu7bK1S0xCaolAwLXP7uIbc8OAu6Js82Rso3/y2Ll8sqDYbK4sJ49Lyt6F8b
VDOWfikVFAUJvvdot6iZtCthSHX5CeUjx2IVvE59uoE8JC/gzYZEolXamLhb/9o/3FpM6uqRZKDq
jbWp+TB08y1yPGOaWhD2kehExN64/yQ0389Yjuxo/p2J3w20EvRx0ErO0uAYSfGkMz0q4xcM3Jej
hXvOes24zAs4iAHOSKRJLw1nT1qHrE323VQ/b/H3TNNVUTuQgmW3GVAbuyBp9Hx8ZYG/FvDoLj83
KQqNHot0tLMkQt5ME38DzVC24P7lzdOlTJauyac8T/QwECeqU8z4TWbTpM4MZkzKtzcT9kVean7F
uepOHCBi5ptDaiVsC67+Z6Odcxu0SrIeHn3FoekbdRYbCHZWlFwtJmKDAnAXe83G7Q1UTKODRo2x
jOiLwZAJY/t1GeRH6lk3agNWauGBBWHrmr5oBV5jrx/pmN2qh+7ygofS4xExeV+nrMd7qUr46+dU
AxksAduhi/D+UzWRuag8l9/wwC0PVBOmtCa+CJxSdr+d4oGdDJA0RfMbdCBDmofJtzTgBBsmNeLF
TFeAPQqVvxyEWCBvDkvQQ7o/oJA0PyqKicVMpCeGX6QrRWdMEuQfA1eePNh0nJ7Y00Jq0EuilHBE
JOmb98CIUPoWU4Ugg0aKucpF6M82oEb6JhDVqWj4UVz9GSnUtbrAIM/No9884chm9gPBBXmJOSQF
bnNToAQABPIdjgiepv3TVYjauQsXxIpDvpujDR75+nfgXSgIK/lzPK9zR4Liwy0huBl6B3xdx1gb
2B3ouWmJK4t9jiYkogMD1QDPAZ2fh57Y+y3pnENfF4Ys/u5nSrHhC50aiiFqxW4izHC/JIjbITHW
UWqtH0qvaj2fRFBPxKd7nmf1f0ocgPThhjU3zbEi+dk7ctYJaEADNP13NSGNb4zI8cj3DOiYBuQp
JyrOA+I/kdfXygdKZoR0cgItbhrjMQqkpnpj0k0dDH/IefcaiYUByV0gGnpw/26OXrWP9e2h7cx0
PqJULVGL3NOLJPNnE5PuzIsxnuxxdnTDk2rjmCaXY4AfrOH+6iO/6qXhrgdiBVyKIy4ZhKwveN/j
S808eL194yb0O5n6j0xbVxyJ17UwSzRbNN7BCnhVgxx7X8oyoIp2Fo4imADpAMiOkU5qHdMYkhrd
A4wQqspo6sOqz7vKMvyUjvB9Tr3a8GrXkDhK7ABUoXfIRmsscHIWAq65Sjv4tr08NPEEeL9/xsdQ
IRY+ChW/lD8Y2yOm1BOcF1gsF3ZpGC2w1c9e/woldoTNfRKRohUZ8IBoLSAyyNq1ZbNDO0CpweJD
CWHLE1X8VyKNG/wLJmKkWiv1JBX5mMMKmeX8yHsiisbrOek+TQJsqsM2fhZ6I6U6MXMTFeBZVDcg
Ttp7fJU2RGzWxkP7gKorBuDKwnzCza9FyVtDyGTS9WAE6GghBYCMHHN5aQ/kFUvauqE1ebJXJ8dF
2mMV2UP9URzO1rHxbZ4tp1zuCc8IeiVr+wQ5VlySiHmOpFq/4Ib2q+2xXRsIiG9Y7YZqInNphURU
di5bdhzkAaYcvXFt/FCuLd4396JJWB+6nNaLk/r3b3b9lZaT7IZ2LhHM0/LBiLUAGtoHcBIjwVr2
TKy0lErD7iFTfqCqg/A2g5Y0L6iAsackSwxsLHAgD75QsR58rGR3g85Zzt/kcpaOhxBqkaVQHIOF
cqdBq9TV2xTC9bUOmrkpE+saeCciJRDHWJTpkB6g5f8iqBTTT17cZ/pYbfMGDVSXmk19wZNyewDO
diQDpDjJHa7HOZP8iWLaitgOhhnAHN9JJ0bD7uvuqDXsHbJ9vEVH9pdI/w/oQuVOIadhQWDSfG9y
aVYwoipg1H4TZF5y70mcc28kri7KkYagKykVDAZP4gUiLn/YAHvzWUhjt/VCgM3YJ/3nr08+KDjD
KUkd+WZIYxLPRR91SnDBBYMMyQOXP7B08tQbxZbh6uLJC7eumfuyCHgoe/hUP2Ej1fjdwRfbPITC
hLFl0CsdAnx4KSOyabdLrM/QU4LaXswdvPqMYHB5nzcG7xYF1PfPptuN09IC2Tgjer6Op5H1I8iZ
sNhBGKFM6omSdJb0PUObsC903R/qmo3mv4833E9l60pefOa1C2M1O31Syl7iIaIAqJkZR7VADuDa
ljTZIOapO8rAUM5zDIDAVRM39kBLz7l1ZTbc04IZ724yNkiFlGTa13U9+WTgjlqgpKHP1iC51RaH
opfMa0PWQSyH1x/NeEvbbsRjXGFzQSghSZPZx6aYn/I69/KWlSoiDAKv9M8tlJFnvK3Y8/Je+TKO
MJeIk1CTcjmyuRQyIchbLPeFgvgJeHOtKSpZkJyVwDPJ0Ryw7aFqMSO/sjvEi2J2LAY16AYU/DKy
ENK5JcLMPjlQu+Ysa4hKzhVX3gIDmGDF/Xe7D8j6VVUc9tTHUeN9sN4S4Ej4LXGvZWEUCAjFWHyM
Ndct/HTZ2Y01sXd4vnmfFd3OnIbfanCJV/kejTry/TqFlYVAooa/zIHZrNBI5RI8jeFMZRD67QKt
RYwU5vfUyK+2+xqztB2Fj1ZwsN/kIkQWzxP45qi5WrdoR/QOtQ6n7QhAjLX6rnAzbk9qr88g37fk
7bHbPvRlU0yrqaO2/3kp9qi0Zx19fdnpa/2JZf0NlOkMNf5hdj+eBqHK81zc9y5JMljn54J8NwhK
U91g/T1np+5TgFxYw9bmIcbltyAhodYQt5oqkSj1LmCwAq8wZN4HU5tNA9nyreCtTZ0IRa1PU+GP
YbbEWiJlJrHY3dezSEqYu8rwkL5OQx3Ziqtg86j21GFfL77e3Qct1FdZ2rVv7XrLWOkCXi+1eA9h
rDwxi2xaua2ZRw/1wfMhYfu3tw+EjjNR3RNfCkSlFAwzcNlQa+oeikt1K6CwUevN9K15mgryVrqc
qk9z0PGAYD78q7zOdkVpxAUy7EERNA2+LxlMswl+c5UlGI1dqyUtrAcgGOgQJphU3M9ZfKzBZTUf
7bIusi9AHDIJdDabn/ePU8JpYaDruHSXwGYrFdvpxxGg3fX8T3O4EJyG1SUs/lItuZC9+sGhQo7V
J9ZO4IhcSUSojMd4r0VfWzIJ5ZlUm3EPToxkYjflaZfRBbKNO361kGgtHvRV6Oog+OwmCqLbyzEl
zG7Oq80D7wKZorACqXOXX/+FIAWhVshzXBkjHrSjD01X0HXDtg1KKO+CPhFBpiDzrOyILGBth5Dg
cEZuPHbwYPzPJGG3xh6AOXMDuJW2TvIEe2OnuF/1NWPMu6xe0a2YK0gF0L9Hyl1Q164+pW4G12u7
hxjngZofgRqh72mY0dXmbEB7EB3zvzKgu/eE4I1bCN8A2HbmkOmeCW8O3HXwUkaLsps1tqGyq5hu
OvQm/Ar/xcMxpie0OHMxG+4JuMj9Dk2lbr/29E3+B6IFcbfUahdYpaSZLDFKnZ2OsZYtFlRu6Saj
O6MtxNF8GrpUURm19tlIf0HKC3j18ispbjuIDUZoD1aPySMGS9vV7m7uTS9sZfOx2e65nTU0waXi
hOhPjf9IYo+I3KvtBagLlcfoUNFP7L3TmkAMmI9bepCFuj3irgUZKEsjthER9m2F4qD4jPqb9gAo
MaC/viexf41iMP0kzySZuXdYgPyx53paCN7Xfy0GAkA8fgMuGFurSfA8sL+95cOLfXjazzQ5SgAO
TyuGnR3Lx5qvJZ+vSLoTY0V7xR4Be2cwJBVOGDeVOdEzup8sJ2dT6fNpf75g9BNFiTLzG49Ox9XB
k5ZRJ/SVSA0CqRjqafEYyZaCA3u28WCg7LBcBnS+EZXkzG7mpFRoIMR0JHMWfaK/02kRM+wRxFET
Om+z6cXEZYcAr6anU4GZokuBA7jIY1zOadIOBx4Umv/b05JsUlzU1rWVYLY6rqvNX8+mPgnDv8KP
DdCy0XWZQNPQZS2tfR+1sRGgf3eovlIte8j2q369PcOkLEAgVEs3u9yrj0HSnyUH0bAkKqH7gF0q
eEl2pYtZ73eQRUjDEbfZBRuZFjYwEpDna1DHxisQXJHEnU7RyuiWRTwfYeJu7bJ20FQiyET3CwZC
M/VzsHIK32a0h5Jd3ktzbQjnA1yeEpt3apQibV8BNq8BdcG7oXN3ItpfAapYCR+nLqsq+oRfMpw+
tzNYwr4yM29TPJKEAMUvjrucAfQN8T4J3VJ/W09H7db8ylgYb4sOAdI3y6egCCK5UuePpD+fv5mO
o9HGmO37tkxreAL1n3p0eGCkm81be0XHaIO1qOv5vq3ThQwGAbxFDVQXzi+g238X0NTtJ8iXg78W
rg9TdVhBuAvgzdqxY7RMYJzeRK+mdsHwnYU4t0W6VraJMFwWpRH2w5yMraguACrOdYYPHTQEco8N
4xANSDV/PBVDbLlbARJHIUmsZCllHE7UIK/kaXr1mEhyl1KN5tBSGJBkCF0Z3/rr44+rH1ZKyJG9
ZoetkC9HesAs1QsDrt9DaJ5ggmyC0v95YnS58BxybUWDMGUeQ9iSJi3+hIGLWKES1Ex0Hc9iOGfx
xl8Z2i33JXHuJ5hjheE6RjL8BtEnFG+VIe+Aa1iVoxt/wHg8dbVlkroxIsVVrdoZ2YCDLtX9i50w
26FFXl2XeqHm2QIK95rZp/R+0FLB5KHwvhFUF5RB0TmgQZ7zA/pqfxLeHtIMayZrBOxgdmDxTwHl
obND9Dg2GEUXloF4hC14M2GNKrJ+ZEqoMRmUIXGWN70DwqHr3l05ase0psR0Qf7RhjOysEoyZnJa
DRRuRUeQDA0XSN71fCuQ6hLshF91mFaV890mMzGMXd9SSQJxxnd5sm6yOreOlafASbJKOFjcBFH/
eY64jhFKWREF/UwqAd5ORxKiUMGCz7MxuR7rmXzb/nlMkpYzlARcz4B3OYqZiL3MXJiweqbtOYZV
y6RDhTJ9fi35YggDa+x8G6YddKb9QjzACFtY4PuHnEvzDzbMvttDm5QSwgtbSC6tyMmGN8ovSO/o
3yyYI66/nFJmMQhs1O9b3HG02a4pgGeJ08s0dsOrs+R20CmKcjvhDf/mdpHHfvsYraIMx9OsN46A
G6YoVnb+dvBTLcie09PDvGlMljCQrSyZLYFJOJsqG89NEveTw6G9k6Cj8mG5Gyd1KBMPvzkFupdx
ObrxVVCXYhsLsFLqb3i4Uf9llzikI+SU1RSgnJDt07GAvIZklsi8NkQtwuwqW1+PYSdfPCZrp/JK
LgNvUoR3Gv99htxb+/VfQ8LfvX9s3ZGLzPFj6LYWdng5uc9tsg/bJLWBzGQE4s73WxWmucYmZwSv
octyIcPZspA5HjPsGYZukiTsaLamGDq+YOVHPbJrbD1xwLeTxD90kqmBjJtApPy3pAzmA3CO/KuZ
B74QYHsARz/xrnDaZIaFXZDYNlu8i+B9Hhs2qVxsvcAj8i407xaKWzJ1HCX2YR/yDiS11gEjrom/
2q2JVELzJDSHJ2qlmiQlQ3vexHjxDYr8s/A7rGRpjqIRWeE0f3hRmMXHQ1M09uWOhiaimXRQ9mWm
tFPzcH4DHVF4kBWwNm7fxDDgnSt5I0+xX6AZwGf73XjN6HaK5O2da5s3++fViHelq30hgJusGWPc
CfAqQbLHdIpgCBnKQyfwl2O+v5kdF7wQZ/TQDVCL0jcirZULlSuCcqOVAGaCa132GdTM/eP/Puty
AbWYJJ3jEfVYRnn1wvhOl+WQMOwD7ID5XY9RB8fJAQNvYTJXvjBV3460j9BQS6GUwQCTzrPtFJuR
U1IilPEmpMg2fIEkqKoV9J23AGSXkzvUmObQi9Hu2EoTp+EA1szIlv7s04ZgsSxz0aoWVRHdo1/H
eYrMUCRFGkbC8S59SAlJVAMTtJmfY/ENlMZvKt8dqH/MNTwVle2mOnzquMGpbDZ/4uTNBEfADrVJ
46FCUnoYnAAtx8hqTHWNLYfVXf7FqLbqBB+tPH+wqNTOY6qhcllr5gtbSEhQYoVWMhTW4UC+ALyL
VvX/+/Fb2Fc2qqBHnbAD/q8sjiV9dB1CJnuZf6ya1iPXPBSWcK9Cal84/6srwrrIDk6WUCc1FDHI
nZAOM9a33Mwh8iy9fWqcrTRWQGy4zkNDSCC6r1BMoD6UNNUio723l/TJkcCEPBnZPdGHYc3KWF1M
kBs4HGN6K/Sik9Dfaf/AlKhEPoOMxZdS9Vhel8504HTggl29fZwbVfCBZdQuNiSQHNnt8xV0Vlou
9L/TILRWgm0GnNX3n0Nt7XYGWVam55Dtj/HbidrGd/HMJX+U+/oZgoZINhHRr6ZBovE1giRJ7OLd
so2tK5rlOPhAAX8fYMiUdBivJZ6dY/z4XIwgfttx+MTLl0AFL8DpplGbnvHvwFQDpnd5IoosyLrI
rsElEpYUyV5tH+38KXoTFKCdP5zMGPfzxo2RZs1lJmccagHSIARkiODEimx4tTfIrBRwWmgKWroa
Vc43nuHR+M4TCcWx7KGpdhnzxsShkwdHXlmrvgtUm56XezT+OjXpYbS2ROPjYe3mryrE7IupAKYk
5aZDBL8u4Ne0Gg5bcZJ9jf4M5JM/0rJQWUHDRB857nvGPKJL8w+mUlRXU/LfY23Z2isBvieB4jdN
/GCwjLj6eV/pOdto1XgUuv2khAWyStUaPaf2kS0lzs4Eurq/AGAeevRJVq6sRy2X5FVUVSBjqgIb
goo5vouJInBuRJS7OIT8wbo4RcYlv3sVb2t/iZOrnLHkomvaZ8lcrvjx/enZxdPbBiYnnmZ5cjoZ
/FWBdLnfx/4qjnhICxBCpdk/T4LrK3BYlqUsukNr7bqmOg+sYMKreLcADRoSlamyRUTV8wS6xHOY
qcei550oIOsubq7erCx1adRYYafugCYiBtz8IrmhO1Rz38wcuOdlN0fFiDi1o+34DZeD4blyrtLH
nqs8vzlkIhfVsLugJyTR2HnpX4zRddvVzSJHWRWAwZP3V6LNqHi1jmge9m6r/pq80FrXeBwO0Z61
u0q0Mj1svMZhMB2UEiJxNUMj8wgrJ5HCdXvXBTt1tc6YVXTbcN4bk+GVMBonHSuWe0tYTKUGyTK3
xNxdtg5k4hCxqVGoPiOwzQ6f8nihIDODdCbu5L7/Dff8Irop3tKgx9wzpCQDv9BEsHCiyTulRHUW
O/woj4gyyty324nkQDJn2i9AhQP2F0hMcwMIbGKEdGcUNIBD4mJSn7RCw2HJKZ1oFfgymDlBiJ4e
xVjfZ4K0Go2cyJv9wiOFhIWuYkaLOOm+bsm0JDEcBnD1FK0+Lw6VfOgmraCGj1u+JzW71YkI+VW/
oIoRyj5eDUxTPaTVfdGIlm+KhzmGlWVYAzHWQ3ByVVjryxkxxJ/5IuEF0u2gTEjzYPOq0ybVZ+4V
q+BC0I24gBHO8MkyZmXLWEhLCqgiNfP5vRFRYiVaYUzer2dzLcb1i6ooz503T/xTKfmFCWU/J34A
1FiJ14QkZqjvZWmUqCE80od672ZHbjjb/V8yz0ErIJ/PQZypcLK2zZdDlF/wVebYxe0DDwFHB2Jn
mUmWG/Y1Hl5LeCtTyZrIXmbEuJHBGwDOLqVoxWhRiY10q/XeMorrV4o9cZwXCdAYBI74QCYgErBH
EOXhDfa2Udu/SDAkjQHjJRaxpKvSXZZ7YJpanya6IOrhDoZI4G4xlEuEoaKoNULCBrkcMeFu5Exn
5fL+IJB4w3Vlt7mnnJb9iI59H/OBGITszzDI+7KWyMVnBDOb3yYSHkOZjCywH3r+jwQabaOwl7zl
EnTOxM8hjLTXm9f5x41fma6yy6XuyzSyzIaDf7A2GyXTA0YKbRgEAwO9WRwlW6PpEcbDOHgFU+n1
WvLqsf0uRqrA6BSZYvK+fK3++R+5ckWp1ix3Vdyt+QR+f2uPAfj9NHkrPwLWGIQkSWQq9ZgJqL1S
kGAXCHJCaPHC5LXK+CBdMNkKUIEh8oworzcU+Tn7R3Xwy9v9wwgYOF0ZyiNJO20kIX27ZkyEpjUi
Cpoxan55WFa1WntNfK+JizMunRSE80FWOphtM0uKcjnAUp8TYSex+CS9rRC1MT6y8fN9zm0jF5qa
yAq6QSMWJd/did6mQbmNGE7zqv1UXCU8dyGzYr5bFmlEiTMIVVgigLgxyPmemFth3YDJOxdTXACF
8wx8X7XMRA7zh0oB565dN3AaodnyymSqIRKBZL4ny1A3MTKsk/t7orQJne0n6Y8HXxtdH9vaW/nn
Vd8H9zcvbmNUOWX0FnTB9xGsRUYkNdXri8IcUM7DphYT0xgswV9VbAaSNu+sxfiiUv0zaStx4f+D
E1Mfki8KQrfxsoVCvEKcLzOSqPHekLHzXZKU3sez1rC6yDGNyzgUFnAo/3p60nc6T8wsPlZDVIoe
exp7PJpL6u0emh+rkHpiR1Zqdtx6/Ez6yWQiiE2yzQiBNcZHquiXkFVPOkWzR2doeVjM4WSPCafi
ZD6W6ptJopm5xvOgR5tB8DFni2vnXl2urKwHBb2l8063f92Rn4geIL+AsvUT5MGSkXSxBe74+6hc
q4kjPQ2HAxZQF1N6xEpVPLHbRaIBqBRlFHJ+Ez2myaoXAaN4pWWlAhbWGK+jYu6vSiKfLuqWut6P
mB7nhPDBpBJQIcSqZ2bRgL9xVWb3jboaDGrxvwHp5kXatTLF0MLVhrN54N84xYo0eaJF0+c9BujZ
xuvcATYol3s/IHbrnNLBmHYc7oDrkPUpTjBsRXy9mxn80idHDNgFHdcBxfjhoEGt2mp2JlaSpAs2
WbYRaN/q4B+U3CKAkS+rV83xan0RpFLNvt6G8ukMGEm7T+Nmz7RHK/snFSfWbsn0U+pEs3arD8ad
6YKbiNh0749Q3OE6yLex2aOQaVMM1DZ/rUc/cyKlOYSNxlX3NM7aoJLu9pmBs9gv7mMb+muUQcMm
zw7NuUGsbuollW+W8o14ZFhizHb5a6BL81g4acMX5XzJ/CFzHsOnceb4+uB9U+73p3KMwlvyt28P
YWryUuYxIdW2/Y9ydVw/seh6Dcp1p7nh7seJ8+gxJHQ9jiwfuoesJM+14QHz+C6m+OHV4SJZSUOU
dd1P4Pl5RWebOGraTjb+DKRG9sgre3DjC9gUIL14TPbKJDnvLdZye8aXJwqvfIXsZaZHz/K+/lak
YjpSFkS+AaR8g8PlnMOskyTalzPFIV+uYoDZapPFpZuLa9XkFZVJy27fi05rAnbKo1RjYRKXvGnu
XMKOpEJwS6yqGKxyFx6bfwUrZu0gzYhQNKhI/Pv4rvLyPkHY3mK0HBwuh4c6K7zSHgU5v+j6TsEU
CyqdardIiwsC7KPGj6j2t5b7FODAHpxEd3f1PoN5l1g9wyEgMwM1SWfPyXnNhSffi5thYHi5JlJY
7ulE3M2n8TBXv5StEkyZHbxyqs+FTcN86UwWMBN9zmJnY1npY8N2t/HwKFCKed0HruFGpxNdH0Ja
ojhtqAoUJS9ix9P2VkO0otF2lYCeehslT+yfMh6qnDY9OS0zqS/gxyqr3/5lTbCZR6pB8Dx4LguQ
GPi6Wyi7gwnbodmNlkR06DCRab7DasHLzr4OW4OxjabseD1Rc2VAVsEuL+Oj4Nj4pAoCKY0flnJy
9qdt9kFJ6lQ5PLZc1cmlKBH2VApAMfJAGWR1u/8CN/kA9qt3QFKHKKG/I9JLQz1gwBHqYRxT56G5
hzTSueTXwe/UiJiEqguU4SfKDrdckyYFU8aYKyKPmHIQO6DgK9q0WbHTBRmSqXtlw8HqplPu2idn
g+HLeBvmeRHPSNIvV8JGqXwPRNZo/fJhH9tiG4EfvZE4FB5dLxqW/0nGY+TPv42EcrT2K6Xvaj+C
VVljnnzP3WMPkLwCQTGYed/6+RB4QwD8uDuRwHmA1pv6CJAYx5X0CdSKhraY5m1C8C/0uwJDVV0Q
SAb87LQ0FdxTnnnW/Ml6D2NcrnIWZ6ZoxppIADCU+yXFz3aRmEnhAkpjmwuplHsbq/iggfzRldIm
W/5lEU4T/OIWtAiPFDKjj7OekUuyy9C6ShIaqjEmCRT0FbDYKehASjwUFtG2zJcxFTHMEnf/8I9s
1zpKsgDtvPBkxJYwPqpLztGvL4LLLSJFUpeh/1T6H/vDWysXCtctC46oi+jiCtQnwwCNJLyAgrj6
Ham6A3OdbSpvC9PQJnM5I55Bsg1cqYaWXXOWzmpdu0jGzMeP/YDRE99Hu5Fr2f+9RHlqeSoA4CvL
WT+I6d3lrXdqeyxhx+PYg7xGP8dVwXaypezJFU6Q2xGbtjyI5hwkcadoxXTwN186G+mlQwoMW0uq
NLe6k9xnjisfoajzoQ5d+kt1rJWq5EGIHRGB8y9wr8nUzQ0WUKfms91Gio93xnefqP5kelA8L81k
CO2RP1Pj12pnwD5fS8ZyfxbM/4vkLAJhzkG/sqmoeh7IecZbqQrgGpaqHr6/PaxRGyKrbdDcWji+
nbpn50hQwSelnFlUko10mrGoNDmjcGcPw07VLZCG0A89aXiWkrA99XI5qp5IgTVDts4Zl5z1eDIn
0UOgU94oXozrVmf8RvRytP214BAisypEgROgI0Yu5DzFYlAT4WeTfsEncVm01UuL0ziue4rKkqkA
/r3LWbBqc8pXetmYboPxIR6qIRG2JWHyDmpxSoAXLiCuSu/Iq5OVut+rPsWSn2BPd3JIjTQ550B3
IFik8MGZKrTJ2XJJhVE7MLoOFGnA/5CRso3GLMmXO42ykVzUlGDT/UiEDMBkFUTnAY9Vc+uadmnq
LWFt9rRb3faEy9OqsfNqUVVYtTlyqIE2G1qOlyHmXdBHLJAb/JHop5plD0oVJ11TdsetFDpvccjN
60Je78zx7vxNa5U6EanM8sqx4pzXY54AqjDbT4WUL+jlH8FwJbDFx44zOTWZ4PBsnopA1RKKDXlG
/1bJFW8d+XSFfR8h6yzxveZ3JZqVDtz9TC8mYgoR3NUJ+OtSu4vfo/IxEWz5T8ccIM6X1k9txhFM
+AUAnSBZh7Z2mfRExx18ZmTho9OohNb3kyGomibKXQAZAzau3RKYpH2qWEQwKsyR9sAMY5geKrcF
gEUQqL/qIqjcwcK6xPD6A2r9aAtvJwXbdQXQ+isCLK93E8E9hvtqOFaa7BX0ScAf1AdIzXrwwN35
S7fAxsGJ2Qu+PBZfruhdKxCvw9LTntfH7KUMaPAzZKW9arJh08ITy/zLYK0qdFy0LUtFVrqPxkQd
iRHL/3+7kmJxLDH1tDmiLraaxGZa4CJ9F6NNWrwa5RNXWWe1ku6UNau8uWibbx1AVxJDk1gJzeo4
tDRjnGWle8ML8zab5Gp5xd6A/MmFDqusnpJlXLSmsS/ygEXkX0CoA8VpkedWKeahWjcKYeEIIjOl
Od+nP6vaT5kYz7IaIvor77r3qE3ZDfv50pVK4DfKNSVOZUWkt1RGXv9f7+ohsiwYkPsjaUT0gwtD
2uxOIaOg9rP9cEE+q5oefObf76ADYNWwgWz/aDKrpCmrpbHzS4SRwtWjKv3BSjjkqD8J/nIKi9Lw
YNtlTJQpxjMVKLTMzHMGAwPWKGls1E3k9QLy7MyXGVqDi+gzISA5YmA6IlAj7+EmulyGOtRChxgZ
BDan6A+6CRFYed7Iw7Yu/71iSY6CwfIQ3YcnLmDtDiMrSlW1cylcsPl/VydDigZ2upuoEafuGjah
8p3+hDXs2/pvyTl23vwzx+XblftsqgCaPs5z97xDgKmzzIA3Nt4FQi7IXO7Z+preKNiQHPs3hmHy
tzFYfRdK9Xzhia7P+SmgFBccwZ9XAt9cgbjC7ygxSEm8DbkZhFQkZtqOyRy2I58efuwu+xRITWmV
LpNe13G23M8KTyfDQJbdvhSe8ELrU2+bM79ZUoYhSlWm0bVKgnK16+I3N5uQZpVZ5N5gUTIz7lMY
3/CXmEzn2oVDOVoxPsazFGoABcC76AjmOVAdV3267ZSeE8bj39iIUe9lT0I6PJetUnE/1+1xjm8y
y2EFLHACFabqiXQ1MQVUtfxyVVs1rPRSY0/SGF05xCr613I2Cf564bJnbSJYqZkBTl4yUhTI9aH8
ZPRgpMFGL9WGXPxtSuBOEX4Ts6EXDr4CXg6vhvABhHcHQ5Yw5xq0Ggo+3UwKhRvlbbNL/StaSQfx
bci+OTcls20mMJD9GeUG4H7bqAEWT+t8ywXqGDK/EoLuEndtqQ6xPCKsns4E2oK4mIhMntbAp1tF
vi39WuImzzCnIjqVQ3+5yN95D86nBgu9MCy4ASZoJCB0FXyOiK0NBJZXyODu9ho0VQooXqIJAgHV
jRvn0GkT5tLrQHkVrwwLzCtZMARjP5HyZOUu3aWzYpiEty1nCcpIKpYLiHtmCNSCxP0B2Or+RSUG
vYqudrLz6DuHyhg96EkJWmtDqhL36Zfvtdij2ZnyzyV0I+JPqt4TnUhGUUgCpnPCX58E3Ghe+uoh
ClAlRbrhpZyp72h/axsOqcmIijohVpfzeiVsBiLoMd+BhTmHZqGTCr2dpQyHFGj/fdPw0V6H4PuF
TysJN1rgKE4iNYM9RRafrhhopL5YBO8s/wNUA7yuneFXmhfyBZIMQcPcOaSUxgNYxkJCqilCHYJ5
AXM6Opz1REFdmYcXV1OBXie17tk3KQLQqma6q+VPksV65m8WdK7aSK0avjZaF0Qv3q/1ryyHh60V
BUUQfnws+cCosRSutQKTSVHnHYv6PLgOHdutvp/A9B29ocbfnf+PD9OIsh6lBbICYt6278UvNcC6
KwQYgolC7S9jaglvvjLYLeAXTFm0Ofj8zq9AIGPTvYeGOhkgNZsixbw9X+ePp1Sd0jnGN4XKzF0J
VFsOa2duAp2WZeeeOhZ1sTxAwuWJ0Ul3KwLGt89C39aRPvqChLEBejYqY0eJ6FSFIh0DdEyNfCuy
9eIR6UdXu7ZTrXd+R2Rw1gSLw3ZNZeyuTkpp6MIktKXN36+ULy6HEBfKE8p+KjUZiELn26aNjqxS
fYeEMjZZZUj3Qs4lDJ/Phry07I6uy8QTKiPuy4JffNoPvXsoMUpT2DxCLgeAKvtPz47hKLuMzSU7
KrlCC7Dn1q1c4KcNpi95ZK0Xf0/2dP/y+aNx9wnK7TyfIAuAl0JupNpo1cAfhvFYIUPtR0a6zxMp
aqUStsXxw2hK0EXfOi1QkOL94azJQaJgLvargR0ns6ebTCV7d2RZiM8tX1rSDe3XAT45WvZwGeiC
4pk6YALdC21j1/e1AoxgmzufC6fEsbroic0gs8351BpBr86EG6NNmJq+Jvuwd1OsPwoT/Am4oZIW
2d/pvajg/2g7wKebWzsTmfGGT0q+89hK7n2PfyOus0d0aAINibC6ZFvo/J+uj9TAPPN7W5AAkyM4
XTlWJnhj4TACSgCk16FeB1pPZwUw5uBI6kKJNgrvBg4rtaTcCuGHrvjejRMlzt+egRm+t5ny7y8u
LDRNUP7ixDAaxFfzVhCCXubZagr3bNSXtkUkHTLKgBCZfSf8ppfxgghezeqG+5WVleAwvBlYEKdS
8eT6vJnGcClQUd+ThnP04DWar1lZJHRkFRKFhutvAVpy5Pa3lEPKczRD/UsJpkmGh5tdnaLFQvKZ
PDB55WbSY3PWWq48rjEvlyHFf1i8a60y7vGy3uAeb9tjd5vIofPcOYsB9KN0RPfj07kd/HEQOWM7
Dg+DFicfIwhQp/oqu1v+5b8qmz4JNrfBDHLAFqgVMPS7LXY88QY6OLv6HojHKf0mIqaZkJoeunUu
zBvfIx0nEsYwipPt1zdE3pREsIYyjef8L3dyNyv3MOqfSvl9EC/7veAsh9dbk4qT/hyaXADL1eq9
oa+ftUMMdeU6Hdet+npjscQyGYaj67MwygBNWge7tcWqpP/cFDfUn4HYgLFAum0/2lvcCELTavUz
ocAGFycsilFM6gV9U1kaXbpguaHtAUe5ujohl0Xl9w8/c/b0ktdSwMUV4KxLmtkA/2Um1APbRfoB
k5oAbGT3wfI5FfIiu5ZfWgl1rnWJzwDnCwTidUdzUIlGN8BruM0Bb8w+qZZoUiw/P1Gkzi6QtJ+l
BhgdgFc1fUyu9Lz54w9j8RO05WU3u/oFfOEN1i/DuYEGMcXnMnXwyTA6VG0PbJ8RwP2YXgW7NArM
K/qetQMBoQPSzamyXlSlwPbV5JYSoIbsXzNwsA8/YuiRbzTvNSE5FOuChJbeD6oOsAqGomAkCE3H
YOzlgsZLYR+mhLisV/JBb7HsHsZxjUsnuHkfUDMBDrfuf3z9KjMWhnDmo35uScsUQG6BLkEL6ACJ
gYMAh6t4kjWIkCUexB+4yMxzpDHiwP5bDfKAI8eONzqIGc4IxSh6VLj8ab3s+bXy3Sf6IfBkTyUW
M50UOWPpZIJp+vB1WpORLotYbWGMhrG2A686IvgWrKxsjsMoDVCtcp1KEeJT2ZfxNNFTthbBNbT5
X3vRtRKiz05uwyNfgUAs7tkOG0ekZYP9x79u6Or6zaEcNIiZ7E+pb0OBOCIIkRU4C+4GxBjz6HED
dgh6+MeuoUO8aREju1g1C3e7ezS0nwcy7qJLjc27IGHbVjxAr0qIPUq3tNGEz8azzmN8rCIfr/rM
mkGOglmlkIRMsKnl98EiSvZuzeHsLSNY24knIJLvLD8ZF/iFJtNNOu3pLpEZJmbJR0BTaOt2jkTy
bPBkBtk3KIjLa/Qp9P0ct7S0IRjTD8YawL3uZ2yMvDc5cz/VZBgFTfisiwEhuKaNsN9UF0P2FdfQ
9A1umj9EgOp9Vf/hBtOUIn8pswoQxjU6jWmSUyNpfBy/Yl/4cnbH7bwxWHCvRj6npimED4nULqSe
JSFdHwf4jRvWTEjbllcWOg+/M5WytkftSph9E4Ij7UTLW7nxhGX1YFmrKRld+vO14exM/HDfL2IZ
sSnXAI+GehC+UwhbH81JltDKyuKzOF8bkjwUUnNtEp10579FzlidKHAcuN47yc1ee/ce2ykSExa6
4Jg14QnJh9yW3Qk/Yrr8L0nvLsgNNs0aKBP+TnKwNz8eSojRWhIErsLyxBQhfWtA9+Pj9VPJIqBn
fXVvXQJdMsuEi8mQqhsNLAlxqfh/nV3d5XNZNGc5ItWyOV1dLGg103SziCtONhniE8iQI2dCxfxo
NFrmLTfFikvKra6d1h9+FRA6L7xfSWWRn+ttnpEVE2zu8YbG8XeM5wM2bZowrsfxcRhY51EWr0eo
bXztyP4Gx1mL7A7Ou1tHGyaNGPIr7Rupv8z0/mBqgCmvJo81NtWYR92EWrgv3LJk/UsRekLZkYVL
cTMMAEPGJIg9F0kYKqpX02SLoSf1H563Zh9ZEYqdTxlLYZFIuoGGYLFQ+zLZWiCOpozQAB+PXVCn
d9Xf82VVwVUpmaabJr7Rk5Hqm2+FirU1Jl2F9d+nolFgES3vo1EVBD9vVN3/vlaPZUcZtF2epxyO
zeivbZct/2Fb6GL0UE3oFqThCG+o6CLtbP5iL4H6EGjIsBNJpA8WSpvuBnSsbk5ARIGdCm0bcubs
ImMQ6FwbVc/ANZRey5MlVpTuEFbky2lsZJQfQWwCkwaHjZcUSnWUhdV1i2MO9RN3DpLqCXsCgiYH
aBBJx9zVMiQPK6NCOCzWBu8E4hbReMRz4OToe+5jsbDuYJtD13brDOo5ORS9mzPPjITsAOf0pOU7
MWibXBuQ7HGIcYuuUmdLySd0wYQcxmvt8lOm+vHyiG0ScjQlRjPN+24/wGfHxswG8q+2WCyZE/Dv
Lm6HnzaMSyN4AD9qc5ziYXGyctciIPdl7/CYN0Pkd9PrvjRi+3ftdQD1+u43dg4iOTqoGaV7F5vP
RgnEtgAHJe6c5yqe8/4g9jtvJAs/gjk0qRrYWr1En/z8K9dBp7nrxYTtfKYMiH8hW1GjEHg+i4CU
2VQcj2KZRgkrekEVfr1sjwe2pbCrm/s/qVUUpCgp5fQwA5EB68ZqKJ2yvehClpIH9MOL2/ilN5yg
IKYQKmkscKwh1VhsiawG+/Zed8Z93vVsHO86s/cqWjZEAt/v3xixhAs3Dod1AThw0d4XwUgz3wKq
+RAhQIcopIQsdJj+zdrUXq6/ondlaqWftknnN2mD9GyPvtE8du4+tDO8tsnm07kRiswBBzbMvzt6
lun19FKO2jN7ZxXvafqWpo/5ggiDTIb4iucX34NE+zVSOy+n3e5Bm0Ai7qBnsYGiL4I6eXbSvjQP
Vu1Aw1bEGbU0TmFRp2tL0CMB3R+T5vK3XSjRHo3W+tSbJHQsZKVFOYQzlDjnlLorxQ+rQ/Wg8ZeF
vWG73Fm3acVfkbsjQItYVUAY8MVuKiKAauVHZvvzlXyNMEPjcd6/ZmP+PcGxy0L9d9ofozqtv2T1
mCRaJEyrco3m2DTU5JTYoh+0QxNXuDbKnH0PVSgTbx/rayTr0UMU5apIFJtafVRr7NtwVVUn/7GJ
RwWoUgkv6rpLvhddkS81JcZVWCy71kveYt9JEgiE/ZCJedPCi0s3M4/bQTMbASTWZQEZPwUHIjpl
qVK5gFr2xefvePJ0CeK8Hw1oG5nM6796YyYpqy37TKpwrfhLlXu9RlI6Boaj3uuJeIGVS2do0dnZ
5NASLSY1d2RLV6IFwyi21/tt6qwb6ikr5co63KeWjXrVAs5fLceMpEl32t6K9BIsPPNF6NOh1TSJ
Izn2OlyqLspbdiKLYUzQxSJTPdcRF4VWLvtFFJQ7kQz/aPJAOqQvyLlwLDXxXqBnIVS0D2pMJ59d
v5bs2iAoythirTFhq7rASbnJKERBUyJDEcrwCmh53CCoxFTWS5zA0owAC6UWEajQTEbN6VJa46Df
0QH0mypIh2EKdzwCK7h3IfJm0sgbwBHXaIzFWhoyBbOEEQzBQ/TdcvqqLSad8s0mWEM8gK2mmzcZ
hUcagYLh4Nt70DXUXDNoCjGYWebYbmWA6dzP5jW9tgsJ2QpiVFD3qaa+iKdj9WZZy+focVhowq59
f1TPEEdB5cFhGdP7sbkdUlF734linPcQNhQaaF5rgbS90bW8YqaiPQQMOIc/GKzVpBojGvxIP2jc
6kGufrbgT5rbUCSRDsBQAykLmPfZwH6IwpTFRt6GSG6bHeCXytKslAu05L2ukeJgm2POSd7ndk/i
b4uZvmHymfRPHRlC/fsT0+b2HVF2UHhNeM24x8w5HHEie3KMZt2BMF1t6AQzaMeTe/9jpoA/RJtz
qmqdZBQj+s5+DRfkSQ9648V/bLU9seSISV6LNjSgBov11C0qwVOUunmXvyM67XkWCX155ts2gz/G
2z48qkllcFxUYv3lCnv/Ihy8Vsu9iA9nX+pOGAz6zM3KzRoera3Yig1upq89I6f0v5uDyfDzDZtw
OdhZVTJPw6SCVruSEiZ4n+c71nbAQ6f5OvAP21U7dJLfj8+Zx6/QZJNtSK6cRdNRca1Y6yMBJ+Ot
QOh+qbdbJ7uPgNXmhZ6VYOxK9YMUg5v3NT1+aFYCFthODxlThZZIVUbSxgHE8Jfn+CMILIf1+Vxo
HkY1S33qIN4iMBpGjIK1Zw0EVJxUpjXef3Qde5zy+ED9OWTrVNju/1JJMTTQYcEYMeg+L3lrzrpJ
Uda0IGz/AmbkPo4ktg2LqDBz8ipi+luLKI1XWThF/T3Y8WSegNQXAgT3jt4sLYVJTcNAAr5V1+cz
c4MwUZmWIpBo4SnFbgx2SfbLQlSXhgro2lhxr+9qjQrzy0e/oj2p5+NwzkdBYJA7xp0PE8huY7Q/
/GrcrB+HvI9zSuEUb+6Udclgn9aOb2ge+EfDaKNfDcw4oitduH72WmDCy9Y77+VNWutJt/oGR1s+
nEqsobUfQbRuidd7KNWMtLkgjo9mkqXa0XNZGUpnSbc6HRqdIwdEN7CsE4dCTMq/BQnXKHMa+/O/
mkZcTzc1fwVzG5FMla/yTWMwqq8Ujc1eo/qiasBfnEO3RU6lBbb0SWm0AwGw8cp0EKsZjJq/Em8T
ujivdHDadZ2ie6vOQd4IUHdi8wrp7xZ2Qi1ywXdXkqN/xb4dBWEGUalWDz8xD1wUCpX0x5b2ZZZf
cXYYuyuMLGvE3SQqo0ylWo0Lb7N6qeJPxokcQxkFkBrZV1bIx6+w8DQ8XlC1PI+sQ9hhSiTANahS
ZB2eMLt0m9sl6HDiAlFrBx0d59mB2MWgULdgC2+vSLaOpu4BCZ+x/LbwiAaPhj2f6AqDn5Qn1/un
5Jl62rAQHaWBl92s4O9xysT91i1POuKB6hmjHdMJ0uRdLrnYnttMV0TpK7CkEL92yccWxqEjNEX3
/auPe1eEx18FHFMHvQ5N5gABHk5OSCrvlriRVgmf7o8hS+QCJpWaTtMK/fCPZrHjGv1e/f6iui0t
p/WrwOBLq6m7awZIcG8vXJ7d11c/kQKoEiarD5PzX5y14DrfYYgYxIUdSOYT67LCVQ831e8//MEb
26v4Dv6wD80le3uOiwkQFbX3TWsxqhVZutrVnW61mLYuKB1AuEbb2PdCgtyZBrPabEb1fteWBJar
syhEKbUtKMTUJMiz1UFlDzUHql61pEu/RDwsU1qRK/TRPpIPm9gfMMRay2UckBONfk4uiTJ1WLXS
Td6clt+u1oeT2eLKRI5M1/aei2AibSe8fd6vXT4ekB70Kj5YhmoAlggYXSBegMkTCxojzZhtY7jH
vTz/qLg9EstbDdibHZ66XjjUAChP9RW0xlPW+PCB1NNFuDWnEBfT1nohkEkKovHAjwN4++/dbDmY
by2TWoS3z4nk1m1EPJGHUu2CLel7VB9cE/tdJSc2t6i1QsJ0Ol6l7WBUQQsGUW+U1CkpTEZjWgal
K172K4zXbLl+UUrh46HYbM/Ku4yfDF5VRrf/lSB95j11WQRvnihyOAJMU1AGSv1tlr79GvV3RisM
EAaz/b7SBchZN5yEiRiVszLNEkLL7y7A4axgDkBmkqFtLEK4tqfJ5Ch5MaRYL5JPlSz2IgSsYrru
Tr34uz9OPo/1V5Bv9OVbd0hZr/5RYKKflUWGS5yGV7s9ZixsIZVLZdjgECKzP8Ylks2CyWHLNBsy
eD12iajDqZCMRGasSxP2oOFChaYnfCiO93bC7Q6IY8aLv9r0Y1nW0ookozgQXnMhUxyR/2o9IXaZ
GK/68eNF27wDKK+dlUZ1z+nLEhOnK9evAbRcOHr+pKURJDF+jQF9lIcmSmhTSw8/AvuKM8B7/Ve8
N+zC6jNVhMCksOIqfqeVQyluLQ6pX5v7yN9UotWzjEnKB5en8gMEWEwOy9owWapLQ4veKNhG/1/n
3Du1sp+6hmz6n+OCg+hyIV/ZxMrt2mzGxCK9hTavwqtaSOswiFUiINKe2Ws7oU2WAm1U2Lpe3TmD
cBq/aV+ZFAR9U3xA6dvq6c2nNxxboHhlMqkw/Wg4ixOKuRY3VYCD0P5ccV0muHkPj0k2aKWAxX1q
UkD8fpxuRSsP+dsZau0u4s62ZzzX/WHOVpXMn+QYt+s6cY4EcAhgEhxjJd49ohtSzzhIV/Tafm9j
6/a+YunHmG8rh6xsD29rz5LjWY2v1iTICB+XfIJTW7jbW7ROb1Uq8Zu4OndVwhqurwYnKWOX9Jg9
W4kEVSS56cl4BLWSU5eZPm6xih1N+uTT0nC9wqZraeL4Skx9++T2BTW5sF3A4DhB2nKZhSQTPjPt
3EOVcTwyqwOTxWmm3hrKhZEfpCho8bsY3c7owyNxXlZWv3EEhXxuEixT3niuYH/7AmDUp+A2B5jh
pdlw1eHGzdAHRVp89Yh81TBaCGLoAtC502gI2JGpR4OXT0G3NhAYsj+aI04jpRek94o3tabsTdro
RvZ1PHAR98Iy3paLfkOBCOjUImy5VvpAw/4xGJrNPxH/85X63xqa1ZULbn0jSceJm39kDN18P69N
3RIWihOcs0GTIuBkilyBWF1tBV0HR630VpUQgBq9NrtNrcnWIAisOBt+qQ4DNkQVTQxv7uxQtak0
TtFLT8Zm1KfiXkjyOg9gfG+gHaeBjLGfWLazJmWQ8i9kGPqUd+BkZbHgZz2kTwTQ+R3jj6iMw+td
ivA/EUIkw7KfB9C8BmzThcKaIvZBPyQCvtWNau5KlBSjP+kIr7Y25+YnlTaphET/eeqyPYW2rXes
WbW4Pkf4jlVRG08KR+dRrWQ6vfB73t7Ck2E+qGYalskTYaa4hfh/1p+UMUtGEJSGXKhlsk1WOg9B
vERn6jZX8If+kvmLuio2PybGRhWrUddbUpHfN/ILsMakiZlmIsWPiDlHOw96//jxtgKQO4UsHWEu
VusmfP4nEhoykdDGyOTFvfslth3OBR+HVcNkqQLPufO/aUCA3eqqdfO59CChYrwJbaQsfyWKOk6j
RXEZcZ6ExfZnKqMaZOdFlmgeORxsTFfXAPtUspIrkK0I2Kw2n4XVFKkV1AEE/Ir0yRnbTKOL3eYE
eapmIX6uvI4WvbK+SHI9ufOomVdZ1b6YGVQnQNtomFxA0bVv3RCDAZ7YcYlcovnZEr5NdjYpFvWO
5vwh0szmPBzMYSj7UiTxu+Emqnj2HMgM3y+iT5aN50BgFA/9R/aPeK4nPiIDl5xL1fA+oe4cj7Dl
5j6acOob1fmj1OLs5UlSlKED4G0xYV+A6jUqhbMLTQvecmArIUQJEboxpvl+vRvCk7y87xIxUtmB
mHOFO84vlSNjdhCf0FXx2mnSvzbak0PTNZJ5jlV5Bga+b4Nk7BWvD4Mp4rrXNS8yE2dUltEp257o
L/LOOvObx65ahBL0cFUbTvx7hPbTB2NrrTL+pHs7hUYg1g0I6HGP+VqF02V4PN50Vq9iDjnZkZgD
0cGrDMDo7knOiDnPjcY1w8zlgSWhZpw8PVzqAAb/jXJeoebMzvy4rXDAW7bx1iZjQ3olgs9sj6eW
4yCRCpRtLm8Xa+Shx0U/k7edhTeBH2uOZ+0Z/RT9a4GhyqkHWTnqfrBUH2GMOQSmiydBjNeehw2l
W0Y8JvGGnQ0Zj0DdZ/jfrHNKBwhfZOyS7IzmHozmDPqh+zyg7H/jyc30cFE5hk6Oc+ffLIJHrGB7
dMm7KfiV68SDRaXEKBYgGSlP9AlAwk7tVoi8BwhYlKjXAFTJD64TPO8ZL3WzzE4iFsMg0Vej0LF7
D6QfEjKaBTNbZUGPYGTwvdI2Kfp2k+SitBc3ynXMrfSPWxLwfpGInMoha1t4Qbzs6t6t1NdkFkAs
a6c6SsJ/A30L0AZGgUM4qr7ayRYOsyr2kWGLX0pFQEJVgrL9zGRI9eeVAtnI4BExyoKotusZhdR2
0pKN8NQMQZaM/0z3Ild8AqeppFpJhkopvFbvH5uUaH3TB6YG6aKW6qEx9fJD/mewjskebc/2WvO8
LLcJgxYgnK3qg/wMgzl3xZ1EoJBorUSKxvx2lyL/nV2epv8LeKsQY7upLBleObHBNpJkyiQnIB7v
MYq3RpZDj6mhgi+shOPdsbjuxsSR9Yfr9MqgBCNavu3Qsi3W0DHi2CBEN6WdfnxXA9CSlDiMMJY0
mf/CS8Tk06rtDUqKvvD71fWaDNHKb+V0vldGKazqMKJs//N794FgwHrgHySJHY1QXbpAVheEKMJ0
rXDIlY/N0xKMAlWsUB7OGWG6o93jzZL2bzP6MgXxuPA4c/7iOhSbjE3rrC5xGT1k1lL2IwhXadkA
FXmiYfz0hF9ttZVwFQAqunOLA5S0MW7VrI3to8iY2y1/WS7cw8v/KBnfv3WCMoyC4dNSdbb0ORjI
g10Hpmab3V2f3gL/rLxqG0qHkAEG7txjHUq00l94fUtBiLh2Nxh+lwH+NHAfnPa7WwXeqffSKmbY
64pI1saHspvdchIceM+ccBdozyaEbjCxwMDC7Nb5B57vZSNcij/ULtw7OL3c6BTB3nmylNfmVaNW
yoQqr83byzJvqT5iZP9JA+0nTKohxvkCHMzyR/tmstGHJjB5bfsuIuBueAxYDnTgUzTeCBLIF1zp
zS7rvJTmZ65GXgAjJSbJsYSD/4XsSSUnZipaamvfc1qbJTA80FBPeiePk2u6FgAP3vuK5sg8ja2/
X94F8LjMit1bYluTAkqupys6xzSmjJjCuu9aLIqk4aMzCsCzapa+gYZsA5bSQHpHMN68l4in8MFQ
JetkM4f+1d6+EVlxzN4pH/a1jplCjHOXZlva2ReM5BqgiuknQzwmrGgmfvQzGiur8idtcyNbqnbJ
Q400OHtib3xP29LIfGtNqztW3jgSk9/1r4iguVwt711RryK6houLi8Fv4hcjYA7U6Lba1FNaWQMK
Jd55JXRAqhM7/k4QEWo7R7xS/5Z2rR0OQjFxVnUwAWnAGtnv/yQGQFOVoZnB2mpaca3mLb4eSlEz
c0ENOVvrEIIlWlrsaAnR84Cf198t7NrmlatJEKuACqLExSH0KCAzhooZ8z2NE1ULggGXriz+U12e
aflRBW8PKCdrth3oY6XfR5FK/bHz2AhbqvRHLM3gnJaPuv8wb5CHjv55sin4BQdJsjFfRzbSG8wO
UjORXJ58Qz7ENwxgizxzPB6bSAgjQVCk331AkwMiO6rZ55ofXm4tL2mVtpMnebUO07XyTpzfsy6i
e1+u+PCAooQFgJqg3vXIpc2zBFaRNeCmGlYpzsZ3Mj4Ofma6gxLlxxGS9HtmfkSFHpw6+MWxTb2+
gwh0rAmuzTNzBQnJqJx8S+bQLZ3xizk2Pax6dFodMCstQw5jrVM1Wjv6R7ji92bLsWRZM7p8mIgb
X9wC62IxDfMSkXfMiB5gv7a0WuKJwPZIcJwxARjrVSKE3ydHuSep9ZiPunEyIs9YJjfwcAcM5W5Z
9KsGvPJUl2OPUOhH5bKmtM1x3nrRJlMMR5FcwPud3+UBvjGilCYK2m3Cvh4588cci9B/N6nQxG5T
z7xSyXnqDgh3XmYQ0X9iVWbXcTOfWBhxQkx86Gr7BbGYeTd2GjA1cSArb1G+c8hqJWx7ln7DGXLM
l2Pyg8hjN7V5YhxGSSxzj83O8SSJQU8puVoJTp6l7zMyoWC3DnrN6n9elimNj07Ur8FhTjPAOFb6
cdq/lGAGdjuhcEZHJFQrLkshwR0rR/pzxQV6u0EKN42uOrwImWx+sZOGh8ISyzcX6pRm57AQbRAi
+XfbhJpgaEN8dpOkYje240nl+cSHpuHJUCu5x09/zmIxurY1gDZYzgbo3SGHHaVRgnrVTwlbu+qJ
VnNA2Jgmzf4sbppI7Mu/Et8gvlldvdSQozPtZkfJoAWxZcURpMoo0yQiEXplyPq2Lls0DtNXbiPb
3Glx9+ZjkTtrpRV+qVXQkGEWoBIQASOT/6CkRP0ZFMSE/pZ7vd7oPKSnf702zmFBXHadR+oVajmY
pwvsbI+b61xTVu5wSfN3Zluws3A2O2+9w2XkhHXbwN1629rMOY7G0a0WzyKjOEQchMuqcUDzLtgY
E3FB1Z8sBoXyrwODObycqRmwv5VnVoE46MkbOhjEvbaFSRAQlzKpB40fj26C17QMysRtmMa58C9t
gfgnkHeSiig2EqXIRLQS6xVz6NPs/IWw5yyd5l/N/pNVI45LDiDbH/oWp4rvdYiflb6iU0VcZzoD
7Rp/C/ZZyRWTjcNZCI+Zh7eo5dcsNh7QAtZ7feLROUHNv4toWJFqnsA3Cj4g1DwvXr5hjF+vdJ+M
5jjRDGzDQ+brxSMz4spL4O01+YRI8UY5BFHa/07fAmmTwHJE9rk9tMjF8N3/sF06woazoO257s/7
KdLN7VLtd0ZjpfP9z7CmG30UDFV/8xqm2EP/eum7g/rZu/6f1wO037imB5rTGtgy611m+aHoZNMC
cf+7Xg6Oaqf5qvAdhXTf95f4RwMCARpB156pJGmSk8IR8za6i+gtXsOOG+vb7fi8lUBulw4yFZxn
6AIcgtkpK3PzLOITulO8J+oC3FW5fIeL4P+/W+fXJUJ9utao85zpovbkVc4CSUVUAx8PQxq0ZSlk
cyY1MZwQ3CV9MiNw+hjI4/ouh4YzHWe+gA1vchssxlIFH4dDI9L7k4T9KvR/J7t3FRkv2MECZkff
j2hyVtKQbZf01znUM4bgNxKYuT/TOQxHprMHVpTVadChb0p7RUp9WB5mYJlh8tQ0eyF4Fi15w68i
O5UOf1yh4S0u7ZnByRUr5OWao4ZXe/sN2E/bGuRGWdgw+UF1ESHNgUGzGL4ej7PWzs9LqKk2jKLI
ZeH0OQMJvVo+vmey8T2H4HZCecSf/VT/WhISavLo8jFbFe/zL2D1G27W+sdmzN1a8y3jAoWjO1YC
4rd2TyAYwe/RkgKJ7FRzjffUxI2NToV2BZn7E2t9I4wW2axVQAVNdg+X1RigvQUeh+Z4WqLf8eV/
YiTIjl8cIa0I/sY5soZmPRU6jdOn1eUS7DothLzq0O9iQ2VLbJDARylFv5M4FcpYTYXLursECGZd
4PBVU2YjK5TWJ+2IMpz7NUi6LwjUhB39MxZ1xF7zHpL0cbaIE/57ZNNlcweBbSaA0mF3LUPsB2tM
JKyMlA9W/Oi54O8fxoL5OqCXuVUqiuNU6Zhx0KTObVL2KT9y2Sz1q3MHcqW1cfSXWh1dfs75UUaE
szhAnYS1g9OESWiN0j4shm0mxETrs5IW2abtsAnku2Ry/1Dbg56pL9mKie8BN+GVCvNQf381o8sP
rXq2QWCP4d0Kh89o8XCbSmvZ67D7Shdu7LQe1oyIaHMhAgEP82fLvX+bGyatXvUpbFD3+u5lac9l
YHn80GADLOY/CCSLJt9Mp8jgij2jOc6pL3cduu1+FWHUu7oz2Sdlh4qApjAh/dKKDVAWEzdGFE5/
gjpAUXXTw7f8QzPB+2aEMv0Svr73/Z7P4TJn4EP1AaeIuQdnf4Vqw0aFnBnmu2UhFPGI2Fo63tRo
tM6Y3yqKJyUHJz6PocdTb00x9tqb686hg1hhs+nJUmOp4nG9/lNHb46idLle+HWh5IrdN81P1Qjp
v5CgrnVIIyZzPQaRIO6DZWq1xYR7sCsnWrr0YU9PSCHa6OIqeV/YOCyQGSv9oODBCHJ3TRNhCh9M
QUb4T3bmGcD1ypJT8JDrW4DNPGJvZGJtyqLkKOZp0KaOFvxLFrIvjVkbOJZZRbDpWyGueemweNQH
Q5O4pTnX4b4tJtCNsmCx3gwyXAHpVdUMAReoZsf8GuMzZVWnDcn4PVaM8Es5WvRP7LQMmmLNcP+x
b5PRuuUhaYrSRPUu0C8xhNMTIBJz11XUTbD7jO1A/QX7lxE4NdFZMSxYM0U9RZMZb/I8WCNHiDaK
5aCPdifV0aaU3J4SGIgMSi1mAY8chVw3xe9q6rxm3d+IvNE5ZSvRW2DkZ9APND2J8phjPvEShuz7
rGXWkzgJr/Pz7SJdsDoUaCpqVCiBVd8vo98PYHN3sCnnZciR8dFF00BkyUsGx3tnxpA++TNClwC2
IR/nqLLDkdkSjS0IlICoVudTVZnT/ZrHE9p6BIa/4PlfsKsd04EiJZEKsGVXZE+1xG03eR/RGQss
9fCXtV9qmknooCr4lXxTqQPslCjanx98Stz/4XQt2fuulbwI8pVzqpwLCRI7K65MpuC93LRVxfp7
qLlPxWQ2si4vXr9WOSVL3R2+MPAUlznPwj2sheQSj/n/zY/TU9IbHSCqY5p8qsZ07e4ePksrgLoj
8OqzJjP1azmKL8k9cricl2yQ0w7u+69ISzXn4faxEKhOtKBuaElEeMsqrwMovg/T4hzTb+mrIH3c
10tCodxeSTmb8g2JqaRQAJLI0dRMMhNcM7Rjvx7GBP79Ghozrtu7a6LDJ5ILsyG1K4uwkn81E6vv
oNYWnchv5BgF7J8WU/Tz8cwcy8G+UETWZmNTuBpsArTvTln7WtgVwGwP79rxSYlGKj0ilQ5sNVbk
IbOsF053YdRz35aE1LQn32WVI7Tw4Bzap2Yz6yX1jRafuXGZMjYnr2jPrEQ0nefFamViunylFIbw
cl2YucNQt2z6L7aWp9n02MnPByQOBf44kQRBgPksCyYhdUJV2f8TscSyf3tjJbxClQuiHBcK1Qtn
XD499k5RqqlnFu2vNqRb5WXOKkGp/ogmJr65e/SURFC5YT0bO56D2NgQjr21KT1I670lSTIgyRCz
tsvfn3yaTDkLObq7smnrQOBhX5GXvuSAykU+jv0toKkpMAVsCHNM154FnXttXMalZizX3PIii1qE
9G4qNUna9qkNlc8KLqkG/WNFDFK7OGLFK/CstB/NhtG0WOdv0BLWzV3zm5Wc6EuFGPq7ANeeuFJl
PNdqYAVx9CoH43cvP6IMnkNEWeD53OUWWLmjMebPy6rkZ1pAEeVOgBe7+jfSmSOypcvbOoHkh2Y6
tUGBrU054OOARagSMET+NX+IMp0Fors3kjqmMXM8uoE722BxFcNbgN0JWK2YAjP5wqgSels79a8T
cM91/ZO1Oz/d5bBe0ZQAsRJQGisxBm+lnuBg1Fi1+NZ1HZcLVTo8KZF+ISSu85MtqlVf+mcbI+qd
3iSnuFIKJrTV/4cCwaPgD3JVrCCFlZSSwbYzg3wJJX+QO4a7CYt13s9O6Crcr5kxYaH95ozh7ecp
RmeCsiJbnkC5KA3Vt4XIj4xouPfwkt9gQoOMd1TqlYh5D7h2iM2lLXSPx0f/7HbQ1d5TNpM0HfIu
dqOozHOZyVQ2A4hFdubEDDSFjL+ygP12n7IUrzQj3YpJiR8hI8ARYnMBqN7trhog/3Wdq+rKpCCM
4XuxDFJiTf07cJRG24qHyDzRCV5nAX3bVGGhzwJrhJHMcnj857HpPjFRsYvSjFLDklWir+PE6U6Z
EJ79gnmlG1devsCOTv1f4YgfcDTrz27RousRPg6/2DpCBbkyQQQMIpJMkFGhqX45p7Wtr5bVvEZx
thJISqPJc+0Lb0OfRT2k0B8/7HFtPkuM8ziEnbhO2NLO+Y4eZULSGCmUB6mx3HKJ2uZX7hzeL0Iw
iKQcItDHD0phf0En+WxAUznjRMB0ygxXLB7U446cfyUHglGD05BWBIHB/HXsG1mvinzQBh96BNhs
ecgueFamr0ctSTm5YU68++uFTNw+16H+G2oIiIYaX1OAg/3cajPb6t7nmL8LrwzvGNP2tbtJbXyS
N7xlYYScoI2oxyaFbcvaSgBiTPGIsIhqNty9UpMXVlYm+KGg6gc1aHxFpZPLDIJwE46LEyyaNGkm
wanRvrnBYudTpGVVo6GvzDi0v7lhlw4oI4+ppThkBjnkw6uL+9t1ODyjWc6kOEg8eTb8AJhacS34
vx13WZd6FUw8qux/FWJdRC6zzCd0oj3ffna3FyzuY+S2omR8noMZz+5bi02g0O1hYeCcNarnob56
4NEEGpUtaqd6qtc2sC3nUnDFU95LOo0b+39I1+Fheza+sFjtRqzl3WGF0gdS8SLoLunPdbVPWvlF
0tXPrVf6rLGuwjn360Y+p5BSM+icOuQyoyRSfJFnjSgWwzRyea2STsK/ebh8z1JT2spQA7HMHDsP
S4TnhpqxHcW5JBaIKSFvH7Vm1L+lIYHmMjqyl+XuulWsIrLcHY6DQghMb7E+Yv5eN+uSq9gPjM/c
MvETDtDUf3pIQRNVp8DjGdQyttuXov9x+u+Sllbasc6nq8orpRDwl/LTNlf4kxqxaauGNEDU+huM
9zitUa4ZDFd7+T1a90mseTVrpu0z+9PXr9m+Gbi3gYZaimJpKfIl8ErJCAbvMB1vaXinNkAGsz16
YS6asiSlTY49xlHAL+is5BKuS1v6077Q9XzwcxgR41AwqCSCaaJHJTDWdZDBgfKDWoujUFXqa832
xd3fZQa0TKmMqbUZjbvH1XeMtGuGBwciDiIWrjm955XD37hIH1cfZV0IkysudS6v7c+ohc102hbn
cgA0NI+r3tvvy+YR69F/VfP+XFaxtMnercsdOsfugloa5IeRWMwK0EjQtewmpSXQN4/U+On/Hmd/
+mkAR6TtkTyHyTLg6Bcsfn0DHemDmY0f5aq7aX7p6cH74njtwZ+E9nuIcJeOXosnaUgnlChcqizI
ac17IVOKcJ/i/DxQvSfBVzLiNlrMIt3mzqZ4hFqnCJwJAQlhoS/Z6nvehKD2UcTDXw8kV/r7uUIi
vHlf9TrbbNxW8PCsg7EYXEnSli1cS9T376pvbYu13uoBY0+xqoP3jGDunWYCneradctUVrtTodza
QCLtq+q2uWCG17shmcwCo7FBawJsN6rtEMi7wAmcMp1DKRytwPkKGFtlYSiS+WSJ+jBnjEbKzzI8
riWz4911Xh9g3duUMWcq489WjE2w7g18iOSmTproTMlbdyIujn2JjhIOcBhNje1Ay7pl9yzMUKgC
S2mFyrjLLxWMUfIJVH2xk4J5DvHeehSbdYwA9xmAz2nC9P4CaA206qxKpdTAxoEJEkM9NeiZ/c8D
UFPwvyj5e2D6A6MZlseBNRYagwpCheHYpGYCTP6hUM50MCUgz30nremvJCOjrkBSqnOEOss0Sxu3
4SHnfEsFEZNjpYztWldSg2WG2TGj+iiVkIgAj8hyQ97w3zxzD6DmjIBXXOjCLf+pmCwNKEgv9K4A
LgWXOvC5Go5q6zFflySszE+h16RaXvegj/5OdfCA9rcYNcYPSqrp51AwdDEYqbUZtotIrsl7Ap9O
KxeZg6jLjzi2w/1eWx0QcEM2vTMk6P6QKaSoAFZzvBMhmvtwkwSJAda3eRrlPcnw/KgSqe7GRzFr
9jQJoq6FycAOnPu6eQPafUwzNzN6Kk4TbAFZifQaFEXHYZJOJpirbnRbiYgG0BjagxtCSub7phRi
+7+wAyhQgZPYIHLM4g48sQLewLGsjysqHtBeoCZq0d9mT2VkEi3wUWFUhvmwmDVOmDhcIBJaCj7C
L8UOLAkvUTqhP6CyB317gUpD2D/ikYwokGkxyaW4XbiUncaV35y7OGCSCOAU+u5nP4AviBS/Bye7
VN7iqxPPK4U6F7odPx/qX/sFOKHg/wwaHE9vTh9VVYDSQET7DOM6njrgJhWBSIQNREKQ9zJIzYZ+
X5Kvm1bzD7SyiOFaKLCEjoU1eN9V/KYoXW/qQlxS6Jwlpa6KE/Lao+qgSO0+iBWU8IpzJX7gFHb9
ylPkJ38G7mZfkq/uA1FenO7hjT2/EoHEBBClJrDAoOw6hqbmPJ9Iu2LArf1hHabmB3vvlmWWVGuu
fSuG+TtqYJC8IH2D+wtMiW+cG1eY8uceOoyVaX+7tjWKDXbNb/WFoRsMsUaGTloSlAha81oekiru
8aulTJn8iDHsKiv1QSQTHNzPwnCoD8SVdAQI4mbCR7QJalaFlmp4fwwf8/K1++3+FjFTsIdpaN32
sqoZDgDL4nhbT4u+LmmnHFPlBBv4qWjDnHzN+wgKQ5RlBZ9AZ7vmH5Pr0lwE/EWkU6hWzfJ2zKWD
gN2LQfFrjJXggMIgmnmkjo1FvZaY2/hglhbmo/iyrezv/AIFkXZTVZIR8TdQQ8euoVTxdgbJ+jrb
8R0Vgp7d2mzeoSAApwfbH0NyMj3JcDQf5JEWeQ1xo3WsWmZZTjKKQz/C1uaTYam4A5igbLgN35Ud
c88j2CH4wTeOw0FNlBNIpEFm9syLxlaJxN4H9tGaavjruvi60hNgc4Ovp8QoNaYbRXBIwcne5mhw
3FahJCj35yT7HCOjvmFl0DJvrVdZVHBCj867YM2WUexaccX5tmki3s20K+nnWJ0XKo1JEzAt9jJh
7o2b35ad2hqxenlhbDQaE/7j0qZE0oid+0CWSDux128M1PAF7rJLDmQ4bvgKfbDDJcsI4E2IPimE
vjwQ96GeneZRahoEr3CJFQ4EX7OG/dW3u/eQJD5yxzBP9Ee8Cx3h7+jHHbFu+n803Pm63Wdmm+Kd
dMSEaF5ykukSN71id3FhrHCbdH91vh/kS78mLhSgL2B4vSqftJ57TNEG6/ehAKcCfd9GtQYPslmF
I/0xX8rleqVl0MuKAi1s6VQNCC+OKmUgBV9IjdANnM5BR9Mi4crOUrRGWoWs2ID5F2gY+i7e41ev
INCN3gbAg0kFqkXDUzDwO7WuMWx9otZmHzANK0yr4W+jusaTqB+4kbcbMxWcuwbv3u921LnmTvjQ
Vk5Gk+VKidQ80JmMxFusV9XAwzToznhZzTG2+MC0fm2b4OQkrH5o/ES5PMvJ3AIm93TPl05ti3Gg
RVgNQ8K4o6+GrV2npeMIIe7P4xv9Qqvmk0QUnuKUqIiaXoA6HKZs3jd8I2prQEPqui5+Zd4DJV4d
BiwPWE3YUqR3S7TDYFH3AKD8SLmHsnUU6HZhzp/wQUcCP5W7+EIy6rB5Tu66I965dn46xSR3Q2Zo
BPPhFc714J0/NccZrnQVhslRodNp3BI29G4pjDv/UfQelQECFOidUul8i5/MA80ofrBQMPBMFEOK
M0pdVvnNQx3Upiia9xzxuY1YAvNCklMuDKiegKzV0KMfkD7gKUCO0ApTiB4OmV8l0xB3EaVeKXj3
xNWk2JUutdkQ3tgDbMzDGl4dPuNaqOG8VlSTYbc2Lw9I7TqUGAH/ZealiJXOkul5YkCZ4AdHrIGA
3W5nzsQTtQapp+HI5xjdN3voP/Uc6q7qqPdaqXCL6zSU1/6UPNaSNrM2IacLnS73GhMAULG6XnJV
Dj2K/p7yGBr1dDxMkNDOxXhR0kASgaOCRGGMs4jLKUsOf3Yy1u0KCUnKQxnG2cl5JsPkCVkZjfdL
a1kWh/Oa8yJq9+LKtWuSAWAjbm/uXKypvOfIQbZucN3gxVdURNGPM2fd6s+5q+cDvzVaZxzAqSe9
3cMinO/P3faOUP9I9GGt12byuzkR5B7y9g4UNsftC7g0ECcC/dF9QEDP+T/3SK1m0hE79Ty3Imkz
WzBwNKsqNTVbNJivulyzjTMIcOL+HAFE63/SdG8Jusn1eKUI9Q9RkIrQk5E75dvcjUGHhImG5iEx
tG2lXBIpTPMIpaku+DeZtWzdvib8YhFL+Cgr5e+VCoL8gFPQSvePcN/lusBnILhFEj1TMH1Sk78w
MyTX9DIUSeOWU+QLTihyzPRHM4tZhOAfzRog08alwsAMyr3vocusKO6rHiP3pI4RbbYfArrgSBPS
+EO15cELGPVK5bLFmWKmkMdyYuKT63lS3t7qgX93Mmi4gP/KqtbKXMK4Zmy8laGF17+q6VmSl8F2
/jcZTgIZqqGuIfoL70hP+8YfBbUSuThJdQHBAQZ0vUGTJjOfczwrgzIvdqcr52wWuc/NatXqe7Fk
g2znuzz+TVN6jxtnGw+dDTA4Dx3D3ZXpxfuip03/DnTGaQJWFyihgj8zETcIMEqGZKtb2LzMNm9w
kI+JMfcSLIdM/m/Lx2HdNBJfEgUXO3NiKq9TkhtX4W6IB4Bu3qZ95GJU77SLJk98Rb13pnLxN/K7
/P20wbzvk56A1+KCFgFwCmBLnXUf5sc4O0uVeG2vxWGC/VTTBHiPGSOEcbOYFOjEreOSkRzG5jsv
6RyPKEG5Wot7HL2oDVBr+yZOdz9QgV9AO8zMs0Q+hUJn/U+YDSYo+SVvvTUvRHJ0pdJhbWQG1686
oEuR2IzWnY6xtBHjQ51ynzoDJcV0dnW/4Jif6IPfRl8Q6fHjs8WEdArtgUSFU9xuj/YcgjTi5GsN
CQRRt/dMBchK0HUgUEAPrVBmKrr34JtpaoFpaUNKRx5bFHjnz0xA2EdNDxESaQFzO3oj3byHl0Wf
sVFitgmk+AFAyX+Yd7yV4tIzjX2PFtu54EX61lYohdAg771s+deSa1vWLDkoXdOouzjnZY+loVoV
nCD1vQNbWeQgZX1gdBiXBk6ZxI9E+XtMXTj+7zhs8zrGTp3lxXYvgnwrd9WNxAYC9snOhQqmlMVg
TDZwI5GFZv29c0+Vm3ce411NGd0nRgq09ucgZfnqfMFMKg2ydGp4p9ufWxiljbQ62aupcswLtZjC
Y2XZuEL10Uyoy87UUVoSpQy30vTBBJacUZ3BSRFEt2w6NcGOK/J2ANLA+b6/wYDlp51Y6EY+huSQ
apVMonQE3gfqa+pjGR8zpImjhnhdl4XtI50YJAARB4Xv1iFjpPP9W+VaOMjRwMyrnAj8KxEJ6FF5
tcr84+FcafKFnGIp4FIzhl76MSVIdCcLzpOd8eeKXZvB3mETdRiiVfSIEDmrzQAcH/DqMkT4XUGM
O5YtVlvyeyFOomDkgsvmtIYM6oM3GDwchoI/qFmynj5kU79JYnqJzPcMHnPrsPs4/IO4VdX4aJ6v
cfVSo4Yw84qZ2n9dl642m/tJwF0P/kZdTxVGH4930p5DiLF4XzcxiG9KNd8ty8tcQHrROFdx0Zwp
LA/g/fuDTVqEK4Vzsq5Kiwc/h0BiTPdrauNEB0lxSv623WxWUXGDrG07QjF6tveU4u5vptghjrkK
QXswpnjdst5tMrPD229xoUfO67yHBKedJxKdkhwkjjCfwxyKYN7RZzNYILyxu+es6y/cuZvVtQ6p
1+VLTn3HcJse7PsQ67TiQfLK/+JQKSVmt8n2+cvuZN56L+Fd93ImHIaVk+1Fmtj4Ms0ALyfkIttE
7s9vQW2mke4x/DMotJDZkgKrauwsE/WhH3+lZha/GG9XIsxxTYj5tubxO/25hOquGa6CTknOoHqr
eutbmbgT0fxsVz2H7sscNfSN5ewdn+MhmsaRfZeIK66+qZLzsXha15zgJPqSoUuw3RCe7czDq7+o
rHylwVa9WOPhThgm6ouwyNdabZjADEjUmObTap1+jTGGSxXvO/G0PT3Xyx3WSN0JQSXwRznRxXjI
DPDW+H7WZP+wh6NlgwNpe5BfJ14oLa9IWA9lHvyGANmH8WTqu/4yY+1Ia6FRnmm1fZG5dW5nHrwo
avks63muxnKX3dfxNveNrstFwLSl9/z8H3Oo7mxXhNA0U5pZk8o4gjtgGOZ0akZqSfDXBp/j/4RH
tppaFvTAkOKZAPYV+MYN6kWYHTmjeqwlwqP1uYDE5YMbzQlmlUANHxargE0gNZvd+2kb0/AMQXHi
n8j4jGEVSW2xvx++vmZtuoJBCXW7iEDp79i9jkRK1PtgyMUbu7oAmHhVTCNsdGA9r9d/2320sBzp
9sel+xd1GQOXJCE8u0Y23v3q/30/lh8V7uEAISiAIgsBUpi/7evW7i5nCe8vP4wTYD5Ue2n2T6ls
SF/xBvtOsOsBr77ooIPDUewBxmb2ERRqKXOZLOLjzxqIsfsQd11dEbWeQ1NioHgrvLlOE7HLNsU9
TfkBs4fCX6n2ZPptzpvOFyw9eBbrBG/w/49ek1dbhF329EnBjzGYSHeK8WnboJOJcAzayuntmTd2
7O/8glvNDK5Ve9aTf9rH4NQGk+GRzkVahcmBInDb8yJ08XxYBujV3+3V//FAFQj5KrqKJcRpaDhC
GJ4ZEl/bnfqOMOyg8k/8ANqEacODE92tMQxfT/M39i1xzLRe7a42UyXh96IL3MOPxM9uGW/Faejn
RpTe+y8qSL54BDK7Go3ktZepMQ65hc1rpuvCmzq3EPZ8UrrXi5UBFGeAYsfNUEy93OkP7NIK8+aP
vlzG3fHxzhG7+RkMeMZQfkZ1A68zxh1nJmzUWU2Bw5ap9pN7fM6AkGxRd1Ga7KcooHwOe3ILGjVA
EPUENzhAy8DMVpZ81PPrnid0GPsqELGH1g5ZKxXaeOkp1RKf0wKZl6/MSPhODd216hCpXyUMKxd7
TWxadrumHhqv/z/KWN//8oubOzC9h2lyBUfvrNjs9tvZF99prPmu6Ca1Zu7ah+qAsnr0iGYLtq+I
hSLQFwllNtvE6JufWRd8clzusjxWE3m7ArQTawewfCPmuMFJFI6E6nUbZKLXhZf+Pwc1Ma+n2wgm
vpdu820OivPnfkVTYFbxsZsZec9CzqjPozjg6MiuV3s0f5HkWUDxSgiIr1NuxXULV7A9+BiTIOn6
1UJgxXOwHK/UlLzcFMc3DexTkxErk0xPPTQzuwaWPFPHfx9c9Csna3zBTBtbPqn8kQu9jB3tPo8Y
erKH0XsapJcayiaXJY4U8orGdmkW70O09mx3x8TxjyPMagKa9Fwjztn9DHveKEur7tVwKsKQUYNS
QgaDcHMTaC/BM7osi6tattWgmM9DzCEZzDtagRjFBR0Zb4KLX7MSFvaxvhDipiJu/yvqmnM2LkRh
FxB5DVweA0Y5x9Hop1ABTFU+qg9FbLbwFBnjoBcQYPj8oduEfvP9Ull+twIkZyGvoXDN38+h2rcc
+qsEeeDMXufSvmy/+qv4ZDkpktwAWDOinvo8O5UP8lzh1c2Jr93wpq/tOnQUPfJPPi96Ht/96Wlz
DzlBn5tc39lBrZABcvBEFYCmuHXqutklgpu2O5c3QJkb7C+gTkox/JqzrhaYvASsvQcKMngLMnk7
N60aFQHtg/x0aJyYHrormw+Kur6WgSH/necXUstVBwxxZzxhM78iom73IHjhlhgJ/jMzhQIsh0kz
+7zRrtpUbytvpSGclnYUHzTE1cuo3G6ayVCcrIcodgRqvBwk729aXjFSmIT8zm4E56B3YX3InsYi
DDjFGKd6KefkYoSqF5uJqYTY79QOMuG8w6qjiAD/NbFRvr98McCPxvDaelD+s3mlFBy9rB+F4IOR
IARNhYIH/rmfVtJ7kCC24jSkr1Hx+W06GioIqN7c/gBkX5b0pml1KEGLsQW2LgbaDFR0nch8MuD1
0L3RHzrWJYSWGg9r9+falH3SYC4B+jpLUkV0ctW8nmrKqWcbJSxbsxUtKmf2QWTBHxUkJ2Lye3R0
ffoX4JyqaARqo+Hfqqtui79waE1lGRExmdOuRi+HkKnvki+M3UeFPYxGddf73+MFwke0BW+RwE4T
CDLvVWuruk+kzI1X9VgPi83SFXf09+4C058ewwDaX7/49C6Oo34P8YjLojdt5rKpF/tlv5JZWfos
1R4R/OU8ErxA3OBMQ3jWiy+u0gzilLtczN9UP9H7j57FufjXZK+YTSLaT5+DJb0skqY4b1OcQYdO
GUj+JfNcX+0RHLVSc1QmpZYlQwAEe3opZzQVruc/ZBf1+xFeTSqfTiX+VaeaNRDfNvPokXcmYWfu
PQaOR6KfsdlMoD+FHHjSgJauId0ymbnouqm0oPYrBOPJfJCovVnn1vLyGXo8SZInAUz/Bbd+HDu2
6mxlJXHE9bF5ko/NsIKnzrwJY1myEZZprzh3ZaltfMy1fRM8CHuYeu1DE8f1zcHJjsNptilWLYbb
ppWVfWgnpH/mVi/SisWod4a15sLtY2NkQTfjVAjdP8upidmCVfa36LStuQKSXUqpy2hxMz0hGTRf
VSgHceXxeRebfRcVwJGfH4RoyKaVKnhwYhwgMBnnUsuFJaBM3wF8B9iiAjbFfJ6Fo1bgw3++fQfL
zu0BAghSDbNy5oxVKd2Pk+mfExw3TbXXlchUbjgQESn3/AIJgo6yQx1RwZx1T6nejk+UaR+rhjU4
fZxSFxcx4Q6aTgqFVqpgJVNpPXtgbxwsRtg9DVwonhDWvqyBtZmJeCfVSw0GmGQgPy3/RQ/Wilz4
/rS2IhPr+t9DFrnQiypiLrdAQAonAC4mfprxQmRvx39hWnAJwKOqCF89k72Hng/BDofDbpuZVvVH
Zl9K/lPHpZSaBE9CCIjdM3A3+BcGJ8VJhZ7FmdVK17W3fJpFVv/4xTrA2YHyLA5ENQO4k8/YaX3I
n6YTnvEE5YpwwLw8n+mXrSOK2DtXn0BvZGJrP3B9kFTvTI4kPgMVaEn/9/emgPqTnV1cFwJSRiVE
X/oPx81zob94Pb+vBAvPBAnvY2/cWxT0jSI9qRwI3g9iojcsfHbyrnSkY7FcHBhjndErxaySwuWw
XZ8C+ppt316wW9t3vOgC/dve8YNyt5HXf96BIklSPWVjzXecAb3wWO+VbGEm7bzWgm63neBLvaeT
y2VHsUVj3/6Fo3GN/f6KpK+anF2Lsn9iKC84pujnOXgPbAmkRWOlXF0DE8IR3fBCTmAC1r65sBm9
r69+dun3JG2eQKRUjDUQ9X/2R6cywibIOE4zcGdP0csw/LiSszIaO2rnO7MLfouz8X52l3WNZ98h
yNi594SUGI7Qx5iPmguW0op/dmxKPAHEG9YyJBjq86SojlUcWVudHU2OrCYHnUmJzlu7K3O+YwGq
hbaXw2TIYK8LIyvTMepyMpkj/qH1IVq/yiSnCueIl9mTLtcSSmNjNPyYhewGmHxaV0E7Hnskrozm
8I78PBrFUgmrTza+pz4ZHgwajfejdb2rmONTQxsuDsabKgi3kMVLBNdZxgRoNEOMYv4dOJT0Q9bG
/NpTqAgTvu/mTkfDWB3obn2KPIM/FXY6XcTe6KnMwCmYqCnslLBWyjKawDug7e+ZGpP5hq/CCom9
nhikkkuKex6FxB1CUAypLmSHZA2KiCtUNo1J8C6yiUhMU8BM05ST1K4wjejT30GZ1M4akqdCyD5o
021146DoGD6i0T8YREArCzRNjscXQy+8s6McNW2AnCRqvdVTO9+eSed6HxIXMG2kXWeHxOSUupQi
deMF+LrMW14SHPlZanFSnp2QasexmD2RadtkBY8yZWdW5lYiOFb7IpxzpbVRnEe5vgTmHdRPD1YY
xnW2m+uJ3NtHRbBAC46/cEcHCHHbOCUvwxGRILbkhJUTWKVwSwmxDQ6RA6+Vemv6dVPU6xSp4MQB
R58fB7c7Tgo9YedfImKrIjP++Pf+HqTmIGHhRqUa71c5REj1TrLasP5ouhVc+paQU+8OfPQ8b2uw
3MgT+0jwPwxqv3QomYKyev7D2padkd6yoMu+pMbUNcfIE05ZqbRZGr3/1Y7QjBzJK8u17OLqbjUm
gBjkaoyczhwND/n9dCR/dupw/de5XHjg+X7PtjDRU7DBmHU7OvSgkPAaFa4JUWlorPXWLaZKUIH4
KLkHsJzI05rrfZ4Ks5v1ay6oKP9LpxVKL6s5KF6+9KDqljtaH/DN4FDqStpTSlFenImgn06heq3G
Dd8HMp+hX18t/Nn4CD3wRLYwzjKYpxNrVoVN5Y+T090RBb64v64Ctd96isVE1LyU7m+E4DKJpSl9
9Wy5DLqfEqhuvkDTHyoGa4r2BAuORRdcrRWRbcq2RXsLCLUt3nOL/N3lTWJPPdol1+sAOhUq4Z9B
CT8uo0+pucNfNIM1dsYzAldILdl08G3TkOISxJw7JsMiMfr+kFgWYkGNbCQybugIGlSMJ3x3+zSL
9V3mf8pfZP49/cPlF04v3fUxXPnjeiZ+73FbT0eSGZkGNAY+Awi8+1YdALMRoM0TGtacbTCzC5jC
BOGnOtvDFmUovdxmRnTn2o3ELuO6PGoMjxlN59UZWVvMoZsSe97+zhS1qd3b054TTqVnTMixg5ic
YvBzcScyAAU1Cxu+B1XH0PMuf+rY1iS+c4iKZN0jEKylhkdAdXmKwXBnlPiQTT1mbhlTwnP4ZzAp
KyLT6tvBOH2lmy+u6KjS6c8WDydBVLgPLUbKOao79wtMTFx5TUsBGl4/rzeUSwsWZcUIoQzUccpB
bhWGU5FODwBa6ACcfY3xirISkegJdzXrzvroW48UFD+reYGEUY50uEpvxWONtkXA0dSBzxhmj0bV
Qr9UymKIDWwzcYckuCD24qPr8UCJRK/I0GR+9cBHyaeUqSEa8J5WU7nNRZQ+fNKIEabtkZqtWwZs
ndUaalWjaC3qB6nEWH/364fjgIRF4duFFbjaRTBYycFWR5qcZQbIoVQCT2p5x8uIaf0ZxiXapxVI
eo5gASHCvVefelJKbNiPh+303pTmqnoNCLqIOb+NXzsu4VCHMfGw30+IyM1LsSUDCV92cBHv+/TJ
95lI9LbEPNv6s+JsqI0VlRQSchvaU87uc/wa0wRDFPs+oFMBD7WVks7P/looOUwzwowLQkyygVN+
jHUKiEsnm7AquvLqNNjTqJl4K70MZ1Jp1FH/Amb+uVrNc23xHwojKNbbcklNnbgmgTBFBJexnOIT
/tB4LxS7i+YTz86c6SxHRHW2itn3caQ3bgSlQq5PJE2yN20qVDapbXQ+eqK/r7IFjjQeevJRIRaG
aFy5ps36r0lK4lqDSeAnd/0fe1CeZh/BwY3Bvrr+1Smd3TZ2/7yqCEFiSzwAB4Kmrp6Hd1Qnmkpf
S9hWhz4c/A2W+jaiz+ai0GrLmhxmEMN5SQhELUmRKXHbdOLu92gyQkgqKx3mrrxV6Bmvq1g6/vAQ
7V1RSUVrwyH1kb6gB38OfmX5LN7UOT8fvi9OwFq8GVyW46vEEk7tZ54ReQFSa4468JYoZHe3fxu2
3ZFhOD606qhX/EbIEAsPTuBJMHXfUhR84jmq1Co5mAGDeTxCE/dmYfNx/1r2Iw2enU4P3QGaBphz
BOwgs9yB5/Q0bfxb3POoEZeqNsr9WRS4XwR4Ir86LsjHwm1Jv+WPBMboCWBteTZghygH4MFi7Mpb
TIPtAL0U4h4x12FPny0oTXFlL2JhsDmktrQvI6LHKJFw6ypgTi1kw+QcI4Kplzc2Rh/MerZwRfLj
kUNDwBFTVn43hwcoW/NCC1wVYbL9ZkihkANbxGCsvUttt/LqfhFPfPvb0nG6PH7Rlua7LrC2qgBx
idufJIiRCp4d5iZ2pq8t0Xoa6cnPOeJMoQ7KJnXw09vJrgOZoYNrV8Bw7/WFBVJvJhttZgdaJAYH
TGmY3Gzg/TG3JoFbbKT7krtgrXUoiNG7opWGEuXeczJ7pzV4g1PKbpyrYSAJlLv6sQ1+iProtea6
LI4Yz0bNBc0Oo8ER8bb2pYbgl1ihs69Babnu7nedAFBp1ExthvQfmhuskpf9O+BkoFHqzqNOMcXn
NlumSHwU0hpUewRP5ICUouENGy1H6Z5oEh83lMLONcuqZHTLhx8jkXmnoO1KP1jvJ1HDAHQmhDin
C0iGFI1UbjJVHGeeAx43RfzZdtRQafYHFNt3z97+imOMmiuD3bmlEafqIMKSNGPuH82RZvwvsTlo
1I+VBnWX9da2r5kgdOJE5eEhRssgsdO39TF3NUXCCE2Sl/qZcz1qxzPvpxucDR6rCIkAQoS+fSpd
mHjJqwgSSw1+cVfx6Ag4jDpMkggfTOd4ogkvqBhYp7NXoWKviw2CbJaO7P/dKVtn/fqej868/eW+
349FUXhPFxEVgMCmxUWtypM8YlhRZM9qGuRXZi3D8r6088pW6xr/UIq3GSwvSN1gdRRenVzuCoi3
4VRKZF+dv24jttCC8+1uvFHZyJD9hEstf42MtwCP3Vzy/UK44u0X05SyeakawNyJkhiS4RXha6Jj
WZNCUMKv0N4JPpchS/nl6FBFnBr/l/949FZXrffDcPiV5AYF4Ekof7KKyTE3NYmWo7SOtTCeloC0
Au63oFjoBA8K0xzIBUBTQ1ZlFkxukUB4rL8g4SloECpvCtbcHRyRatzauqBda4reoqnHopmvwCN7
Jp9vyPBUyrGdATk3Ol1Itoc7Bi1m+ecdoIe1DLgmBMk8xAba6D5sbeZqzYCboCadyxAdFAEocSC7
QMenr5FlP/pjSNk8W+Oy5gWjHzJJeqBiwafBOfkzYOnc2ulTyrwHAZQKrJ56pQdoeLkDnCoVGpCH
Ul9YAYOVTcTfxionuprhFphZprXj/pDD2GvidPBiAXRBvSiSylFM/WciCKhTfG8AFqHjGtD7Tf0G
zpBBle309UVvBI0NMueegZybLjv7p8iE6mbTQD3naAWe5NbAWBql8Kjnifp2Kkgz5ikqtbH3BgDJ
Dg4NF6ypOANkXnjJUF6ekwK7lxYw/mfZm3ZRp07G6fid71HrYRcTglO7yS7K4SGosTTL225zAQz9
jIoX6BO8FBAWnc1hg821VotAcSQ3xNqmn9uDh0nVQ2aXFN4zsRW0jKD4ySrQI5Zsd5IAi8KeGNBa
mx3+HkYErdJQwwFu7bnvGz+B/2Lo53i4WZQRDVRYtMIF04iXddVaXbHeRRVj/9eHHIzx0cy7LBxN
I66wYqgLXadRH0aQ/v8AWvtzHSCb70cN8I/NSI8GH95Hl77Pwhr4/HEMu/oEFjHrAVKCJGlS3zjo
pQRrC+/aMQ6rlCOn81yWbSx5k9GR7hXqtOqxq3U+OPipQbIij+nmYBmM/CsyqUiSdwz4Oygw3N8B
j5hCVzQ1+dZ5gbYjz8zswgtW2XFxz1h6+LLKiZGWFBtt4PT5OUkjoezvs10T6V9UQEzmALAqKLQp
XFGm71tIXQYcE0LzDOvXBxnJ0iwvqjIV48cXZD5lMVydsapEkpWszizsQT/6TP3zHNyB9MiVLPTj
5NklFtpJInVdfrmKcicKIWVKSrehqqvO78cknvzfgnzDD6oUvYhvqm1cEqGS5UXx9jlECVBnCVKk
qaPHL50P9vICv5vrbm7360e2EpZpSsE2OfWTFrlCl9pESXFvKOehnOe0e9BEbo6UtEwSMXb4D/JT
WehxX5HxCaFNJOIwMSD/vLm/dypm8v51iPjGd+aWotg5J2LXUkUzY4oQFGcmAi6C+D1NEzhIJqLg
75fKm3DjiRhiXbHF1cUs72fVdziM9jZhXCA8cNtbfao5BY8/4bNjLwYHCHNwtr8ilxeRRa6+jRO2
fxEtEHeU5Z2eSlqlXHL85V14dN7fSATTJf14OPbFRqWi8UL66MfXw/uIJYUEXovHODe/p5Wen/c9
OaYemQE16tqyeV+a0Xr9hFccsedc5268wG1V7D0BzIkD4M6QCn9aR08F+cE/wWWnMMIxoibsjpk6
e0sS6jXcD+PE/7eWSFUchZzLWnntq/oJi6bC6nmEtDauRrVZAE0wYezUjjILffo8YS18UpMN1j2A
dbc9+50nkqoJo6Ph/8JE+NezfVcd2ylJbzw5wnRcT4rCyXlcPfneERBu8ImViTLKyZ3mmH8qW/T7
XmSK94U2xLR1CDFNtHlEUXoHDFEHwdX24tODMNeNEdmcVffeME3eG4EJT8amtnGkcHzRKsMYeW0Z
iq/BbB/DV7++L+NETEw2uBcjAvNk9hex0hKIQxYCIiywLZQCsB54o90gmfggB5JocvxZSzK0+qp2
TVMX3m0JvrQgZiCwfNL6lkO0e16iQrWSSAf6aCp0SvsRUsAyZgpYnuIRu/XmkmwYPIIH6/Gvi+RE
M2HlSrxIhWjcABOyymy8KWAk0E6xjfwqIQ84sIpOADkK6uAqfGSX1jWq6NON54Pwdyuo8TuOuSVJ
OTxsclqfTNAJ/8gnWq4Gb3aNXO2kc8gocf09y5KQsqY2oDhQVeMe5o8G154UCOQUgli15iEPCLei
BA5IZ8kEUJj3qySYwOSDfkIAcbTMi0hAkFRIVm/Sngf8HhUaN8q4K8uQCzEmLGo9jt4KJmS0GAgI
gebJ8sv/qvXkQxbvIpqKTiZoNEroCJKh2Ht3MmCTtILG9Xkt+N085hvqin8CKWLC+/jGy2BtkOPM
RTH8w7F/U1LAIUCFUixvixEFWiWK3rKgiAngnQV3lMcohRbK2izN1nsZZzsVVLCPd8A7Bt8Vm9DV
ghL7lYtodbnhCba0TqUsQzUjK+vWctfwcRJteDqUV7qgbji5YtYMpBraEPRV89s44uPMAqSOi+6N
Ynrg7TE4koQrgAn2XD9D0NRI6VPPAoOwMdbj/PiRkhnbZu4H3vbL1SdxuE+iUUnxSuu7yRK1eS2g
dkoEIB/AigPMRvOH+nNzlsYmKY+HAgzTdQQAReU3+DHyzqDKe4dXTaP4Sz1/7LW4T1VcKTnecL0i
E+Q7CJcRwcg9yj3Z/iSK+0kyANMGh86aKGW0IWrOJJJQ/P2fuJBIWVQKiXKXXgXHWX4TbPmGkN2F
Ej9DwmxCPLLlhgoZIfMu4Ttd+4NyTHFt1qQ0Y5W1/FQ50KdUphnZACc0MszWn6QJ1lcT0h9YELlr
c3pum5+HXlzhvVBNtVTyXeNmk150K9LhnjM28W1I5QBhsA81kZgHfxmd7BuoNROXnkrP2Nl7dx06
TrP22Bwwzehsv1hkOVOuHobPd807unO32TW81D9xsERYdYTMGDMyyzm7YdE0aEhjBMukkGWa8ZbV
44NWviTDQ6D00sGfpKlNbaLjjJEgNzdm/UiqWlK1r/feZx4nExdpsLULdE28Rr1Y6ocu2UHhzb88
37n4tqRzok482ri/xvLixbNM/DX/5DxcCccXDtR59WkXzL1u98Sm491wMg7QfiE1Vt9Gs19+2t7y
ebi3UgQPpVLWCjTTvrAMjJlJq1wRwidJX9gyuHOh1x/S1YlJ8cY3EU1NSuRCf7TLFRyrLWQWJp5E
7MWVthW6jleYTdHKA2ixK0u+hhD5NsNuWDwqYWEF6ri7PLGqG6BMPLJ8gi0ZdfNV1TYtIDS+0FYF
Z/Gc+/PS7lnU0cFXSdDhs5amR7dA4KMRsk2yFK+UZcoh1Lcw0+h2fvdf+r7KSyU6M0Thbyg0kMJ1
Cpzfb4vGqAM1+IBFk0C5PHKSGN5DZ6WVDtxLXIp2vk5X3jK5TDx9c3JOR/LasWPOce+O3hnaPURB
BNaV6lF0S3/8/DQeWcvdhirtPlfkkeT+FKYzBgzY3ehqIhEgvpUSJUmtUkUxG2ohyhIT+jaB2s9G
rKY0epy3Q25uonzSpIwEttVR5EDotXJr9kPZTIAudHtlrmJwfbrQprvM17QpqhlinOHD5iBxxs0f
/3S29uwVoUkglixMvcrOZ4mOGwdiQDyQ8HkPJDOD6iSm5FeD26ItNbrgxP00AbAg/8iJusF2xrwz
ci4BaF0jSKrL6gxvzZHuG41X8/Mlnp/MYL9CxDEUB5NwvaRbysJgOC1Pxr9oYobmhu4yQuOEc+sZ
Mdt1CRRXVbPnGwXCBNw4vkoFykOD+UFdNHKyRZAPJiF82paVXN2Cr8RDr00EXs4mkb4elt7Gd6SD
iZuCWpyKO+ebZH/E6F4APbdATXBcAD/aXV/l6Q0YSpJiUa6DWDFVeldfjz4G2h2Hxd52M1AlKQbd
tilA61aPU0DfHKSOQAOARAvwo47GXAF0OXR1lFB5L8B1lTwCKLU5zUVOZtSKDt2U426JMaUHzMtO
ttg9MD022bjJHQDQD/5sCVhBGVmS7XOrCjylzQLcelbmWj3yXKAvyoka0+z2Rp1anLJ3WM/1fMhc
U6W5Z5Siu4bePpK9HGeu+s/ztTz/bapBl/IcXHmdXT16rsN9S17TgNGg/25+RXojI+cWHeQl6d5D
3+i2jo0NMXRLx2e1h5He2jz4bw4Q18XJvCsPGuGfcy7XmzgPYiaWia+jVhqMubfbzvHXHmlcN6gN
agASPll2S5f983calqaChGV6ZhzWQYCLwb5xrgDGCkDZMbO5/VJxSH62VD0s8GejUmso3Mfp0+UA
9g1VxECAVfFN8uQlZTnxQZNtN9hPEnZvfIdxeGQX2WTU43NomJ352p3j2hgX/ZDKsPItosLfozsM
fjpWjQe9cNCkzXDrqb9UJst2dB9Btdtpj4Hh5Q/i8ZPSIRJmd1zA2qYSHl6T3D/7NUe9U7CUfmxd
uqydnMdBZhtVPi//drqm6hdbWBypfi1mzhaXFj0cxhyIOrQUJPClrwE0Rj2UB/7/DGJL4TozEL5R
/z+6NtiO9lfsOFeqisdW3lzi5VEN0Bo7rqsoqU2JrZbcSuH9ua7zTg1JfwfLG3n8dtA8CA3HeNzr
JWuXoH/n97Um8mU/34z4FaVMQSDoauP+fCY7aV7tA3WxtsWn5oo4/CdqTOGifs9G3kZcEGA/ut84
j8XWLS5OBPqEzA6Qxw/FWzi1pMeuo1gm4vYIAuJ3xIsAk/a2LOtzB4jATGkWMZ9W0XksDcQD8jz/
mWikCWKpoiXIculAvNcr+W7hqQs+s4+bdW08RXe7o/+OuKzmWAyLcL/2U/2I9g93J0w/QQZ3N/eO
haAHFoOOh03sFAak1HKZ/ZRZZNlm7SwjU9H/kqBGmM7VVocKKPkR9WKPvGuVQQScBj5+Vg3RnOJT
bY4QvaBOClZOOGhy//p5Txm3LJfz35fY9ri5woluJF15XDg2dIIdkGj51zzWKoSQeS6S3nAn7YYU
9KQuhSnZIHsUtSPT8M5n9cCzF5csPOynFCKlTHIZxtTT3l5Q0H73pQrodDPejVuWsOupdA4PULMh
n/Qlkwe3/vObFCo7gP0kk/cHImDqm4OZLIceXg7s+aJHTCOtg09LK2mmW94Fm+2pMNG8xT/X1cSe
+tJjH3udjqFlS+yJdPfTshdfh4OgZa7nBvk1B7QNQG0Eupy1BCDhUhVGnpuZI/PtTjb/lw2nm0lI
kTDk8m8cVHcY3KbqDgdCWMNaA0WOPVDai9FnlGv0bnADftg9naS4Wn5hxValWRaqDlDiokfq0Rmj
6ABiGq00hRQ7cvG/imr037rJAfzQ2EJEI7QWoyYg131knr7KemysesZ4hso1bVOBXDKnMAH+0G3s
06ixxm4yPd+IkXBLq1el+4/O9hN4SIIqt1yixPL218pcxsvFW6f4bNFvNYQERbroivfxOuVi2Uq7
wR9Ei8w79a4cFGFtitS3T8S8ssfTdQB86fhJFrpGSfBqhEv7KSoN6SxTnjpZy0PqTsaFIfTCo1z6
YrgyXukyiBlG26/svMK+K7rWz0MjAZNDkOyVmuDFTRR6v1/cXdWvWkig5DJtoMGGAZ92aJI8wE5W
7M0RRVq2SIl0HhUWg7oqDVtDaGFNW7N69GHkmwSjAaGeg1yQsZosTpFfdvqd7QBu2t0Wmtx1QPab
iluLSYresnrL/QDjeLgShVAgEptFsGZxkcyehKNqlLkoJDqwLxXxjxCXUu0R5v85iNeyhnTzNIH3
zO+mDV9NmyNfZoH8uKPqwVVBsw5y6c/q5JkoEwN3c5rtxyJ+brQw45Da8M+QzbuOe6iFC4+PqtuS
yQAoOGGW9Y8vg5qT42pv8bQ5iLc/BW3XFxuLy4c6uubPz1MjwVTe+uo/nWezM9RMnNbw/EnFYTan
MfAHNqYGHounG6AQj3FJuZ4XMc/V+Lc1HvLHvPOosjiQsaRwDg+i1efgBtuAK2H5bLON2JUohD8Z
qFVP6G6DZ9Q9aJlklQTwF3de5OuGIrGK7APdow5PsZFOs5xs16Ee2xTb9stnKNbDb7TRMiDNAhOv
J/mvtBfq+6f7DZNb+7PE6tPbHBBHKeohHiKYfjon9AUmedu7ukkahveP4ScDqYhLBVTlKBDJ7Jwo
GzC7A9Cvy91duddtrcvm8eRLvcEF0LifWYuIunM8XLaNYyQv/TQxK7gEhyguG6my52si7OYAiJem
3yyE0ln/z7h7nN5okapqicMNT2qEq8sZwzIYIOhzkQ1Ef0lqwnnQBgPfkwJU+e/61OBEm+kISAGs
EY1JA2sPTm/wPpwRfNADXDCw7c8z1csMvrZ2YEItPWeuUId+fw4+knEjNR7kQBwWu2LehYZ7yUrk
HgwN95y+/SbjTfOII0zKwOe64GKc7w/XOTvyGpO1eUlZjp6LJrrfqyycRXgo5h1bi61T6Npduk79
6FeMLjgn2OoLgwPLEwuQCmi0znMjitp41eRjoLNVQr3Awo3CDZ7/vhMmJEoUWAgpcR5Ll8Wm0JxV
l0gRxVaMsIi9/nH67C33f7n91bAVRJ1pVt8IluILQ2xX8xpbUx6A8S5I2vWjo13If0nfTNhQg0OD
KWY0WKIsIHFPGbUQ9GPFhVJQXOSPvnP56NVjbGJz7v4WrssCwMJeY+euFLqD4926PL9spRd3Cp9/
BcdyiyVoBcbevwENKwjABY38OZugtewNHv+geggJlHgeOzZhJ0SomM7iZuRFCXPytv609W1xo5J4
aWNSfo9xc68/WWYEbOsstXOblKPKHx1L2+RmsNcPQCskSAI0UlAgIv27Q6vRw11wQnR5m44odPuH
H3VuBMoRzErrFxZshY4ZNlEzXw1J6rdDHre/xakF81PoRyOLoKlUVGEIW5E7SDvYUdIOYxhyDBPu
x17jl8TnQ38XPFIHjnU3Xy3z+s2neZsG9AUiQ49BmNgX5lkYCnxrjVpL6vlOKd6tYzp1CdCxZg2d
QpcBUlBCFUedZFxnJV07VNDQUZ7c0wR0tRbvkkpK0II0IsBtt1uQR96lE0qY/LxF1Nzm818p9kVi
84tc9tmvo7NAmyNvt1SOTHlGq3P3em5XyWp2BxHsBU/+8koI3/om3gNUwnhjQx0Z8tWoBdVGtz+7
NKaSbPqKStJwI9TTtKCeZspNFvnLTsxSi+C7iucm5EgbtziPkVKg81u+iLwS+pRYrqYXrtFW0HDc
mZ1rCHg9zFaseDYPPPGLBG86IusAfbgU9me7YPhQXoblfuqEgcQOCVBhNv8Gd6LHpI+zsOyDkisu
9nz/gcvFW6yjE7lzddRJllwNF9nATB0g7qiPGozTiIsYQjk2wM/A/ktUJ6G+YkBlO6pQZg/4+U3B
AjNHPUZYj50Weep54PhIFkKWOEDShHAGfip3XvnA3C7Ux8KnnWkHCuo2yrPxH/Ozzxs6fWdLTO0H
67zjFJ1c2XVpZCRf6L/Vohya7XDv9P6kh4OwMHe6li/MYg0RBQQKQjW4u8q2RbylO5hvVpXmylS9
bDsLBxSl9ASJlyaMJQj7Iggi98jQQRLswah0E884lo81sEAR2AXId+EpTTUBHZy9bTM+ipG/q5uI
NsdAm5hzKNkZpUwHCw68BgXel1eKK4aqvrWWjA2HoHx+mVMsgu4i+gKtdHGAFHzOKOcdhw1zxNXI
RMJKKZs8pxVRQVU81q2JIIc1i/rrLYie6WFNXdQAq6qnoCjCmN6STXJWJ0OX9F2I3DJTbgZOgx2p
GSlSXzgynrNOGIigIw5PEFcDKI9VLRcCGZKIpSIOIT3tDAFHG0FME86q6NslcxqLFzbqG4Zloo3N
yLPX9bRmbesAfZiBQczOQvoKK6eFpxdV7ozqA06PMJtpQrcEQaFL9QkrYmiAj0gIOcdfBjGecj52
Fbky8ojzy8G6UejvsIOk/IVgUym5kNhcnCO8lbfUTFNk3W7VobyyD+OCL37CcqCA69gTAtbTMJf0
RQMTzfZkA+uNNXM5Vwuht516C67Fxv29JtB5+su+KTjfa651Tr8QBfzBEN5ibYQFHejkMsy6E8xf
O2thAt3THADwHWJVNxgcZRUHBE4rrVMvRp0dVzQJPtSgg5SbGaUmnAztCZnQQNflyWq0K7/Cnjna
1gmTPZjTje4kkD44DvoC6HxUQQrgEj96PcHSPK+A6twTckj7m2F3KiqGce5wwpkZYM1w+zUPVhjd
615YncLbiw7lN3e9hDfbkhN//cbaiGvGAJRTTA0hNW6KkmrcaPEIK9nxBxsrruYzcmOFhuMMe6L+
GbRmKiTTqBWWVGiN4hmIs6EPOxN3UrX4UpZIpb9Qa+k+NvvMHFvgkoPkwv21fSLUubJWmB/UxHtJ
sm4HenUxjVdZJzzhHFUsW7s+exqOSTGf/uaWkbZXVOPujMUdUMyBug2UuBhGWErXVOQzZEJJgI9X
zPV6S1pdPA2LRqCptzGUlnOs+Sw9lTjfFN4pjZvx+3Bkbton2SBGpITlusFF54aKQCvjnnqo+Fsx
MdGwlOP9iQD1FNsTzKfp24BgxXSF02KGO/3Xlc1+n9xn0YRacK/QBtncfP7K5yxZdmJmPDEDNI+4
Sv8Ouez9wVl+n6G7GUUfbu260FcaXDDlXz4tzxndCoTdHAAcepFrXjF11GxN1EaqNjHNSOBC5bhW
wunXrDKnrwB+SGsxedHgj4gbW6WpBPszY6rvbu29hPP7tPTKSA+6Fqof2pgw7Da2mBvQu35MDdUn
qaa97V7wKG+silyG02LS6PgypSkrn1DhtMKlDqJH+yw/DYKoSNY640KE2bbwy1cRb+W97TFjZgCK
F92b+YbfCBHNzxsAyseFUpCuOGEEi+9JNIquqCN+Evg/6ciHzebcJk+ZusykIIfMorrMTo4x9JdP
WprNH1MRmjcASBejJp1JI+3aUpJ8dbRZzC9jDZ3NIgMtPSU1+Yb0CbYyQAB1q2Y8lM4pwsSmKH/k
h4IPhpyUPr+IJpjjMW89eHqN3qOLEVAynZ8wb68hn5NDNzpVVqyUA+22LuwWE3PbOACo+qb8sz3/
0cuC34rj2aFm0Aw028Se2g9h9jdVVDcHhbOItDkKO+Yeao02eEOmE9W0q9QiSF4cu1Fc2Pv9FDR2
pCe5Qj7oL6U1/CTCelGHwtM5HTHqGge2jm9tODsYwR+wYECDGV932+EJ63ihWcdx1oyLcZ527blp
xa5MQ3bwgEYepX2YLIpAmlQNv5B7dfL8PlHU0oq9XRkXQxO66/2kf/1qWfR8duokjdM8MN63aMo0
seATDeQueWMHS8C+ewUIB6IcmOOMp7djIYW/xbkTEsE7YHLX/wAcf1GqqKiH9KFSkv+L8x9bE7iB
hvKmgNmXpNKdQaXD1LTX5qe5U8nC1E7gEjqlfHhdy7pyEfE2ZqOw3sCYABiQsjPPU2EbQYnCfxUx
rNWTFk7S94SnITci1zH/+tG6AEpmqu+IvejQauqnEXfR9uKmhvdK5l5DGP8PAQo3rX+3zfUlD8mb
YIUa6up2pUKFuAaxYzlcsXmvmx19H3UZxAGnSGSnloFhuhuedhwGJOgE0LmM6APSnjL+HghpDO7m
b6V9GoXyLR0R1gvl49vjW02ERYGwwT/7+jAsd+jeP/cqpQrXdXJDJZ4vsM0RqunbQTjcwTCtLUYv
LtGWAmVZ1xiBNvV8/oVpeKXJFNKFPSzOivbzzcX9y9AvtaSXtHl4kRT+wtGgkQMHrOD11ZO1aCJl
MyEyJh+k3jvr4Zj9jfi/I9S/xgDDfwMqXIPFzvPv+9deIfham8IDUnk/e7ulhvZ5tKGfgOWwUdak
aczH/v2z9IJUeWrVbbAgEWEsnj3XiDuj4IGebbw5axGJXmbR7ty8MJ1XGkTceWGyjegSCags0fu9
30k0N0Pg13Wbq00jE4SAxySO4XrP6C7VQ9ne+Sj+FlmgQCp2lbDx38EOnSixAVYcncN2yzdiD+sj
VAIr58rV8Kj9jnATk1MLMAX2DO2HRqwejFiMR5cETBP6okDU5+Ql4XNB2K/EMexLBdNABM6o4g7x
wNDt7BrZXEWJNVNWb+MndpEVA66ZJcfuLgI97BpeGpJnnAxSfUDxeRyAfpopw7GM5mVoEabUb3A5
Zay/VXapBPUclM0Ir0WnXv3nhVEwEtGTyA9Yemb+pk2YaXNqXuHi/9DfgE8wIxMPrbMkZ0TNw6YX
Rov9Xe3FEk79M+CNFcBNTn7ri6xN3ybJbFQDpky/1jr0pV9Ih5p8w/XCuS+lEZefUQ1mp3oIe55/
6aXWRCItVMjQQUCatcQ3oKTZLh7xGPc1GqL+A97PN1VNWQoUfrIa2TJ0JPza3TVH8ht1O5SriI32
Mqc3JMdwfAri6a1OIgin6iTk/Gnh/0/ZRubR+OftTpskmz9NMZmBQlZKzp6gxn6KlJxxFIBZTcGy
/W8kxBBNN10Fll0r2m1Pym0n83+AYVnu2xRgtP6h5RKVq2j2eQXkmMtf2s2Jb6fz8V0Y/lu8hf9Q
dIxZ5QGTpCcmojIgsfZTDL4r6LMKNaUoRD4pGqB/OkFqdimF4CDnSCinL5XeuSX45kPYYdbVO9SG
AevkmB66bt7fTu9naFqQKec86m0mBvDEa3L9IQijJuZKEY6R7k2x+HdxGL//sxR65kTbSsOS2beg
aM8nz+W/si/YlgGjnOa3lWyjg2uY+l4fNeNGwvHA5rgvGR5jeG4cEeVRjAJdRoM5nvQCV+XChnuD
u7gUbrrxM9KZCjLt9GCyPvyekoxj1easfLFFSwaM7hRhwWIL0fiTTGkmB5QRfvI6CYNBHeXRcWXI
FXNuRd3qa8BwS8H/+x1DYZJSIgCOX6j0KeuZxngEDa2dyphoSHUB4rCfDsxhqIGGb3uvGM3JR+JS
HylBf3PfnurQDG3s2E/yEwUiAVp9Q4ykrf/GK7SmIorOzvtWhghPFHjBdQBowqQ06QMhGmCUlUXa
UhB5Z6RzhCpKy0cDBxMj5uEwNzOX631Yt/wnn+nV0J+4LD+tYOPye6ku1QsTmu/Oja0GupkLvzMh
LTEuLq0QCs9nv9dSy10ANCP9+J8wGIy9Mzin5sjdGj4+brl/HeK7a4iGosZcCgr9PScrqmWf2Ie9
xQ8zqwr9LP3bWcYKyhXXkE/USTKzSGu/ThiP2kNR70r9QMXFqqEqWlc2X/GJUrfBMLW29wY/vVuR
bIU42YWwK6VHIXv7HL67N3Pgd8kJHollLoaRimelbjVXUZhE+KaN2KJggRjyz0VJs1CTtrhRamrE
4KDyRD36hS7VKwxQEpi5xFDMtA//4hHlE9OuTB9xj5w0LXIrOsJ5h8AvHA41/Un+XUGn9TtFFiTR
Zw6YMs4bJPJyXeKEgIY/+hmakNcN7SU+Z1fF767g8vx8oy9zEto/zisx+uCDWwXljUG4AbXWDrZe
nTSHynFuztp26mVmR2MuMz49LZfgKoYbAGU/nmSfuGv2RYZmLq2FCyzTZbVzMCXH/qraXDTWRhDd
u/kAnhfFsdeF9aLo2YUMu8WBS6gmT2T9I31wZRYY9xUKAay34nVuVP039CfWzHUOUazavhlE0v27
ddWJr8c+SrYaizO9U/66nAgGXzT5wWn+jo7/W2AVHESypbRYbXfHjGUh36VQmRqTdya35S0mDRqA
Hu2s8q359QEQ/BzlCLIAE/JL7XNUXv9NSQBy02L/5SJZNcN79ellFkpCJ0G5v6pRIR9/tg0w7OYn
zDuKyGQh3ySX/hKlZ1IoY83AYAgn7haiZ4QSNlWmyrcLiO8WjOlPgL254IyWSWOUOrS5gEpn87dV
JXwbYoI4bq8zX26W+MBUV0DiTxH9z70gVbpx2wQt/MRlJp1Q7edWc20JdBWbk0R77gHiSngTWBTc
z+6P3AKf41GkmLsO+Xj47ToBCjqiI5kaGIdSLbYHy7tBpVBKFKqwlYXYHCN61uhl9VmU4B6rMSiW
sIUnDhimw5JgLaxsYNIBA3pHovsyYv0ATWtnxMfndSo7o1K/EKCtIEo/PDwYg2yL0G33PrXtOcu1
GKjq05cu4TCsJ7rlkCA+DgCO6fsdhZmm1EOdaOdPOuT/6ZVX1vQpB19hXjZuja2IVpvl1uwewL+e
+jN6Jv86yzs9K9Yx0PQpYxaEVb0PuQnhcJi8ZX2PUv4NYksU8r9TV9uEmgBhuwmf/16zn3RVXEYo
1svf0ySXM0q/K4O6FmC9l/WoW34ZMbZEckZxAown7Q5egP9QhwtIaCGfXcgHCnN4OM6TTisCMlmg
r2l9tiKU5c7XID4QC7ZxHTB3TPtKGcUulassp3C+u76Raxg67sPRk/ts2mGUcXasry74jyp9odgT
Hg8aQ75ILrnY6nT7ZyPFq0tb6Rg9LpBn2iA7jLxGv8fpQWJhHxORAB7DnL0YIT8Qgsn03UHKvEQu
4gUKIYGBeJE2np5kAf1iZHS5dHVX1bSjKgG5+Kg44gA8JeaaLuBF9KR6GnWYmSdut/uEouEdprc2
tXzznVc3UhVwuu+qT+NdmBVJIh5I8qa2tClDF6d39v2/Hrc0/uXQpK88hm9wDK/pIUYn8ZGqwtlE
TPpH3xNIB7EnYeFyc9TSd2AO/UThwi0KilyJOHf5/SZ693viEgAXAiFBP20G9QKaU8W565ADyu3Z
PxlN3fmPEyJtdHock7yr+pcbjOI/O+P3rrBE0KrFeJUEb4V5q5Tc6MWCJX1OllORbl18Lb5ONJVW
vh1V7qF5Z39XMAol34HPA30M9rgkZKMSQP199tCQxftX2dI5UttT8ESW9MOhelVy++5nsqvFf7u0
/a7QIMcSbdLbYAke/qUe/fnat28Vg8/9NdF3GYy33DZS95buzzIe9lmuSboR3rPSddO0YLbZc5aH
btUqWUnXPi9tpeuMhtwG6hebFXYqbixYSTbwUhXZK3ScDZfy+FQble+Qrx7wy0/iJZkJiQDUnPwH
XQjQIjwpIyujWlPyIsufihf2ljv4k7xqAc0MdjTook3D+JQSZEffAXVlSnxgVCUK0C9t9xMFc3Na
r4J1rjySlHQonXP49WrIoyEAn5otI5zxTrlzX0RIY5xIOZuqD6f3hco/UQaODx8jaOdLMCoxnwpQ
xrnpk8RoOecJzggmgkWVBo0uxVTt3f2t3dkAQw2WyL6mdqeAxvkcEbLqKEYZJp7gJad0x9c59Sct
VPrYQP+2LMSjv5R6s+YBwOrYSSWWN1D3l5bTUBwNbTFAjRrMk6vwqSAWNmWOtyqX44gR0sxlL4v3
acv0JblDG4Jg/xDmLPTXlI6HYRH3giPXsMQZEchmuWSrI/o3tkyPAKR0gZtZG2fr+Pb/l+wAWQAC
4/1B/PWRGvwWjoD/VuiVmhZWk+8TjcLYWiYfeACO98NszAcPq1VOkyfohrOoI7dyvBZp04WIf1gp
MFIz3SDyjKsdl7FnlHgNt4CkMBCiNyBgsCesM36Cjlo6H1r2eQr0/L5d1aHMX4ZN9QY4+xwis8YK
SQPvmN97c/GEFPNTR5duxTYihtSWYbgjHfX4EBzUy6hPm4T6E0cDrQutOrRocSAZUhT9dWd8ggOS
yqs9c2E6ZWgTAzFy3vIfgdPH3JwE/wEMca+HZSekpbMNiFgUidRgSO5+aHUmefkxv1bkoYrj2V1W
kJhSbTwvPrtbdFLi+wzWPaR6XugmAXREP+ghsaJhOsblqNoCAk9+rnX7qy9Jz1uBAjBGOyMn7SI1
62qvBt10t2Q2awE36Qe+/mYoSkjtIVGdX/ZwUVU3sBtJD+3vYlrCrHxmLoD3sfdkVcu987aNkiyx
AjwgEAV4frlqZlaJEbBn8C5Tur9xgE99eVOhzNoAApLukO4vfhkmWF4w6D1XzDFmKi9iks8aEQxn
PK9wucIrbOMmXzNnOJY2tIylMdrTuEyPcSPTMwm6PXB48j/PUgiS6+k1WlUs+QuwobHWYwxXL06N
X/Yczo91RxcXKj5xK7Gp8X3tTnVaXP7OQZB555gx7i28wgs4n6C7TRaF/UGx6x2/JFqfMCFg6OOK
x1XJTQV9YHxlrsq4FjHqkxBoHpjhuHn+OVdzZKzoacDnWtsMpQbHsZFdVSl2d83QF7sZxbwm4JCN
oaAwkdeiNKs7T0nJXTs+hC45evCWdrzCI7+CqUH5vNzGcecP5oWBFQM7v8BTwIZ/0/BFwUCb53qA
Fv4IaYPXhHekfKnFkvlS+0Ld5XhB1DCBzLe6c21Mppo+H7SGCuZlyJ3m8vfWu0yhxLUVYahEn2/o
ATJ4xfBOUuQ0epJM+zcip9CLpEJT7ESlt6PPA32kylMFXBV/3cDHIuxqr4QSCXFmStQZ8v9F1a0f
bhFz7eI2HvehGdtOfv40au42CUL7z7nQwe4ePwusXTyWqXHq5ojYGnjN0l7RNYKadsYkXcgHbWF5
yYfqTXc2y4sqARlAY/gXRxfomuvyuWxVxnr5JZ+BI4hnajgS0pD3dcwTVFTfRkRmWkOcwAeIi3bk
HlQ8JYQ0LKHY4V9cfA/8GDV+7DAW4m2eqyxrVEXq7/lcQyAK/Qae6YXblmikHXbVmbzICu54RnJg
IOHA8YuuDRTTHisSwSxsUH+2iVHt02xDL8X/XRzEd48tqVzGY0SGW4/V9YF3/ode7JxQjGLn4V65
UCO/HWhfpX51cwjtro4IORUy6SAJaMPYX/dGCG3CR9wbjuYvgRyqhf2sVnokZZ57Lzm/T6snU8To
w8brSSkd/sP9XnCMydrQT4PrPHTH4WRx1+RL/XFr6zQLrXD0AoQXNBNR/UE/8RH0Kgvq1GvGmiNg
sQh08HvrCT7BYG4tho7hikjIpFvGLGyA08wGz3BsMxjfmTLO3NDBvQY04IaxD1X18xfl1FBW++8b
akpY7SDVYq5Qdvmz3kW2pg73BKGCE2gGVCdiRkmoLV5CsjaDI2k+qe98fTL4Hny/+JP07IRFX33v
4dLbOCABqjZIjlB+ldQ5sva/a3N+vvBIVH6I1aXEFNyjGkulJJY1MLzhKToOrWS5nN90Q5rHXftH
KZiv//QuNQuX2wm5ivCsULesinxvQLEk/43AIi9bF83s0d9R9sBiNFocbqrIeA2RmP7CGLWZr/aK
jkMAa/0y+SMzZ+XJKvTPgUv7DyD4mDzUCg4LyO8QYA0uX05cyx7EZ8xSljH9PLFxmYWAgEWaMFXh
6sldVFwCBaJGgh8Vo/ZwHV4cg26CHQQC6jBhnx17Gb/tm8/BMyp8tL2TBvnqIQEC56FOA0V30v8T
pK3ugRQlCx0npeyzP5Lxg9e/86kN0q0b/0q4mG1egzD53LHU40oORJJVhtp8RTYG8mCXSv/Xx9hF
EU0vTqCzW6tiLIeX+RoDuVRz0mYt4te4LGNyK89djuYnJrG7KO9GVe1w+gpWsYFxPnmMbgPUOHic
jU9RCyqSHAaQ3aB+zsPUJQ3JFFcTDCrbh2uScTNG6subhp01DeE/xYVmUU3QHGnwoyZ+/G9Q3ZKT
QaXSlXD/0zPtdq+JwUHkxg0HTQQSd6HX8Z6cROkpQ5toX+KX06skTog6dAkJ6rVM4NPKxHHdO5nm
podETucOVU3WL2kRzr40ODJQiy7s7yiyIjwaewzxLCCesD7RaCRNfHHzWt3TMhbnA1AlLNp/1K73
MmjS4ScU9dc7pJojaxeRkYlv0jUwtWtGJki30m5MKVJGxIZo7vhs/KtOucGqR89zQshH6mMNf59A
PBzgI57qs/EmSfgN4xqQk/ft61PBAcQ2qD2N7bd053gwqnHS89sz4Ot1iUBsBFfWFJkNBaS4g4sJ
7iU4dgaP+8lVW2FdAx5ak0OBOmXkRIS51AYyNRFDkSZzWDMjwViUNv9kFlC30ttRqeQESWVMUzhI
zhnm4ClREGlZlJ5iovF60wwdcqicBYh7F6mnKIBJhCh57qea9mnu9w3wmD/FJLSLXH0uts3wW9ZX
0WxImYYKsQEOQy8ovqkkHGoqQhYHO9C1HyWbD+ceW3A/m20iOFb9UQwmix9g1nuAew1IpyZC8xXX
ihwbbtwXUlqzr5chj5kGhDqXSJO44Z65eL6Ixhdp14VKq7lsmNBXPkE0hIWV7M/g8tmIhbDHYDfP
hyVCngKnRwawMcsoKD7fgiYavYh+ltYBfGf7P06GHsdQ0MdR0VtMlU5RPK639/kzdjZCjrEape/w
ZLyqhHpdt1sWrbljo+2WNhzDj+gwhC2C9/A9A1pP70b4w8VT5YmftBxhHqK4OaFQi2itErBpPJ5c
XQy9XaZy+mi19PjHWk70idfE4bsybenBMOjZScbpKLyUT4VMnGWnRWTRnAfMMiLNMKpxKEqNJ+Br
YCfDKPao18vMWLCFEjonJd/HwNVAbjQ13Q2wEctJxvbnPNdnPJnJiHbL2JsSoVxpR6Hlapi1CKma
xDMabqi2900DG51QtxxYSXKt9W+ejiuuSUv2i7HGTL+fDTiG86+4QDoxK+1fTAzLNNIj1HuNgAe0
C6kx1VXA2ym9EDseF64cbDuo0GvJpQQcTKwVmzi3bBcvoqVU4ftigIJUtr6mjLBhaa3suznncxWb
yMYLpY00N/qU0TDArUuMlUVTCHUFkcWGX+FkFqS/6gFBMf/hj51fIFZCBqVzJ0hcWlT7Msc38Ctn
2Af4w05TkPuR+tE6FFhrtGeCK7zyvJwf0QxGSrpTBJdCUpzaQLJr6v2egch/QABpQkyNbksXr7aF
HrvJt+NShzP0vQlcXL6p1nkqsJC3RMaQyvnT3qgpS8jy8CwdILpfY1U3alASIlvyGGMpnZ+TbkD6
nxx5Ey1hbUivpKPogqhkq3Lzk8o77FXdnBgQYm/5H8giNxBQwLBxqrJptN8Ddzgn6gJpooI0Tfv4
aZaaj2oCaGiQEksD1XIAHg2g7PfDu1RSFfOWo1EdP8ZwpTJPaJzwvSeW66OcxvTgrzqR0o7SIscz
AK2dowGXOvKEkQf/RZ1ZF28IvH0J2K/HrdNqVXQvUAxyTgYWhBpLUdnJdnd/O3sPHda7+GAP83Rt
LQHRxpsFFVSP8tKvY5WKijao4/gdPXpBcvB5Jql9GcybJ88UkZXj2jxjUhj7DIYD1kLlAWP8aiYa
frz82TSREqOf5++AqvnvfZ1O+cHqPnESSo7PSPrBMKIEiEnD4GhNbsa77zFN3sCecDK598ferLUk
yDygAqrSgWLJwWqc9Y9QUjSCpkqxnSgEsxz2DDrhZX/VMmiMj+vrM1QN+d9x2W4UGP+uxtH2cy4h
XisLMEMXPYs9pt5/RbMgxP5CMqmUdHgrNMnrtQMEYkNVPW1xUGgo4GujW66xDBjyQBIvR1US+tDC
B9G0gkxxpAhfTwvDa+PEzsh8VYQVc91elbEKfr8swA7WZ8o3bMmuvHCMayzrqW1alD4QLM5hMWTn
B9x0bTGBZ1nZUoYuZqisgYsasADTN0FfJTBa1dJ9jb5q8YE4Ixj462HlQ9gaTOBrLTLqm3VxnIY+
kg1zDAuNHbbquN7vVBG6J0Fa9rJQ/CSzEyK0NPa1kUDSwdXHsf5bW2te/kVf7XbJpKKTKqHK83nZ
aP/rcGhwn7dWK2WzkfoJYUx6G9p0sGo8mc7KVsbtHMsCH1UFSBXiYWahkH5y0nxSQ/jkf6SMG241
NhHnaxZdukAq+P1MpsMcQ5/diNgw/DvvF4FZfPY3iknLkv74VMAPvILrqZD5JKm9wjfA5CFOcdnk
91y2HLUNQ/noXoXZLJcJxgwUahmTZGRCW5ZR+qUZly0aOHhTVKNmmP47vCZQq3gv5HZTQokfFrH6
3gd/oHoPB3TnOzSuV/d57kBwLZc/AhLzxdJ7+RRRJBycmgZHCypz8FE8LGnyERiDOPs3ISBqqdvo
ABoIuNb4xEJPrYibyyGV9wfhCNumXvsf9554E2flQvSiy48XGmn2V6g253iWp0AcD0+oI90/HqE8
yUIeeiOFtatqdZk2XIixXZHQCrPGzaYBki7LA0AkT9NB+xJae3w+CAA+mmjFIO6CLABOqcoC5xrg
x/Tq97MXd5YIdi97fNAxW7Espdgamvz3wXz4NY5K3OyHx1BFj0FWA0xX571i+sPa62eCNN19ypWQ
I/W0EJo8CQIRcFLtw4+ieP7mv7HJ0KeHZL0jy1Gu2Erb/Wf+k6Ge2M+kM28gwKveun4Xsp7B1s+0
oBREaJ5bF23Mr8A9x85gmrHT6orLiEDwdH/j3MJKDlWtHVgkROj/WqaIPqgNT54sEuxVfdiArHaD
SM7UGQnMtakYP9/TqRzAw5Fa7Qu+g1u552Czl6XjuWDf5u9UBIf0urTAiiBdfXtWC2+Ywk/XlHgR
DUvedgcLzMstB42J8QXHX6u5Rl5KnGhwZgxgW2qDtcUuBNPes1lrO0lMXvbujtxU7MEkI3ngGSJJ
Tr1aGbQFJXasFZtI56n/Hb5T9AnLzT7x9zvl3vzY0aletk4ae84MDYhi4/tKXrpy7KKL2YpMgQ5+
wUV1vvs7iTOLSi97Pj4xTOJnnURL52gIl9mzzDQ3oOEvfLRnJFJd2kDWjpn2te1dhRPLxI1QpC+F
zM3CK/tUnVCdrV02zYwl9YeCenEPAgo0Pw/knolssMyH+nH71LPvjUCX4EFGREy0amsuIdneTJa/
Xnucm1ejV+CzFaHA8zmcHX2CsCVqZGyE42ilYTz5fPsQBTfgMRo/HOWAEI/dSX7ZC6N19CZCsqHV
QWfFN3K5cz9KTv9oKhGNC3zn3ly8yrYXUkImIWs8z4ui9Kmzu7cL3Fn00qryIfQ8OYfNtqfCRQuB
DuR3hBKKV7NatIx0SAgvjzpId16C81BPqjMvhkpyvKkwp+BmO2WyXRkxpkBGJf/1rv1l9EBdACyl
iww5ls52fY5R9v/ARanB4AaMsHcyM/wqjTnu+gMeK98D/8ivqv71AojckGHcG2mPi/x6dVxOHOZy
BguGEm0kcQJc2Em8gsP+LtaCRzkcMcjMRxpwt0HQOxyaOfV9Ii2KLIS8c4uxkgJCHD0VrViGKSQ5
uPY+fiuDlB2nXeP5/IRWampc7AOjocTLrEf+xUXdzcBxvu5PZ8P1gvFX+Oy8HFVMZ2pTVzxvhrd3
qkgSoHAY+IveF/mrTHPSc1vxTjaK4OLNvETEKpSqQjAISh1a9BGrI9078aunhKHEuZEJ+NdjZTdw
UyPVeuw0m4IUhBTCYUJdZts6oNmVHFRAeA4r3QE1xvMbSpmPhafUHRF2bobwNolr8vWRr39YKTrn
wLBaLfrxopeXAbiOkMbKSoRzeHwE/bBLJs8CEOyW0Qz6JvAp6gr4bmFCyQBP0MGmFWeRVtRUPHPM
+CFVf9NCfCtdEOhzV4WGedq2rs4sUNAI+hCtkjJTA8+jCrsb+L4n5pbDsLkBQL3aQ8I0TCI0UZja
v0rfs2Q2QUN+3O+ALNtj3maEl90//L2+WKbbt9bREFxLGnpHJEn9BQIHDy7XNd9yQuq1bxxDQ1gW
Ee8nrHdLeEjS+ukQGhopZ+KWWrf0J1j9y7jdcGgrEmQaqT/y5+cTbpoexTaVkTuDO46idUx2V2Z1
xLZy9NfbOZ5dijK+Jh/kGQ2AV2C5v2yXIAZuBbDvkVD0XSiLcJmSgfpltIuDibmybQLK8ZDQZecP
iR68vwj/ML8CDeDDOfnNenOpFWbg+gdbJV25xemBRwsQyb8b9KM87WaXGGUr4pTziFDtcBVPODLq
IDbLpl9AvCIDhR/V/nqhQC0z3KE8onHfa7CadodNWPaJhGgERq/Z5CKtQ3sAblMx30i5nv1tSKzP
NYPdplYHL1UDSXxsNIc8LwCsmJqnRTcXy6O8Ysmc4pXJt8/3/xkSRleAq0Iy6w4+KYTn7DuBM9qt
n7pwVlhu2ZZ9O84izObykgu8Ws4NJeU2fF9aBkxer4yleNNGl20LcqiatW0GibvABIFlx3nDjae/
568vxyLDrG6e35iJKCBnpEow++DmVivb2gL0R1mn/UQ/pf4qu5liAHjQNP8paLeCqbhPZ5apWPMw
fv8Z7iluoOLknEbAOuX21iznTEPqf+TuBS4H0Rx6l9KB/sO9uVdbGRoTY8SqxMPCc3M9OVCMdW8M
g10u7QeeodAwif3bbzKwiZudQUDY0IREM0/jTafq58UInwhMWBAbXpYrHVq89ExV1hmkVk6hmLn8
jETlDEDPUqhY+hbHbSr17Wumc3+PhXvXvK56eG1BvDiSLeVhqH5tzdi5gZgXmURRfmYp8sceXRrH
3a+jfyQ/KMsbT8FEZ4sKcOL9VUgUGVSZ58K+aL4YVg4/2hZFd+7gW9Q0EIopnas4FnExYSSEucrh
yWWplC/GOiTv95JNG6FmKe8ERKVxRoufmUlWkYm+rZoF+qRiL2WscTMGYW+wd7lr04TvJnwCbvRj
s5jTv2+9QMTDRyyh1ZfLRHv8SudojqkOz2AI15HDv52VCe2Y3NqlZpczyCQENpJ+wXHRHyV5j2ei
v+fQUmgot3u8l9K7vGLsKEUjaNhlHKLClUCdfvVsl/OsUtERjdKlDAfa6TxWzCaWM7o1WbfAzLCH
23JJrn/8/CDKPuBUImRgC1xHbqEwihjKOPgw2Vm9Y4KfcbFuyOlPF9pu3/3p54FijO8NkTud9Y0L
sjuZ4ySmQo1DooH+CtIJ1lpCmsUEivgImoBZ92KOV2Wu/J9KwsH5VRHMoq5+Pvoslac7IZwEUwFQ
R+ous8xGc7g6AQ0E7iil9JfFGvsi0CxCZHiQDhZbqzNqprnpsw/S4yWvsMurNYV9LxPJ7c040ZJK
NxnRBV/Q8EEpQCOWELOpCRPm8xwdG/L3bqsYxk+Cza+bLViG+d7TaL7ILjzxGIP5T/1aJcDv0F+1
ARxeRYcUfuH28u4Rf3zrpbiCi+an27tAwruHLmifsGRzaKVmE8vsHCLFwQQVu7W8ijdyoYYP47jn
bwdWr3ynKCDhQsXB3Gjp719WHNei8zSG5B/Yvr3FUnfIsh+cbbLr2T0rb4jwHJgYnkBMQHvqG3A+
eaKy3hVi8rPoMvG8itYSxUhKgAzKpvNCQwSMUgSQpnw6iwZVpR9YPGl1Sd9Xf76g+DBg5o5B+bLd
aifyn8zq+qSF6a0CKebPmsQPGUW7fxB+8hAF1AVkm+91Wu8lY2qDNggoZPTasaiWhV4+bMe4BE35
E8rcgMgMgXJfmk6y+Mj7YWVch6JbT/CjgJQC1fIerr01iIrQsFf16waG0i7PWQtzTMAWfFoqElFo
JG8X6X13GxIzkf+9R/rg49gXwc/KGwQFLvOEdBinmHHTBlbmLtg4xFjm1lmN5kREEpElj7zE0I4N
0n3ygIarmHarpWuaXuYUbWqbye8Iy4WBbWNSJ+rOKC0kPvyns0Ik6T7cr2MzzygiFUod5AyxqQCR
7++qw68niMk0EuInmTuMjrSbL9jCuzwzbUfK00LMBbTwEKj1Z4TKiZrxliE4hRaFJSbCsDx2zd1w
YfwE9u1h/RjvWZSCRCQWY6ZtomBCGTf8Pry63Bnt4ZErPIrlaLW75C8+X8oMI+K1uxJIDcS/Q6Ab
tlrAZBIjZXNccfZrAFcsbQg6BcbNdgku4jgmFl0ASR2rPFWI1Lygjuy669eeFwINQCxMeIWZf4LW
2O2A9LPHyHyiOe//U+7YMT3/s1P1t2z7AXX+18LvHNNCTnCyL+OJykFfTG9ShebgotdeuJa+8r9t
DDi7VFXt4jcwQ9GlJ3l3mdZ54LPKdGsFKBUsItza+g3emLs1jK6RyA7XrcTrfaLJQ39zYQc7e5gR
rfmtEAmsujNqxMgjFVVQPR2nprQbDE3h5n4sBEq71UNyN82u5Ef0YriUP/FS3xmQ3fg2pLAKR9iw
AUucnvz4wJaBgivKmzSdqM6EdWlb/tsocW7zBk/MD/wWcFSvlqJ1uTjwcVGI+DtzFVSyDa6HqWzT
WGKwuolQdeAOFwAwNPuokxYJo+S7P1LGanrRrsEGoelpsKqAbYgP50mA8zswghZDQqyM+WdG8Imm
PVQaHIFaI/pDpn9RQksc4DV7D7frmN8MNljAXoMI964jmodWCyueXND4cvIGEMA0Zt4Ue/1XqCyQ
cSVGdg94gSPcnTleQ5O337ZXmOI7x7NSV/5Vxm0/jfVJ8Ds/wRNYbKTIRjcuTw/ewGzMj5f0OVox
4SzN7TD9S8lwbSfd/ARr02ALQS9ezT0fsu/nww4xD+1IEcIOQGhko5VyimN47x0USQ8ScXiSkXDP
hF0ZVwmDZMLafS6nLmQN25LLxljON+weX5huGhpXJ1CxBt7Ahmir3EgnEzsV9jajHWSZAOeMyp6E
RBmHQONzscDANlYZbXISwyp8PC0UKvs4PaQXwrGr+BUdm2D48EBeG07/ggoRu/y06SgTdwaN8UpF
wVoA52WOGj2HPbnQPY/dmwZ9bOUu6hRXTS5r+OP/bWy04bs33BCknpeuM8ly1fSo8kDKLGNxBsRb
dHp3WAqh37uSjVPYYD8CXD5aqW1mr1rX0wx4YtuueOBz5z0bdNgUcm4rmXfTdz9IpBKjgdJWtnyS
+PgU0KRb2uQaQg4Hg6A82nE16QdpdKeYxsVMAwpQqdBWx78WYdbZTEkV4N7+3V7Sl2wAeTa1tk3i
kBaO/5egdLWkbRNO2YUoFu23fLMRC0AP89Lmoiq2U1AAe2QzYSmHjTkYHtm+H5ARWYp7dLywdsnl
ZZ5yiWuHYEj7w3umkX1X+pC6KgohaEBxSiInLKZRMdKvNAVdNEEkUbpS+wXBb1D+YdAb8DYfQaGx
O0vhPrdHiGJCY4BOqr4IoLn4VIhlZSdv/ogyII9l+bPcv5zWcbzkpg/ZxF76hg7174nW62Bpyvmy
nlJkgfr0ITPB5ckvVwrzMzci7JNb1dHt5y6cPud4aXAq8y0okKWc0M3ZIY1PDUbqc40x3aeDT3yz
S6GmvaPYnYhEAg/4iMdgdXX7w4x4rQNhjZlaFor/KBMgaKm4fLr68LPKTYOIHCqmMP0w5pQnc0aR
RjwYLBm6xCWTLTrXrz3dk5wVAqSoNytWrHWEYt9ob2VThPK+e6oXKNehD+cx5t+wV7gau8mKXGUl
eaRbX+jC4T9r+34WjvjIaH6Ww38hq+A7FFoJH8XHWUlJ3zm96+smU6VCh0Ien13GsZ7ZjHY4kXJR
gChR1Gy2GWhPyvtPXn+ytatFtRQfVX+dhF6J5mVhpJFzQ1q9PkqE6ikwdITpR5KXub+U09CjKnrz
g/kmA8gKY8xydohhTiJwn8FLxZFKlW99exCrV67brrqbM9RRekD9rHqAvSygJpGy92+EEDws1B5e
Inhu1ySYxMOy45tc8asKSaa8hDHMqLjYGzjXSA8UxM8jNGT35B+47YY0+w1r8hNPDpo5If72bnmL
04A1Ye8wtE6NX5YlWFsjwG/9wSz4uZtwkPbnYM22CJ0afrjcQf24CHuk5ArnI/gLBcfq2VvfyZ1V
1PnrA9EK70OHqo2rMVWMffHlvd6k6MMi31nEP5SNDvlhrskPVqPF+apOIfHyPsZZMR81XM5xhRji
Ofmvhxra7a3HiNuErgHApc9hzlMhXJ0UKclT6viWr3OdzHUXURrK9ffCzHdERxVMoR1N9acEHSyc
jNhdiK0aEefHr96hao2bN92706fjvkzx5+EoGlxHslC9KjmaGvUXsyfiVu2kKGTcKSrW7+jQIwLM
3y8oYFSDmNLmsWU7nJLuRRi7j2q77FjIRH2dZHdaI4l6HoS4MihZWpXJSGS+U+QjXLmL+gwRsFaK
TIpBCK51xxgzZyCELNfPC04uFXO9Ob9Fd3VEmr1XemkUGmFLRoPQTzsqILtwTEZnr/n02dpRxP6Z
g9A5FuhafiWcnOTGYFcU6+Jd8EdaO0UCezMJsYdggKOt+h6ZV6++bhYtQ1UW/ZrFoyT5k38Jb1Tc
8EU0iUo6BbNOd1kxGKRyrfiS/cdbbrvlFF9rNX9L9ejyYxe+53N3JE7MSNCHBD9nrXEZKiE1RfEf
rr/1LmLOJ9FCCWMHZ82Y58nIYAQQjXjTbXx9nuaZiMN2Q7gCPLDnF1291CwTVMGxMk/vh4rIjH1H
svxewyRSuOAgn+N7FOsnRrwsmE+UXcoAt/BK0M+qqGWPt0p6+4uViweFpitEHRcUZEGOIbANQz31
BuF4amQlLKRR4Kl8kTBqxrmS85Lk5r0dxFKgOmeaN2aq6WeD1t4DbUGAwKR7BymuN1k0wptROqsz
18v8r84s/+mJcY6u0YlEQEwxaF0clM4cirbceUlxuwQoQv2y6ZatJ/CnTX2SXh41r7LRQwQSijN1
49XqWKGT63R0llbZEcjlIT/5Eh5ELFpxThPybR/6zcXLAeLpdNqBkPVLsKCGKs2G/+lRXUju5/ne
aDdHWbVZkeBt4SxLRqmc+kY4pSjXFIaFnnoWkgqlzl/LqxhUEB0NIUQDybY03IWvvAChbxUiUtrE
vjhbfPTF9Tt253K+L9mdmwdrUCr1BkAqgUFNJT8Y1tU4/5CcDLrommjCeFnqR49Xqj90DcDl8MN5
F8GhrNLuKKVNGYeSj7tO+xgTycmV/2SVpZJ06unTloHhf3lzM05Qik7QdVBTkfRw5rubFx/yPZpr
DQFuIE2Zm20BQX0s0OA/DjLvylmckIiguxmEwcQo5iaUjD+PLusnGavKlJoWa8luPZV7kJ71pzzK
we+svqdVjRTNDqIclpSBbWemiGnFf2iLYlErk64m5loB+rFGNE/dc5Z06pfI1HiCgEXmdNSjfCyq
+3dI3fWVuWDseZZI4qFaZfbLc7LPN/9SiZ5vPkQaor/RVOZmKohiwBfAyZSk/dFwin4Nf0wHMOhs
xxXKulckucXznF7Yw/4py3sYFHfSdZ9MRMhRhSdvczejq+GTVn5W6iB9jYmY3PikL+Z12Xth4AZC
t3Cdn26vyrMvhybLLAXt3EI23GyIcA/RtYLZz4IdHdRAh05V3jcDhU/Dhe1XLIySD44TCv+7sHci
s3MRMrAGEcEbBrCuMXCEfIk2jxBuJxhaZB9XigWarER6gQuvbeP/pmKSVzpsWJrgYzJOXF44rM53
PEsQ99lPk9iy9BMKMB2loNVTU+3lQJcNuLTekQkVVNJykW+VrUMVgogOQkCz0AVLreggCLJeSvix
4HsPXYY76Lgs3nQBToHqnhbJrWlTbLOypQNkuVB0CKfhxfpoDaHgPMVd4CKONtTL3VVkRfS7Id/i
paNu2lhj2pKJb6vIjm4pz+4GLl+Yzcns4o7EFeEVuCR2r8YWtEkwzhQETKshtQ1DjVIROOo/riJS
3t0aoNqSwG2DGj0M7E7kkBXML6Lf+0hVlDZanuqcNY1rElM+sbiO6EJpGPpnx/3OKFhx0tTjnMed
wxduaq00MvwqiWNP3pFDu5XiFdn4Q3MElsuo8YCW5jx+z0VLYoF3RIMNeu1inTgsxyJEO/d3rGSt
l4Z8L7XUh6wEalAFJec6ZgyeTJcvDTPGN1rP9gzBg3c9gGArFDZbNwTvTkJ6UdkLYF8ilZp1aQjL
eydOVX5qTKBj75VQ+9jj/o0F1ZOQ4wC43hYd9QlkwACyVb+5xJBM+0d5NAAr/+J+B3RYbpg/+kYT
WVWuTFqHMfZZlj5zZzOS9j9ffmM5P/KpAb+g5ZgYDWfl29d8UvCtKjOhctBbLc26yIpxAD4vl+lI
zgGSkLbx3dDAN4g6apoRRBIJD1Xb1JFuaNl7Y38zF0pU1f7Lk4fl4xYq4N8aM5P+qzjRCUrVH49c
XiFzxi/FNiyxkQbZiGGz4oZGvsUd3TJrXpUInRz0qpkpDS62Q5wWdg2wRxuPyVHfdNOmxakCDaev
4n9hAASkPCaSbCUkrhzBcHOSXjOFt0LIK44DGu6ucDUGP7bXvszbKFldSGlx6VnIVmsmeNaYygvW
PS37ZhqIn/ctbS/Q4X+v9IrSMg6KKJ6lK9NrDQXAMGBwg63ibCzDz+0xtEfxLn4ucgzfIxqSElsK
CydQoIXhNNyUyj3wmgLvOAD+12t6pjSXfmIOTPvdgC1Qd3chcfmc4fR2poVCCBbIQ+fJqMOc9d9R
s4SkkU3aNSaPfHSgTm5yKrDugKuLZC4nsdWM1JQeAYhLnagOtZKV90P10NEm+k5JSbgZ9wEs2mpX
NNpQyjwDJaLHSN9dJSsbkB6cccAuc+uVIquhdVL60IGlwX/iEivkvPE0jmtscOHbAD3OEojNpKIO
u95jvshiugw7uYzLyzqj3Q/CiJlKXUBe4Z4t1Tq2t/h3xVW4KT/Zgl8ZfjbkIzAf03oXMIy+4qRT
9hTEFxwF79sK201lYL3BA/nsqJn67z3/pDDnKhRbXzuX1qiOdS0OpLc+oY/U4+nnsMjL/q0NTd6+
YMRO+RzN4pMBSLKRVIaCcWymdlqx9ubCLbJtx5f4z6brhKY89O3Dar4Zny7+7/PQeG7dZWkoxKcS
tPf/ZsI3Uqe0MF6ce5q7GmKYWqTJx4/wX8YkwQo+6VZNAFtHcGncmSgBCzAfeWdWxXlQcLk8tL7V
PO0GFcEO3cPi2YloeGAF5VIjiaITLy+rgeKhApwkdkSOAwKdSbSexmDHIrvvVXTEBCgZVlbwEcZo
TLedh12PTXJ6sHa6bJAC6j3tMrvvisvQBxCn9/9ninIowHtJLMqZxGP7vKE2POBWJ6h5gAeW+OYp
li+wSDUJhb0eCdshE6CXLL/UXNs1Ikb27cHLfBvd2/l8JK1d+afZIUg21efxycuoe+FnrtnUn55K
ZMrOypXB3KMG3jR4g/xuFwIYHlFj8ovDlmn6GSn+tI1VjxGKE1b+qoB9rDRTPdEsiPdTcqcOMBsz
2sogz7eP9IFLygJVavCdpmMSB+0P3ywVBeyT02NLjsSTbBXOnu3pXD5bVf5/Ux5p48IsZYeu4BHF
12YoJwzJbU8YQXxImiwn4K2zN268+2yJtPtaziH43FG60NCvkfTeEwlGQmh5RcuAaBp5i339oqsG
l02VOX9VIdbMsezKV8tmmIR/bSBiv3uH0rf6ibkL4rv/Z9rAgpM2/kboL0VHbws3ZEIXu08ANyar
vpq3p6bihLFkx3LgpgJAwFaaarUsiTRiK5G6m0BAV7JtV1xCA1FjItt8/y2FDyy/h0XTGReFoVPx
9ldNfKyBfy4DRVQ4rTlemmPgqUt5FeN5iz3HLieAgeJ28rd+TcSgURBUS6ZI0mh3Gao6XWO6XdUu
78MyFkkKNc6Ct0kvl63DOQzKNj6u9jLgL/90+bkJdBx/KuvNdBxdJuQ43N5nnLs+aHM0tbaCZtW9
ZGE/96uq5Fqneutg1aA5vgs/7X/PCtQAGYo4jj1KNsVLuDm4PWOLomnHssG97HJL/5rwZ2Ic7EAx
rSShisvaWgXsZVwjFm7vjm3ICGNus6CGsclqdi2MpkUDAnW2zULFKTS4MLb3sdh4/2fUsluyf3yz
MYaGsu62d4IBANYd1v4KQILpMS+95SfxHNKju58iDhb0/A2RioUcm2aem1kLGnl2Uhv/HTLoKay2
TixnhTwXTaUsZBL13dm94sGAdDtc3tW5alZ5znKF6OndOmDgVcvBwvOntCCCxinuiRsFq99+KDzQ
Ss+vOQNeC3OqgLMDLkdemshYwcQCG64IzO9ldpglYCqODbGOvhrlmqLV6CZXXnu0eN3zkOcZLOSC
fI5OW4xjdJW5iD3TEFCjn+ufngEQWL2kvD/Y5R4jivQeEjvV6Y8S5MQFL/etQCk/jhddir9Wh1qq
BVFcc34rzmAtAJ2HMXgYRUQEW01e1ORebpqHcPnoZQuwnZgz7xohQew1ZABDWiGPxMBrEomL04HS
YGk8uN1AonvlCDcallYGt72+IQRvNfrI6LdECAmfX6CdZpaTv9ohJdLbA2aHVZXUnvvFHU1P1WWk
EuzliTKb8tW0Tc0IjyNyfappXxvfpkGNV0HEbesfvGI5EqrWi8IaeNU2ldlvPUGAxnNOZcTMdAQl
XetDu4ugn+yjDpwQ5SsgNDlGT5GSY8QawM1eZR6qlOdrRHPi8QY2I5zvmnjLfLQvQ2Fb8Rdgof3P
O911T6mLsbZH0y4+LZf4+qMCg7Mw5WsNy46lmj6NXyxDpE9n1vo7n/k/4k6AQACtirkCJMNU3l3G
UOemhPXum+96QtzTG50to/y8lIkU39CCc5NoyXAuhhzk7zLKx0U3wAYVkIQuC7p8nhq4Dwdtn1Ur
EKv3eIvv9EpIzBQPnRpmI0TJeepWANQ7LnEWV6Xs3UddpReWR8OyK9hPdJQSQ8pahMnheLHDUT4u
djfCYI5rhgzxRze32hikKVfDFTfu5vam7OlbejSrT87iX/M4R5jQVqQ8/3aIpR5K6iu7hzGLAtVD
mKlg9JQ5TrJO7HJD46OMbo4SCx6Cyuq/KU7aegyODNzThVIhbSNEOZByE+HzeHfxfZOmN2SYz0+u
rUnyjzWLcivJsmIgzfBcUWpijAPYV7saeLMlPMUPxfjSll+EVm0bSdtZ6f7JcGQMxjCcg7beiD2r
mH1N9/ER4AueWx0C5M3fVVVP3G1wyydxdiNKp2nIPgb0UC89dePGbq+84Cyd1kSQhrhM+NrVMdUU
0p9Y28dNEiSIExVbdT9xQjju87KzKtu7xT0+ujmblZYq/nr7jZviqqvvFH92RbBSP8AyWu/gWh29
oin/b2b5pUhN5DGgptZx5LMY10p/GgPlVAj4ocWkTYESU6YTeAsL0uh5ycjpBb/wmbNAwvRcxAk6
yiD2AYThdY3aqIDjgmoX2kpTHWsZhJvjebeMUeOix6a9hVuSXaXjGu2D6r3ppEifQ1+HqcDitZTk
ya+xfQwajjK/2QeopjXym4/427siykvLWyZ48gHGW8hUi/tpf8GfU5CbxUAHpEtMYgkwX34GXXD4
H3Jb+Ur4KD4vRoUxIfhOgR5ZgeSouMqrhr+8qceBPri9aDiXAALpaOBPVYQ3xpJ8SFHMIXWCBdf4
QA9vUYV16aPmA9kX/XHKK3y18I1fZy5tORy65QOAFIoPrP5y6PCXKmfUfeQWkTLknr+jAEbdNa7t
rDgOZqc26RF1UudySUPND8VI9R0KFjpKPCbAv2NyHXEH/cZX0lnH461hN4nXPttnXnHdZfmNGIyM
InprZUrMpPRYjUAipWjbHLzBGrc3oQdsD1163K5PT7uBIwRFKJEkuW+NkKaNWN0TEDCcb7Um42VD
1GTfCwgzOAIJWX+QtTNNNMnteI2EAJ6YzVzf8TYvty8l0GGVhCIeKzyiQICFA+/F9sTokMUhTaBC
twO7ciFE5HNcQQ9QjAkUn3tnbTmpGcHV+VmmADTMqlNDT3wFdhcrx/HxGyE+nv4poIfYcNFxseCE
46u5bAl7eRCe5KmHO4HUHctLinbV4TyZXoGQaNHR9hW+PPNVwRt3xD5GBij9zv/vEf/FcVm9fgIE
GSzbHeDtMqmVAlswzI9LVsa2c07fnGtXGIYNKtnR9IFAVdFoAvCTtnaS/sU8QuLgGytUJUF5SAKr
4rywBVLYH2zU7TF1s7T4fh8vwyC8heq6fYbkyzPBna3asUVnCtGm0yseWlEkV9JL7N9NT+r+/cnV
Xy3c8JfXpgRkQLsBDy2LtByN4zYW/N+GdyMZ/GTOzpTFrCeIqo1QmBD6l5UKFJw9t7VMct+eHuu5
isT716fgxoSu/g093gb3BZzf3iKvLW82Y+o4S9PqfDxgvb0qsqwNIkXyIuSvEZow2YIQcYmHMayb
8/ITXsIbUGwAKUD1KurU+3CeaL4qy7qAATfi0xCdFSnZaNX8LvZ4Zs/jWDHjjsg1vVoqp39u4Abf
cpTmGuXLCeAEPoUJS6WBplRC6gWl/rjgsC05NimaB7N1HppwjhCDwQtqn+d00xvD0K6IMag3vzkc
LOdUQWxS7GG3jVKiOpPKUPmyJhi8rOP1w0v0lm0EH1bEUT/Bf0nJ6LHqFceG78ebnhf7Y0rds09B
7yjU85rRp17K1im3n3/RwUyM+yx++2szYaXcesCbprryBxT8ZU1Mr+ZvsVAqF/J+DOIVrI8JkZa/
dESKMtHlRs9xXgOC/x5rLd3LecwlyTRL6+J9HMYiOlD9mytCCMFx4T4wFY71qGcq8FjX7sLGHyv7
2l++ZEq2qZ42Am07kG45RhmZbqgEw4v+jXO24GnGGdJjKKHPkBRHKZv9NTczmjVhF7alIJ81R81u
bsWTYoYUv18ZNcekgM662rBWmkDO0SHMSTrfUaWUOIKJlRamd4GGzXIznLVdOG0OYxZ2ckTSs2NY
6kAEZHTejEKck3EsvMc0K9CfeFI/kUKWYUDEqy8qqckfJdC2uFgFYAtktEV1Zg/5L0eMEiTLA2i7
q92Xfg7IAn2XbXqQy0wmfg56g4m/hiGQvOyHfudTPreTuT4hr8y3jgbDf9orURNzWUSmpgEF3AV9
GPGg5DH15ncDKs2LUdN94IYOws6OwrKFymTcrLjkE2c3LSSBxdCP2Fm+9gR5w85ojgC5am0r5jk/
oGWXjEA7RDgfIgVUYtXDoN49aNnnAAFVgnCKHQl+mqW6OlbDUFxQ1p7nDMhmmQNuSDxja2ZLtsMc
NR309RjhpfR8Lu6dDWMYwsl0uxzr0gEVokCa7evc31Dwsf1aRlD3ZdWxR0rz6Pc+PULG+avdJ2tw
sKFj+/QhJwdwlQhWXbHSd/k0nE14eJgSY2AXo5rLBtQGbLqqUG2DwI6EPdOuYQU176plyr7HsjLJ
Okqej9Hj2Ex/p5FXngFyzoyfOjTz+kAzaXgXDlBXSscCw5WjkceWaUJq5AePnzdyaA3/qbJI+jei
OvxzQuOtaIAV1E0T/JAAp+1EzZEeNDd3fiBmUHGDXZ2XaqNezWF/n3SmrQ7p5olbKaca3UmqhUmq
GFzrdknb1jV6sI9qrsEvPxwm66Jj+ony0ODenHDA2FLsl/kGsXSMV/zdbfu1rBtwbYZ8MvlAq+jg
l42aTURUF0e4QQzIuKPM71FpwkUBEF1+FhATAISh+OmEyitgSnFHmcsG22nmQ2rQQwi2ZeCYqwxK
atWWu8UBVICyLlbjg3arrq9WamPZJglfB2/CpC8sPo3voFL7hU4RZQGcTxGQqC5t4J6TkCaVDzlO
F1TpLH5a2wk0WNir34KbkGXrWr81pB913tDPM/FwKY9vomkifNqt1Cxiyz0JJcy4GfI3rZEncKJB
esFidChmo+WrdHkBfuEZ8yQWEXbbE3iSFflxz6PylI4w+0+qO9skCvbgrEGCLuP3l2NmYmMWRTy4
K7XDTPKETSVytmIXb+pF3rTuMJutNX0P/dGUJia81NeOFgHmUP7V9qbkdxe8HiXVS5sjUuM/ok1Q
bwJncpyAmasTdmhFtQuI+khqRfQsCpj+07+PyLCIcytvQxhZRHSQPqTiOHRcCaQzcUdEjCMpbNac
Yg/79GVq9GwArjHUgzK+spAjHIxwDKM4HS0tjLGUGuJdT8hu+91eVOwjPQRnYE6j2Qqihz8o5AQ6
dm/YNhHRVif3ebQp/TNzXnUZjFeSJoUn7uHHscIsNespVh55nX86pCEz8OGmu2cn4asfW3owpQqt
zEQwpmVsCJ6BaqOyYT/lOcPq10Ka7gx59l2gpky+1NWAWZFtNp8x2JFdF+zBsxUaWNwT2k+Lr2my
OYCmVTZdl+qUyZLJnMEw3BIB33ouG1WuKKDFkJvjrkbSyZdIORRtKLXsb5RTMM5HE2QRx0ZMUAwb
u0kYjFlFd26iY4g7k6F0ILO/goIXWDz2jn4g3XSnEWmhWg+QRg6gmGLHtYpBrFOHj5LqlhCFbyyE
MKdpJrBQ04vrmZpL+sLbK/sAcze22omyM4emdQAcyJlYbEzKSen9PK6Zm7juayGctiIsUzXgWucG
jVLsSTrDKH4qrC2Gz0DsGxtZmnZB61W+5RWL57ZT53MGOv4I31pl2fdMmIhbwtUEJxsNY/95RKZP
NvZa7EuDNtC3sy3QTfzFOPWmMrJZqVmmn4u6EeexHoHNeg6opoBhYvFMPdzsbfTKcPcuQZZCA3hv
EVMcRMcT05HYfeW9+x//I0XwkqGMLikZjw6jxaYkFIF7s5WwYnCcSSZWFB8lnuAXvr1gQOZl+Tev
FZcBKxlx3ld6T4TFEfaaGvCIserA3shtc3OIAJfrOdGmQx48BhHjm1pENm8XjldsEzpDhG954MWN
VbtOCrvYdYeaYc1un78zRgROYwEkZpzL3jWpulKV47uUXqEFO13HIIZaJsw7wwszJbymDhT+xnGH
f5TKPcmeSGIPFTEC8m2YaygVv0AAR44E6p5i9ebJR6GWtEx0jEbKhVADpO2avBYvgVpSLzFgEeR9
DL11qsmFToSiHML7a9YV3hlcEdMYK5Zgbd+dnr9KFtt8QAcsHV2/e8q5XUKLnc0hScxtp/4lVHb8
VFz4SkgyF4tCZ0nK45PMbtiJIYyMS6eCt17Vo+nqCG6fyKowsugdhi4rNTzJU1WXt1oCq/Z3FOmh
RrJLXriUmnd2LE6G5uCCKbJxS7fkeObBAmq+ntnP1yvTc34AlwM06fx40AGJWaV4LBedFh0SohXE
LD0C3KyfbuX+0TW+XZj74jGAsJh4GH31XbCrEkbPBUkjlgFyOaL0PXYwvbc22lM+MHRwd/gUPwvI
+d0msPsMkeCb2jEabXA88j9TUUKyWorbk4+pyhFiISf6Dnb+6FKuVNy7VHVL9Cr1xVkQb8+MVtUW
vxtZtWOXkwH5FpoN81+M/zgZUUDY+nCU6CtB3ARMIZCVa6xep5kOudr6RAnXNE9LAraPUNzHll+t
iOaPwKcOOAY+V5cr8AiVhLi5imQyWUqzsgXvJtsDQ58Zo/jwdJb7/sishc3WmcjDLMC+T/TuGAeE
IyA6gaMco+VPk4QuFvcNX75NmEVlx9SVgpeKop/MdEy6bv1h52mVMiBZtUyv45cM+mz0BVCjlMGC
RwIW36eLpUTTFNeeJWUy8UIHBCHTaz/r+S0OEXw+ZW3OTB1fEyEgriq4YSm0TiKI0Jqtl12kwZTe
S16Yf4eZzKNoUuXPdJ1lgJM97BOoyhKeu+3+3R+afO4J+RriczuZ6VzUHW2QTVlYSm+t47syiYLE
55GHTDJgF8JCBat194AZTxN5xlyVUsZIpXqIw/6+Bm3r4HJRxiPCmYtCG/VQwU/bHZXleEJYTBii
X8J3tGNFgk2map3kjGuODH+dvIB0G1zhe/zRSs0yweLM6wMr0UMwnT2o2hFxjOhLqXqE77r9ZKlX
8DLs4GTCArqNPPId3KY2AoPpFFKmrLzQXqi0PjfKa/W4vPboSDBApqiI5I7ZhB74nCVI4xT/aKpw
OvJqtFUrrZ1gQNukTaD3ifwXJxIMoGMcoHUuL3e50AnYnUjfTWT0ktlwO6oVjnDRRbKX7aV1zaD5
/tcADQg5WzdV4dUtJtPuaSWa9RhMg7mIQ35+ZhqgAtZ2AA8LO3SsYgPHv8fQyO8QkUmzNSdznVaG
Jgl3ojppUCObZ6beT68NUet2/h4ieFF6yLSjd9y2OIrnCqQSErzBEh1ibuY8A73fI/HcShFVGTmL
T1cD0/Uo+V2fiuBankQiSiBZFD94/HCgPe8tvGUPLS4cn1W++EDyeEXipw8T7m/34JDqUFjQ8jlV
OHgWvCoraGst9SDPKtp9SjC38L+UAumZVXD8+RSLOh7cLUwoIue4PAm1i6ljSeeYyUHrDz7yjYJa
x2nucyYj2nv35TA/5wALX+54quHmN5DGk3ucxNzy57XfNBe4kPRnBjUCI8lzQkbFsUzphQqV6U7d
l4IM6qXiAQnBn0GQQv0wUMXUFDAm4pVRgT2IbcpsF2zA1q8j78BHiWi6Ug3M7PIMmzJftzJ20cbS
GoJQsa36zaYvrkGLGtGdlix0An5EAfpMWW3CXCy83kMEApGRyPebm678ODPtLgXbFSRYi9tYa+W3
sX+Yg25vF9/WExlnELU6Vd1MNfStR91NB3DYWpREsZFnDn4OJ69khmKVgdUJrRU3Vq9IVLiW4Lj3
oS+DyQzkY8Y/z9ZD2RZiwYl+E8e0T+H1timLXifGRWAfcQfD/QjcFhpdkZiT/WqVBMUmw02RjJrY
ivO15HcFH1gIM9i9WSl0eEvz32DzhC7EwtqLpSKOpTFEA+BtpUNG4BbpluaJvburQyJNvanMS8ow
CHGCpddBv/RuNZWYUsxqugE86rX+AJwtYLDyodFrvfgWXVYGF6YDVowmvyzfvko9a6TDMEfB8ox8
zfv9WCqOZTcq0c4dzJkJd3fGop8JxDDQqSBKE1s/xWspx/axeWy4SmzZqpyIFhDkSbG04fxAAqVh
kmSmG8bNC9qtzs6jIqFQFxIwVTmCRJElznknrvu81M2mNhTwHtuxVhf2WliYicr+BRIlfuVBgdWm
iKSsyRK52+9kMKWugMrFAZ8KMhUYYPStOyhV2CNq8jtOHgyzQOjAzB3f9wurlD4G0Gjn9NbMmwX3
gKEfdD7PdhKNmDbmAYdbiBBB4my5w08H0wIBZoydlC1eVft3Qa+E7l/DTKlfNmv1yQPxQhnMqb9X
pj+CzmUsvOInZuZ8u5slpKsQ0WzCrYzUNo9KY14JsJyv6/Cl/OSqQgNFfq8QdO3fROs2HelyF8ss
u4TtK0yVzRhhBIwZOwqUh154O8/m4UCvoigt8puZfbLhjNQGlm9Lb2rba/HfGt6E4K+BJKPd8xKa
BIL010USo6kdHRmaSA0Hr1bDr+ZTlEf1TXqRgYZODkuM92dqZj+2Lm1IAX7rA1HLWpOTMOR4SAbT
liB8nrLmXtEcwzzJTzQjGKR6OwkaFJomgP526w/sv3Cn8KxEKMzihOcYnW+Ri1fNm7TGr3mvXreS
wa2rsEb/PJ372l2CS+qYpC4MtnrVxr6F2DcRp2KpJ/MGstm7quEpZBUrlvCNs5r9hH2jymgelkj4
fGvLhnTJuCpd7lO6LpXUI1g90aONZgTOStF/GwY8Sux5rFHiVEm3kVjWVPfSwb2slfkbl0Ut3qtZ
rRviVOX7LCQYEs8lMXYkH+ApJFAqaMIQayf1mZCNAKzAeYdFP58+cCflD0UR7cMT9wVfP+Stsve9
6I5lWY6/Dn7YWbMw2PpuZpuol9DOhbU934Vlnk57eTH2wCOUUzVNSItYZIPp3b+7XzygwiICtHb7
YOiBaQOJGMcn2smcId2Y9qUk9kHlLERARfrPwSIHuWxmZ89q2R7rbtbsK115YZrgAR05IxoTBm8F
TmVr4IWo1U7UvYg6EwsxBzzsrCinPQSIhzGdTc75K8/0eGy1gcOV+vZ0NfIkYv5jUouzdRBe3PN5
Xn0ehGWKXD6PueBDd0nE9bw5r5X0fqVfgcAUI74NmtC7075N3SfigonhFhS4sZ7to1uy+6SbJa5Q
xd7DVlEiVFmN2YJYYaPRugsHrPDNP8g4KCuYC4wPp/tV1ukxCewiS0RWXBgyuRmdTV6VmQOo+7bn
ZkqXllxAnrmLwdzgOPlzafjpNulUaP78SDw24wRzsJfDjm1EzMI39eJRkQK+IL2HvwRPl/evI430
T0hEkuysC3NBimuGJP09DtXoo7Ky6vuqHwf6Y09K4TmprcpvLFBP0m/s3wOPoy7NYSboIt61SJQI
rU+EfJs/LrkB5Gv4uyKDJg5r+Nx5bnRAD8uvEk52cKKXDzEI4XcY4LwIY30sxURODeY1eBAYc+Vv
ZskkMWlgExnyaKuda3yVql1iVe7+iIuoU3eANSqPHlafsVPrOk21b0DOeF/P6nuGKaJ/n+3R45hE
6ml+D4elMnL2NKyYnwXCH57m223EIhOslrhdoQqrcQ3UjuEG6Lh96CNwohR4b3nBpxvMPTGz7m9X
MWnLz25TRQByZTs5H+52glOu6K+tTi0klA1GStP52VfhaIf0PBTx1QksmH+qfPoGnyVo6mafDj08
TiOqi3zNr/1hJn7x7PN43FRt6xoJL/4UYZR6bruQBuzcmfLMN2Xtz8mSVexnoIaYLPa8f8wwV6GI
RzkNPqh9qy2Q4BwlYlyxXJ+WvH4LcC6f2R2BE4SOve04Se/GsomNjHniSMsUP9o0or/64TjLWp24
SdytDPD3XSzOw/6CogoMuL/mV8OFcEPxKCPVeCZ+xL3gXBGpP/NGkPPJPVykYzAZFtWS9ikfQOaj
CDPHixaxw0PePC7bizpAfLSxlsyWImQCVATKqkuLDSuS9wS+oQLQKU8bRsVLTg/dJhpoYas6E39M
XqsiG9/O8P0jzdpktzvQRzC0bF0e5iovQMvYmadMszf0xVlPbmdHyZpksjM/fSiSVwAKsJFzN2nj
RK1ygdxUMwoMXxOm+eeosGAkWxjmiV4ENNZXNUq3Wj4tO/D5hWshnY4IE8LPQo8V5PyfzYOMtflC
UQTVMsXxMTuKkEvuwwb2xv3gKpg+h+XguocbMcWOlZOgWuz9PhkAHFKTu168xYl9Z8+KcuQpj8Va
3TNX8UIDOik5awHlJLcsv/pjmUB8vuxrZGr1zUU/IZHOqe35QgQx/H/ZdjFqtDqP+39JUhz4obCF
4uAfwJHlkpvVzHzmdQ2WMUH8j4WNUfGdMUEOm8XePSm2rg8Nk4S/f/87ZrDmLNoXUN8r1CIftvrV
JA4KcauwT86wjeRFVo9x+3OpzRHrm2o4yptQva5dhnL6om7tHCQikmt/JE8c7175OAxExmSqVWnW
6gT+kYaaq+BdJwvkjQEr+qjuV1wh7J1lGquAJ04WsI1L5ZDJYXFFkXbOSR6WhefFe7HetteqJe1l
gn6dugmzh+GLnFxaaIGUD51LtCy825bpNH4P4nkF/WnIPFy1OyNcz2Uy47dxHxuhUG5UzphUbUA2
7nMipSN2JA31thqME/A5jSho6j9q5sR/I/xELbehxeyVpVZFzD+zHBtxkWrtYLtBJVJy3Dvp7REO
sarimGx+OWnDQQxHUkfbWuoPlwJN0vwWmuQQhK20o4HqRO1sg99r4ctIKTzf4FsvGoERvxVo9Oxd
PDmE13remea7VzR1QPdZtdG5yQLpppU18pYCe8FWYAkiYNqzT90ZIacmz903ahABSlBhg63MHlnt
qTv1YlXpbuGtllGGkyyz1/e3fOkeYiRiUvoqc9PjmaKX6doS9UsIxH+GJb/cqmfuBAi73db2NdrO
w48Za3lFlisQmWTLKrar0BEkOIwZOgX8g52dm/9DzFqHC+5zy74cM1RH3FThhVs+DTuuqfXnMqit
C1VnvGXt52xns23RHqjkAUYZyUBwJ7rZTq2G9gttY/x8t7b/Yq6UJtMAsLo8K8EO0sNsAGqUr3p/
b64X+leDyw8gR6rSMxLIxJcxrirgj73pt4rs2gIS0cNpjwvm7VjU/dCi4abVv7i+gdRSRNaVo9AI
p8UeQBkykLbHzseGdfiQPEe+QwZ+AKWjbZcFHf278XPwutYQQIQHP0IjYOVakj1OLIRWu0MXkEE6
K8SokbFzg0Novwsbjyw97lOAghpUNFoNQU/v+bcP9evoOk6ZhT9HXSd2yUhSsfvrf/T1lc1QN9xp
pKr4m5gRMSzEj7ycXJ1icshSqbMuyBvbccHLibSQJjoim/SDEOZIXwYKc5DmWRXboBEkx5fj838A
ksAUeEEGZXmVvET83xLObeQ5NrIRDrnSmHa2BYLMCrxGZN6NsW+8ukXOLtS76p4g6log8HR/g3FU
W2bHXF1o5A49l8QmOMArTYtT0gmph/1ORW+FZE+q2hA+YeyEvgZCfHgEIaGMRvnLjXi+70uSHB+j
wsjXzl2yYXTJiERm5eKP1KwMIC8zumMz2y4eHN4WhTnA1uvTmYF/MNi8j58BhWy8TPftCa6TxVl9
NlzBGYsCYcjFYoidgonEC/13xxIktBEPa1KLwLNb6A5fx3KITpm3DwY6YLdqx5rkjkF4gfru2O0H
ujddqB35JvWax6MdY1nIvCDbOo+Jd2qcVLmMMtoNffL5bmz4RIwTBdsDn44bzPFcUKCEU1S+EiRm
nGosaDFCTJ09wWYP88wO7tuCvqNA4cBM/M2WS0PLy9MnB/oQ59ar8q2RazJD0exJzsW7gRd+pjL1
IJrDv0iN86QLAz2q+tNAd1SllBFVELRwZasSrrNN+SICCnHA9D7sg1fTPvb1IhFrMkc3eFFuIoc0
9b5EBZMgpCW9igpqHYjMAk09YJq3HBaTIMPpftAOiIbUP2N+q8roVkqg1iq5ssFzytYH5KpP33S7
NgokGRGyWDXZXVUalGxETqtuWidDWmyZgRISk0wdXCb834+HLgLrVbC01fJ0eyZMDXDxFE7HQIxU
O9JMTXWeCeYSPvltlnxMsa5UCTVMm95cXt8mmRiOHn0q3bmg4/8e8m03EcHPdBBuTonsRVftheX7
1p40ACDVwlOdTlN1YQOsdO3kUjuHcPC53fKHITpKu5MgLVK/hocK1d3W7rLEDI4em/0bhw3vlOEu
jfiZWero+q2tcy8SuuNG0hpBCoOkdANunO17l3aO427QSQt9SPQKx8mCITB+xRsroblgtHMZhCbL
WvQRc9Q9yUAxG4W/WnKueG68Ulvv1zAqtqInMyP6ybYvPw03R7RTsEvkVYbkNlu9ZFNThn9mZ7wQ
INZFsvn7gIfzJvG2OnrwoYJ1OvU74djKTf85rqU5ohr0mmVlY6CP1eMqSbklrBGas7mcIVUEKxKT
STnolg1KAjXcVAK2pUxXSZw+CWKfnaFcppi5M5TKSMWyeNCauRXMnYLNS2bGumYmuWqXOa2FVuN6
6Zs7yO3Gas5AehC4RX7/TSjkWf5T4iooNFu89UjRHKm36ZGzqIM1jxEZXQ2e5COQEHJw5C6EVskq
zBnvTSpkqI/k5yPd50SrInv554S19Hj9GVI8xshWjOB8DRl2A37Io8W5eX2jQUSuDRoUP0fvexbS
1DhOOYNFS/R4BzxR3Q0QK74WQSQuLfZsm/piXaY5ScePj3rpT2J1XJeEZGdf3176TmKKFYwDOWsP
gLpzmZq3U4r6mDxRSgUZu6ALRuPYuyhvwzQEzdK3kZRUaTY0f/xcJm+HiePEmLdcn77cKSsLG/lt
7iS2JPyc4ut/bQdRpFFGaSRS0zx7+bAjEO+Jif6ZyCce+x3VMKz0rnGYaBg0F0NFxbfurZXtgqnA
CLo4VdkD7HqHDKOExeQY6Ed7pcp8pwmHcFF/KUAGGCYPY3hQQzTGF9xDZA3m8s0bcgKiz3/oDIDc
WsTE9nGZEevnpZiv0CjRbLdrnkHfiy22v+8jOTLfNl4QOfvcPE2TlHH74YChxd/XeIjCSeF2Le9Q
e1EptJzpU28bJhdHWqK2+Dr7dWqihWZpNf61NNv5KRQFimYsMD5+EE3pKzcTWW8qOUzJgzyPyBbK
nQkl2iutFUGgt+jL4WHvZyF6ujIUchAjRH0rQasFHOS3dW6DywPnE1Q4iRsAgmOn3YJP3X8tbUdM
4MHQMXO0ucwoKFUjMaspQDEd/76vvdM7Cu40GI8iLwV9ogNhdT79QBoyyUL8h+LWIblUfoW1N4aT
sFWZWWGlr0KTSxZBfO1jcH2oSnxOIAJfj+Ys1QJL8Jwt+5MoOQS09SWCk30HB8zYuuQII5Kt0VrL
xWoDPu4wVX4LPhL/s8H2Sj0mxh9fF3P/nrIDpE+eSQtvOUMuSPdwa+rUDZZHGcOX7Kr7IP54zobb
8d7EPDdj2Q6WF92a3LFpaJNtXh6dsy+ilLPYOx9Z4QP3NkSVPNUHmb7zWm0Q9mf7SObZ+uz6B0h4
AD4SHF7wJcPpJyG1bQXLPQE2PFPdzSqMl1HQkkyC4IN8cdYNbfflW+hJCheI3IGYPQ9qgEEmiv/m
2OTX05UlxMj8KcCiOXEZ6TSwqEU1eZY7iFmciMy30bimqFJNElbgFfcwRd0Cjj1XEYx2cKtOMXFg
8mjB+3TrdQYjg2t/uvMAPv4jXx6N3XUE6uqy34awxp9xnyFDXmDkgwGsg5E5dOtJFLljWOcWtv4m
kFJEn5yJJPXLr6B5jaULFGF6HevVHzybnVeFFIcvpcmO9+JPSEReKjBKOWOE55/a6+jHnc7cBAIx
0Ltgmx6r+4KfTgkuA/a8UO+TlTll3xBTR5RMDX+0pbYbfB1ondFCrid5CYpt22gGK9MaJDuskFGQ
7cO3+lfj7R6JcI/vNlaBxeSVqBdFMMd5O6PtBlq989taDjMGuGRM5gxBItPPm5qXAwOZDuxPn7pw
FLcDzf41Msc4QgtzBuMCyfvM2Sk1a51lThKjBK6KbbP/vAwjKvh3t3chCIPi9ZKq0GHEZX0ypSH3
6YRR8PaA7s1NF1bNjo1BHfAizZM1C4by7sWVeaOwIomSNQ0mm4laZPMoUz7tVi1EVP3hp0uAE1ST
6pwEyWmopRv/0i9/DgPKsNv+pAMwWHiUGWU3vsZb9XTg0ORLM3mPg9ueIYWCB23eI2nbVNVTU+W2
/dvLuIzsQrESr8rUm0Iw/NtU7DVHN6brGxGW2fHXOrK3ZCMBk1vssChQVvSBJ1z6RQA8M5DJnHlF
qcA66siFcohL/G3rko4n1VXy37qNPsBZA+eYHLr0NVfFvPjfohpv2+cTDjPwb6ZMe66txf+ea10B
nJWVFwO7n6XnlE6egRjap5NB/QQxlRQdbxwDZ8NTJ8hsN34XkQU6TPUrp5w0pgCYa40133pQ4pqg
l30/tr1EOj3xOIQ9lCAARR9VMtfB+2f9yB0qZ0A7zEh4FokEA6PybgfZ6hmbi9iLkspruoLLY318
dxTAvh2p5zFeD4mfuJ/P2nvaYUQYPqrC739IZiB1p+qxZ7fI1CYucqgqVOCy4ewJhJwNSQoPUKPh
1GtDf2hEq/NrfAM/PmFMoaI6goEW1WMubfw6Sm/dEcy+wrZBt7+Ro9tFWcDHWkP5k2eymG6DF/35
4eGS7rfQwLMEFzdWjcVbv0g6YHk/VvPFEkO5QoBCrPuLzx/1W/ZWBf7uP5gy2cEJDJf5vFk7G4SK
v3oi3pfEFVpGvfJaiNDhSRVmsOj84JeFQyb04t14Cm0pGpOmlTHI5u3HO0GyvbgYQYdk68uTQRX7
L1hpiyx3YZmCynIYGFtXM0/ZzIgIbEYipWe99YiKB+inWUC+HEDDmOUj6Fr7YYXB10jW/sdA97ce
l9VOORi6F5kS1oUKAucybHj6VAPfmRAvR5162OVUaN9xTXwAXAN7vQ3jIWIqKf506SLuGuNKUWCq
TPOF4sLRO/FfSYVVPyecvb/4X/GLhdjqFxPkxF5j2jTWgTFtwDu9jKuJaAd6uZeNPx/IUiJhHkHA
nd+wQiXuxYzmq7LKEkJEPtBFFH5VpTRx7nTDJH0QIlZrEwsGB9M2GNGBhExfD5n8Xiz/vB29mbOe
iASZv2dU/6RXbPMvtWF9BzEvL3NZ9puzEaMlPGjA97nykOwhN29ggUzYRawVyJtYj2Ek3G3/aqvW
CmuMvb2fmZ6A3PM6KBGe65qsJr20HiqSOqTCuPMfXf4fh9fFASvWxIwgtCIKpDoM3NxeUJWRdqOk
OApmEmfY7lf/uh/MhV/AdjL0TNU6EgIJnK1emg+Ev8mLhogzxnButpRQsf8eTfNuXLCEb7r347Uc
F2NdvXZNSXOKeahSGfkT9fT0hKFCS73q+RBre/0TpsUh85mXe/587oyyLtTwk9UeJJiRutCegGws
JUGnWz45gLgUNTnKP93HJX6oWBqbLDCl41H1oCcyUstvC/5gXz+bdKKeoJ2t8bxQJCxTfQP1ntH/
uchxRA0hZ55APcl0uFCME7Z8DfbZQassH0Ewe6YAHm5ATregh4CFj8JCVsVKTBSdPUrl95xrHn8q
Z/bW1ldS3LMvADndjbkGScoOW2BaTqNnEV1xLCV0bKgSG4O2IGsygncJL3pzEkkiEX9m4lRCYnIo
ZUoczmW+uXMZ/uNBHQ+OttU8T3L9wLTFhULTSlm57rUAfizuDr/wpRORKM9XIGG0Quif3vGdza3i
ESLitS7Cgj6tZhAE0GD5dZgPt98gvg5KBmsMUUHhXdrugAjRVS4utF+EzZuiYyLwFKjczQK9q4Hd
Mb1yCwpfhWKf7W5iqYpfs/iYp94XhvZfR57bfd5uhukRWIU/F9rW7n4lM7Rz1EVGUGTu4+HiT6C9
Kqzfld1Ua+KbxXg6Q2m8fz06AxHDl67pkhzBk/kxn2zLITrUyB78KXRf5BEzD6i8C7OZeo4mPrAD
08WHHfxMSxRZp0P/F89bty7GzNonrTZHNQUgHLiIikXHjnfKcSqT8+2B2kAA0T+mTSNNSfUXDdGQ
qk7l/1/UCpJvladsN4HHBDq+N5IxrfakQgPyC6ss7brvLTMoDeeFiZAUNfLKkc3D7eKNhbSwTv5Q
/x1P7PP+J+r+nLsaInLFvtgjneN7x53reWatoJkQnZqis5qGQuMOM6+6M9ZoYra8L5mS2psKnIim
nJhxveEMzZsxjponP1Rh+3fUOY/LzFZJ4zB8SzDpLuf0d7E6Nbakox0C3rrai2WLxhX7CoA4RqyL
R3YpjP69KQrm0bnzk6L/pjiokcXBQcAOo6zYUKO/c2VkbcQXYHXzxDYnCH+p/Cm7890HLAVZham1
nVrHFg3HgivkDSETb/BQQEsN+HkEGWSAdvrdoMe36m1GMRiXtUyPrUJEEHySZsESFzxN4DAqw3P6
g+LUKQ83mocWwS7ssAiUaKA3slVf1tU/qHGean6znMKZANrS9k2jiEBsbFzLi8z74JNKJv2YI2Dv
ccj3LnYFPRvkfloZ12pzOOzZkEBxHNI+N7u2nNSPNBM8AfF2UVA5YkUKPCW2xlttoqHh73URWzyS
WM/gEZC7+qepqLxy3upUKyL3pYtGJmBSTIfeNJcaWB9YaaEbq0tQlPIHFpkscIw1mwfghA/FZYrY
fr1BeWNa6Zt2C+B6T/3V7bG7h7ql6rs6m70OgdzQPukDUsXOkfFeTSfGUP5ix8UFBU3OQtORzI+T
089vvmYbDNDAORRbYxl3msmGL9zAHJIWwXmIanJcGy/WzBR14LOtsUWfwHgqSInVfIOeIIQWNzbG
UM2eDeFaaGBt9mMmdfEsm6XprGXDibSTJgmtUu27A+TQMbMm72f/OmY8v3LsQEkv39GYzHGXWvUM
7tCv0quNixeLUzZ8qGMhhGvLCvPSqeQXWP5E7970cSBrWC9zS+ONuEOY7bw7j48UCwaW8wqcWZzR
RsG2eo7uT7zvTgQspolZdw26szdVAU1ucwOxj/bN8yzpopN13S6WGPzfgHaNfoWF/t9QaEnHn6s5
15b6NnStlesNnXEhUyP9bJkKF3+SgljqEDffbfvxEtwJyyOZITrTbxewpgIm577AeLK7nyJNr2Mv
4b2mCOx8bNv9XxHAVUnXPqH4dU3OVQBA6dT2cL+xI+OKyI+mMpea8zmK+D3FbosD10u1nOese599
4pz0Oz6PIVKgIi0BUnyZ2cnBA2WqouN4Hjhz0ZDQXYPEUrmBD0mqWKUpaSwPJ7JSLvedctB+pjk7
XAI8XaxVtMk1z5GFu0nQtBKARbJph+Szo3GItnqnlAz8l9qPndbynkHZK8vxUPLIvGuaN8D6Dy8w
ZWUSqGShKsGEISwejkTDc7U66eqkWUShdJPVVQL5h620n+WRv3UR3q9DQdCLhh9d1o5dGPY1759T
4v5a/uDxqlxKWwbc0WsDJpq4pWAGpQZx5Riw5Y0yxg2ST0cMwgWEcQ91M01X5tX1DgA1xCwKDogS
aJgsdJB3+kWSUbKqcKMvd1UXi9CxswdyotyS9PYq6mFlrGl2Sgfb6xVqYDHp/8+kJ6SIdJFpg2mD
wL73Bqj7StTYU1XcWDQb0QePUEJ1MEYKdfOvbBcPRiO+ov7OlW+C341w1wCaintklq8yCyzUy0CE
61wBkvivlh3sZNVUpEXe7EFYCCfLhsasVSv8bSnuPOt1YzfbIIdgv9iEZzfYGVuK/QKWrKL2uGVz
AYX6UZrhO64A8UZfocoNvsbqDWHY4sHeJ/hXTHc4M2DruGoQLn2Sm3edy820ITIEn4576HGQ/hpk
6DAYihbF3h8HCLiYGwR/fMUS85wCMQwJ7tODNY4guPo7C7BsoFqI/vVLpKBUvhtlwPhbJL1d0BUC
nkz+/ofPnM+xz1bId7tU7TyrYJu3jLrPvxZL5dZDzEpPWY1koXLBUME4EfUo2Gn+Tf7nq6IGyzDV
5KrKy/24vcQ+FcFflqZjStsFULtGXw7ZQ1S5mkvZasAPzQBFUC3B9xOiS2n0ZIReX7ZFixxLG9LA
6Ux3UO/slZ0cH9wvWBXG1iys16Okqp8TIjjOdZEFRDjdzJokK/8N8DtP7FyWC1r1pVUXIhZZe6tT
hSJDUtb03lvVh2C3b3lKtE1Tf6sWQAAulCFT48VUdKqS7e4DfTfchSWR+9Tw93BWX69scoJxDYL7
+z2K62UQNnaPZCI74oNJ+90UDC4+FPvTo8d2e6Cq7kpKbKxdv/SqwFbG974Kd6O2TzWc0SwWgHbx
is70WGPtn/bM6WIlPWORyjtzf8ap2J+MSlySWs/mMmvCzJlNHtir4CvDIahAm0XS5lxYNGPVR8FV
jPBpyX/ZNWJAE9LG1SQNJBvv6j9Gu4d79H7OhtQmlSsRGEhPhX6KZavTytKbIZZGCR9LwA1+EpnU
Z6M8X3lX/o+cC6gJUZHfOR+1NLaLB3O7dFuZltWAeeBjC6CZ/jhIT4KpdODI8bY7Wq6xQxYdyu7P
xC/49qHnNoL/yCidIgc5Vr3/CfKOOLtxNboviOCdZcWeCI3+qI7q8Cmf9u3O3hlQepltDVPNBH61
y2JoZ9/ky3CX4oFTTPR2Ph20MOnSJm3Z+mSZzliD/jQv/GEstTDMp+5+ZAaSFdRL0aDmS5ypAxwF
SengZmjwFtlsI3A8BMSCpoBrGVcpQlaSwlw/CDsQKgX7acQgiEGx9xG2PJBuFlzCSZ9WaV5t/5dm
qO8y2JNHqmFS5RhCdhGoboi3Jw5nApyhpFAyW25sNVeLO3cTEo7xJ5dLs5+usKeGgWl2I+00kot0
mz6ooi2BPvn/jXlL7K2iRIrDBhU7SyNhrSl4Z87mbbx+5oavfcB0wDSEfS7EFgW72tBLm5bfdYfI
R+0dVUWzrVKM2VNJWnAwA4axg8BUYhafDwa3iSN9qFxV4JyK3TzCaIaEA0/zTpiKoPvlNjrF4dq8
2nteQez0qTaeYlyg0l5Y+owXotGnx3vdelOai0sKK++3iqQvQKSbQZt1lm5RoB24aA5JOnTDASKp
OEDQh4fITEPnQP+OoHK/Yr3JNUDHYG/lIIn3bKYYJ68UQGLTQ4+xJrJirzabTNUugOgYW/AiwlxJ
nfE3NSZ1gVw0jTTRxhatPUaPAN9qZUQ6e56jSZMrEvP7ubK007hkdO79OzDX73jY8F76+Wt2gPv6
vQ6XyNzd9crD9tG5cCJZRCTrxgVZpsNCA6oqpoEioR8bqD0kJte4CO1iRx0RlIoEjgpDmh/6kcRR
xfrMp6EzSahEi8rhvvmQhJIqyPiX7n3DfxZGBAQfHmpBDIrgE5G++kgAqL3N2xff5mfLUqYicqV8
1oFjuvqFxwmzCAiIVPLjzteIjfoI6CHT4FP2kT2RNPBDVRPghKZyTdnh4JMSJjsoSNbqlgqKQgrU
+yaZpnM6sTVs19pAuP0UwG7iFey00Psw2XSM4Nc+uAAdWnOoXYwBUHNSLNmbXhWF9tM2GaFpIXLo
AtOfO0P6kmGeSmqZJ3AaLu0MvKsYFahTswmtZQDJU9xiyNGPpKEl3h1mWWYi48M8raDifUkhA5G3
DnCgbOZq1D5/wEqOxmQ4WP7IIT6n7kTXA9bl1Wu+QcY4oxdAy+61ZixZ2KTikXIcISJvl8LaAj7u
m9pcQR7soJHboMHc/VMr5wK6ZzE4p81vFmrt9ICbtOccSS5eON7b7V3VB0ity+iYzPj43a+qqY8X
FqQG0lT5Oncz5i4j+BcE6ep9PHuBUaa2IYqDc7QjDxM25ZeZizq+pnxCRj5ECaAvwlzfZw9VaVm4
bi7t33+YLgmByJ7vuavy0sxDewn/FKMZaJjfE2WVYxsDXzZpG3sVtnS+yqC+V255Iu8egUketgNb
8bMO7yh6/RmyoNUzbIE8flgZQoIDlB+X1YQ8SPLNfB2OGbaPgX5lxL/Au8XT42SMup2prLWq5aZx
gHUdljoo6ESrr60yv3HMUCYUEzd8huxEAPt3RpYfkq5OdQib4TexakSxJmPNkANG95h6wk7gCKTx
3+l3klOtrGXL2ynmpYpwtbdifkX3vaC48+ovQ9Q2n01Kf4j2I63dHNoiF6JvF6yqdf59hfqH9p00
YC3RfJUBqv3AS6Wsqvf8gTfUcm29cxLydO1xQ5Tc948Pi4WTWrGdLFtX0SPdIyJy05X2c+LG79AF
NqvBOLrbmaPdGbcIrQCqBBXw9gi70fkC1vzsJgthqtkdokA6ZZ5EN1r4frG/s1EcH7orGWDgaPwa
JfsoHOqVsUXYV8UHcmcjGt1pHH7K8GjSUoG4GSaNgZ5SCmsq/vxirYU+4+BreQ8kTRhX5TL/jOEr
pELiDjQrJFpFIfXxD+RoRxcyFyPpbaP8H1u4MQw+p8QQES17UrNz4dQiHfwL5xjPEIzqAvdGq91i
uPqL0REX3GRLTb9CWk7BLjmoa4WjL32t8pZ15ahlKYt767JXFvy+TCSQO9d0GvHPyQQocpYJydOA
++qTHwa8DNLvQ2W3Kz4jJOhbraw1wXqjlaXnC5ihSHg3RdDrHaAIkTxnjyVx6fvExPefLzgGY4+G
6tPPgC2qc+ZveQypOJq3zryv5Q6SbVp04dzurJF4Bz5+yI/aV4YKDxjNUTvxcD39U4DvYG2sz0ZH
ZqALI6FnPvw02iL4sYi8+waJFyrmR9ecqak9v2yNy0s7/vT7ExC6EMSoUHiTf+sFVcfNixDaLU/l
PfeH0CNAyvfgH82xXUQfm66WGFqTUDQCS7AdbKF6A+NUrCPGeC3uuRJ6lPDmuQ4mISKB6lX2W+BC
BVLMU6yB5f4uegILNf6IclhqfNq+ovoX1QqczacPCYL+H4p9XqY2PxQavTqDZF73Uocv4nlFuwkZ
5nGmYdvpnYhvFr10LWJmjfAo/xboNE1u7V+9E8hlFvN11d50vBJghDAtCknA9Vl9AI+991YUeVL4
rvVQr0Lyw5LW6VuW7fDiWxUx30uR5gMEWZNz/1hwRcAho81rMCo4qH8OQ+yoP1iG1NAQN7EOKEEa
NGa8aBMIaIu5IIU5+FnIj5I6mvDEZLxNfhzeT2ktjmQRUKerwesMvwa4prGBz82ofMH9Q36vacbr
UQGbte9yWyjrt+iY5spFAUwbvlAql+6nUYp/LmeDJCq/54fwm8AVmAvZEAcU6wuyLKesaLiP4gHi
Y3ZF7CK6lEeaAZNqKnzzuX4D/ERfxVMgXVa3+DIIhYqnJ4KxjXmxfoliDa38yTm6TZzWdcYwXy3w
iuOk863Lit4+P3dZQ5Z2qd+3ev2Jxg9fsQhsy1nF6TDH/WVEW/z3XS2GjHLR/fOy6/99QqLc3u8i
FvpZjl+rk1bvbChgqJPMal+dQEjMAECqJiCEKLd9ir0XcPO2TYi5AYsi2qWOWbqD5owoVwxR5x7f
gG3Wz/gaf0OyTFX+t0J0K0nIiWnbEHkzMCLErC0eKskcUPIVdd+W09klCgsfIvcRET8c2l779nSZ
pDf1e35I8ELcoe3n5v4A16JnkcWFBWYDRQ8ni+1WLH5kLa9UoHVSOqK5cjb1xWvZMo1BWL4kwtCA
qRpIz+w0FHevN52ld41VZt4N79mrHYlKPR9Krm86C+IwK8Q8gikSz3QEVgfOfIIgOsCEOLYqLqOT
1QkXoP1GmKVPNlET5LHDWtCGg8YzGNN9unmfU/QIErrWtz2/TT7RveVLgkuOoANuPf/8UaWLHMHX
O6gIYSJ3aUGceFtrgtOc0iw/tqzLuHRT1Q4buw4V2ii+nyDNV39n6W+Wn3Yz3PhYR9o6Oyr14ZhD
9r7E3vy9eyuwc+5+iWu0qJ1/wGY2rwXBjXnwkbN38B0nn1oezsa6CU0w/oCbnd6MSQt0KyFYJQoa
gqrGefWMov37Eed1wn/AU2SF9H8xe5J2/SF5xVLI/UAHZS2GLULpVzHj4qpe3tnYJMqC9uLnzfzk
IhkObSH6QwaaoyA7H1GVX4eOPFyp+xYP1TRXpzHAKOotKNFpFVfNMduAonj498UOwihgGpKFTn9y
d6kflQxxrOgyRcFzy0Ukbs1pR+jfgPNFMA7YdqQ5uHY1rMNvBQv/wDMWOJlyiQPLNEpRj9bm3M8g
fIeRU9FYlQgY1pn0PzqOX8erjnmg4HhH+4Y/318+m5FxJwgSlqxdAoDXVju7TT/aJUHY0kKK3nGW
XTPt411UEolRbQGtSpUeKToHdTO/NcvNRb8oi/BULZHn2UmK5/vXuVrwq2HtQnwCjSgAlVkowlMM
uGShdBlJge+AUBJVIsXDDzZMJIgH+/HlwoeiR8OP6Xl13dsfynJQ1ffUNwoP5gq/0zqR5R6xX9Tg
+DRHwuSLB5OU2XkViewvBzxRzUUTai7/1BvZduVIMqFAvGbY5/W9BlXFGbYaVzRiZf+Hhrz9am94
ATPvtcdI/902d0cncPczoT6CGoXKKRRdtmjo0cHoqEFTz5NEciwcZI1LBd0NfGxI+K589ZXdeEbt
aziUxmaFfjexCE0Dt+VW4MhncXslETXmWbWWn14iyDIhjL8jKwhBLZGpUOzXt9PnqcBzAy2s78oM
y0PjTZsr8d+t7dDVh2wVk0Z4ByEYUX64H5MCUw1Y0TFpQR/PloVKSbwPGVBy9UXogUmV80iRQDTN
GvDKplKqqFetftSsyt2IWgls9hvqX4JwSmi1UX+rDbGZnGnjv1P1hqd6oYcgcqvkaJfz0MKSURlm
teTqaejXpNQ6AwoGA3V6xIPMTItOjp101KjdED4MERs2wyopX1OMtysQeaMhc+tZkrkxm+mZAT66
GxY674BmDZpFDVgLSq+lbdP6tLgi1V4uXm3zL38pml73+FGjVuWMdDZkHYqkYimu0v9V1LUdowsf
JaSrmKpEAg1b4nCFEoyPmd8UpY3T/53640F7QYNNeKx0BxCFfxR8Kisk/FhHnSJZUoADhCZJ1vqO
DYGHCftfSAka9a26NMJCXUs5i5WqCW09T3YdgN2ZSqyrmx643wgBfEwdxEXWWxzK1p9MKScodIHi
VOPHWyH9clJSLlXtAc2TbkotvnE1W8nFiQI+0d6R3e4OPPo7kyZXiVdEkf05aOIqVncMJIoyYkKy
yGG60gC5bZVuhkXanyDv61MXm8QBjfqiXlHLiJQKQUlw7OwnlfUFVBbdi0Rr0mvAyJJSfj8Oewc8
Vp8cR28YdTpW1Fr1Mk4z4w7q9Q66JRsrd3IipcGp7r64S0OhZCZLRlZEHWtuZqAqED2gpXnbmNv6
5N1F8fYi39IG4Ohpzn0zwvm1EbU5hwMNUz98mLWLEE1d2hearTJ8yOJS5ckUZBo7D9b44AcdhsNh
QRdVQaYc6o2Hrgw60TySAKEOWn6gAHPzKnaCQvEQytXjUIDvcJiRLCxyeCQd+EIx/lUe9goybkiA
3ckAYt9JHbV5PzKKJRbQh2B0nc0yIdWU/1KMqdjYmwdNYoMOCinEU7OQjw/P7kfwxtRO/hwCKjzA
VmaPn4/KnwUUKIcVV3o32mMvRIMJECK0NR28tLg6PY2VPFbsx4a9kNktrM+eh2Qk1hQItwFYzCaR
yM3BUcIqXjMIQ+msgJkqa1+J8YDaeKgNZ4Dnca2Xe1La1vfwlIkxKVLd5BCeAgSlQ0BvSxyRqXed
k3SHlYzg7bun+q4ZNeHt4g1M6ljQH10nJJroMru5kKmwhQS3okkEJPvd74+vxpDAbvlgdAMXubmt
UaRYRb80r1Bm686TNcR5mskIs0n93o6Pf5xByBDoqPGPH1ruaA4dkiQp864S6Xqg/3oUqjvWwt7r
Aqk5r9AxEegKyHmCANsOPUWkq5DfnVTrfXHCPGsuFcwvw/Od2L+hLTKMBkMBjAW/kCQGH1LYDr4D
+LIe8GVfpG0a0K95fGbR/2kAdhqPa6MB0OLgldbKUtqqpwbLXPD2H/uEfJ1xt/dF0nLoQV5mcd2K
GBAsr+3DUqM0GaUSUWbrbx8UzMwc4WMdBLNfml3DJNss36HvIwu2mphLQNYv+kR/WMT4oy9u3hN7
CThr4jf1UDCVPGnMHVYhOAwVtxUS0SFlHnwieGBxKY20XdrflfD7rmcCcreyocfQqaS80sYDxap2
WCSH9Elm/wne/Nt4Bc1LnXKVC8YmlRVhl+X/pw3brT9kMdYliyIS2CRTRMJDcMMmNmJbRo2OmmEb
WPnhaHRGTIA3j7kuvDQX1xz1tX4CRpbQdcVU+67CyCawhCqcDTcZ25MCPnk7UpmWzNjgA8EthdLw
aejL5Ox9uX5ZJZ9It1Er9q4csSkmRXcpK9jHONDC4L8Pnfztfh57PdkSEbuk6sBDJ2xUNiMyMm78
+udrWCIfhPHxeSZDeroXH5WrGCR4mz+Nw1zH27tZz5fv/itsdNDxeDQL8I1tu/kQDH8GLROsx1Ej
AtrSE3OyhDtThw2lWClCz5tdCqui3aZV6dlIEPQThqRmbSI+x7PdXVW7cM/Kf9QHArFRVHEmoGkw
6eitBEEy2LTo42qK0onxeOWxEu8WzA2BBsfYdVHpzU2so+uIpEgBrgzhYEACPOmhYdW77hQnXPoU
R7lCZu3BCPU0vM56LPrhU+/gD9tAmMk7Iej4kX0RhzGeoMP+oWMll7prN4YiGoglHxTkeesy4mS4
neADcwt6dbcITxsogc79V7gExIKzoGDKgRzpSWmTKsWehTWH01merS9XBweZ+iJwBQK3IvXsGdRK
e0hYBg7vs7ZVr5kLPnjKJQ+ZljvnmLjaIFhTdZ51zvmgtAc9LnPpcpzf8dFSuFZXI75bNPJPOc+C
2huvorKbiecmHLzrmLYLt90YYF/AUgk6PQpQrB7Jv34yiQD3BcWA31Q6wNplktqc8dwI+D0UlDPq
UmIN/GHxHIA0OpTD3USBDDlsRzr3m0NScbsYYMFyc0FNYifYluWt1biTX2uLpWXNGP9J0V20Mzei
O8+2hL6/Ry2+vOCFAb8oUm2cri3nkVy48Qx+WAB9y07K8qUHDAeoNbYCb5h8tWGIO7FsY7te6tCg
ZQR4GjUdRHUi/sFQqsXSZ4DfYpvf2K2DVzYl3NlaZKXArUmu3K0bJSZGOKHG23poDiEE+RLZyDRD
Ux1PqYM3RO1Nf1VefTRK66ABREm7sCNPu2kcsYcmRoTsordynKqHXI437wOF3eaTVruZnWF2XxX2
8uS0HseNigyUyylOKtCr3DjqOZNvH/jg6YyYmJFVT4xbFrMXllERrrZ8tj4QUBWQre/hmTeLQ44F
i6fIjG709cD1X85eZGqO8i3rtTlL+14FCa+66KTpDOs3D1dcsiPzEURufai7IZJxGxrhHT3m3uDe
p0m2fjZirmqdW5GZhQlXLKRG/e+iaIBC9pNZhuTcAUwTzxea0BCm1QX7+aD4v720eB4kfozytwcE
FZNwuUqlQn+USPb3pwXy7BAG8veJx8F5nc4/Vgq7sv0uivrDeCM3ks3KX7uS3NfRNkrGEqOdfDi3
eMUVzDWCxhepw3TSLZyOUq4sjkrgLKTxsu9lM0BWFd+7lL6vdIyv4z20kHN1jwW+J+lubWoVsHgG
dCaE5YWgmYzk887y/B3jZ8TfZviFJHYvQWWx62Gna8U518PZrFtLdCTajGRFXUm95QYe8tCm5Reb
Bj4UmueBmq1NW0TAn3pT/KkWMaEZUk9ZUzmEozNlKprHegsUoVuojh79zwlaiJDkwq7hy+ZI4dsc
CfMwNGCos7GkPUnOVoSTq0TgVMNUPIizvLW8o8kkc2BKx5fkkX0hHuBGwMN6x0MH6v4dIRLa8TTe
UFXC4DnaUdQLm7gqXMd50ojpKpkpuaARRrD4ZdC/SN4Z5hoFNr8hAXswAzcD5/4zwzN8opdIwJBc
nqZCt3JXDVad3sQ3riO6lx6x2hY+S8HC94CicqEFMZMgizQZvAMmo4aUV4AYZ6xmM9FHr+/dfajo
dw90IhgfW86hwhho0IZtYKPfHTYoFd1NtHIOnQ0l9ajaSi8voi3h9Fw2k1hrtnRfC60LRuaUzbRt
BcVriHj2rYwOvDYqIRwUErlU/okF9Jr3VSOMHMDv4we6w66zsV3JA1OnFjZvxH8ADrYW5kxrCrn8
uMFa7Ftt95G3xGdKf897Asl4/lImMZdQKqoCMty+ZprVOqOk2c4t2g2sFJWxYuuZS/Cs5dc15sfa
Zy38qx8Emd+Pt9pP9lxKS5/VAJ2BUwLJ8R0BJ+lBMBYwen7LCB1yvGrU11ccnXpeJ+5hFJnDOs3F
9g0qrmZelZ2rO9/Ecg8Imwj/xdOvQp3xwrn65DMLEH1/iQ+xY+OXKfcQS+84n54EE7/gvXZoKRyz
zBEXsX9aM+mnoXLJD+Ee1ZoHkWaaOEOPRM0OG48yHkOOSCz3f2Adh0H9GKosHFE+62Qto5/BpYqu
JAnufOyso2+BH1eui7K3/Ria3zXJ7ru1QFLUtkFIJ8PJnHOFZIpSTgHl/HX3gtcgVohyeCV9NIQZ
P/Dr4cpQM9mxdB9Box7FZ7GZhIR73JiCtLDI8s9cIFE9ruhmc+AE3jj6edZuHW/aZ8hA6DyHto1r
OBX4CKLQ44PREA39WTHOqB3gFdqYgrC5sGciovChYkfVGlbI+W1Ri/Cftwh2RBTG7639xU3wmFHp
zCpCC+Xq1etxuyTnfoA/c0Ob9zGarfmq7yExhcQDPx0ucyxsCUZjW/jNZAHLdzd5Fx8ucGGXbzGV
FK4cVtAhhWxNPJYsS0uEs8Jkwk2YK/DT2aSVQ95wM8IsJmFdTXQI9miRNSflFXxcKNZV7Nys5/mA
C/1QZyTYn57PIOUkClrGHlJIzg4j7mQG9UXw4eJUcYnACWimaqo3qWjAL3dMEgdsZrD6VLqbux9X
wSCSqla+e13qc5dpszd7DGGGPgsFRZsohfgghZbdI/672GiWDdU1/pW1YWxSKjgGzNmeywvDR0Xf
s3SV2ehFoT5hMUv1F3+SzacAfxX0jYaCPLlD+V5NPEnA08Y6QVLq7AcvKEBLIEFfHj8RtzGDPUxT
ogMXgs8tX8AzmAQWtiwy7LySuq7mFH1ToASQfGazvFOiEOgGi9NLf/aRR2XYHpCpyNRRaPEPRNP7
hRH0VR0MUnAPc9oDx6YfzqcJLu8mTs1/tPwJKndgCNGlCvQZSXLx7xR8b1LnR7qaNravp+Ybj5Xl
32ltvqHzRrs3cWf5GtsaEYwpyzmAJ020Tgb1QDB9R8l9uBp15dxGsGffaTuPBTTi9u8YwLM+UODE
LXPetHR+ttaITfcMjvxZQHhfhfFO7zv+aqbWnyH/K+wAqoc9PEDlyAN4KUiREqVF3oqxy+6QBBeR
GnkPSZmKyPDp8Q48r5AvThmbzO5F5TZRZf+3huKXeKU0pQ3gMKFfW6IRLBb89fqmwdx83reF+buQ
6s9eYxBiYJx6WZTJyhdYTdgc6QyJY0qxLIjbqB9ch79IY092Trn03O2of+blvGXdcqqrr0arVTg9
te3dBOn8ewlttribs4ChGqaohm9ofxpEXqh8SfLyANlZtbnYaCs8ZTFDvZPXpXAWtNeiXFOLvdIQ
yQkn6Tq1n56hhdzKoJzFGeC43eI9tRgjQS82sWoIzybJ9ecWhoGmmNhiG31ogNdJWM+oBbRYV7el
FjvOT1isbXiU7CQ1FcxntAi+K10HJK++B6xJpr0SnJgWeqG5Fg31PjXpuMqaEUkaCXMk2xS2zR87
LIFjEbgOj2eWODs7wkE7FjEsNQVUjH8PqYCVVSSPGew2u1Jcub2J+dkOv4pvIOs2oV67/D6TIamy
O/deZdV2Sgr/duN/T0XfN7d9fcs5mLd42cIL8eUxlGTFOmgezbubWarNL0BeuaB64ZZ/4HI9xYql
LwYr4JKMho4P4A16hfQDRPtA7kQ20c4yidq/tn34WGDy8Doxjx/2Zpf2laNsHo8vgrrHYCdmsoN3
FDn9/4DE6fNEhyEQmfmjHWiMrkZj3b+fpX/6ROyMt+rSAWQBDODA7kv3oYzaC/YX8PD2qcKBmfDu
YI7XzTHJZ6+fhZL+rBfhqCCECY60GoWw+pt3oFz6IXbPM/pPS/jTw2d3GgNmRruWXeTGd/0agywf
YPWLzOcAfEi9NM+ng6zHmDMA4WvnrH3UmGoKbRCo+EHFGuG9QpHygBoRTXLKa4GSYPvqOUH87puC
XhtKtlq04bInZwHVP1X62cYHMAMr2WX0/NEBSRxmb+iQ1aDZrPbZ1X3p2vMUgelw8acv0pRx12MI
lL/Kd+avHjXirs7tdNh7k/3fvHhPWYjuH2EE4fraDWlurquPNrZj4BE/K1NqJZVNHCdycfMRMty/
X4z6uKrGAsuW5auaU5L6JFnW319UnQlp4hTQPwH/kbXSYLhMZeOOegcMUMM3grcuJJBWiMjdqaWh
sGcFnoZER1RQeYp/rCg39DVQg/UJgBIkQVuJe284cZ3KrcKYid66Ql3yTcWzGTyMPyeeRmChDB76
AkbKol2KTEHH5tjiZuuN7j60iBPQ5IskXtLgZr/sMbV44ykNiw6fvwaD5Yw//cYkXlqEAuO3/Xbh
3N7N1uMK6P6pL9QOfgCnSXZNR1olvyX9MJebquFKe4I8WB5H/TGmxo9IHS1a0q7o7Ws4JAZrNNvS
ROWHYmSgK6PbfHUx4IEgZrT91CgPTEB8NMD3+bvMuF3hz7XLBjUthJBpwTTvIMyg3Yl1KtdKfHcw
sM4yAXcddZj1ky7FaHDilm7udomj1GrCjLDxPPfzY90q4BPWcchYq/oB1rNU7RwZ8DYVmssynOxt
N80yPleUadA7XTTmESe7FGaKfX2ufADnaPDIrtQG7AQnf/SU+px1nIOGYBIM572s68BAVemm1UxI
Q8ZHp7gzuPdXhbr83loCi7Jq9VZ3PPO+XSJYfsurpyUPoAYX+5LTUYOE3nOQqN6QjmJEOdgps74M
outeHylpGwKjC5fdyWhRNbWf2DxYeI4bY4Z543EzFk7XUwCi+NmSymW49949ckXvxEnYN0fejin1
gvTP/cSSfxgJQIsLw8TesrlKt773illk/WyDBkivtB+++cxKthKWGFCsF3JDV4CYTIc56g+5vLoD
5PvEJWb4xtgdwsf0fR7VCRzFu/MKxn0uvwkv248hlKybauq5BUeuuycN9+YkSHmubJRLhPLoHXtj
SACwo+EYwYrBYQpdDeaxTGd6MbTAor6QzmY5M7b4aFTFNY0JDSt5Gpxd9YjQ6WAguiIW83tOFsKT
8ani/PVs/8HehVSIPOnlKmbLWfx7j6EAWHzEwhDMRcy6Dv4cApFGV4GtIx6Huq696XGgtIP79MAp
grCcgvWTqplnHY2fqXBzukffK8yj7g3mEtQk70obXlNOjMv+KjfID4W5wCDtoI0x0SfE0BL9FhsW
wq9G3rINr690tLwHfPG0nSGFB4jkGxFWl4j2ajhfAZXBdzr6oTGJPPOSTY7EJSEo5p0D5axzHads
PErMPkD9hFUNbOUnI+vsw2OKAAj655ceJ0ecFGguQGNOhRHrO6xLEGFYkaoEvT4hyCrhuaEpaWQJ
lSphCHwkoWENa3m0u5gE65vjGlJ9KCpepoYKZrBr9k7veGxNbwhaGW2tWHirilaEr3Mf9kht14p0
LF+ee9R/0O24vr7J3At85xtpzMG5a/skVmkFI/kjA0KLceUq8YzALzSTNev1lJsV3Sqahb0QVjwz
AbeXMxMYoSMii7F8RFjOQnC/+/KfB5zXHgwzl74IOGTa41u8H4AE/W9CkTO9fFn1woNnKjnmbu87
KDUegNmoOzQAEFRIuZ0qaLYYGZs+MojZ4q4F8PSVasHIqsT1/k9snNMjNEUaeN86PW3KmCfGd8ML
7IOCHpJdMdbtPNg8ry+urfD/ku0FO8LfwMujuFZb5WkHLkHuu13F9sTjGAg37CtUA1SMw5yG6sRD
8ecxRcyoyDPUCRLhgfcg0KAAEF3hSMGn1pAuCgIpOao7hznw41ssPEYLO/uqc9F8HiGB+B0EZOmz
ORf81jCeLXdqXGff4zLCCWKOo7fWM7z2CLHAzHRBxwNLgQpnBWD3e3f53Sa3DY41E3tGzjZbXeT9
p7ZNNl/fT6pz2YEV6yTQmVHKHfrwGB4Tvi2IwYwnAZ1Gpx2I4KDNp8f1/45oRiM4Hu8AZdi3+RKQ
nKdWVtlClbt6hbFFbGTuCnXVMLxrJgFzs90qSMVhtWsK8qPdzOcZT3owja2m6v+GCnioCX/L5I30
SmT6kgpEpl+/ssNKPTwGt3BkfKL0XFZtRsoiMxKXHhEwypgYe9xwVPnvXvIiH+2zEUvbZUXk+pgA
Fem3fhqlrLso6+jAqurwB+GmK26ChGbAUpeDvjLn6YBHJ1TbAOX2xZamxZOZ5PgEaySxtdoXXTZG
5+4Oe5nR1ToCpFd66B496pt4z2d+09zORRrCDcMeucxBkWoysJHlSoj0A96tz9DdtKuUelV/h4x/
wfIZtVKkYLHzC3tWgFe/XML+mpi/KG/ehKygrSRLur9cTiQ4Tb6K4KpV13tRW6ZiGCsrb0sswAde
M1pveN4nzwdRWN6S2MHWd6EAFGBTo/FiC5OM49TObQYyf9/wzmm68ska3R+/X8fcRUcxmSPHXmJT
zciVTjw5mR5VG7e/k7i84SGkr2TppJP8fqEGKW+6V1v7cytQOr5EDpbSO4xgrCld7wjfILH7S4Vb
VyhfpigmFKTgUFUctZexUrjLa6z/sPJzKcXcRQLBbxauW+y6t2xFlN0TOp723GSOy3P3jiP+eTeo
AhMabT7OWPRr2dCovrgtEHJirjw5KFDoRoJLXzb1zVhjjglGXlD5NkyCTMpuISfSHVeF0Q95v300
gZ43rKhdu+TM4jATTvgQk9guHr+bq5tV9vSJQZFkSCwBVpYwmlGReIM29+2CzlXP6ONe94UMw2GN
jBbloE/euu8oOPo2Vjtwbi1VucHIfo+KrtUhi+xnSivEgkddoOOGWZqdS3j3laPxptbo4RTD77MG
OPitaqhQ7HuK/mTeLddv6SGEW2S8zUbL+dNMoRoPdO4DFaa7KHUQRkNzPCfM9mKQM+NolUVsVnoy
RZd8SdTxUsvsfpyzsk/ltiv/9h659NTfE5zCQKTILzAiVA6vJ9t8hmcZtHscQ2uOyzYdiOFGNA45
GQOFyB5/Vu29tZgaUcOSxrFPsceSwSqxbJgAC1TShzLs8TBH5cFdWgr86qmfrJKMT6NkYc1JSoni
4ADlBl5TtcqlwJcLGfjGhSyZsElJKM1WwH6Rfn7HBAuRK2fg1X4jvklQt1CasjuNqFVhG10zTaos
GFOYVprDNPx4jQgtcZA+hUbMXisMLcpLMYzwtg8FtFFFNtFIf96TVvFIodtZmNNg/T01iTKiKlu3
V5HBIVS4P1/V/UdBss0oJA2YKMaaSdazsHESvt8o7jHGc2ZERJABihoe774aLK0SHlsT2lhcEKUc
/70h/cPti9k6v5LKUoqlQo3i6O/WBEflsOJ219WlSt6mn0YesTcbIB1JgoGGQWpMXlP0UOubDzWR
cxt1lKdAYOAv//AEskLhmai/qDOuR+ypFEIvIIonqeTh4dWItlV0K92lI3A7B82NDjIsYbllkKa/
bMLDyI6mkfPUbgnk0p7+S8ga6b+yyDL9dLRtAtrpOyHH7RU0v7ohaU8RAaO1vBI+3HZLzcRPLMBs
oEjXipOApw/dtrKMAJ6Jh+qDm0oJ1npZGUP0zqB9s1Gui6bkXFrHGCKHqpyZyiT96tOifLEisgeR
vNzTYnlhE5MV+MF/YJoBVS/tyLCZ375r5WQ/9OqGe2NCh/ulJ0LUmjdojyk5+DfWcZICYDKW2uv7
VB2/KWmkTMYipZxLJYgFkL9PIl/FFVScGuGSyRFEfmyfClMbeXOFNHP5Kb6rANq36WE7TLbiIhLd
KOziYbn6sgktcyBzjoEhWunnOQKFsTd1U57j5hcIekBnKac1QANb5b6t8rvnY2o/GZJO78BK2V52
fvjU2mahIyGlHK+lzyIHa01Ci9EZK+7Iw6IQtYA1H2v8UBYpfdYxGNqGaVD1lUB85f0Sp7mT4PHB
bTc9TkPI9A5qsvBxBpKs9A/CLCNPwyVvG9hgV+0v1f6ScrmUEDNbgy+ogo2rbdvZSgw2G7HBeLmC
culDzHlIJe287i2djuXgxCEtz8/ebm8NwQXqgSapwKQwyYljxL6MZzJPbQgavdAa14WaSNE/tyPZ
xI+9jp2RHa7qHfazmSRcVqm7VbPcFkBK00C8i6yhqLI7M7ITmxZo0imxLlcGMZq+LDTG0NnOdSDN
lg0J9oYAgZikEGGzd0AAWWQiDbzaUMJNGI+eYtIWShJHIlIC3yhn1q1DQ/7j65oEG4t5BeLzB1s2
vEHESyGAfiEDjaYRGLoSj2dDDaWCuCPUKfZtp3+CS2L6f/E4aL1scg7OfYLbccWkDiOM5TxgUjPj
KITK9oeiIVHaGSHCApDO/Vfsc/6cNtHMoPQXeu7PM93M1BdlZy7FaQiNNtBeMAyT6i+HuWSjOOIR
YlzQ0eOWor7tdxuvEWbaa1LBRwKGRwRjwivu/GZKWvdBCPC+qgcZrvKafc+6HhzFkCdAElSwrPuB
ydQfj3vMpLAjdcE1K9M/GuKQpQ6Z5s5/MxbfRlnep3B1Xx8jj+FnIPwf81Uy4qScsUldtAYXQv8q
E2zxKfPSGSHgvIS7LctPdPi8e3hJ27fWYF+4zTMLR3a7h/dzNtiU8VlPCcejaf3iuFKcUNxoHTzA
GtwjoKddpSLlJNnSq2xR5KChaQKN6ucWxjKT26xUFogblvUuCOUy+HxwAOLbomJdIWxgubc1dbxz
IRyPIaOaOgr1fwCXRGRmc1WEybCUniqOthiBd+qkmCZ33aLydFYzV/eEPrxKp9uEH3weZdkNn+NE
xWlVX/5tXFYYw8XiLLUBg2AEHQAsgT+BHz6V3+NR6jMWvrwb8jfER6DjAG6my1bFvSzT2YTqJvMF
t2bXLB1MWJLVQCaiE7me2ibB+UlcC2WiB25nQ4KcyHpBwaHpYPua0n63xOD/ztO5pm6U38Cl7qjh
1wwzLUCFxTFi8Z//8FdS1dE/2aQH2c0XdST8rYMvWwi8PmPyBOtBnHpsez0rEfQrTvWQXFu4kRT5
+/MVNihW2nv5rslHfH+bLKxl1gJOql4Ck7WhapYUV05fbQEUBl598xNzm1KkyhTN++7HAFy8Azyk
sfP4FYZcvXfnJv+Gbtsvf2jvOgiKyhoJc2GXQvO2lNjOO3D19PCszerKUhmPAlAGrz/wuaTHfA8a
UGjlAo6a5IsnsL+fiLVLdfK9lxXqazxhGsZ50FODgzih3sOy+QmWsZs+pRdkcpjZG7JazvbU77dD
3F07aEqZycOeM4nAK3gMIojC35mTN7aMMiM1e5Ssrpijw8JwymkN7LrLZ2HcuXh1Q11eAH7KBr7p
Sw3GkhvNx5dp9nUXHMwwkaa0qHZWh7h/rPmAKp52I334YC1/XMEb5iFgYUG6eb/DVd93KC9atCxv
RDk8WCmqpTUWsuep34h9FyI+3dwkNH2DJMQyYz96VQNtac9/YGFaz2Aa0vugkjCBepUyrb37ywEm
uUzZUA4f5eIspL0c9EJpVIODW5fHVNvT7YioQvdX3khrQXbk/eI5tH1EIioy35csYlxmygxpX/R+
0y4H1rjwUZmvlf8Vhi1oYo8LJCCBgMO+hkxURHjomcBqCCOx7APBgEOiqwqPq/EdFiqonboSsipB
5EpF/4Pyo4eo8YD23gF+DOrcUP2QjMmCOzjQ9wCbBYx/9eeEx2HFeoEAQSdKWXqFbTaD1DQLo7BA
9gnshgygvkPhN5tzgGEcPFMVSti3DrEYTby1B40cUdgaI7xcDQMk9o3I/qlXt0tVg7kjNTXhqe/p
qv9vqWHpaAkBzXlu2xf+qXK4nnPAJpXurUfoGNZoH7OSsFdgsShmhbI67x+qlHxQqUWls9Zf2Rih
qHMdDatsj7Xl5Y/Ww6/bjDLsvCeFTZQZpIAMLsSKOhgY5gJWXNCZFP8fWzaG73j59xA5Cx3pqqr6
b2mffEuC1nIj8GE4R6zJlcZc/aB/cJjgnix2bZWB2w0PdB96zwiiIURTkchu4ZPwRxYcOvoCJaTQ
i3dB81LXDSv6k1Z2yR83gjwvmKw2/zD0fGR9FySt72VqHrqqrprmn9qcAzE70PWO+2UyATRPDO5a
XwZ28Q10oCTsRf6SnqVLWuIOzd3Zb2TxQF53ARewDwuQE/KM+1wJ5V6EPhWvfOL5GUNix9057p5K
SEwV1cD7Ia2tPXS95flkFi3AliTh4ZXcWN1WZZ+pJlhQZymCKhWMy/8jPQdGGsOOsTFYJngIgZJc
CdbOrjiZmsi2MgcF27otWCTZhhHxdKNPyOl9goVrzlTBUd86z+eCr57JYJo+Ittio8Gmfs5QrSzv
zn4czOCl84NNTMMZyvT0mQzk49Oab+CEGmJQbDNxoqOAtY6uDSqOyf2XvtTwXUrMktJq6XFDG978
H2nmFgOp/g25OID1csQez2uixQQwGk5bJjk9E8pZgLsE9FZpWt+EyPrjxQc2Wm3EpOd32igurt9I
T18mplQ25jZ6A5ETBga5xmHNtJX1FouF7q7i2nLGzZ9ZRvBPbAz/jvzaHlteX9CJ5LDzoy5MdePk
8JqwSOUwC+qPZX46xKAA9kxI6aTutGbTP7oG+moO4GSKVnyNBp0+SFt/4I6JggmnM4GxIC930vsU
GcWU0MBmXtrfFaY7j22rGrjeQMYwFsaWOX63vHMO3FIIst0X0yLSq1otrt0J6QmQu46vs5zi+kJN
M3HU1sk8TsEXn6CFGMY0HMAfg1IyccBL+ElVz2AB1HN2MTDV5pASb4oIc6jXVmsGrpUlvfoQZ0K1
47AD6dK2mY0FTUK10Q6kHBalWw+Ixakf7SHBaFsGFV8kLvBKF1G7BZhaDvwETSq4csehXkwlKGGQ
Y1Vo2Kpuwp6E9EJ1rWHjEorh8julfOVW4stSZeiro4Ym1e9r3FxtwokD6D0JkTplYLFmBYJlUytg
yHrqd+DKXddn3a7Gg41wyGd+bYnsRXtHFt6o+kJUry7SLh6/XwwqYAKt5coWNRPL1ay4mFXhg21e
J0pn+6Svpggo9ZxVcrUnwy/w+lGFvz9OQASWbCkLJDowNT1ov8D7SOxVKE1ojNbQ0SC/uNax3dD4
MG9q5kTkkot7wmqdfaolpgvTcHcR3JGlIsNYK7cN5tKQ+M9FUbbhvjZiiisLHI0a2fycMxbsG/5R
PO6JKeB9qwP5eiJl18OF8S2ffjzr7HYgHzecGmqCMdrdh4gTrb6GGoiExLT+1TKHTM9p9sa+2BCV
qFnu4i+ibqvk738oW56s97rks8SSv0xr/Gf3jIhOB6Xlomopd8JA2rmro/acJ4OYlS+01FSlwH73
5pMg1kdr2m/pV9jczRklNWxzI/1yD9kyYnsO2q6a8dPn62MMY6HlitQxeggY+wt3M4FrBDA1/zcB
07S2y1a49R8kcjmWtfpzGaTu11rxIVR6KXJXljRcplh7CPBhubCZVuMZ6vbLAvwhtUKr6nBHcFLp
0B8gRtFeDu7frq0eNDFyqW4lApNgWqo9G1b9nN0NrlMnIHw6JzSFJYfq6XRsrKwc5gXXvSfxlptw
/t82PEfo5U1qqKwsh3gZiw9jpTlmjwLI+o3DSWcfMyycZ4dVQslUQQNpXzoaEtFTZbB/CYzVg0Y4
3Rgw/sELgXOl4nh2IpB6jGRMtSfAD/bu9KMgU2Ufe3yOggXgcjkwDtBDmNBcmXyD0sFSJexuY+Pl
sapso7qIpS9hvD6/iTcXcRu4J7GIN6iO1+2bPtuSF2ALSIlHRthzndx9mgZU4uqXQocWqApC9aNf
JDOnZV9KhwXKwV2oVptx+I2kUtTzUZDJtBTYGWmlUWNll/0cJGPemRBd/Rq+9mQf4ePoPxS+pF3U
vvqDKAJ9flt1tLHoiU51AZla61wbpKj+QSxSMtduX7do6MZ7oME5mjwGRYSVQmILLyudviOErxau
vxNVhHm+YoI/U6KsMfqnrJsC4MT4U+jIsohVMCcoa1bt0RKTKnwjBPro4sAkdD0zpcDI74LSCR5A
NutDt1KZCaiZYUPcMYa9ZDUjagvWnOvJo//a/Tdr3y1i2v049KPLpo4tq/BAcJDa5bY7fu+U1aos
+7a1W2DuGQX9pJnkgfpFhxjz10yV/oWIyCn8CV5tRyzBovfyU3Tp5oUd0S5pSyZktU86iGtoVXUy
P8hRPapp152cRJORTvSyS/yftl6jfnLJvIFygY16f+1LxWpkIhENeGbO24rnNaaL0HguKT2+VTHE
DooxxutaRlM0K3+nySTK51b8rff29iWua7SBqXYfLGS/kXlTrxgLZOhxr+PHdplAE19BHXu3Vygt
AEdDuGEz62y123pB5ggyKQlGgkL+G/V+PmYUmKLOpHeqNcxeSmJkmWROvrlajjTSvF79KLlUyZyq
kuoEEdHH6QqGrE6coha/x2Wvx8MsU6c3zcblnVxnVOi9vIyZHZPZGEAwy18XxkwnW2THFl+Z28Sa
1liw6e9qGXD1KrL85/NTwwEi4WJoesCF7ZIZT0WVCttqLMiYZ74rGQ/4BXNmX+YbYWujvPcvVnu6
+kendi4g+syI85d0te8csJM4RQ+o9ZzlXooSFlh0yTbVtbCG7vw0ga84/khxKe6dLjAukTcXobqE
Z523ze4yIHASCU+in7G1X1src7Y9rXTeRY71sS+wCr1YAnmQzgptCVQW/7JPF/FVn5JsOkKSZRWm
yYo/ot+3yYHUg1CbA+19gU2sCmdXUwDcsP1eBD+mQunA3Tg/IfETWzcJ53rfkQvc+u9RRU5epWhi
x+bM2qdxhZbqxLl28H+JzZ773rjXsy9oRVg0nE7ZEyilCQzIcrVLxdO1mHwphti+52EF/E8WUn1X
ph4/MkpvI2oQj6Y0LX0yftWSiQPPwQSrmso38fZn5WYqxS8R+x18bc3JI+qukjicGb6VGbzRHy+3
pevwX0irpDcsaYMDL0CE+YF/G+91VMGw4XS8zx5GqK5RNo4zOmwPP+z5UrkSUrUrwxdGiWpRBxEC
nhnsXYdIDQgz/6ualVnfveoQVsv7ZMfe0WyJfuqaWZpA1PNbMxGYosB/B4gA41qyUpC44ACdXT78
ae1sZka91wTcQ5H3MFO3wbeiuqHM2lK6q0vysewaud4Hyi8eiDESBisAvYK28Qka8yDzGr4JuXjJ
iftHBQxLzByfXdn8ZTQGO1saVpouCNyQ7ErLjqaNxDYIqbxY2uplf/21PvHqFEnn3Qky7k61IgUu
y1EfKl5C/ObgL1aEojRXATLA4E2E0Nq+SAZfjum0YQPsGYg2F06h2xYd+jjPRxRY89wo37hIg30I
SbxpNC2nHG+nU+cdwlY4IJeycT1ZG8ynPKzNNqqp0gJLhQKwiy9ui+8XB/4RrYGsFxcdhIlqKZxp
D/CGlI+YpegxwK9X8EHx6BL3sYs+sj92r6MzZEFkTBVHVY7cNwXdnc/41qKlyb4n4aaqkqEWgI3R
xlKEA9dBOrLkyFqpayZ+r99LKRZElt+ldeZTvQVQMW5vzKushyVbHGremcRCy8GTIKEq7EA5NapS
00su8bqX4+gwCvVonKXXGVHaJrp7yvCXarDTepWsdTcgB0hABstScC7nJxsZb0XDv4PKpB3rqO2N
iGhYUokOrtofpl2tTWfK68F9lfxnnxePeFC4YIJK1998h1ODLDLCpvX8SppJS7SNjNrU8sWyWTPh
HRJ4wZxDnMv9EgE4CE0CN7Yol00NwdvgNgC1D68UmFligvcpVNgoRFfRAxgA9q6Q9C8xsfrij9py
GaZvb+2Fh6Jv6piA8IB2UJRh9ujmkzSo2SS15huUsMWUEft3N3op3t1vn2VmflR/I8eKCGIcLht4
z+NeoJewf7Jd4lDSE+uBYTRrhiePOG/JxK4yF3pgCSgd1y0JqrF1FvCkFVl8inuGtKhAN9JBqrvy
uqrLZNn/2HhUI1KGjoAe41BRHc1GVlMDPApR8ogbApgKSwPlLZk82SiRRwr7kTnsj6RVsvTAdGVx
DZ1YudW1osoZph8em0FRXpDhf2EzAo9YzsDL1cr5hs9FPrsNvHK84yVBzNSZYugsVc+0Bsfm9yEa
aE+idJiV+7mCxTamhoDWhIQgv53foQOY1R4UYMJho66OhwAjCqE50I9WVJKP8BE6W5Lz6gR1Q8Jp
qPH7HCkmAZBds3pKLjuZDWTPP2937ySECCqvpnhOpizD65joqH7EWTQ7AUUqDIIrsIceoo5Qf6Aj
uIJfRQPITW9wwJz6QZWssBm5Vjm1Q4ImtIHBbxGyfiFtt+x6BprUs78i9XBE81nxeI3vMXVMazaZ
4KplYlrCuV/qxGzXhSou3CaPYEifxk+2q/Zt+g0C6iSV95X+1GmF/8z5J345Nr8bnHTOAmLUwOj3
uR890sBopIDuIUkdeMx1RJOnZKefLIocw8bp5q2xW+SJ0ru6lyjwvik3yj2kiBS1OTYLSn6dvrRM
F17qf7kQYUpC1+emaTg4lNBiv/Q8fV3EqpB9ZjCD0jYbE5D9HfoUeZU5gB9ZFHbNKRDqMT6O0DNL
49/ieVYXtTq1lzGUZehpT6W4E3+IXbiZmcCp8dLX8ShOPd3M74huu5VzSDpHXRdkQCxxtFMIIFLc
Qt99HoJRyMGRw9aDpvGw4pUWuyJg3W4Lh9mqwNg1YXo1eBry2WEXC6pQfss2JFw2mF7j6MMqGctn
0aW5WUx3Zpxxeamz/cUMBvHHqtxWUT07ruMb/5x9giN4Wy+AJSwpIxdDrpAZxYWBkDzN6p+4HGg6
SVUN3cJci0J9MkmC1ra7vwVNK5Y4USA485c+zh9hLva5FZC4DIxw2smltqGDheb+fMO/1AsuhRmA
fz8EOY9L3hhYyMRYX169S1PTXOPKFjxhnnogSjRHNv2j1amdsMHoMYcr0rPqJyStfG/hxWdRXV4G
sfsU3cQ0sC60Lv5jbMIIFu2SCBTpAxJrQMPA69OjGf8ZACfLZysopw6WNymHZB1yjP8rsaomkuL2
G78PSLgHgupy/jV0mF4bGTrCoaibeA1w1gO25JulmW+pggRGZwC9EOj2UPAq7Bkev7vGhtQ0M+JT
VKZ2xRQpAV2CGWGXIjNrYyCXyJ2ddYmGpM5gkOlzGF9rOSLwx8eScbi9p7YG7ACk0owa/vSEBsa8
tQWHkdBmhGUWS/Wp/sps37F+n3ov707i4edmLwWXpKSp4K1Ce7PRu7JESX7Z6hDPMQ1igV2apJG8
v/mSglfnSkX08DP4xfNfzf/jz/hMyX02TKl8LzCfVLWsSdeFIn5MBpTlVOIbRKrwJXN5bBInfyYb
MKBy5KJAkeZgwUR6M2/QeoLVNaaPYWglBQ6M5hpxPhSkYfFrzA84fVM/9LEWtlOLRlEzWxtM/qup
g2GWhQiakQM3zLUJWkPjTqYx7KF9RbpQ11bjbXbtyKxlt2g5Gaff5GHzidwFFFtw/S3nHc+gzQqQ
nA+uzKbQt6frT9TOpAGX01bxQFnLNVTts9QNm5llI9zACb3lLaECFWz/vJwqUB/eT51uqMlGcfnJ
AFSIb80X/i4gLSWuv9aVkMqhPBsr965C+MYf1iTQEMeuMXvguLjIlIAtZEqR1wzf/41VryrlDvrC
2b2n2keiFKCtyVssKwlexV3nm8vznJStdLOoBpA5LCNkXYLcV8WY0NGovMqSZ/WP264ltY5zzJ0y
iAgfyqRGuWaofrUIvIfngCs+ZIKC+0wSEy1bwIF4tQc8LENd45iNc8yJ13F87fUscvDsxOWWeL2v
dcnffYpZUSbCyfTvJTRGA9WdHjGQsrug7XMPe4/VYCXrd88oWxk8ygJKHpn+3/w3Cvap2ZzSrQ+o
DhBWna7XYF/bCx1nT3jCNuAFqM2VsnyU3bNSl7spTKyNrhKIarm3xmiC7hIqUWhMWLtaAS6w03ml
T/6SFqFB9NQWckt3mjLvNyXe664FIIha/ADNVA1LtCVqzAyHXGdgqf/ItNhsDTbxZupaoaSI7NBg
1hNyq1PL3OCItXjD3Cd+9wuXMkhD7ldGryBHsIdoVLY4fWS1EKo4SrGMA82n6KosdbIMe5Yq5YDP
XzlvvltAoMN2Xf1w50KPN7EkEkNa3477gYmycGzHww2c1XK7BFO/wGKWnLBg74AaEgoo9tasuitR
LRqyN0UDfZz0KPJhPOF30D5NOdWDsNN8LLYec+rTt41c1Ioxd9u19YLYoWCN1cAavFAOKn5OMQag
1Wu063LtlNoOW7S2BBwfQYJJUasPWBIgnk+CUTKiMeZfE1AhUCL6eThj1dJFXIxpjDAddLptsCKy
LdxtR7cWP+atAaK9CGncgIXG9EYNiisb+zn6Oh7VOQL/Op86RQazU6S3b1zwfPITHeto5cfZ1ktn
6PASLZCLztkCv8VB1IPymWrju3rOdkjnn/7r3BInuLf/1orKjyn/stMB/n3zinjrmnoWn+iW/EcZ
gs39jQOpXkRb99l8qiYmjzUibJyP/PRAmslEGg846SnvzAPP2j/c7o68MFR+HaDaogKzREREM/5I
ufeEnI4JocISRRqdQrTn+f/IG5jjor1QBiupvHdrhNkTbYpZFogglNjytWegARbqRC3vb0aoRAnX
MFIa8I6COyNpOoKbD7wVwATHxC3UhOaghvLb98tTmVf+hDtCbNVq6UZ8TfTcIWnaz3jKnnhtjrJ8
WBKUGZchEU6Jp1gUe8RWqFsBdS8FUXXmbfFFN6YMUbMrARvgR3xKs1py00yarJwh00gGNUZYPTTo
HcMtGtHq9S69FAuBRIPEo1k1+cYgAjR5RLR9D+HBhE2qtI+9vGkryPbeIg80PxUTzxFQZgsTwmo7
a3cKzRPVPEiB6z97U4l0OzsJxOdNeCSIRgc43zgxyN6yxmQIuWimxiOY1+OIMfVXl3VTpu/rCA2G
CxO17fY4M7N2dYUnWxJA6J+2skk2DNq6yINc/0/a2NSbCagOL4njdIOBKhRVmNBfQWmBdUKBgt9K
9uihgdOOwN0H/bD0YzJSerpY9ODAooYjDOEb0kMZMY1ZG/4kfviIAcNCgOTPjF81XMrPFwPUJ2GL
gkWPqHb6iQjqA0O/uU6T3cNYGAyWBEHRclffaVFgQRh85RREUGXonShta7xI+/tuVmZWdRn0Ttjv
k+4IBrBh3hqFasqNDcd1Crwk9lVjcTCubDoRKEuNXbc/++tAf5rkmXvZTpSOwXTc458ZRqCkrZ1a
GWns87QWTY3iNTEETtKTn4t+PDDLT6z5kHvy4hay+bkyHuEc4T1h1mGAkPwCs1ggDPhcecRvBF72
7bN8Ja3TrDHPuFoK0khkGXQVvvC6x2pTyvDFcTK350DebrIRJy5Cdy2ghO8wjD2gZ2MoIW8MpTpn
CuHHC8Nq8c79pDxlhrXKtfHiAVdp70MVp6bkAWKDaJ4TeRYypRxtVAO9L4LcIhvl/FEV5eDJyJsq
sjG8GJ812SCoE4akaWDB+SSxMknlImr/7zvoE5qpmf2CTZ7gadsmlI+dnSd8xQZYfqRJeWwvEcG1
lFI/ZUKBr6n86KM6HKiLeWx3hGVQAe4DTcDjGQsuyCdzD/PmRhFYSGZj1de9DrtCiOTRggeSksEy
hgXmgw5oQcxinLdSYOK9q8wKYOBpEs3Gyl88xeG1PQCYfmuuD/LNvkOO4dGRFXQuLq8K/1WxWIwz
9P5c/r1znulVAX3jUWL5jQN1/cFkReV8xrHxEbcCV5OIxwbyolwT9q/hUbl6f6lnpO3UInWBGst6
u53kkfTtmB0uy7STzYSBzqkC2rrAphlZgyYK9QzwRTfKW4KjjcQ/iTDPBX8znj5OqMTJ6JiEcbR+
vmEqbVl2ZK5rU2/ptrG/F0LL2me2ZkHMNII34zSmj9Y6QBT1TFFdhKER9QdiYcuQT26zPs20jlJ2
veiSTrsBgUWzALYsIw6eyXio3uwDebBsr7+xDAJqfEFCygLYSE9qvJmK7XemW75HTtC4jVFG2TxE
9gGXF/hkvL+qAP2f/Z4zalKagd205Vb4jV73XpdNWqcp3d+0t9NzZtgfhJvbkxfjZ8sKqWJznXFS
lN9ASz4/QcPLgeSqdSrKDdf3N25O6MKwtTknfwAPh3bQupl1kWG0N9wXARRDNNxgbF7PuJfF2LKI
4o9FFR6WlnQoObdO7YVmXBvSHkHFaJqSsA3feWXvSWlPsBOr9ZZNLRPfD4l2YmqD98S0l02h9ss5
8xKX59QYu+ejZbaJg/HDY++1XNh0G09IMxPFrPHZZrXUzr0okm3qIHFhC0J9r2aVM1UECueCdnaD
ne9eGOCzgb+fZb1eGKUVxldLuLiGMEkG2q5ThJxDudsKMgU4P8xYld6afmjzQylj13Z7QwTrxLBn
alQCvShidvvxkPOF1rVjAb2vP+y8jyVqTjgD/N1MaW0fvAWnJi7DdLxCbAVTXZhnajCmsGpIC1IY
f+pdPFZ+bR31M2tRXFbTToYHXKhuiUpEfe6sF5jD0CMDx7Fn4JiT9BYceufP1gc3BiSddc86gKn+
4I4o2lvu8HMFDz3zufoA/nRatEU5Z+93OHGD47Dzq0MDFil2eDKkrfMKqeAaZgi+sNDy0GQOacW5
pM/nf2F3G9ySJx/d64QWV5/UyNwGSlhHMIZ2c+Hbz/EpDCzCml6lnlqqvrMUr/y9uZ9luopumZSi
nhxwd12+0ZK5BAD4VmYKHvi6v3VaKOK9/MpSF0IE5pB9DytPeAsClAZ03ZR7vZjlrTckqwCkBa9S
+/+0Da+5UJ5mhob4TY0GiJtxj/21tZDQjPVUSq8czOPIMqZ+LFuzf4iqb28bv4B05PCzvY2Cuu6O
9eBgk73r6tGk3JDKui/akiRzxNYi9Dg4ppqFEcLy1kZo91leBoM3s29uUG8mQhQfRr7YobNQS85D
h2dwhB0K3Ye/YtNZsiwe7t9hwrFWyxXqAfcsiJ99RfypK9VyGUa+BSacFfVJ/6bzBqzPtEjrJGRZ
md84tySbYiz0a0mdm4vAUXT2Jv8pqJwNLZ+8T4v7F0+9W+wakK78UxbTbLMGuQfe5xZZ5zwsVmNZ
eyvYIQwJKS93jFG6SsMZIcPDhmWL1wrhBBqE7vZTrSh1lA5g/p7y90V+Ux9wouCS1P/KbMfOlIRM
u6J7WGKLNjs8xQMSGAlWaHER3nw9fi36AG3a5T+nslkHwV/8jQxJmfULdv2e8nVIDAkGK//VB3ZK
F4yi5tLXVjjaSfu1ZezGUbEpT/nCiUSi0AIlTAYPyHlL/Uf9M8r+PtuDMxSOeAkBVca62KgA0l37
RG8t1y+fiE0OhrNQXRh+j8gJ8GuQGkMNOTGyt5aDLL5F/VsdHJXQAOmuTfa8eaUBxmsFYPmKxV7P
fJtwWvCdFTNd70tP7sZ5erIbFT9kOOINMP3e7LP7Oh0PwOA8kp+dFnqdKpg/FFDlGeAx17Rb7Png
AXJVVe1mnZFXvNZDy/lVTzRluUx9Obzt029TEWb9o6MHtbp881eez5iM+l0zLF5/HosSOsCFKLC1
Ttbtjl2I9dd4RI8DPTXp5jLMqbLl5votObscwjcJvo8Wm7m4nSBVjZ5s5xzh9/o5YXFtFj0AfJJo
cBkj3kR+32GG4/pFocOoLyetfJnzthqWTmwXfVG097CGXqPstTo2NNU92oZgasHrwSk/SyWtZcRP
TibR7F5wnph58tmXO391BG+84r/Zz/HEfMoGpOqSV/eeoJWbCsaIckwfl3o17qMLgEGNSYp+xj2C
ViBvK1/5uFdHIa7snJ02Jx+nylWZ+0PawFreTXXZgTW0P+ElzP5YBToW2/jy+Gr20t047q86aqdN
qisAJMfi1WEqrPjnmFV8L7aQkrFmv/uIcL1ZZwOn7lHuaAK3Bz75tKCaXntFTCjGoL0PofmMQzY3
khW7pw0h8YZLdA+Jq1rSRHKncvG9U3/hmVGUZwWMYAiirFDuYhLgKl5dV8jIyllgl1wCZLviKRHs
N/MaUkF2+QEw1a3QwuYebyUsoV/3ioQBJPq4TJFNz24Pt/zXHi5XG5hrmMan5C42MjEF4tpzEDbI
gf52Qn6iF/1tLNCb8o7c9XXPR4UJk+pJSYWVC4NCPRb79TWweP9FSfHw3XwoDZangv+uQztKvLHl
xB4iJfCJ4aSUF29HBynSyp8rfXuSGnjSRxZq2t1DjBaTTcJm6vAB4tefQ/WaLcNcjvTKKi1BQZfA
YSaVLDAvVEj2e0zPtlGtF1w2R7aYrw5FHgs21HD1bo7IZ0bZlBidA4+5h21da5RNMvr9aeuSmzkw
plfqVamFWpSMmg50bsg0zenjAMl2sxwEKxzwlpYdEaP/IEdT+rRiyqFoMEMA1nXwvllPQJyPkZyF
cLPve76pCQ+BwCIF9oCGkNGrBWkIStQ8jAFkzc+K0Jscwe3NSsqbTqRN16ffnwYxX+NoVAcVSKQr
OiwFzpTAHtrf+gHh1jPqMluRdhTlFHIgRxC1RDraSBLX6t10XTPM4rbY0bwmSZ0HhzVKlLaMFCvX
DCYT+BugLFYcyHMEUyKjX2ZPeIvPBaRbAWQ1f74eEPpE5mY7S4DtLqraxcogHkfBdqYlJWhergw+
CptmAKUUnx6GdEATBIqH36wQpJKyWrH1T5aXMgipVXbnqTkNu989dD1Ey6gTnzGe8LWk77t8nyOc
AzmQl+E7KYO/dRoA5hQpLlWI1yMU9zx9vGXecPzv3ekgUpJ5Mn0omoFv90ObhOYKiGa+QoAGKUKy
1asTP5QT2M+2hdEMotiDzfjV4pCnWeP0bhumczV1QJjJe9Y22/8m6/IeS0Rpmi6C57NMfKwoZFz2
r4b5xjiCSbyKG0QSxdxe8kj1iaZicELXKZV+UHn0Vl/Y3SDjIEBnyz74XmG88CJCHDsuV81UG64J
GaUYv9QtxEUYwpFmMcyy7SaDEn1Lu8E+22HTfJa5BjMaStKLngjMqngUFt16WEZMVwCBTGWiCs6D
qYxOIGO5k3GFwzzKctqZk/yEJZ8FevIZRvQWQDI5slD3Icq4qXpF2Apwjtp2ynMMhc0LsYeFcrv2
FYusVaRVzJv+3Q0gDn2qqeLyZYxQLZrU4XJIKMEx1G0ACE7DtzHYfnabZDB1q9f0HdW9L6RMLaIh
D+8Sk9UwLBWPetlhiOYWp/z2F8Mtcarpk98d3DYrmtqBIaZs7YUI41qIOGcGP56Q2ci7AcM8iSNN
ixKiaGgDAHwZpZnAD9Ia5tDkIThIKvODTywPnK/8bhFSWMXzJX7WKdzwuQJPFVb2Vtuy1bYSgeWu
4LSu0L1oXG4sSh6ovQhk1oOo2VGNc7tBFyxc7wmjsL0ixKdAlrrll2z4fCufrvhyEae36gItWAvK
SqOWqkNReLrGLif9rYbTH5hc8L99SsVZYMeREvIIS3POZEgu2aOXaO4E+XpkbegY98N5JSgFN+mM
z/WHCH/XOz5AYR/Jb6jb9pfG5ttB6f2dRRLOtDvLJ7k41/AS9zHGr58OkP/Q646fMiSfKIeG3zol
qgECU+/sohvw7hjZHABHkbwDxZrNPDPttfT1IxIUFIyYwJVUUX7FwI3mAz+UmapfW7fEcsfx7Dox
DunM8A2pRLrJYX1R82EERBugDKOEKEOy5WkLe806/vRZ6OQqnCdVNY528NaZsr6LqP6gKobtSrdU
Yzwh2yuXpN7j0aSwaim1rrPxT5u4pwLTQGzKnzaGHLNI+zh4RmMcVD/87DunVFAtI4qVYF0slqBS
V7UtWFNoY/tCGzwOg5IuGQRDtvGwnD/6RsfnK/KSoX4v1LR94hZkjVyZgqwHuQbP5tvUJKvGiltU
ZJuePmJMzGIrUBUCJfsveYIsekOzPXMbbZj2Q56VY2JqttridQiwGy/zManwefMzbNeFaQ2/sMRB
sHrBQw6tV5FuHqArQKgg3Bt0/MfCD50OEcrlFQW9Z24IM4bFj6O9FigKPPKGLa/AV32A/wxLR8fu
MvcfribNuT00Lh59sMziVClBi3pOVJse5PA5UtrLPkL3s0GYSyR3YCbZy47L99A328zbnGQQiQSb
by24xEXFZ6T600m/PAP3lwqke1RN1OoVYCeS8kL7Hsq1Ts+I1F68Lx/b5Kay+UjWjhk2xTNtzqGs
kHxqjaqwuzcE9tm0+WkxhU1MpTyMJmy58bBcQemXgZ+0pWVIYo5Uv1jYEoFuWA+GXdEaZ5OfWhZu
vJltMpI+kB9j0KVPNDNxvyKk9biyQqBDI05vWCF9RybN4zEntGyvNgszDg+BpVvgHQnMjvxWOVTQ
TsLKiUzoHQLEOYSUkb/4IUxoPA5ocmKpjw3zMveAuJoXdWp4a6XMZITpOd7OPzBxY0b+PPVzLRnS
koZOyvjmwUsdJniFhjnNVWvPJRo34J+YvBY2nmmlkc2VRfYkVOKpU+7dvZOIXQ+CSUFocTjaui5O
ttY3jZCOlG69t9f1xMZO202YmoPv+A5e+xzvTqykQsBV2bwMFAecpNs0O8QOrE1IUeEUjFZFK1PP
2R/0OqZAtaxTKEtNfE82bqoDCX+dM3VkCtS47kKmyAyDerZP/GdU7lS3GQvjdRYJXtslG8kesogL
sA/Aw3t9L6a5U5EXB+luB8w7KGBGRYKRSjbP87wZ9FP0tBNXqkjvCSVBVlxYQD9aUFGzHmA8MWI+
Jm95VQzpNuVYngPaKu7bb+beaaOLAIV77kNk/nqAEEzKGSZMmsQjiOO80q4/QwzzdBxCEkO9mG3S
8fdrsgYcu6WBXB4TUtwXgVOJw4ZPGlbd3zWKxvAxbOP4W6XbfEurW5nMwYi6y33KkgXkx67NXbQt
i4oMNnxsqIAX2e/YBaO2NB0jP+gqbbR80WMp22w5BxyhuBKpqkXFgzwtaFtGre/xszaZLzi27nIw
lI9nuKJLwcpKEvS1j7JqgjD8sovn76I58JAwcsH1Vr71fIBmbe6u+7VnpsyiAj/RFdo572iqzsIn
a+6N2xI8/F+fwDbgkQbD5qAM/nqD0R78m3GXKmLqjDLIjfFdTRbR90+zynxEE2u21RPpKIUN9ZwU
eWZvDAtsBqY8si01ibBbg9k75dhNrCmyObowjlOMk3hok5f2jaC7LX/cbmYq/ntQItNKMA8LZpAo
tORuTlkqwHcmZGnWr3phr0icjGQ6+JexCL5US0Ecu9vkTgLG/ri/AXvP35//dnbhw7gv1VeVUvCU
clPezBn2L6kHb6/RIJ9IZ07oD9uQrFjINHpBYJlMkkoJh6ax7T4r2h41GFPoirryGlmqKl0Wk5+r
JdailRhrqFJUuG0+8/Gm2qVgBQkAaSPqhVJgvxPuCTu6o8FrAkBQt6VJA5inbSF0ZDVok4Hfr9b9
uyBfugQHhBZ5zT4Rr1/ZaeZMm5vamq3pOk/I9rsta5Swf71qTdjJzE3MsXtZO389yVeWl1UgJRav
YF1G959ZdYvdQ8Er1zl9/MzQc64DsH9P0vkwyM/EI1lfli3k7Nulz1AOm6Qb6mwFFdjJmbHcZjia
cdkAJYgAReQ9bD9WEN+dTrzf+kth7qCrxEYZJDT3lElo6kxkyG9B6A+L7qz847pg8+Yk3/ZrNNxD
nkpXdkHjpRfGwzT+LA5RAhlAS7tv+Xy5yWr/ayoyYDlXZNdzHSCVKE329C1OSXCDE2wPHNgliB73
vf0aC2yQ7aiFkK/OnRRJ3UI7lHPH2lH7IQ3q6tTaWsKMGIGam95AYYq+xma7t6nDVhS6xOfUyEQY
3R+GdMPx/Mx9TfhYBJO4Z/oZlAmiipTk5slXHx7uO2jFufnWS6SdxiWyQLaIMFGYN5Z/ri7bs1DK
gTU/CdF390Yiwo1og9dpiOL/r5MJC+D97dsY2j8M5bwIRCKILQ8gOuOGu9yK4GslKhsEO+sdJCEc
UUVPXe3bmk/2CBFqmtTUE1L+blUvjssxzm0jKf1R8KnBSnbGVW0CNDwn6EFjtbZw8A7TIkSS69YR
/TP8xcSZi8hB2xFG4D5bWyMCwpZFjTGtq/hBZ3VFYyK4zrndmhJ3I5ho0B17Ac0gKb5NRn/E9xvY
r6iqn//JR6XQxsXxQP8Hdesq80fWXwu59OtnVAHTzmTa+YdbMKyqkrCktx6OxpldbqDqG82wHLR+
vNXDpaH6SWJyRKmhq17lPfJbyy9iT/weHVpXra8qa706gnEqArOhN/GjNapK3BMMGueYKrrH/ARC
3dCUYhbH2onSkH3gw2Bc20E/wl0GYh30eaW840YaE7rH1WhNtF6LyM6TekGvmYvz3MXYiCaeXviM
8vt5FEvwToQ4guKlVmTGz809bZho0qknONh9CxgZNXtfrnD+ERhpH1P1exWVxqYmwPhkgCOgaagG
P34KgYbT9uCX5KSIheFmDEsrHsis5VB0ewXwixDcT207lSysNGeFNv8md70l3RaNPXcTWxQxqWWa
nmDxAd/U9xlxmoEItRJhbxOHuN82UR7Dk1yjx1bbspMgCoKUF4nQuqTlSrJ1usAgHgEPjLaKBFNH
++3lkHX8arHR1sPLwcDWdtTncu+tyH0S2VCpm9LQgnGr9jOfCTix+vud/vTRv3tY55dSwCHGgGDp
xCNWL/NIVhuYKPcjziysnSdKQPeKdpR4g/OeM8+/n6RS+R440jp4qc8yQ92rjSO1VWKQUJxrhVAT
/LEpBLXAbVk67U2JcruOPkYrYXitjfB0mGNhUv7zxkmHLWCOykVXlRSymuP3SRWe+p8W6BSue5lY
PetuQJfLlPWPMmPgNCzMW4oE5FGS6WxLar+j8zYIMmRxBRAgnbuXIJwTtgshH8jefjvy0zkvMC0T
Tql6jNrJF7SRAbGe5MJts4GZGT7adpEnNvGTCwxBTEXWb4Nw7HZB952zNCf2tuS2A79M5hoI4g99
Au90INmf4YHNUo/stkz69IKfrWkpYubBYs8eqMIHO5PrbX9Z7M68cMWy7tvuXxcSaimzz3nYY4dW
6fkAERDA+9YAccNTycFjdq3WEi1mrEBfjEVn0dPVgmNEYCrapRpSbSsfPG28ifQ0WOhAw+OALDQb
72bSgp/GSI/D7iT9fYD6xAamS61c1gQkBCiHPqwKq1j00I65BHtwtBNhYuPOw06PsaLMK3l7B+c8
UVw1dyzqKOE34r7mPozGrSRtgCtgjV5HZI5GOLKJj3QqkF7VeqMtdDFrhzLHDtsAMPeL9FmoUJMw
huk1YZQFzqrA5M6kx8OvTkZjWGXdTuQYRUPGqTPYDXZPy08/gQMbx4i834um/TIqSFCbWOFA8w4r
Xgjq9itFAXR5EVyNtNNvi4adg6n1UMOSR1qUzQZeTCkBB2rpuzbzBlhjWO0Cb+dINoZsOQEv4p0g
9n6LdUH+mHEXnZqU4BPEHvFvjwDeRwgtX44/k9ePXhCL/Re5anAbdyDtsuzmsJmJNyalOBtXft9i
wwq4hKqQ4YofBB8t17Tj7DeL7qiUGzPu5QiICIUoP7Mx216GfVuQ+/5ZAZ1OBNswDfYNEa7+7dAW
miNQl4Vqta7hcQorFQz0xsUPG9baLalyz7adDPIvwYBiXa1mHNdX2QkD3TKlCQ+Bg1gLxLH4acBw
95sU2vue8GcNeAm6njuv5MBEeL0y9SKEXBbyOfDcu+92nT4f5co/6rFBu7q5jaItCGnfupO5tnz1
gEmpl7gMcDTsfJgt3SP7XwH0VK60+Q9DusZIKW+fkRmwyVcyk7CvdCv6IACD9Mx7BGDENvb/EJaZ
NeqyQPbWiVWVzsnKSLsu7/rP3N1EZLangyURCESpFgcRiWU7ZH7RFQ0Q8eq3unuE4d+/qQVcR4xV
cbSVEoo1KSods/f2KhgpXDbyr8UbfXYN3taV3D2zndB79Mf2nFyqsyA1QqTu0ec3pE7H2T03eTMF
GYMc/YJ5qCm7cbMtSKwt/TFJeTAaIJHeIZr5PrPFhnlZU2/2X3cVPoYWVJpmvJkVWs36tAIguowl
avOx5xm7f0y+UiJA3Dw3cshjq5wfAKRPQVs9F34MPaQnBDQ+KFBzCvZkBrL5qJoi2AsD7YI4x0TB
04rxVAM6R/z70FWI1joDzYRF1U01A4msfc/yxUD3NxFFbD2AdwZGVgss/5Lrco8IErHTrA1EVb1H
i1ND+37ojAlGXDiaabUsC+5HUV6hygnMnN/Xx6c/VeyUdisGkWKZdnUHiK4OxRHfh9f+Br0dUdIR
W86elUb4w5hlw3uHkIyudPP8EyWR2Mh6Z9ofdm65oALpI28TgGZRigeB89nj3mU8lA7IXT+1/gxT
g3yumXRlBZfkL76VwQm99kmkzJ2uK6gpQSzQBV+qJV/bRUZHPZNLbpND3PnoddOYYFGBHXX0gmUp
gSj+CFoyrjRkqw/ssaAuPbiiRWTdTIsMnz7AVd9iTIv6jqb5wXjUhNgCmmltvbAiN2kN9g2V0Liq
xJbmnR7Msqp/EiYKPRMlKiJlFb21JpgfuqVmNzzwzN4qA+YVT2M3M+hvRup6HHzsrNvykwONo+0r
8Ph8G2pP8zeqeyV5U6+0+Xyg9pbHQ96p9SuKZDHhDJqBvXy52fSPuAbmc1EQu9ZGICIi+ASVRakC
nqZ7IGr8UnOawwmy2dnn1fRPGwFxdDsdrbX2o7+4udJMdlqusuVBrT/v9FdibWeUH92tUS1V4bZf
kdC3R2795klRFfdGhu+xi1lfj0d6nJ06FKd0BGXa+2wtN1FiY/1U7Oft7LUwYhuqbunfJTNZIfvq
dAa7Dc9x4njlWiaZDvX8sKbkrBk6kydEF3Doib2d7Yj7+qVbqv4M61xyxbCIyIH5zgJRPfiN+g1k
e/mrYB34/sh2F0dTiicezioAdhnkhuQdoDhTOgvShn6iRjeIKK4lYpbNgOFD95zqNozsv23n0ss9
OfZ7rvyZMEB3wdPLxxcN28AQW3A+oxMVmpddbUSeZ2hDMorRvBd9TfaEiswyhekDoHehsZD8iCun
Qxe8Q3MG04BfqkkGKPayPNG4sypn3Ew5z0bav7tCtC3CJKw12DdrGouGbiyq1VSRQ1yUSnzjvY+Z
4A/liHpXb6mX3SgSj7AuUpQpzh0xYSrquTQgi83m9t+TMUz5NDrN3wYEQiT5nNiA+SDAGMtp6EEU
FNS+1FbMXoaelJohelE+UME0cRDSbRP59J/OvgBFm+bCNE/gRt1KOCwKX5wAOtzyh/dE5MFFTq9Z
pMO9vAT3kK8MoU6SGi9xaGZobzhWJEfc7ObUp0I6HtVk/ZvORKTRQ6Yf518SF6Sg1gqDFenzUr5N
rcIIi5tIuaj1oYRFyC44j4H/BreGy1yPGRj3qNN1Og8d6K0kJetbFpxaKaoVTsboh3oR08579rSY
D8OSPPK+hyM20/McbydzTgebAFt7KyWYb4P8H1XqCcawtf7Uba3CbRYXHpEzKspzLmBoffdGLqer
MvM2LhmxeeKAJxZZAYNwroKCr5nmeQVyaYXEwCQrvuQyrnrBTDwoYzXA/p/7sWRl4Fgq6J5VD/9E
1cMlxImCXIglGQ9AOXN+5RZ1iaIQt9U0jFy1VEH7PXHD3/qnSS4pw9dLHAayceHkTY0akQa8v8Na
08m8CSL+2YNws49fSss9Z2hgcnMBSCgoVaa9CFJNMLEpXJREWNyK6vmUZeqHElH9Tif9CQppvdhs
R6XIIzIy2Vzxra7opPDPHjgWjgACeLS4hfO5Yt1pinupFlQZy7HaseIO8MZiPZ+xffTHQAsJfcO6
Xlr++C0rKQxrCWcJ1OvBwffSzgku/ZVn2VYKTZTHPHiyJ6MGCnMPF3G0Dz8lOEma5fnUVd9SuTs7
NN2t2Di5JBuzeDBFM6DJnICredt1+hphzh5xhPpfIGrGF6xReGOn4oOSMKOcnKWrw3hhcRtPAGtR
yfdsIwDmFRUJQzO831z9YVGT3/fVTlWsmWGymxTUQV1WjrAqFAsglOtomnVZvLmAtOLRBp0d7ZZ3
pUyQ5H8cViEF0akAqQPl+iYi5oT7bk6OQ7M/nn5QFO1Q2vEZwtbIPbMHQR/Za2hO/WwukghMn9pt
11bB8hO4fBWULc/CD7+coDtb65q3LSL3Z8KBwPE5VxQxI9wVldACLy5qU4QJL3nBPyJa+qETvPs3
jf6O8sePMHruY8Qr5Qfv+19WZBlL3kVKVpULVMgk8P/t8trQeHu+R4w7Becq20qEfEXKxNJIghls
8M++l0c8orFH+6aNjenApSriMYE+2D1xs54/7PxoUlhzZ+eU7ajCQBqc9kD7gNbgizkfPS1VHXTq
mVtHIrsTRQ5cI7EbxVAvdvt/xrdbYwoUJoJSslefUasZ33On54KtsrI4C0PCRwDvfgZ/A/eOa3ez
mJZJDZGPqPI53m2IJ9Yxb7rP7Gf6fabZXZGzYJKWgmjGDjn5wZ+VNrub8BrFyFtToo/RbKYPUGbz
/5cnxmH+zS7t6pGox9lFrSiNrd+3sSUYI5O2DeUCDlmaWmTww9ozEDpfsN5n0pl0xEzRjByfIJlR
BqAuf1C+ZpeaXva8Kx1n0JrbeN8BRaUxiDNxDYrGX7niPgShuCDIHi0UjriJTEbUOv8dqWdOxbIZ
95XVIVkprWO8WGJEDCfRjxRRx2Qa0fxc/rQpN9ImSfZJTiMWJIepuEhGiT1PPMfNJJIfYBeQAcOe
0NfBmPVqTAgq1TsCODeIwyi9WHV9Fqfu2599oJ6vJOxeM+K+f8RhCYw9Xww/4lAIJpIc5S1M+Bzj
/SDqWlR1PbklEoYlP8YuJ3Y+dPAqDk/vzFX4pdexXdOfe6kgD5g2luSgPms+CMeu8ylJtbB30Oxl
qNJEFFlB+QECEWIEGc8HEuuGzItdtC+lSTLoArHRLoF/KBB8PD08XKebY/XTYHzg+4MQt5dOOjcG
bwVkQLhdMA9wcFsvs1O0vJCQjcdrDRniBivdNWlsXzh24Fx07WjVv9kiUEdsLEdWOxNf2lzlmFtF
xTaGKehMP9m6TsMJYr8O899NKIimBTIvkdm8qFl+c03z6sXYoAMn45kSp4mw9xQeiYEU3L6HHqnb
PoFOs5EKJ91VDnPzxlkvEucj0I06AkXGJeFOHJA6H5Cvn9KMHgaCCc9DFGsqxMNYmM8O+GjojQw5
7SwEqhNfvH+mIUDG8qPoGVbKRBYdTRVPU3InNUhOqCcjy02g/AYpbLCEUzuzrQIbPgtrK51b5uoO
EBlIMh1sncLVup53vKAt8o2+nyldAohzQ13ZBr01IB769Fzp4FE9LjYNpnmwnlrG8KEheSRZjvuk
w+B0vqp7ZwJ9DzU1k5xAMZAI8l/NS9DiDYT8IF+gDG9N5mM7Nm0qFeChjCzG75OV7X/luyvN2TOM
XiWRqiK0p1/gKd/evFEpDmssdqT0Ww45aP/V+HwnjHlR907y+GT48Ruk9bOs62DQieiCKqWk5WnZ
1mttjxu60uwXflGS80ExFRZHxcH6UQPNjUIEMKgRawMg20luKxczlelKbQ6Ho1hk34yYJ4efL/z7
I8XGVwTq0WFi5xeCtjMotS85r8OUi69tksy2X4yHtWleEU1s+a/wau0/nb8E4C52t/yHRFHNrS/7
qTDR3TnvEYzjyffHLDCmTvGfPDzFKhKGnFbLR5deWfrKh0V9mrTDMB0UOc8vikZzQbwD9Cm8JjLP
tdO7xrod5+F3EEq6e/pNN4DMfY4FH1WV24YiZAV+loX4WozzC6/XYUiindGx3xQoAXC27Lj00ahQ
fqXuEsGeioKtRQLkCblhJ40w+AeMSbAQroDg/G2tRh++XK8f1oEWijalBIhXEzVwEq+yUSJScpmn
gIAdoywKSf9JegjSptRBSGsclmrVS5uRZ5Q0PuqQR3GgkkK2KC0uHsP2nCCeR9/zsizSp44TG/pl
5errkMs+TUvV+xIBdFLIpjmpVIUEOksArxGswcHBBSyx1dvFubNg6CuINhaxPEkPRv4WnjGO1umA
02+3tFVEMvJapvyoWr2SwzrYsRf6iOCR6WCOoX/C9w1DJyMZvcVPMslC3iutJoB4LlvnH9nT51c5
Kt1YnmCrublMW5L7GKG8KUVR7SdXfklCJRoDbJs8fgWiSWa2OyvHnYc7G1eL/3XvkkaZjb0PN8OV
Z2+hgj3kX+0UW5lwFjxLqk4MzjJEmKGFrr/+YT8UpJbSiYw463Ltv/Jl9xDIkL1SELfpneEuIsEu
JQRlRiHOa1CrKjKK+bb7YEeieDZ9u53UtfEW8ZJgBMjTwvo0qKLeCcFGyLuqsYxI43eXy7kGrBwa
iHOp6wWGQDLdR7IWUpPPRVVRq5VozgFfjhEn0mh5GY4pJa33WT9x3pf1Vs6mxsoJLBfbip2Q2rgL
7THl4loWBsMCiKPicDFLT5tP2pS/l6kHb3r6xCgDItkjinNPwwkEgagKmRsN5fSseMoNW8QpG2wB
S1DH30mbxZ0T7E4nLVs5+fU8mR6PJHgsMOiQKlmbT1U+xb+U4UpqVl5/idFXl3aDm7jp42L1ul1J
3qCShkeveG19RYdrjkZGVHD2+eGzMNtX4E95xiKvlZSu6XfKLW4zedmK7YfRBKtfcn84b0JBnuid
Wrj89FGbvIZE4Xyb4n5bTqpSdNIroTQ0OIHa9Opa1Vj4Be/kyHLlr2Soh7YPbut4rYXmUEMhKNCO
80JDQJsXkD2ZoGz+mPUm2J2csbPle8/Ka3wO7ZcQbLJJhAdQ22qwY36nwpTWx9qfOdGPze1wvSqx
k4vYhu1ujq+WZV99Bl6RcTvkQwOz2t2ZCga2LC6AtKwsQ4u+takVDmZKFR6gz+WYwNfJYBBJbUBV
moLKt9Mf65w0WrVELkTN0rWN1FCDvWVHBrvDqIlag4YEjAOsYi98Cqg1aV3NRMWoxwSqkVqn74Bh
itZH5M+KSU4K2/D20ySmszhuG+Ao6w6dfP93Y7NXpivoHsqTahylizHLikWY3R7l8hZOereXCzz1
um4REfVWf2hlXCIXRIisTc3gpAft5HPSDqDWHNmvCIk3haTVogg2tP89/jlfH0oVwMpSVIFsRf9r
JNejZGCpk6ZgQLis9qyAA9t5cU3OGT+lh1ZEgMW0e0QG5ZKAlnM6SNcRosR0O03xKn2qRQ8oZtah
+u1ZbDr8wpIkF/lX52CH8DggfRCaeb3xOML37uId/VGcm8Ijd7x0LZyRky/bqS1iwbCYcqNBq0JF
qdGgsZGNn33Zk3+KOOaEBQswJN06r9YNlTmKySXQny455ZoUhyJ6Ec5+ugV9SCSAWXYHpRdQwiC4
6xky7464PdznJKIuZDJox6kZabJ8p720AAfQbt14hDpfHwfNFC5lj6XeKamdYSm3+m/9dSwaV6oA
P0MZ8pyRYjcqjXgllVfbxGY7s9KnmLPr6Rdi50FoOLV1/ziI7X0Zm2saZNyzaPKioC98Xaxgk2+d
7MzTEuZsShj3vr4oHRUqIVmiXuLc9HzFoEO4Jt/DXn783IxZr0SnUI9y7xPPqBTcKgMeOnz1ev5t
HlxyrHC3AgvJf6fut83vCOutqw2jiOTzglCIsr3V41cWEyjbWjWDSOT+U5Ks+YHhsRKDNc4QvPzM
kG8Gr/fLnSO3NnKSqxe1IXSfGrVU+P1Y7R3iaaOkNjOre9z2FDhh92cMotC1YbIu71JQvP6lUtT1
V6CWP8ayALCj35+GlcoBpwqwGDBrojcwXkf85RpGgDvgYLGMkpMvHEqCs6XIOFSVzLE36oCIYFb2
URgblNex+ZsOC4xhC4wyQb1Yv52zL28k1LdVyEwWeRgfX4JjjgsH/0WRX/NYxk7PDPF6rVrjTWyD
IkspzY8aOzSETOm5FTbc7E/9CqZHy0Hn2yodLPuyBQxuXvA7EP0Sgud2SnoDmidGAiO+RnCL08ZL
Y1g6dCf46OE71O4hXS+ehavckvylJmmBy0dBLXOKjtjPSML9rc9Y6Bfk+swJwcT7FaoI4+0ljVNy
RwMfTLg12EAPIbLCguL3j5fDTeFd21JckxZAG6IvsqC/uT0AjQUhmOKzRnl4VmF2wclajWhHM9Xw
DG6PZyro/HsdE5TOVTwnHfAOhIm/RR3XZlRFJ2re+YuVggJl9Xoi8OLvkYeBkxx3Esjbl3vtlwe4
m3w9ZiqDeFRMEkyM6BplY89WxTCol8JPmZ94bYmkb4vavJIKjX2Q8XczW9w4IHC/s06hqZoznmoK
kaDchAbgqGaAIHppHmEH08FhKPpGY1v1riqwdlKwYG3kfp2hEs008qJO/hpmp/YcJWWkswa0doOS
dKjvhOvAPSDRHJsGmeGFu443KWcCynob3WTb0Rw5xaHPEMjjxOuyyuea8+1aEcMv/CZP/J5zHAVe
b/1BdtbZXY2T92iD52n8O75N2i6c170JGAKpJ+lELcHyNxgcO0ZHTWjyESV+iq5cfBL579OmbMmI
zjb6OkPPyw2/3s0u4B8x7WW3HzaILerzGnoX01nE7Dg0k/IHgoD/vZAQ+Krswh44IsZR1OLuU3Yj
dIywJYEsXU8JVA32w6UcnczZA1eKu9cGba5H15XcjLwhV3qxsDufNvYOt5RQOJC0B8+NJ0MWSyXS
yJ11IUOEuFfiNr8LLnJsOkHbzF4FGDnFg2Xfl+rEws3ceOBwVY54yZZ8sN8UEgQXBrz1SI+dsGis
8v/NC2g77fu/z1uOta9uOmhxid6FSZ8iYsSPjIzNPnHEIUaZcf23g0NlMgjusw5xwaKO63grbvWi
8p+M27E6KyRWgOtXLxZJDi04T7UTSDiOivJFemioGliZjxbo0nll1E/5AyDDcBxG+RNKcw65qQUo
Jzd/oiWNkUdQycdNlSmhwMNzH9GKDsRpFCJR4aBdSgtj5rXU/b55Jdq6QeGZWvG6uajOveodgXlN
FF6qcYg3n00QwqSA8EYYTgRYxYdTbF/rAfQMTLOgKfF3xiUy/qQ76DfyaQKVC70oTVkf5WotIkVM
W0sjr6uwzhaVka1DCb+Rfc9TVVa+aNSBK5j+FUCq+6nO03t9XQ2EMNbvSzAo4BiTczQkiaZg80O2
JYJ5cHEjQDH8KdIpWK1XP5uRJ5iFvAM4QiLnflQLiWw19AQNIAh/a9/qAnyGllZq8mPafKRzI6Wl
B/OrJQe2bLftdUYkMNJV0noNzRThfOLUv4w0Z4dV1+mITNaKYCCkA/CfXmchayXXYyHD/c7X3O3v
pd0OQdCxZgXmjw6gW2joAsIpstg/c/4JlOytU+jdz82BN+OvnZWqlNqdRJKnzXQH8epwXvaih91T
z4f6TfmgzCOnICp5MIf0OGB1xibphorsBozfpqoGebUj1SEsU0VKwbTg8JTTfmBk7/PvFjbIHidE
CAGjdlzlR7abNCJBouqVDWNc8/7TL7TkWh14gKoDpPGBH+B7lNr4jLENvbCA8d6l6LQlp14lxgN6
PoCvUGh7KGRCCIDRWXg0laGCrJElogT/fHKCzall7SkIpScedJsVLC4U8YwrFzsOWHoKy+VeoXvj
8TJYfEDOWGDPkDVxXF2aBDzD5myZWACVJXwT3fwNR1CuQkQp6cuR4+qMCEq4LopoA+JvsJFb6grU
EdvICIr4mDQS+BtC7nqqKWSBIAR4DvcQSxlJXwcKB5x9595yHw7leu9OXE3ef0ObQVPfETnTtZuN
kMTXaWGWu6kwtRRZ1UD5pd4iXhvsSUSRBMx/94akNAiVXpljf6HXOBpLULSp9LnGorydcs+5HUGC
jaubPZ2ovTHOF5UNtbUOQSDqBaUIzCDzJ6Oj7aNMEUCwv9F6d/unGP9vjF5uSungYMU3/NJ8kNEB
aKrQJLmZ6DDJTtydC21cGy0BHtNzat+J4HrNEsDoEdX0jZQAV/l5Y1ItkHetRpz6lkkMkKFbjkxs
kaq9GPuwfqYO4OjXPqD/bo6/4FKss+i5Rz1uilOjj7C5egtnbdAzT/l90enwdfzNd9JKlYEGBrIR
b0ULjzhetU8wQxjoDoePE0dQeVRLJB6LzkPAiR1AxRk0svY35UbgD4XM581s3msSEgRasa1Zlesv
3Gv0lGA6fDEnEKizHzru8UTY6sGKlMfowFUgMC3D4VjID2M6GNsTF/bXtMDph2+24cRUBsivtSOP
O7g6qcL5gKfy0POonf2LyJtmOVHhfjUilJHJyReUzZOrp/XsByYBlOBgoLIaBFT438UhJ0vRr7NM
sroSL7boUd0iPol2kzd3NcL0yvynRyyOU/4uP30XagATNqlUfv0IcLivqAiJRIIWbvYTexanE1jB
icvCCLazzODcrFJ8ZL61Y8GGDB6hw5WSYePzQrEPadNYA8flE9DiCBo8lR+60f4wXz69yhj/tv5x
ba5MWMkuWtYsB6D0M0VoHTN5zO11G4wTQzJtremCW07bDVBcuOhlCU2U3hbN+PGTvcVFnhM3mh1n
UqjCXoK+1wN9WWDEgo8BoNkvpZswzffBl7oVvPrDz89VKzycozMF48S2+gzepiwcszzWdR+oNOVn
Q6s6DGMha1/xOAFQ2HS+DOe5a2heYFbiFFWZGZgMDA/yuUflYf4n1ThiO49TcKmOBSX8uteKTRjh
IXG3/OI7JMj2IFnPFTExWEEWTs6vUoskNXwbAq686VWzZ3jKNm701jA0h2fuof4raApeyNdD5TSf
2w59eyqyWiPiuvQPRmoLBZl11UEYsAUoHS75BGaBXzMYAR+53vdW7UUGUW7TJlPQvdoTWgVi3R59
jASafBjksIjJr3ArTo14XRJpZn6zmx2jJ7XYT1pE+3tUPNJmMrl0HnoATmQiYbW9J310xQMlq1Kg
KZS11bqwzAaxLH6e94hbf4dtN2XrCYrgC47aUBHKsLfnD9iM4Vr2EYiTeSpW1dCrmH/SlcN2Hj67
jKw1SM0f2qt+dlJLgF2vMgibl33rFm9k1Rs2tDkVl2BwNbUk97sf+Ym45BcIzLf45yGDolLo6voS
w3y7XVVowvNZjnHJMDyv3Jf8EYb5U5psJVkOQzRhp3m1XgmIBxWSoZ8i65zUKD6cC+DAeJ1fpZxt
Te/JGJZIs+pV862cuLbLzAiXbMTGDNdCAKYOPRr56ali5mFd4vrQV2t8FZiMFVQCqb/jUKbiAV23
q0QJQRL0peIpolWhM4inQyqT7GWUWOX5tzrhVUhjnaovzYqam8tHy2yqX/yFOQggOc1LlZ4n4IYT
aJZ4Db0fzLUEIUnJBJxZcpJQpdoVRvH2I0eTO3Rs02za05JJO7+4WQvb+GdiZs5T4Fk7gkjr5bur
LgoB0ZDL/XL7J7Y/QnoWedacz1QBKbUMaQEPHdYbVhCFkbyVSW1Sb7ILh2stTMwKUg3PX+/RDFzA
PwMbqLVf90B3Tw+M2bmn4SQzXra1sFMOS22kVAdkhqdv2a+TPkAez4NaNrZ+w7pD/0lhLBFKnmw5
lMW0UHTnH52PSTxsO9Y+a0cinL6LITQkxuYbcsXucApQ9uaoA9Qrhdh+pHu1Um24/7Qc+Ub8GAts
+/hf4KbTuothSwuVabtU4Ozq10+Ofs+G0bXZaBs+2OTy5AynM4Lpb4Vgy5nX7phptecZ5/6JxNYF
Y92ySIDKLZS2aH9V0xIzEKtElN1opw/mdgPL37TNVi70RQEMuPX9tDu0Z884Q2FOAoAUafgo+UMM
vbu11nzuGEQuBgV3uL/09XROBU3N2/0Dx8CFMQpUar/Wotl4kOPZYxOzwFeXOUNN5Xfvgbk23zyI
29IvS2/JCgnzA3VMKWzoAdmxlvHCQVOjHxycYh0dXjc+fjcOs2oBe3+3CCuKY7lIDl+ftrvtEaxQ
FIBBFx2nKSEgGKRxQ/5T9pthbTk/iXJbr9IOsyE2fwOYRIE//r5btzVVJkxYmR75YCeoFvgBisNd
RoggLBMn0HXzfIq4J4go9AIWJBcXDa9X+hVK1nz1ZGK0SyfOp29uNJwDJNhiVf+Nc9oRrWOLkIuh
0CUJB7gKa/RlcI7CDTFmofahi/cOS0osPjKPGnoentx8RP7rpmeAc0pqzbmpNGj8yEfjaxQuSzBv
x6O/tXNSaOZZuvh3J09TXlrjluWIsq1Ljk8+HBxcsJCUSF4CzHiYh2sgF8YBinQFIC4GI/ycAMbt
o2hphL6RRMK7Fe9+0c4MLg5DXzCPEWtmxlNN9MaV7ilySq8k7arG24wLKsdLtEaUuoaX9Xmo83Oc
4nwCKvNPib7cGdYndpF+5p/8T4lPiRaK2JNTdO0s5ik4JJ5tHhQVBjqopUn1Ezdiak6bjCHpYNM/
5htUPZIV+vS8mBAv6LPdaYMILTxvPTruq1RJZhCUM52jr6mE7DJ8HNV8o1oTF2VatYVqJ15Wmrir
7n37t+pC7F0yi6PoTK9u/YnOy1wFtw9tjFxHXceqH9OzeACdYthCgaVlTyouhQ6OU8LgWzDF/2/c
EU09xIHGiSa9w0JjVDuPzNm2BTzegNSK8rZUQGg9WSXqsVKmDenoAdfAD85x2suvepWXXX67N7Uy
gY7OghQzPlUREVF15T5OaxMlc1vL385nD5ywkCcBiqqB1M/GboGN9CnLh/lyUFLa4se6jFsJDUzP
C7cqV6aBF/n48uX14CEXYS562fIGY1zY04/aOmeVr0n23B66O3A3xd7iQruuU0zjBelrSAzGquD3
4ICamA8oNJmJcuN9XcN9vdDKVacfLLdRA06pkjKlJ5UrImmie/cUlIBAuOLgNOZS6x7H7nvmqqKm
EBGfB8xvr9PbhVa2Q5ax5QtaSLp+L+nXOAW6ARjbX13xGzZmGc3yjAzklKK0O+tELokhgGMM+iK7
LH9m7pjFj7xfgXXd7HAxuo1109UF1ZyWaM9lEvuDpIFr6o/p+W2sI1WX/re6nTPiCmEtKHlqpBjI
l48uiePoqFrSn+zZPxl+zomimn7VsIP9OAoM+Um30U4M1YTvbx4k1Hb2ilFLK9EUkpcyVeqMAujy
pTYh7Z0+qjluyKwkp4FP8N2id57SO8FlhuousJ3WB2nnt1B6eUdF7WOc9KAkHZRTKIty7Z2X+oXi
lYVQFhQCw5Uath2tJR3qQ2gh0SsgkVHFJFJa+f5mkK8Jn1aY57oo7NFWb04TqQiJ1d08Mpg4mGda
x3UbmKihXruhdaVib3oLiUjJxenCyyHqvoQ/v7zFaaKgp14ZXRnJlE0fSuMwLAzUbAD66GO0E+Z7
LNh5k+6NxycOCNiKW5GLpWiOUx7Xp6BZMwYUtYA2iKZ0GVOzldMBww52cuwFOnuwFCosxDlNZ/D6
RNmYPTV+hzibW8ALzm3Zl997lj45SGPE2stu0+mRCqu4zFFoUSkmfLXStxYJ+/BXqwP+fM3/Xo94
L+euFfv+2lBefBmYaCj8Z8hJYUUX6uTznW49Zig3WZ4+K8pkZAyBm9VLonhsgrMj06PLYBgm23Kz
z0ri39e1ZpRDekd4jz/25t0pTRDVyKbunLJjwihGzkjTUuau9GJ6TYtEJXomFtYKFi/h/MqkxbIq
560CyX3amcmcv2hd4p3H4oBrtpN+ZYYo+9VuueItzCHszdgSaPMN965lEX2SeDTIigfQ9GJ3sT2Z
jou5I+WW1yIzFvMUvpkXylrWS5VgYqJ6EvrBPs4PubbrpEUYZBttZEZpuJF/ASKcI+sYl4mJ0hgs
IcQ/lQ+FOfI51TpdBOwUVR9iEBOeMVHfLhQ2OU7I3XK7Q0/LWb4I3hiZthxX2L3ncgEAj3AaFa8h
f30ziNHenBnV8IWLo/uwl5Tw2hs0DF0XPP7oHtd1RsDPn351StPy4IVexExIuF/JDMW4kKFOuejg
oUnH9aPOUhvr7foMs0vhHqX6ZVRplfkmpSIuSRO+DWWBVx0h8JFrYC6D4SKVwdyfb92IzNfyhhQH
mjucovzecxnk9Sz+voo322N3G4Uly/C+AbrWUNjnRzbqKqQj5f5qyMpTNokM1yf09Kpq4plWhpfq
DOfoWrR1h4lD7Z1SvmPlY1ojRoHiH2zFjbJKMPCAm7TREWex93bAbGOcQs6HAh5u5ydCMD6IlR1r
VQdjmCdpFt+rrAl6kutjwyShDPlaNjMFkp2Kl0ZOGE4UqUWUB681rXWLc8hcH9n19C1moSGN0eTo
O41LbLbqYHuxTwoY9kLg7aM7kyOEJO+M/+Uxu64W1LCVxziB34tweRq1xSTNfXq/de7/EZH1/Ebj
QcNKhIEtyjTLYHW1JEvKK5kflxzJxYizHLVR9m2QZrNa7VjbsEJJMT6QSj4tW90AVbPZcD6mJSsq
MAOy/H7eG5KVIaolfYUxQqYlMIP/JB7zIX+bhOB9foHwaxgzfUA7uBXSGfzg/zUuIgQD9Bu26+Be
p7uVjKYdu/6S+lXZeEO8PIOjhhcIZreV/4lcRkaXCROwk1NdYlTdA7Hkgrj3NVY4dCSUNMZa9yIj
L04DYPqXsOX0oDkLeUNXNIIlSKbtxmiGOow+eBDQ1paPQn55BpKXah6+QLa/tKqn1bxZPRubsbSo
AvzwJyt/VWzl3+oMp8tU8jt97G0v2jVBHZRcUFdCtXBPUTiecAXdLgZi/DLC7VNIsXWxim6rd7JF
f7fKO0XgECDQfDFhnMgGfPvaAdy/+mvJ/qljdK+kY5NW8xjE6XW1zJN4+wAcq2WkjEn+f2/JdWYh
ciyMa8Dy0VguPs76pJ5ePEhECAPN3knCl0cwRlG7zTUfKkCwa+UkmXCHuQlx5lDN2UyLe+PDfgy3
eOjCj8DZbW538p+I8b1Mcl9y6Fs32pHVe2S4PTDT1IVXqBjBntfbjmAz/nP38v80rq6lI+mKYxbZ
d+IlDnyEo7Sh4SNQNIIIoVs+c9uSm+HIGVpAZxH78KtrzuDWoQcRl2Ig8MqO3I3EACF9AkgrwOkk
Cd6u3d8eM/gorlLlRSXXBD5KeG51laAE3WFA3HRuGyxxT2EGu6HFA2F8GehbQKZ0MtGm7R7Grnwi
f2Fa3AC0R6Lixq0i8SzEfXLBoIQEA4aKZpTls5DvDbfvaiqH5LjBMt8Rp/BhbV0QGZr1WiPy+ycN
KcnwbGzgnNr/aSwHwhqSCuQwjD2lfiZzsu31zFT4Dmw3bih1kKkMQ2pDVFD6BgGV+V8FBFRHws7I
xp8ZbYsLgfRaascr4ihSsWMMPgMjPQVaewYexbgGp5Sfng8RGsAIy3mxy1R09BUaqTemkUiybOF4
yJ9ArIyADtaAw1/j444C+SSTzHD9sujJrclHScikW6xUxEAcAmkqw/mAHhZNs7shssQXi7VbKdBe
Wbt8X+cWEe5hNxAvl3C1kNLfA7JompAxhbmgQNZ+udZthIFoJoVtABrSQ8xkwJcc9H+nlGxcEmBJ
+60W/rxjVv+9A70j5uzZb8fMETrIInFz0wjTu/N/OjalNp8Wy8fMx5hqrUerBNft4AqBjdzNy2KA
nvB2zDS858HkCFVDq/Wrqon8PTqzmiQc4GhduZwMdJiTXUImPZhhh4qoqiYGpuWWtrW0BSGGruaH
CKXXxEQC2kVAMSXqEVGISty5cZsnGHiMZND4Rq0Ii+Ga91jaUoBmXT2/P2ENHJIeNxjg6Lh+HOWN
16Spor3quB2bhjPe1vfi9bcmd6gPPEBbRUVT25eQVv1lsmTXcI2JY2ZoiNtvwQAhyBDFnH8UYymP
Xbz2DIWkPHB5yKeSoHaUP9bfOm4Bg8oYo7mRftiGrg0NjKk0DQMgtLbYKkNOr+Uc3hDSm1AXJxGs
RtAmYSFAITx3RWTGEXYkPs57cJvGtqGBNj78kF4s9j84WRxBDQ3/mkGDTz7guPj1hFAKn/J1nVig
XjiPKC68Piu3YN+llGWSipdASeA7lq0bTvYSxEVIpOrhgzyhYXNOGZ0wPUNzugIiyQRraVt+IDpD
TKFDTbC6FxDZiQ1g7ds2pZJ5aiI+5jQSdl2yFauMswriWkA0/Mr4ZuwwJ8ybFK4fDIlDyTEcRKHk
MNAoiQZQ9+ry2TJLf/rdvixTK+cLjz+5HdfkRbCPpjcPxNFkCOsEDneUUhnRnvRn1bY78lpIAc3T
+2F7DMbG5QHa57IDGkZcAQ1POvUta2HOl43RW9uJKj8ACe2dDm1/bfz8fz7JM2Yu/3Yq4QsqUrJI
jcdQIzyGjY+PNSOlKRIqyEUJEKiaVP/KbJJK3tfX9Yk4XDNniHLf4w/ApASkOs8HsbuJlySi4S9o
ZCCXtTvgBZpEc/ZQVfxoV4lAVZ/ARS3byDM/30dKiNGobHJbZIAhQaQbAW8GBo+fMFQ5mzthAb+o
r0N+wgX8wATpQyO/cpXiLW3rM8Ip+dFzyJIlo2386H4hYFed8RDTud3FvRhu4IhZpgsq5O+yXWN6
eO2b9XVxXmDFx/dIKS4gJjDnohzBz7gqLAS6HKFVukSqjNiz41mgU5IN6L4X4MYR445FU2CKMxeK
5AWlZqRx7g+TtyIXsOxA9I6KC6NUG1IbNjio01bz9+iS3LpVRUFzsJWf1oayLgxBwI4Tmooyh1Mt
0BiSG8Qgo/CJGntpOjcpHSAgWsmT+RQpsbi4by5ffCBXA8kINhkPwf8bps1lycmFDLCVDaW5ejpO
gRhz/Y7kWIExIPQWebpIwDMj77wznKUyMwHpngZm+xjXOzgP05cnCJRfsByoxRZm/5wdsYwwvmNl
Ltak3AhJHpE0/MdVt6YT6s1WtCR6U++rqDmBHe3appLr3qUeMQR0hYkypaDX6SQxAuu5zO5UM9Yd
fOa1eUhy3nWol7Xvy4DMBo5RYXGLyE5ZOZ/XgPI5YpD4rRgF/xQTxTkji8h2hAosX2dLOgKD/Vsm
Njem6OYy9Iu+fsU2hMryIdr5xZxDMZ9Dl5IZsYcP8hsZuHjFwsMC7eKX1XnMxyupYGkmdWhUsG/E
X0forfvGlwVjbh7ntKM7c22KWNcKeBsJs/QC3mYRH9/OMVjCRYj4cN02Dq5ViAuxBbb8ogE6thuK
SHZUqkFxVzbLdqKrDFFQGiGYJnZl9dICBpaxc8IwsqTBYYbEB9a78JzBfWLTwBbNOO2KeKj4r0jw
/dtzIaiSPsv9utkJWeNLn11suPwadb9u0UG4c4014aOHjTiI/BnfhUipAFifzepqUlbbph674uuP
0px9GqjiuPa5EpzP1CYuyOLKQy3IYTyVwtF7WGqN3mKCtcN64+V7vPtVnZn4EQZI9rYFUF5ekal1
XTf3NPcDojBLWGnofHJklzPWklC4YDbot8c0xk/ECMeKZkokDyMvpoPmznODCYxQc1DU+HjFWb+I
ZpyilJBoNpP7ZtgEw6zf3Xst/pPTnCIRKAg3fCSOTJdEbGlgCn/XBaciQCeVmd38BU7s0vRDxhXQ
+OvojNj246TCJOwuXXog3ecDIVO7ZpcMB1sRwUFlsC49l10v3bCu/urBKfL0uS1KCcVJJVMyveRw
Ebpvak85mEsa91pRpPEnpl3PShqLHTS/vQH6IaZjGl1it38497CY54+HiVKC9xmpF77E0WvYv53G
Sce8sr/TfXdNKJlyLBMdJ9LvlQ4AP88KwZowvEyYYfcUvRrRrMppnJBOEd9SL3/jpSochEugs2LD
02yfSeUftODEXN76ut/ef2EuQQyeD49eteZJTF3HDRkMZW3Gy22ZwQq6+5IBUKdHA478DB9JWpsv
VVwKQm9tV4pC0vOqipiiwhdDcwHRjS89aolCqWsJ/ubPy0JtAZJTIrhG1O2HdOIgCN8ge3gMzHOQ
iNyYXzzLMx/k1dJcxrPQ2bLlCieQ9oSRgQtY6L+aqaWJUn0voSHXWl7P2+4gHu5bTvaHedLDsmOO
wLfLafSFwLYXgzU9Mq/8QewlgBykzf5Ow6t8YNIw417T+druAiDMayt2EBjyH8paePweUqiREiYf
CgOnDHqqIJlFaSeD13hbMkfCQkrM7j2KHgTD5ADqUddb5e7oxKnGcwQsqI+96ZsPiQy9tlho2Qs5
LRIN9NFW0e9u14ZL/lHMLzlJHMiT9l7VgCN588ErHaHhh1+sBaIzZK7YJ2habEbPm7pMXHkJLjNW
VEPwe2GnEofuhXn3S6S0YI+WwC98rPXnbEu8xmTlsq+u5Jg5B4W3mIz76yJBLIji4HwUSQIAVWPV
nPm0HbZvRkLeSzrwWV+Ohva067kmwxeWlP7YvcLDJPNiGuUJf5jNznnFPIHUn6GQKyraK9i3ZgeC
Ab9iX+rBAAFv1KyTHDg8HcW9p0h2R7qKjiKpVUa4ABvEwiZp806LpUgQCxKbibLUi8/Qr960tUKU
CreoP7mA4zwgaOst1vGIajGqA0iOvaadI5RaaSvw3B4iVMwfvGAp4TVRrP6yzGbS0x4iro2lIdCd
seX8ek0y3HjBk/z3bvnYb8S05Nj4dfoe2yIY8D8CCaV9DHCAoblNRn/vsRPYekuahq1YXBJ4cmwA
7yOFFyAWJ+1uMjvrrf/70lVRth8iFSUYydRsgkNCVjffxEkU8DQEIaSma08ZhRGbEUCTQzWTPCtA
RbmPQzvdltjEg5uUbHywO4Ob1wfKMyzoauxqNGZF/ls2jc243gV/YtxhwXTA2kXkhbTqyvET5RV4
xtzKkndhkLSSDSMXP01wrhAH35ICFfSP+DQwjVpZ9NRSSlSX297x/Ibj52FL04tGKXZyhojFHiiz
97eS5FerhIBnLz3bg8E3F1vvZfsSNHEUmrQOAO9sBqLd+3e2D1MzpI7Dew3YR7uMhOx4L8Jvbm1r
ZgphJXit4EOiHr69m11zQ24R04sZ8MnVLat9ef8VV/HjYfLdVCd4jaMYyl+efpMr1/OJkHzY8oqJ
vg36gd32zAb/YEJ7w8dGZVIIDcinrLNOqfbjRBPB87PeyOM7FrIpL1nTZNtjsQCa/oYAQ6qPlrvY
PyP7U0UwFUSJl7htCOtF7U0XIo5YV7k7Vdm97t0cxilHWx7IgD9w4bysV6Y4rC3GHlMYeDib/meU
h4NpurC2R66dLJuVGYDdsEhuzfZKvJKypsCtnuRraLhDXKJSRlRHSJtPCVQD7g4ouBHYKvRxEprm
7gM2oqvuLNEDFhEoHP8ZhTtVyg0uktlxql6lHQdHS04n0L/aWEGdIfBNpAOLYJwidOhPbubXymmV
zCzFM2afxzkt9ywUAEuhnDSNeZ4Avpwpyl+Rh+qm4H7iMlwcvx9j7a/nP/QQ8GoZvuiT3Xyk8jo7
/9tBHzrWPcWZ2SqdtO2n82YT5dbH8B63liiu/Edx/LGJOj/Vz1wQZ0Vtf7Ni50tc9LoHSIMnuAf2
tOvNSABwlJUhpyAFMptR/Y7IXJXbbSXLQ85U+v4xUBXcI5YV0uLRAHRoPJzizFyfjf9BGDSTyfz9
9uhREM+sY0XnaS20iIkKUp4D3FkO2STL3V2i7JWe8sUbFkxQPqDV0npgKZJ+dTn+sb0YOWdyofZZ
tcTt9ehJLMrfTmbLD249L49YUGTQGN0cvfJaPLmE7tiyHKs+7sCuHmv9KtBRwdKq8/4prQALYVa4
jFSd+Ioxp0mXB9w8QOJug4h8gVnGk0ctS8QKIhKF7s6P91inUoUcAYrHbG11qzeYCxHOtqFcJ4GH
ayzm+lK4RuitlVKbXL9ULs1ErUetbSZto4wDgyXepu1wbqNH5dq+s+trSqpyHfhPLq9o9owZAYy6
hhV588FcxLrokc9avDaAzCJGhY2ZPC+hY5dHNxpMXQCpguSCdoZD9o0pYvcx4O3CfWTa2mf9PndH
x5OLyGVqjEqgX2nDI8kO/r6czFmejsjiVpwKBxf7Mq22XZOzqgmRSmciXpaf3HcA3qQz3fklAYMb
hSXXABUUQhexc1kLBESYVwdXPpiBRTaizDNh0gNRCeCmHHDw2OuHw4OVxvEu0dm4u8Ca7Uk1ds/a
awvxgCyq4xkU6Mk2SkZwMTazkJDMsNrF93EmoD/Jod0wxdpITj6s1vYDv9XsUVCk0hEVAglcyiOz
IxsbRwM26+RkwpgSMPl6kkcXhTmz0l19oDHEJtuXPKioraFkdL193v+RhuVAAOBlT4lTztu6GrPc
mh6hrygJxxi0EVrqYS6MW5VBYHUYluykLT1E85GEO0D0o5dipUQd6P3dNpBq5BcpUpWfXIVe9Epg
lmErEZBmWX+ZQK6KDmoXhzmYqYJALljQ4Ot4lQcCbBXUt93LBDgbokOVyOBRBjLxRrhbPcmvpPAQ
vjyBtmjYK58bXGEGHkIwjL9m5ImicJHNN3JsjpdwvouZRqe+W5ewc7nfsCTjAFb2Pzyh5t7QPDlx
RhnJuM1ECsEWyk7ihe7Gu44XjIDERtDpvaIWl4VDG2xl+JOeLZwDENFTwjRApdhfs+nhUi6GZvwq
TDEDUtt9auyRe75TUcbne3fEV9olSpHx+qcdIsIjUNPaIMQNIULvLn6jNRkF/k2q5m/3FOnKw0Yr
103DxeQs6iCGiYbhklp8iv3+WPSMjY75uQbMUeZnKwD+9JTULUwCksugYoA5WA4NjwIyWxQTs7mr
JSrcz4dN7Xjmk9LMffKexi6um/qhFaWcTykPSjHVkR6x5OYw3ja0UHzEaEZHcyfWWoJ/u7/2Q/CJ
/t07xMu15YIh8tn+2WmXBg6zbhgSYciS5YpTUDVZ0miGY7A6g//nvsdJISIuw0bWSeZBPxTghJOn
nfH8xmorSQGI9Ka6ityNz1s1UE8Avjwt5z514JyrHjrNT47aWEhogput9UQm4NbUXJeAo75TGVEY
45eVPbHbYGdOmocvGrUZgqMnsT2kJevOG9DWebu9ksiKYfM00cVgL3qgk4pnoGw5E+h/RQ/F3L7o
y74wpkr28sCJsUCoSrSbEzsRqX7CbQ7jWaJqBX6iYkTip2FuruK1DEf5DmQvHaYBUTeyczXatt5l
58CX1JZXoRJWZiBO59vf0Zc+3sTq6ua4SXhl2pMrQPOA0/ENofNi1ThB7QdpVC5fMCrULLGbdkea
mT37byHis7SGlyG26B+/NQ3lmFUSMhD/vxY9clwUMBAYlqs/p0ue+uh+oWD1eJRnWQMJS0w9cSzD
Qjc0yu1sU2gCkNUIYO4pO7JNF4Y54/MSbS4Lg5P7qV2QdUlE212USoI96D4DDen5s94g4jP7JXRW
s0WGBsES+3N0s7CRYKr9XrAuWbWIJNq97uq5yWKrf4CPASLrIrTe46HoGUb9ffSqE+H9BWev+bb8
XExdTEYwkDNXNyR08OAGLOPvCayrVo9dfDzP34r/2T17iVqJAHkc5+/rmhSwX90DBTG3rxonJlAh
DRNy3rpzxZXxjElYA/6nZCFujmKSmAblTOs5zjxrbotJkp7/NV6rBwQLJ3beip4MuWa+nkSGNwM/
mKt8bYGXNrL5xLUpVdF1sOGrwoOtQ2HvoJTaQsV5riayo0suc7CPFJdSLLjCAmIcWfYbkVYknKEX
2SvyO48U2doTF106LVRZ242k6xYb0oxBnI4ux3a2kAC/7WTpCEh/dcufuSpx+VSkP3A9Y6sBJyL7
EvZEnUiFLAKEjqYzpHJ5e1tpgFqkVyDcvdfUM8Ckkpa2CCgS331IrBgboeXxyNqdvw627uRSBBEs
t8970bTjEVyYnQNIFcTcJn9SdMMhucHzYGo/JK4bFGYr7pT5DueHwM4RM4zhc0jHMkXW+Q5sjXx2
cqi5d617IMjB9JuHTKLPiIFI5COcJ/BszXe83ri9I3S1JlEEcPKQsdG/8ouwwm8kSOQQtjHGUJlr
VpwG0CTpl3s8jcJaxiPKPr3bunLRKZdpG1SzEY2VD+Lfw9pEaAXmWooeQ4t+dH9a5t4DK+Ca9xH1
Ci33C400U6MbcsWAw4fAtQHcQcd3CvQBw6IcX27e8TepCeApPN2rai1t81FOLz+jKg7prnBNQjFK
me2c8IB1sqnGYvAJH6uaLojFkqoEs1NV1gDnUaFDgramYGuRnoFYS9ho2Tk/tQ5ittl7P5zcKOys
q4mIviuZGtz2SLsFGRH87pR/W5PmJoy4+JiYlG1V9HGLePx16PkN5O+H9cDrvtioNrPtlsWQTQsV
qJViPj9VzfbHQR3fWOjj59mEF46dmJaLMnQe2E97Shylv7XxyilvJ+S2E69U5Bos0NntoMhcaDXn
nYyCGKk6LDqYnzvQOkmdCvMYivjUD0Wsx5jdYoLw9voghJtjiOAyDI5MfoJ/8ECslUcin3iehYTc
KvRnJCurKzadiIuK3yGFE6Xi5xaGt3lfWyL2dJpzqlX0ZGXv4MD1SIz3AnlAoXuUPP0v8TqqewVY
ZvKur5vTXOMKcdWuREfI1L5j8EDSo+7ozsOIiz1MC9/EVrJQnuawCVl0/4LTmscgN7q7CuPU3NUn
lO6HwlFSXgAXcDWSX9Wft29mh3oIeNp62ERBDg/v9Z76LmneJQMfCiokV8Pp0JQFM5GfzcvXgtUD
TNMh1+4UXt3SA6hOvlNsnBBZ2TRdwTjCwPnlxyPvreWrzFKC10N0EDb+cdhcCqkvEImNF7GC4kY9
S2hnfR3ScRGicg8rH5hXdKJHBFbZjw8i3z/IiJ2jF3WlzfemAw2z1BYU88xvPhAa+nCsalGbpKmK
IlfOKg6mtGIqYLYo5241GtzmwdT0dIPWuHX6ic73ooiZ+P/76gcFaZat34+9vStOSP97qTrIjaqR
JG61Hl30NMvPYw5QwaRjIDIpj745ABqkkHE96pTfQUSGUBsIZ1YJbX0o7PMykd3Ah0ldbX5fCsdU
y2vQfQmx1DtxCGqiQHuxtJp7AWuPuDg/EJ99hzcl1rwArE0L+T/5uMYMdSaTyM+jMmooHErCDLdI
qINb3Vi5hIVajbcp99etMX4CjtVzj8aUFwLTM6yusWRcC2qoo3YrgY+d7breeQt8r3poLmh0POKL
yL/AFzyWYAIbMxThXRuJtz58Y12axG+/KLStl/WA8JhmT74N2zIGxLuBem8tShJ8FkxkuenlYGAP
bbnXIIa1tMYj8wFGQwobnfB7Aid8I/Mu66k4pPPGXkggh3cAGf9dVFavzkPwHxxoqjd9hETFPWHS
BkxxKcclPpyoQLBRwH87jCgVRXZZ7B5gj4c7nA5Nd/2U76EOjCJUIulKdUXqx/jY8GoahMraU2d3
UeTznRQOWZgAtXK/ofWWez3EYLUBdTvxJkgtNkrhs/LnYFquEHvKoGK9BjvlAzidNNs2SI+GevK3
wzXh1I3YBkpMAnbyNtzSmD4o7VqKAoGyEpSFo00iWQqTF7hgwIJGWuhZJXEIgfavL322MSMjPQYI
FO+F2g1UilskHIjpQNkKav4v0drji1i6C5Hzb2KXRXg/EJVizC921CVu+eXq2akt2ENc+KBzQG+8
91a6P+B9HGGNHoMPGs366QG607cSEHXN3Xr/N4J5SnIaJt9/XNBRVuS+ZYQMksl8u9+b+6SEi2Bx
Pj7REXAcgo/jE+bEu4M7BVydec+0XDClQR7rpZ1IfzARiDH9oQXLfOI5d7iVkY/f35Uzn3IEGtCO
Ruu5CEVrBwFeL7tbsEzGIrW4mvWBHnUIRehQq7S9POmxEBx2XdzVc5+CWDyTLSt9jyGZym+yz/Hi
tOOxiL2+pyX8xS00gNyEJyhXGmuoQZXMmfdc4d7A9JBcu+Oap3w34Ne67N8o777asNjzJpK1QSP8
meUKxCYAm3iab5ku75cT6aMQhxlZefwryxvfGDZlnV5y9ZX843nMcIZm7krBkLUW5/NuyYymCpqm
yj4S6o0hEqtFBswMokkkLy6ag9+nPty3HDCQbYP7rRusTZmIzWiXWxp3ixLhK/IoIXp8/oj5ozV3
bwH8Rb5rJzlRErdg129BVMo05xsfYvYD/rXEWKf2eQ436QLm/gZJHD289bhOzA6A0MPhxdkx/y/c
c4QlzkWYdGWMzPnkv91yrDOXaU3oFT1I6BItyw3gaS0dVCfFgXW0hbfGaDGrI4PwWo8Op9tpWjvT
/zCYAIRmtxHFgzdfJ3swKBfg6ocQjMEjIJ6MaQhuTLwz+9jlGMqL2AsO6kCieb9rrnDhWH2/cctp
1zjjucOivkqtWSoGvYiKtXbodrQqJ3xV8fYPTnC3hunGlUPEd1npQfJuY6dN0okAX1oZy5FQnEgW
gZJS5SIgvOvqoBGC2lgB23wEeaSNtRvtly0dunn+nCu7B4sBjLWKQba2mMUjHasfgeFiApNwa8Sn
U2R3mK5S6f72UpRy1NMOKUwb4Ue6krdGLiD6sge7h9FCe1h/GCp+fRmoOWuKwWgLiiiZV4hGZNkE
b4saM1Nqjj7sa2MZEqognu3IcTM0rzw5x9ca2+uf3VnKYneUGrYOef2s97WlWW3ixpuKO0qLnhup
QWnlKi5Bo15BLtuFoXdxMA9YO6ZhGaOWU0OiUBELhit6zQ9EQ4CM/RTlgG4bpiil4ToCBbz1KnI7
RYS7eIny++Wollghhbwwh/f+MPcZWFE7nFffs/YBbaFemsUUtpqssgc8uIlTkeDKBFxCpZpzKAhs
5qxMAQMHNyeona2aa3zD3W6iC5lAPO4NYVt1X0L17oABJi9UcIZbWLifGsTCtXB8szrBUCRCtt5k
Ko/ktSA56jPkJHTN0C38V6hcMOmrHEcPiYJaJSCcBsPRtMXSsMQlrrxomJxu3sNbj87GWv/dEGRa
kFnseSg26Ud6LB9TUB9N/i5RmFAlXoeX3D9FSB7GRf3wRf+7ZCrbXwB18P2MKJcTp7kn8I9xUpWe
VeoSPNzFUL8XGYYP2iieBTGab5T0IvTvB1wzIx0wjO0SrqPcXG0zVi9EIwbPuWzSxliB23935LSJ
o6P8VorLUaTaOt6t2dzNnvaMEsz+XUsA20HKh8QczW5DfMDZ5jdC5g0X6D67Xq+bvTdJ4BcJ/jP9
4Y3hcZ4gNDswgYXGVvQIliwwsotGW+FReIYrDMFewTaNYRK34rz0sOuN5zj11ZZBCwIrL5UrURGK
d4jF9fnZHiW2MCubfaJKmJoBs0JwzVxjX3UWnNQL1VVXo1eo6Cayk63gah3Y64bN5842tFvs4K+8
mVx406w/pzcfRaG//HNjYXXbUPZnvC2ku+q7e8JfUITCWejfOwtS09QRVG2SMLQmoOtCtp5TwEpA
3hnzhSsJppdgFlYi7WEZ20bHkhws3SbhhYdkxGaVDVdPh+cPtgXQQgEz8Id343elqPxFi+znjyJ8
VLxRyMZOJUUGOsy3OXmSv3JKhHpCjoytvtQqjbRPZZfIdaMDz8CNyfEaPnqJZZnlXPS2Mrja1iUm
0gt/5quOqAA2fIy1MD5HpNPo7lmGkmHITQpQTVbIAR4XP/CZXvbx8AiLSlqcYsWw7EWto+TjM4CY
3V7w16xssPi9E85MIA/TknsDrQ25LjzZl8oJS9E+s0aIaIv0SIcHgbHV5FYaWI7BnYBMz//dKmKg
0jiN4Rd19+Ag6gdOuRuHIkGMsSY1/7ZO4J4ZegfDGkYEYvbQCdwPVG0TopRHfQpo0KdNJIt9Vtn3
Ueko5seZrHoEs1Ut8qt7/wiXSHzxSD7+MadopZ7oxEMkmzqr245MJJfH5HYY09Ww1FGle80wJ627
/fEyEgT45NC4FgHMYUktph6CkME5t4JC3NrpaxM6dnYdL65aGTULZ2R3YV2rbfruaW+qt/Jm1ZP5
gEQVtKHvvfeMhYAj/Ja/So+2dx/sePzp5HJD0uMqcFnuUhaJ1SCzjdts77aWeIYosBwbY6VA1OLQ
NdUZbiIzmSAcSt9Xa2jaO0nElX9WN6IEYwpvsA/J1VkuUr6CEt91UpY5eA4SQ4fmn32YaKQlGcZe
OHrW/ha3emzjCBPRhCWtpumYRGkZkQr/unrkG1/bbvPhkpBFRdJ+HA2m0EMYmoJbNcS3vTX+TfL3
tGqtEdnou+rN36xqOKUQxC6a52WjNbBfjA2PHi5OqZPI1SygiNMUYdbVdVtrC/ATyypu3Z6ZZ/+q
YnPyQvzCjFCcc8ssTCgZ7LvoQfPdf48Be9riW8Iv17eoNiQoNGmks7UUn20qtm29ygZqjem4GWNj
EMY3r51iZZaZ7M3rNAHc4+otVRdmvi9/vMOxJXhrT+7taXeVM8y+KFvQU2vBlqXxE7ffxJXlgdlR
/7zFRT0QEjzeA05PFGgw1AT0lbLHDKxV8R1x1TCkmy24XTRq/gJahEAlCcvz6PIPs6OKgbRg5VXq
rbUlgWF0llg1Ew9641SVIwmZUBe4SyFon7guqbDGhntB4lFgWB4cWcnZZiAn4cDuUpmttfHIKdH1
a8PV6tqK2J0aKPUpolsi5eTpPwsgblT5d1eDgjWFVbEdkJ9XwzFDiuHshmnYk+YrRoe6UhP76caU
i6znAApv9dTfKENCTWJ/RXmgMceqDIyg4YIzRpHTYoSwjYwUs/XrPSvKD5obsYjOHwSuNCgdYZkp
8pO6AMVY8DUyE6R9+7p+eVntMy9I/j1PDIueRuNDqG769uejTcWnaMboqo3wxz83W9N3c0i5C3yg
mOQgtGHVTr/dLRgdqk0d3ZSk5kdoYIekjZqLNmlWsR7+lYlTq8ClwnD306quMGPhXipiRRX7173T
xgFDD2qsRfCe3o1Qhq18Z3ivtJosUgkeIJvIuck9F96GHUiygy+tYYboo5BY+Lu76AirYp90ca5M
6olAF81wHBa21F8oeQ4cFUrkGtWgVCK0iL3Rn6hhIRWYiS01PQDY9VgZVYFuvQD22ytw/DcFTt3R
TCQCU2TbbFz6wIcfaTRdjM3nchhU98dmz7VxAlPKYU8aUHLUCqG3FV2yKnfpg5jA26WAcMxreIO4
sSoy4KkNs/MLsSxpwjjttkmdatb0ihyxs/B2dDfJRprxQEaG6ftjSxZE48sVBnklWBm59EiVrD7O
3UPwq4fGAYvDp5Rke7CSdSkmAgD9DXBNJ+V4KxSfZeE19UFvGm1K3pmXBVG2aC5h8IMDQ6iK9Iah
jDbHSxnVfGLzEI1rzLWpuiZ+WQgY7V2A8qKMhzLlnS0IaOhK2oY9HQzbywTBDt8826TJ/sF8arAu
99ds+Q047fXvmPzI/UdOMFOlNdlqe7aUwWK1OwwfX7EPANpasAwO/fXQrBs7vKcL8N2Flw/AWQhq
GPp769MUUetXDqqqF+3UrPz2wymSBWhMSyaDPT4a3p0+pKN1p8IM0FDCz2O8lt4igR+g1tyDAJF+
EO85oX5e1dxqcIvm/TMxkUhBeIQqXW97HX5W/nSJZBI1WFMBnLj2/rZpz6rQuvOMQ1RSCPZ/F8uV
0FfU3SVX07vRD5BuKHVeJwUWFwlgC5mHltXLKp4zJ7687z+A9uaM9oKNQTHhQNvC85BnU3K52Mfz
q/dhzJuwofo8uJd8/7ZZb526R7MQ5kvbwxrPa1Ev+ZTlwlHMm4ntKKPngg4nf6/ois+VqzV2OOdc
Iiep53sLJ51lwzr9qYbLhmDLYmD71cjd4STPiJzqoknRXMCTyty9EomKlkJo4jjZ1dQ5w7VU6LSq
W6JFoCwrZN4ySVVPvDuj/5MbpAh28QpAOrQHSzpSXf/dUD4nrUF908kZQrvuunOejmhAPB4AAqEu
VDIDLVvoi6F3HX01YVMvJ/+m7I9BPZM/bmbHmbWM4HKCh55L5YhLvcMoE7a3dgPutJtXrtNJkKSP
9Z3WV15GHwOILIfA53nBi+D5/WWeRpfrEcxd/EdNr2Ndx9rpFZO7bhVI6hO2klKR+ykoDSTGgDLB
HWEcNFJQPybh8uMtuju3l6cT+v6upu6vdYDrphzbyJwVPHClGcFLVI3Eq8+600aOybe7mSwxegIE
MU2bfwwshb+hgFzKsP7ZY9wML8yEbx7V391TOWQE7UhSKAJxpwTqGxJngC9YY0fctZczI5WNngCU
R7hDPALyi7m0XlWbwMZ2rljl/Cjl8c0D/hY8nxqh3GfDz4H3+qUbJ4i8WL69T4WEQEtFovnEGuBO
uSfWmUuzuwKYO/Bca9k35/5NczpYkNLNHkZG/SQbE8ZIxRbn/oi7YGVYhThW6bwkvswZz/1qGYTz
0jHzwQUd8jqe693PHEI3TRdlQOjctXfA1uHsUhfT24RTJZIxPFwIHij/EF900tLUqI7od1FTY5KS
1bSx/uBNgjfIX/sOXIPg2/enR44fCByrghoxZypXCjJWqQgiD39UdxDxv/0cCz034W4kfw5U2bYn
5dB0PKqpiosKRiTo1NifSRUvNym53tlWfr+GGNKNH+kmyAe0o5e+lnEI0kZusBr/A2Wd42rtWm0k
8WSpmOmUB/HEZT0gIbdv5A5c/tbEKyprq21hVB+xXekkh6bNEsHBV5pgXtpaHOPOOL78VQPELtPj
1j4nK0VuwsEQOXVMW794y/kJjCduefN9DM/1L55U2gfudLE1wMkv0IvdL14tlR91PWPx1FKsDg1D
ce50aB7mHhn6rJ9gNxyp5TGtvG0bkJFQA0koTXBxmyq/8aPL2kF42sTULuBW5YdLmZ0Q7TBEMZ0B
xnMCxF1+CuYMXNHJ3o1Sgp9DJs4ql8YWjaPq2tByziM20gQW0/rYGfunoeceZboT6LgWofpmib5X
ZRqG2AUc99FmJKMqzM53tOp5BBRHy0kPAKO+6M3oCP7Gt16jBnrW6+RdiP4Bf4LyAa42r487ZXM2
zX0QfGzg6n1h3G54US4Hflv0uxA7FhKRzpeI6TSHkdjOAkWb5Ln5Q4ot8yd1k/TD2h7tCrRx4bwz
HNiZUDPJjFol9/RDtDpvXilU74NjFVATI/MPHfFQqbHYaKtS3xmANYrkXVCHev0IR0wd9zxRiF8U
H1N2QZU5zp2vOdKbaeh10FF8UavLRL1jab+5Edz7yE1UlsrO9zCHbPxlalmggm/WuJKUrmBDbhwR
6fdNVlrpV2gghy3WBnWdHpcbL/grWeDCzzHT4TwzPwfJUAcUyRzmanLbSxO7VGK2mm3t+FaYocxJ
bUyJazfcmHpmBwaal1o7BKGyG6kTpd5+VZRAfaZRt6NTo9pReaXgJgVckPHnqvoCXLw6bc2bAD9E
zPrfYojFBkWdJWFJuoGT8cwCKpE29rihf6NOO3ab3WYCHRN4a3Y7G+IlyGAcSq8r/cmX/GTcLLza
29s37Um5SwN9dhTDF599LJiLQ7kxcf19sCnwI0HEH7eZGFT2qZJiCHr7G8Z95EiOJla/22ofGM/Q
KlIS94Lmx1f49HxdRZiKZmivtiDG/YBeBoYCDFstpnUFMSWCKfROhfza6lZcGB12LrXxpyr2AcUQ
h1zRbPAhEOK+1WaXmMYiqb3aSZeRxnzQ9PC3WwZ/wU4jjVvGAtxn7YchGxmE8JwUjfD/ShfD6ogv
N8sgTgbeVSJO54vN747Rqphb8FeYBe3brQ5djfzJi/IJk6HyWpIKluES92mwT9k0r7EiLIRsNXu/
P1bTrw6ItRQOyS89G7Ob90/NxBp3JEu/cqXPyiZPKJlazlZVrihdK4kGcFyOrxfVR32rAC+SUDKD
fJMJq/cGzeAw/mumtYT2HGJdLpF7SGAMonkaAHZ6Vh0dSl7SJ+cMUN2kgN96cWCpVsgB4aLcBh/+
i6yTOBLUlBfuHfIjpGKbKqbR509tiCN6uy6rn4pXJXgEW7XO/2XeS02cC16EEGlU0OEDhg8fMBTc
A1IhSiv1Hf4EmX5kZmZDYlb4MqadZPkKjRFuw7pyDHn2hQZ4AEYvviRWw5J9sbDPxxJ39iVy8HJg
BZjguvXlqRLiNbgtWPbuhUKbWi7wHyRNKnadBn78ZhLGJCFgZ7s/JWmRhozQaJ5cbE0JsYZp37ew
qwUxMTaieAMLBrC48W8yHMIeXoNWoB6tq+R5WeTv1C9UD7cWWjLva09TM7zi5dmtT5qKNrr3I/yB
n6qYVZntL3FtSRRDJRWXevbkxLg5tYQai+WX567KzniGE0S+QFymHCtQ8IcCHsCXqB3sIPdrSc+/
hOjV5aLC6LTBOfZAG/aVF7M419PXsOk2/oc9XZVOY/DVk2N7xdRO9h1q1OMqmGc8Qpdzp0FW94E2
ofWHBvVsKXOV+RHA6UrMRBNJDzx6QmCYsgv4AsBIEqXovoxF+6UpHDQxMT8W6LqbLj39Wa95gleE
r1Yy1rj72+BxXWjCgjwdIqv1/VXt/aO4uJ9WLL/ny8dzT8Zab+i2R3uO0ILzn4iKNuNVGbPY5BZ8
U3f9LE2PFUxDeiAv+8hvUkq6QVJyhKCLCmyOEpyYcE5ajHWGwnAXsLSfEMOEyq6w5Wd45KNlfqpB
OqXd9WWErafoURpqqqhHevfjgF4yzh+a1jT1NUjujO4vAGtrmr/1ZupNSbgEeUnTxPXrFfRDvqHn
Pg4PGl7Ms6HYXTubkkRQUCXOUnBkjPJpUTrtqdbs6uGv2ea+lNdM4hugpB2rL/Qt8R2+2WqOJgKL
I+Rf8yOajcKMw36yLoMeqwwSFkAvaYhyeOFVGO2FLg/al5x6WNE0pK3LiWhOOljWskcPNELW8yVN
+mqjqwc/3/lBvuu7yVK18tWLO3PzBoiQLUW1ZxFBV17m4D6lT9dOpmqyJsT2IDx3LX/OvfJo7kj+
3YN8ktz8KK6HeQH09GbrXWlvnpq+Y3FC0RoF+ckeRn5+oyAY4b6acW1GAE9322VX6aBFsDqM3T/N
tCYpxfE9gHEqn23qBWo3PdjhO0HxQfaz69E+KdNsGVIKBdSb4uYlQv9bW6gccmLoSmQUiR1KtQkU
bexLJmNkXkNqBlClqIO35FKg+a+yzR9eZ7Rq3dyv1+0+0CzYDR6wnmDIpwTMz39RDKPCoj+cc/pB
mFpKFKRCe4fYYDPldLAjaA8vTxIo7EEtXJu6VnF3n+KmMckBuPCKbFdQ248nTRyB3bsxzWR3Daic
jqurHk/hRqb+umjMyuKPiEx4aLgvaSbuQUyVAYpNHz4blhbAONTjXZQECSvW6adnVG3W3/BVwr9a
r4mXFLPYp2XwNkWffuCC/cArlYjdccE1+uXO4qZEEH1G8rIobQf9ptugj1/utjhjTmHwtPM7Qw7X
guXJyAupp7lib6XVfsXLoZL1lF4i+kp9jSNs0Gzf+IldJlBB0foxaSnHZ7BApWeAEAK9z1C55l25
taQYbzgENpOsU4Sk9G6EM2f1K2655zPtBmffGoirJx4TUE0S+/fOSyWXjk8lfE16zRNMSxML5yg0
XjUUccDVFsnGEiLDYCOOO+bII7vWtQLpZfbK//WnFc5pwin3t3HFVow9roSLtgFZpckYGPko8y1P
1tCZd75FQx7cLnKjMOT6W5BcRDmTrNhkvpHwBO6jZU/0M82wBP5DeKU8c+fOEz9pIZHDeN8dWCop
64d1iDe9Y8EtUK/qoyyogug6ZRG5BKZbblO6KN0WkUz37p/3KkbgR61So4sfF0Hb4u3w19UA5NgL
wODF7PJelIRUbKklC0MzkkfFmHfbzFjlrgB664/0MKBLIBtXR5uESviQbcknewDwi3PnegmmlIsK
mm49MohFy+3VKcGZx8AgL1PyoXEpXI0kNSYQGGD84/F6ViX2kDt900kCAxZM0DXiq1zVNGAZgI7e
yhZ8HkUqm/9Ag8hwffJEr/oPKGsB90pL5tMNjkbD6DJHVizQwgpo85kNtDXIvefKFPP+C6fk2tR2
iDH7z1+dkADVfrTDa1NCoWwJH/7rQvcJ3FYXcgqDgA18Xe7BI3x51UM/LaTfk6bYaH0ysjR/3SDE
6GsnM02scGPG5w1tRWj/e0gzqRVPHTNNSqi7/OWriiUhye+Mr9uVEdoaMqkv4YEmJVPkPfrslIud
WChSyRJx5wLSYOoDlzPqyX55ZimQPoTZO97A+tXtGtMuOkjrdiy3O4ufT2rNYCN/+8UxFWNj/DpR
+fX53iAPq4aevRKAJ9JU2OSrcFW5J+250OBKMPlpa34qhEArMil3gkQDaxBF+8jiJuxHbLdm5CGs
CYikJNVrkPy6+OKAvQ3XSLWqbRf8LT3Gp77Bg+OjNWuAUXVG1ydxgsIT9IyvC4/LJ08mJG2zU8CK
dLdJUk8BjWH7KFg9thMJ8cEVmw5r632vtw78lfQmfuxYSqlZ0+jQGGLEQADTUii1I9EY+HBuPpeZ
t86BYcjEQ6qRUlpP4n7hFL0hBh1tMiQ5DSUPY87K14ibbgpJrmDvcGPeiV4Vn1P+P4GKKhr4Ysn5
Qop8PhXzNDy2tfLiv0d5ZdPYvDET5lRxLC+YHgcI3sxrFpJTF0PuDlveUkaSLTT2W/EaryhxILVJ
Dt7pRDY04giB1i36FXkdvgzhsMcJN4xcMZIdEQHqMfLg0OwnexnYu83zdNjbvD36fSgRQ2/TL2cP
dYqepK8NmxBkMMSl4rysxmrrMt+/k6SqtkuofNjhppJqARzBEHiCaMl2ntLHLH+jcYjF5E3Aeuhi
1JtB4rjL98fbWLYfxsBUnZVNTs4Tudi2i7ARM1gxko67g52QhWUmCEU7fDY5ZRMQQHuJgu0Ft6Cs
pi864H7blccOCnyHF++NaNBcq31iG0TPZ7O6PK6HioUpNsQVHxMQTQHdTKrp0gPwhTKRpdwjYbkA
WRUf6EPOIEDiaetvz8Ik8JCyTc2r80yNDsD6oslfReLBh3VtWILBgd1v3q6FMFUOgDKmyxB09KtJ
aP2V2+zuLODy4+f/C6wGVDib+yEfj9EgHM+0waUpSRFzjNMfxYEFIlmzyCp7quVnoWnwkbiGI1qu
/G4/Wh1QYwZRVB47tqt1ZCStJjU8oQGUln4KzunP9zh3uXTdxO4XWkHrepxrsXFo+KOI97QPHKkL
gyqRBGy0R+RJXKq6tP2DtpCISurB3zipW8MqiOV4YUGbbQSwY3ojtC4SL4N6YeB5VQPiTzZchqXc
M/5qLurn7RMWeS+fotG7oWBYcKPK8vZpTDpwb9+30aCogAMqOMqUBK7gWbpeASDmRuzZrirtf5Uk
kGX3IopuV6nJBnxi11+NqFrdCZWjifNIonKQe+7bGWbrz7JkL8ewIhnlkegEihohV6Nlpdy36iWR
Tcn4zE5c2U3IYfwRO3d55ddLlP+ELWxVtUhe+MKIVrn0uu/AzGcxkgbAlrhjwLiaU9gReW8M+Q/9
cQMC1YUqeoNUflPCfMOZwvNCMweciq9RCvFpRGV7VjR7UldDIfvZ16shWgfSfN05Myh4eem1IZSf
qILWHr4dVHgTzalwObQJJM9acEMAmgRHqdxFNNQ3WD954DcD28Wh43/tKJFnctBljAw9TzIe058d
PShuR4S7p8BCeiWjVwWrtYxGJveshKQKLycsayUthXuit5//kkXb1BaQM5/QsAX/FIt9p/DowaT7
pCh5TImT6Vi0WFUXB7r8ZV+8vrsp7OZePgNiKcOldYoqgse/WF1femqKVlIEY77CqPF+9erpO+9t
F7DmlXKg6fdqdOqSsX3XhcizkWV4ZLQE/BBQzRRzSYu6eE1/ESYoNHpA0dxYwJBN3dymMnPVfo7C
L7NHe9Ev28uplaRHvyi3epyQdIhfdKKUCnUSmnfUNiD1kAAkmra+TwzPjHt1EsQRd8SxitkBxy+a
45ifaUuyraavAwWssX7RopaletKfc3W5PITe15ir4AiPLSGcmDkc4PARk/wEX/l4aib3jSpuip+t
Gt6sJlhU5qNYwsylDiTfnlrsnf4XwFaSAoYmn121lDik0cugHgfzapVDdL2Leqa3GrwlYw9a+Bws
m1n8suCQTy0XXksEMGJFvaLgciG//iHh6TCkRRskoOXey7X/VzA/GKCTTgm7NAaaLXBPA3y12LIN
KCTW5CCD+Y+FClfPpi8T5PGCtl0bR2bWluHkLRBfQ/X3XTaGnb+JsQ2cn9x7Y6wyv/SyAmhVuRRK
ospWbQ28WOgyCqtBD9VlwjMfqDbeFt5TNzEBzxs50WxOic5/lCfV+9HyLTC2ZX4Rgm3atQ7M1ger
X5NodL1pXNqyCyL7IjD51iLPRfaHiTyARa82+7Ed0+rG7IxaMW15PhhdP2MEGgecR35P00c30bQq
QWi4Q3Al0ApBr+NpyiFeKpvlalsF6ASlRA/NX0AQa2OIk81Pd0roX/e/m//FAQi7aarQM+m+p7dw
Q6nTKyr9O9BAr/jGZMlPLXEwuJCk5GHtG6PCbMbwLPtVzyGm/sujEpxsn+MDkJv3FO7Iqx/0ZMve
23hnF5P1wjj5EZlT1cdhAKYk98/C6xVH2YTJ1la5B7Dn0Lw07Jt7NGTZKoqJYRdl7MZfWov0oWvP
gHI3Wg57IaenvP1LThsxUQoqLlTg9oniNH9RG9qUAbWktnRTFI4KIRvuFwmd9OfkD7R2w4Dm/NbN
ri6TeIrENaTNN7zZzxqlmMEhvlNsebeF2CogPHP37QeGEMh4H3yvB5TF2Rk0oNEvZrOvDwxN80PD
5ddTz48Jb9KC1uhNL3iir8pk87XFO74ZJ0NTac2fZcbkFL5tcNstrsNXDQSIjhORTo2oYzXSUj0S
uq71AmGKtsrtD4z4jKuBQCRdPj+qGdhGcxKgIx6Q6S2TT4XgHFGDKiLISH9o0FkY2Zn5EEY1R1A4
HqgLlX3dm+E97vBhZm4e4SXaw2AEteT19llN1ujXIGMFzVDH7IbfbpYEmRs8BHSTzi4NZpGN2dh0
BG6ZLDCGWEbF4xHJRBEwuiF7bOavYADMukm+HBxnyWIUmZJkGKbSvapChACzjQt+Pm7Clmf3IAa8
NsAjbYeY99M5KvX8U3ZFIbNNiID3l582L1see8P7OlalDyTxpeHUP2pUyxmr0/LTODZPp61uTZHK
jlF/peyT0edKMsFdOaVfRwi0PsgSn2UOz5/Cv1qMMeDsQrU3dAVdnE9gZKfhFgkQN4c7dCJ9eelF
DPsIIE15Ll71wwZCppvQU+ZEjA9zwxYgd1t7XHMcZZjylxjsRblWEhvqfoDyug3MWUTsTNAdKqTg
XhNaUzZXiYQHLghG+EIZ5XIP5VNtirn2dO4GEOfbUQtiKfR3BjTbGcdWUFt4yMJkSwpFq55Aa8jB
MUgsEON1gNbe1fhVrgU5ap1eiGAU3KxKgfPymtmO0aPfxblEp5ddM7PNRjUZDZ0iL/kxjf1TT/YU
Jtzekuksoimkeze5PbjsUqIMztq4aqFajx1IS44XNDH9v51ilF3Ztm6kQmX9pJdLNHWgSsnI4H33
6Bf1M/1VMHUDKIVBpp9ZWx6jV/Nu25hTe7NcFPDy8+SBQ5oioYH+iXAH34TYeWSXYBsoU5l1acae
PcxKO+oZUVJPM5VO8bk+C04wD6fkR/BXdxWyEmbBVZLmTF7WY31eJhjBBEQTayeNLaQsEiGrI7nK
QpGAGBwyOdqczx3eOcXx91QakvdYa4IDKLnI0X0jbS5mjQtGoA6Fb9ga9e1oUrld9jESfLN/Pw9l
LrmsNtqYHDdpnPizESWCj5vKTJ0yv/eMEZ6hMjryPCS58AOKp1JtDapCUyWl5ESNAre2Um1hszsU
gn5cxSxLbpe2XuAhSCKRLkOchOqmArFXbMqdk1tC/NyFgtJUX2f5IVsuILErZycB0g7KYkbMC2mN
3iwe1OEURtU7PxLD3sNyD/eL0b7Okc0nZaq0Xpj2FtFXJPyqSNscGmvJB3T973PciDt92/uTYQig
7zBYE8evPCrjk3+i48CpAIuuaHNyMivU0BcThbYwH4aGml9URKXrrvKrfu4eghFUwbNBbM4f+ZrH
+4BhDR8JvLPypHIWETrRL12j0xuy5rQImjg5XShNKV8oW+BO7H9YGCLepS4CR1/VSTtUWzpdotAF
69Gu7tSLTyb9p2GMg2tKxgUrA7pQaKXXogNwP4rAzOz0N+HAO0shUWUZwoEaF9l8hAFEwh+Jyyr3
mauf8Enzd17QhPjvo2O48SAayRcjgrePQWbTdX7vD1M322CvK81KefymtYIBnBq3tOMe7UQhupXV
xZEIT6FWUO6KofVQteY6X0R/MZxpp8kSamlXxIIn2FjU1b6iPUBLQ98G+TEG/zaNtr8gRMw0uqJM
3UVTjxllSqOd4+UWbNMfOceizQnBhfO6wSJuwJBKqiu4ThwwIyRIDZdghzcu/psLoVPZFXN6Z9qN
twZ7NMYD39+KZkLLzE17TE/bCeyah5X/EMlt/srj3rYE3Umg5yfdFCfpV/csGtixbzW3MB1PgsvW
OuBopyQSRT2cnYURtcMtN/KPeWTxFikm751AaN8nl3zDR+kjn5Fzjwy02idATvURYdX0B/D12ZPM
7vMC5NNNY8LQkyOgrJ79/SFjPZ2Azb/1UJTxhbVYh6OvaL8WChg+sHhK+0ybptITy6x68xLqFwhP
8SDqw3rGnqLHZE39NmIXsVbCqQXFCG2cQhCQ+Qackw0MYM0Yicch5eWAGbgeSbY64GpMKHekJyxI
H2/O32NmvJbKQNRdAuvcx3ND+blcR/NKDbKDIq6TJpXXNsTnJfWSeEGz6Ddwqe6NgBr0IHsMfroQ
SagrDsSfaI4lCxLy/bJGx2i4nMWXqh/Td9/OjhToBbgjkWHFuPH7VU6g06kUAVZAUQSFtxDyjGWD
s6GeAXw3dFHVNNCi0HTVB3IVOgiHTjnsfBOUG3nAFT4BP7y8uUBSxzM7ccp+S8Lf+9pkc0ABwuyM
O7qZDuWrbFfswyoxeTxcA5uqWMiX/NhotZDjZVS+jqv+JiDw9dALDuxea+qVHOdrApgoINv5KlR0
EDBdKSOL9cIQCVc7HCtwqs0YlqGfsR8ACQAzxcTj46EnBvB7dAF2LPZgVmepN/fmGMUd8FRD9HWu
2tPQMjyDARXgKlq3oEXi77ylqopmyxBHXoW/5ph/mEwzARGAWRHvHYoOW3RhUyIjOlhPjD5Iakdq
GOYBd7GIwyrc6wO1RUw2JnFH4jVl9KVd/3oZeaVhuxlcYhLprIJxGLfIIWne3jZe3tRSyWGlTeQD
hFe11W8TtWgPCY7fef9/r2aTISznz76T+FOPnV13EvC44mCBS9ApsdRdjyiAmNZqAClPbA2cjuUl
7rQhR744fZ7DfzZoZP5TOjLCuVs0XgBxa5Ms0a7GDSJe1p6RM8tXSO3izQ8SpMQkLZetMu2tB/zX
0iBrS1K9OkiayzW3EjmibPyl07/YcQm2ymt//7XeDg/mU84mg8wrnYUlfdh0SbYjYIOVJ5MKOk3b
xii5RnvptMGkloSc7SFWQETxyL9efHXJUwQDP6GkQq7lOpQg4YcfzWyU6Qumf3NYQE8E+cJgEIHi
/68R8PPdUfmudH38199l6ZWIqXGkGE4+eNOyUXRyRk8AipUteA9ay5F3NVdcG1t3aUDmC9G+sivg
6qXbw+g76vFH4wSanF0G9pCDLPoUNNnCw345ZlRRQR4+nqfUi72zzkRjQp112U65unbywleXpUZB
wu6Tlv5gAVXQlShOlCtKWD5DZ5EUPi/R7eYlb8WD5jNi671z5ya949jfT9Em/kiiVUuulveiO1p9
lT6A21Yr7eBa5MKun65yBTAm2QIKH/WpVZphInglQBlFG37rW4rmBSlK3nc7FPypbtbGuM8p4R0V
3IJCPmyeoft+DqGGkKJQBwQkA7L7h8bHP1zfEkJBHBc4n+H3SkIfurNmsWCD7yGmjgWeduvcDZgS
m+0dU03WAJ+oHUS7QKdmIv8x5s+H5GiDUwd3ZN3x14nfW5G29PgIPEp1BOK60VIvkywQ5f2TZqHv
PA/sWzpAgha7NKM3BnCmx011Ji6hc81fBJZhfr+7GXGS2mQue0xgd9q1fGvjfCDLCGGOVpxRZ6DG
a3nOc3Rnpw660fFkfJl0mm7eusUk/dcIjcTszPjl8mKAho7SXnIp6HXyqg4g3LAyAwuq0/Y/cNZc
W4f3fjqV2fejoqRJ5G6cuzQsG1mEG4fbAPsF5ZaZLJ2GpvxA85EipkZdYv+TJ1x4AJJSIgv0O3wf
oGJd2E+ex9ux+yN+x4IwmylChjwxvyMiXDn116hiKCQbv7lU9XlZOdX6yyoP6z8EOnN9JTZcyAz2
STaN/XSgKTAgm0BYG8vpxkGaPETYpqbor5LOZRi8hQbgAiGhk7I75T2Oe65IDZw7AhUEXBiNiQfK
xnBJezKIkLijjiJxvoObVV/0iDeCD3grxZyQthG4SDdRvShBj+Saz4gkVFr8HC2hv6L0Z3Gerwbe
UcktcWkNP8mGZO/P+RR+wRPo9361b5Ol27MkLGcBZAwJyEXEIY2OtiN/fqYuHhTREAI17rJTz6PA
wIMCrjYle/LNs3YgIAKIjLcqyqxR/0Ro7YRQSvR3l5K2FHERF+8uQZYvzO95E3WJYi/S8oUWMrkS
kwMI4JsmtGr9N6zPZAMTC4wa2eNGApzwLkAkc1HVEFLFcXK3P/JvW6sbVPzxw7UkoAn40JrXckQ3
voY38V+MnJNoUqrchfFt7bkGvor05tkSsLu7qE9F38bbcIiSUaJWMJ2AYasR3RWtQcTdsdoLGiud
pkjaZo8bZOZwHmGHlv7kO2i/5zQIaV96ImpGUHaXylYIOEg+t6mII27rYD7VfRtpJqCVnBowyVfq
Ub7KDSZ0WsdNBhw40OPpnlkHypblWCMhvU5VtDhJ61B1HypuZnhp/bXIQA/eZYbxtT5OZtNDrvET
rvhPUO575xvH9CtnWAjgcvy/41KQh2Kae7d1hpx5UlhliKPCbW62+KdQ0z8p+LF/Mn3lsJbC5Erl
4jb25dpkkMNN1NqulVm01rKoPEr0TUktV1VSMkRVjW5JIT9mHPASO2WQX7fOWL8xVpJhjd1+1mYo
1WV7QDVyla+FFcjaMnSrTuyo6vwf3RgUwks/KPlJBRR/h3hVbMN/9TbmUzeCtlVbHU2atwVB5tA0
+SE3tTijJ9S7ViLQRx6B03QNOHPIj1Ri3DelhCzMbG77zyy3IPrYu3SUrBAVvGS3sxS6A8/QdXwa
tRIGk1gKhrIFdqF21hU8RcY8KzwuOIlMz2/hrGgOkzY3A9T8MgZQ1kDj925G3ugW5YTIFnXETeuQ
c+Nw/OIZCu340T7GZWPRqKuKF9Wr6Knhh/vVH3/wWhfCG42F2x1Ox7ubs4gkceJCCJ0OB5LvWyGz
O5LlZ4q+lafg8Fs87bOKitfgXnZND+47PAUlBY1MPXfM1hUsSERawazxsYxiAu0igRj/RgNfThTR
WcJaSn/Ww1vd31vd0rv6g/FAQTOVvT/xb6IkED0+HbMdbpR5+6hmoZgcBgkuaIXP3gI6SXwd/gkk
Ay6jgADsURqfUijeXfknPLzKV5M616hSwd+FMBlko2OvP8u3gwyeJLKwcohn6QvyK60iJnq6te9T
XV29042oOAGIdJtP6b2UvoicnYLd/Gd7hcgl4hKvxFpqTotZxOAkJBKK/ycGFD8tQy3loctRRY65
CpRrOp6txtdUc1xXKeiSNzHRAX1TzQ8UaOQe+e5xZ3b+3EPfraKRF2lCDQTYEnv1DmojiLPKpUOB
U9UsuTMjhrMCZvl9TX1gs0A4vnm8rgpBwQtHReUa3b1S8xddZBUP8UhV3wrsd2mlE9Ik/3RK4zFX
oLV00ig4btxGUd6zyUGuybWnMguFKlt7QA1ZPL/xr5gKseHCnakoC8zsmS5xy1T3YJrd8O0UCJmr
8Imxt0Z0m2Y15o3VQaQ0xt1rUJ9C46DFedPyZgFjBXQc0T76exNr+SfxZ6HAMdHX+51KIW0C41/k
19HPh31DyLder6mcxnJkAztpUWemw6uc74BCemljEiUl7GJOr9xA+WxZWjZ47D0ZdTJo0YFolxX3
ye714JucEPAPpwvwc5QPjWJM/jdRNonkZ+3rObi6QfdkBymAkhr9vHPsTiknPIM7/ksKkc2gkg9d
X5OS1y0OU8kX9e9p7oMXkjXJ/Es2fNRtXoCC7/SMNrGy4WYIuzE6aMBIhAgH70dRf4S0oNOJuUJJ
SXLnjGZzULogP6GB35LRdNoD4jyY+Yy3f+zXCe/xCO/mTHcFpRauhQIgBMoOcg+AaP3J08YY424X
uC01bRe6ALFoYkWVs5cp4YywrrDHG0ZStEX7EnXzLvLYwFdpSsA/WWHTTBEijO2ZUZkrejtKjzUQ
Ppgvoqo3KhnZ2esMzcygjyfWb63vUu+PBiK1fgaxIp4dpdHG53nyqDi12+qu0n+S8dTaDy832i8W
7COVnAuj8se321PZ0X2hEUqf6jiEa5Pbnd85yobDeTfgDtK30UENMUET/c6YKDrTjb9WEp9DuAgX
TLMM4ErDoa2WN+In25hMvZ8mILdQVb2q+JYJ9X+Or+IvcoAVEvPSjJpWsswshKcfQog2usmOMFHA
UscmE1b7QIfScUEy3W72xuRdpzsVDBT2JA/VtdtWqap5W4Etd8VU7KS4KKcFw/m1Bu049YATRg/Q
DbclLU5wMonjfim2TidG1dloRcIrfEURogI3wtd2RskNTEEd12KNId9XmjmJbjJZJtahYjfAz4Xv
VZCeR4NJ9G8uw7VNCJ8sIOAD0qYk7wXw73EKbmXcxONeHxFcQk/SnjT02a60/K+GvURs701i5MCj
+mSWYYFvpD2gRHqMbyIkXDjPr1bYlPuNTm5Hg+qwGYc3/Dzb82wBEASwXwJCXDHp/s58FDMWjOkU
bm8UT5C61t73YJxScxILQWM3u1dqujZXW3DbVmUy7KnC+WWtONyd08GnbdmYqVcwgQ/YVN+IFj1M
3LXbgUVJ9f9+ByxzHfYCEg1QekD0fGqTGlT9or9fGDHp4T1vAHFiLgqChpdJE1CoNZ2llzD3mx0q
jbiq1Z8TMrTgq1SL+/SOL4PtM7ObnjTtdZW2dEdZc8q4CEq5VHst88+TwxfShZ+9i2n67UP2FVIw
bDgvxZGbWZHjGKzUSblF2Z6VjHnhHMSV24sefdhHas+2CAFfj3LDM+qj8b3eFhEDhVYm6W2Y9jxb
eW4mERzpDpYC+fGG1D3xrVju2xVpIVlT5owj3wEoTOYi/cuwPytFtXHEjssoG0hDSEMXbjXJJ5G8
PC6ulZ3hWIhVfUnV6J/wpEmRe6SwqxEVaQQulrczEPMFBZ7mLrpMHCFL5ENgdSp+Fxgllrfz97u+
KW07Zxst4hnxT2WC6t1nkEACVUclFJ7PGeNnCgt03kYh8Hpu7A/IkHmXV7ZX8mjO0twV0R28JEct
JVFt+b7srvwV7ZMchrEBLOQJfZsExuGpz2/hHzJF9LZItl7azYn1CaRz5qsTSLV2uhGjOXZt92gP
5Y2yscS2+eJvl9v1lAgGZ5OaFZqrgMDiyiXdTuyR1BPSsB6TutVqkVSLhqsZvM7SPM+L/2dxVzHx
UqNVI4PtYIxr2gT80GCRfeclTomlaBGE1buzRoNH9TOgxdxnPAit8mx1UnSwQVeMB976sfwx+Z/D
pfdF0Mff0NxJF/MJ0A0jkQJGu+1Yy6rNSvyMz8F8VyXzOV+je6+PP3hRkdgDU1iNGm+nggQNR04X
559WaAVNnH72cmJv72VIe7DJEK1hLm2NINoPJRQj0y2XX8NvxNun7u/0lcW98KJxbxRN0XELDOe5
6o/9zBmuZjsDX+z3h3s9AMVpeN+mf5xp0Iisg9pZbEjfZbIzncAx6/d/srQj1uArEiZ2xy/NwNKx
u6gXBM2IX5SXSjPT0n9/5lDfixTtN+NOFmYGGGcRJJSF36Ilz6CxDJ7nSKdm1JXXLDiAoph5P9mq
5S8LT0H4LVhdFhdihTsui9RyvjV1W5rPjeZNujnDAc4vTBunSWOixdfHKNBtLT9+l76T6xsG6d16
BD7mC71JAVQDYJILp33zh/R9nDomVjtjpc9ojAtGyHc8uTfm9bS2IEtLcC8Qarv8EMa7AOKDGSib
N7ALY76WluVaSxDJNKl6LFa8UOBa2/PFQwPesfBIGWN0GS7+mkrr/2iT54vSSX5E+yjkQvowqhtx
gP0HGyBo/s3xzYittWf55uy+C5fD/Ax2QyvNWdRHU2yE59Z4ytCMpmJnCa5BbPOqv7IBfbyODh7L
AS9wmkglg6Hit4XVVI3oXPbdXqOZpiCfDqLSyIJhaD37ZpJlJ5g0Z8+A1ejyQLmT4B4Y2Unm/hha
xoM0ihRExsADSBpQzhbx64HiO1/zFCpUTU0YWvY5lebXtg5pJPkegcjLK0QI02GQgFufXDqg6uSg
SqMqvUpbOR82O4ef3j21407AnTmnA1sjEk8gTJzcIJTvYL0AyySYNBhSuY45k2HjK0w3Cm5lv2Qq
zbHpl17giQsrUurn1VSnhYBqKT06t/26BOIpxdY2tzPkA12UzqFX02CKPtTaVXUoE8KsIHwz36en
9h7XLK79if4ra0KYHprBie5GAwhMtTYqzAumugG+HLDteN2InP1TCUu/joDUVMKbfNdQ6ESxBULg
C8MZCuyCDd/uwQ6eqdwR9NGzLhx1t/GjgFDPGLbX3EhGZkBSE+nyvQebb3sZDibTNkMoYco+/nBJ
2/goy1EDTAZfDceE5z4hTnG61rAQw7phJ02L1YRb3MpNNLz/8+ATakjb+AYTWKKYNVCdzkDCvlWr
mnMEDij6wXF2DED4TTaiUpRicYhVmqNl4A95lzVW8ZR87x8yoGdSagqMj8i1h9i6NpJ4cr1ITV/m
pIQAObOHPANHs1vt2qtRZwxaA2umqgIzuMqNSlefM1sV4IGQZNR9Qk4HyFmHMiFkCj/Q6JhaVqAh
/8O2FU66MiS0CiwiaRZisgqHsRwOVljPlTr/wqFyzGywyVcryVFWWm9pNplqR3za6y9k1+7FA2q+
EucpJLT8aWADbLg/K/zeAXoohfHPbANBMGoDGpX4Nk+l0ozLmzKLR/OLq1chWJcYO7aWdAo14P69
hC5LcPNd6WgYl0I31gneFVShpzTTjwQJsIVhGDcmt5NUVSPheclzYEa5e4aA90YRnLGXQ7eA0W2V
Uk9lt4HJRSqw0KHIc+jY+cOrH9n7Km7bLxpREb9xQlYi3Rtxm+XYyLLZpqQtHPf0tFYRUzdUMheM
ArvCeMIXYvfTr4sW8PbV2hL2nnK5hMq1O28IFz7jd6IddOhV93Qvrgg6Mw/3PC57mCRIT5Qmd4vI
3Zh9CdU+EXt4VXupzAus7vCA3HuRZKxgxT0i0tVfPUx1VNekbjpPl+aIPCby9obzPoqZauctVAZ6
O7tSM69o2IIvC+AxvcHatGcCu1qm/hsprg17OZhhaIWk9KZHkmH1DHB4xt2rEhAgxg10owcJWW2Q
eehiIhnTkxXMkI30BaKvUQWCMptn1XlMQ3PIKyiwwZs4MLjv2pvWuv7DxCCJc5gSxCdrnaFHXwHc
XVBQrna2jsK2DLPgWssDaoUHWs2PB3YHJ5sIIw1swwNjq5ctg4UG628Z7pvBwWaPd+7h8Z6oOrKU
D7sX0ILEpyaarz/6apEBqRDyicH4p5UVaMyJxiJaP3HS5MdH3iYQffaIEyhkXs1b1dw2JvCgppp3
UTeAh1xiUkYNWROpWyR1srJRC7AGQ60tbCDh0tkPevTvXaIoqaFrdPKmalaPylOFAL08t0R8hO18
h3ei6YIc5SfYmMwkOn4/F9K5+EjnMhYnE9sQC7utdBvt0UXTH5bDr6k4Va/r6kj2HEFU1/dUB8Yh
5uz+3y+I2ExHIJ9O+aiylI5CQYPTZo24UjF/hZtUo7c+uR/dOOwMWr2/CwEL2MODXXxBhl7mu6tj
qgo1lqthWujPIuX5Du/wG8XbitA2tNaN9ekaeoddTXiIi6oN/hEJYdjZOxpLRSYdFrmQo4P/rbDA
H9yD1VxiRCYlkMAKBWP+LOtsHi6WHPXwo0X9/imfpUXTcAHy4e7W5KPw6eTUeCoEDHIhhuPO9qsU
LmHD4rFKi92fL7xtyNaB1URxIprMUawhNtTBR4GK8mkXpySbNcl/oVFq6l+2tru/Bsai58LnEvsX
mWSAh1KyiTqojMkv0aEIf1ajt0MzzAF03muiGy8q+WIJ23SDyB6Cg4DnF1T2OHD0xUz0Jjn8cgLm
+G+geH7VuSnuCwF6MXXzUqiPExrSDAgR7+nTaUC8qfmnR7TXNfm49Aee93kqNF+dv1z3k9rNVQFK
cvhpCG+qDskN1R/eb0EsAyKjhk18WO6lDfDCcuk1ckdnQXI/xnrOXLNq6eWPh1/IW/uYjFpJxHmm
V7O1kPg25S6FhdKDKxOBUF4OkSg1+bolUh4R1sXL4McSdQB3C+JQhAQLwIcYhaNENvqqQm7wTTlS
nP6nVpUquCbZRXoO+m69ile3ka8YIfyY3I2sb/sLqT72N3rSsIai2wnFE/aLMshxTpLBJ1M5nydj
828+zeQBhRlK84B4K3bGnfM/TiG825WgME2g2LClqjIDcPnnhM3SCO4QwV1TpT20cx4dcxS7JLs5
YAcCgqci42gWAr8YROLBUgP7qccdnqapcc7mbtKjNvhTMo/flf0sBZLxEsUzkZgnqIXsViIwv0/k
kpxOQz0ouziI1y6Rby1Bmvqz9Mban3GXWRPzmMkXI5hi6w4PJoHbs1zi3XgsdfWEzbwBA8cG4shI
3gkOm6pBQGGLTiYWYRbZDtvoU4EcM0zBShE4x5iRia/Y/0o5lZtS6wVXPQyNmgp0NAEvo6c+fdet
zh/d2fLWfIK9JAii7H2h9Y0urcHs+K7xdiLldFfozf4AKxH3kqTeOf6IVTxnNPaYsjREVDIPb38k
+Bl97tzIADgqVya6D3CCQ+m7sW4Dv6XMoTE1eQSgjcBeC7u5uYgAk+aIfJYxefIeDYrfnnrDTp/b
QiQ149vCN+n/7rtdzXvhJuvi3jNh1zpD94jII2eJvYodRJmc6JXrXtzHcNcySeTe1mRnpcxWm9JY
BUf8FlK5+1wSpcd/dLet7SeM0Yps9QOrseHABGCTfoMlqhf/guWVFmIxjztVc4t6WS1agEXRodZK
ACGajm90Hg04U5ibdwSDV0oKYbNlzjGHqA93kh9EdY7jooGGdk14Mp9KS6InvqbB9MBfHoZHeSBj
PxDZiBC96U+Y6u9YVL0C/YarAjN3RNjunDs5XmDNq9glyLPLqgDNj8Z5yr3QYkhJlwV63csBBoTr
ePuej0PKA5vXYm9Td2Z5dFYXsmTAcm8muLccFUqyh+gEMH4O+mRyd52YnqrwJxSapc0dPkjP+2cJ
LgYdCYUAaJKjZ6YBhN0N4x4Ad3Z204x65NrPgSFwi+zU0Ln5MBUPyv3/HAtpAni9sQpxQxQUysLU
us9XHcJI8PSlpqu/hA6Cj/Luv9VvhzK3ncYbqAqIa/crhQJqvEpHrpQyPltKpoMF/8bNrwmN9gYi
5G7WHmo+ob2hjV22rxA/8948U0Qer1pUVIZvTqBlR+0E/CnI/w7KprZ0RHq4jE4uyQu5ITGgk2Tw
rZBMcl2ANsxTMlgL8vTBCmhFU8u0YTh0MitGzA/Ivl14LQQFjxcXmtdWW1SDPgKL8RQT7SzrFhBA
QJu06ySR5Il+VYksTkCZ77siHqaXDIRqFW/+PiFL2HhiXPlpkCe/emgaFBH9bxUFZsBPBSBrLKMd
4MtgwfmfTDIzdUq0m24p6zx0N09qHqTKbhwx3zxtyYILP0HVQPLL1/j0wuFJvo2co1JPL6qL7+8n
57AxxUNmZ4Qq2dWp8UpxvibOVS6dNy9cLncMIAH6yq9MQNYy66p70K4WJwaB9O70P556T+GhgX7M
cB0WXq6uiaIUaYmxOCjjyXvY++e3Km9vjbpmEDH1TEBS4FUkuwEUTY6v8+Jjids1AzzbaAUC2zkT
WwAznnhuNSgH/t8Or2pePULgAw9MtF5J4a/i2GXzUf4qNmnwAt5wp1ZqQJxHZGobPCvdGecatlA3
e4r+yfelmyU5DVC7AtQmVIe54J7SkCIcy0LJeL5ReiYm9mX+qRt/pM8JsoJph9PXoGdfRfWlk0l7
5vpjtmNHkKrNIlV4QhlMirvcIucoFuzk07uAUJ055TDbyt10oikrYpaYx9G49SlNAPVOq4lWL/JR
IUHJyhtr143QcssKqFptEicAHyjKlt3Sd9QVDAqnnpr3tkWEKeX9X8NTW8sVTMP+cMueyDuscj0Y
8QfbHdHPE579AadE3g6WLbLdaqrSPFB6FIFCNDZZTd+d3CPQJBvatgmiWAKI1wrFiMNXXLccn3dv
TE0s76pSjVxB8lUP1wMtKtJa0sXguXkf/DO7yShQ75jisxZD/BqITVbb/KufITxzi6fsMH+9Uxiz
Oq0P/vz5TCIz2oi+0Hz/gr8CoZgWKjIsgwCmpJ57YrmHPGSF+AgJB2VU+INY9jUUj/I21RSgEE24
po3R1tiF81JdGD9Q6YkKHOUHv1vhvFgLDn3Coi23oMkcQh++brJW7gItPc5bY1Q5AayAq2+8J5Hj
658EOShiebIPncJnQ6ZCpJkCbqZnUYExTg7nzN+3etVnCcGPbwfq2qO/r4TI1CYWpv7fYCXpFEDJ
+o4LiitSH+vhR26CuHt3zxx+AzW2wdJ1kT+Z4OZw7ZCanXn+XtloWKlfgv91FtSgT2elAbTbtLdm
M/0rki8iyvibbrl+XpdzYhZbG/3iZzsUaNj0qbYn0BwyplJ0Y9zNhSh968psP/KyHGeSeAtoE8oE
8Fdkvo/3hwLmRW5fnY7PTYdGliZ8k4iG+qOIzKlYraTwyhFI7fBHg7czW8XEXUAmuv0Avz0QrZEW
Vezh2bovm1MU4VP+tOmHtG62dtCBaWLvZ1PBcvA//79gJlYgNpAKm4gfHj8soJUnptCnGm5vPtaN
vmXKH0Mq9m7W/SeUfhYmHafLMVneQDotsz+o4LqNLe0EXXAPR13+vIYB+OAHWs3ARgZG/U16iMTR
m2msySOiIluZivr3e5/2cReyePleL41XTc0qKjB+MVB+l0fuAVyZsmKlsLMgxJtNTAGGjRW/mPby
ZYhB2VVyvW5g1khVLOgLGnFLZJN3xicQS6g9004dMqCYux2mL6GmV9e4cRTPYjcYMcBHSepiTxzZ
CrMX9a30uEmDSIbc5O69IqC8DsPHlAe1/8ewYhQhdPUQ+cAXzTIydo7LEqeDHwZq1ga20Msz53LK
QGIncoXBKAFPDWI0zURHsJa95pUfblBvbituRffNXROpJzfoGatB+15kHv+ylDuTNTkrmFWCjg+L
2cjls/h+91H/XGY/NHbPyfzFNJ/lIvN0si7hnQhPCGfu/uDOjrC7Lv09k+FQKROIjBIS5Bp6U3+h
p4tHGddmT+Cb+QaVgP+auPzZnTYPgT3o4XmtfrrndYdW/CCy53yJLnO/dzCQlYc9cfWLikwDG0RU
4TxmTLo3KD6MiFbNjyNfyM1/vBKfdMMDNFLBuwCyDFXIwLBroofzDi1/nVdsmNjh1Tm+vqkUyqBO
vH2OiChS6FNgpD+8mZJk3XvqDRNRS8Y5E0zDgIppz9cMtUnfatyCcYChH6HNnF4aAq839aoqa6cF
TvMWEOahRgAp+JVqhpeKtHIDsEuUHOX8ETxVmg4XlELlQtcCPyx/igjX1mUmOxWTUOcT8B9OodLF
B+2+nsqIGxU154+WEucvTEmOlrD6htXT8j2Bay6d5/I/ngdTfr+jZ0JdbadccUL6kOc91/e/nAKo
UsvIvPzL9yMFEqP65AzwIQoJnkX2GUi4YkXBS5/I4l6E1gFnSneItjYqsbipJXk0PuG5dVQNFoD0
BZN7+mJsUi9PHNtsDTlQfAmwOd6r8B5lVh69YBt5W6TOlkjvkAl/9YEaOheZwOotqOkgUcYF3wHX
moe54IL33XiZhIDVxhs3xx+HpqEkHIVgBvdeosi5jk4JnvyKBMrr5kfaUivKzYe5NSssLFT62wg2
6A1wDntU0oUzIge7Um+udy6fh+Iai2igwyRgB8cDD247AJxarJRj9LlHFnGOV347BqArfnGFgS1q
lj16DJ+fH2A+0PhDmckpTvWCE2lPhXbpiaoggO4r6gRpEg//cnedppzQEh6eDut/TKIt6bLTuyXL
Ju+/35TFWvIuLIOQSQj2RJJLxRDqzGwII/1+06esSXz35rLLo1Dca3/k36SMrnCChzD5jm+17i+x
jlBANrx8SmYaGo6hwqHNRXz38sk+4krl0H+FXWBa9TG8ZrFZ7wlpR8Bh9SBmvEEHY895CSDEpPJS
lgqi5hsqyYBC8SdRqhhYvks37X1b/ETwfzlpWnwxb8+XFj7Mx7N1KvLMNkLeT4Vq3EnK7rypgu/5
SJJ4OL4eqRePAcl/+NVCvK7wxd9RhSASGmbRzsTxfNP01wzwsae0LtCQKwb2ZRwrhjHTDr+DaSY6
lbbVluUZJhVA8RYCxDAoGGvLihS4UyePuaBrLHdZSYzHkD8BdEeDh2sx63kF1Q40aHbdleUPNNjU
6iWVYg30kTzCgXdp74sJ6eEe0Ssct0PDnjSJdAgIpWyuHnsFptJT3S97cN4k3zcEJX7pTaKLktPF
Fa4oZPBfkoObNKsUA2aqUxNimS00ShKc+VrZXQZZ4JLKTsGvnQwEqpu/Ix3fkJM3UtvOP4wqbIBc
ARkMpxFi2Y2zEnxKtp9LFO1FYlahdRYHIon1tcNEM3198wP0r6R20Z3yMfqK6DyJ+5sVACrpdaTZ
ohq5zx8/dqJoDfGr3+3O3v+9sJfGZweiKFFQYWba4We95UngW2mJUoICZ8V2rHU26nCzGtczKLGI
3WZV8eWfL+fMeUEwRLymQ2stu6Zms4/aEMMf/JbaID+OhzvXUdISjbN8FN3jc/q04hSp3J2JwoKg
imHApzITZCEwum8UWxYG1ZD0CPHn339dgDaAkjVKrJA2U9k9eOMRXPfJp6R2g059JYffVte1twMM
VMMwQNyS6J0X5hIcOO/Y1ilSgqIUfWnxBCMLlHAPN53C+d37mbFoIoVzw/hmRJ8vm83ZIQtdW++K
MSbFS76fEP45YYXcz8Gs+oF2KIOUx4KGGaFWRXDFiVx/76IhX9LVL4JQhz7ombj0p+nKzqFEP1iE
EAOFvZBTpcjZJlZpCsoG0LmlM4z4tYHmnuGYsX/KVXrIYB/LlzY9ywvKbHpXMk70D6ek7R6l4LiJ
gqt/MdHWOCa0pSalF/O1+rd5bI9HwMjovvklgQvdDgvIM/MKnnYIKa3kc9bjTCuWh44ZPE+ng3kd
HX+4jSg6UQob4pvf8KdfDx8Cz13u0kLZPBftUm9QjRoMAIFxpR1SNlG0BvzyASBBmDDIEFlG14TV
iefYX43d9SiQHIBAhq4sS1YTIrwen4OixPBJvUVEYDLScq4Wa89Uzc44LJBvpQnzkcissDlxMD52
e8TdrXU8zirnA0wXYtt0j+4vECEtAnOJ5ouVRGh+f6S3CAVhyomQliN7AOLHLITm4S0WlVEj9Q8t
+wY+hPLt2KCDJxPq/wqmSUXV8Um93V83SAx0kMBieLrIbtUYmhZMGE+9SlC7gKUIc1a1WwZlJXkg
kcmh763sMKhPgl2lvHK06pHEfDgHGbSNwYbr8ceEoWgpmf+2SB9afCYrvm718Ibi1mW9LnfqxfPD
gczBzjClq1LgqHkpjG/fDHAzEChKe9MPnmyb3wewAYsdDOc+YU4xEotKxJOePN3rF3Ee2pSajklL
PzP63V95d2g5P13TY3BGKFG8OSZa1KtXamUgCFfKv4uLaSS3k62dX5UdRvVEbYkfK/FGhX2GSLC8
W0OifqxD5iXX+ozXfrhzDvdUYqPnojk9Dnsqno1idsLCmnUv50nC2rnGu+oyOXHtRKmXbb4lno01
T+bRFUI4Cu+qAkErPY22M8pD1IufXIRQiRUemXhz7vOwOSUKFYX/aVn+GovgWzYNqo4wt84luEno
F5KBoOc3P1uEim2iE04KWxSxjMAXX4roI7kUepCLome3/iqtFfJl8D8R/6x9O+ZVBt1OgsGLRNsT
ls12T6czzD/vLq4nc5U88ctqtCckbAehqghKoOWUMlfJLUc2Aob6ZoOCa6wu475yL7ShBOPUfe1E
k9O56BfzTiZNXNzocyZCuEyxxJVqbtmTrpWTTztJhsAa3dYq9h8NugYHHJ1pvNlv/Fn/yV8B9Bsd
nLGjZOa6/EDHLNuodCaEAls8+FfTu8wPiUeDnPKZMBoWs+bJlZU+d++60NG+RdzXcWcKg/PRY60f
tA6WYLr1oYrQiQex2zKgO/G4gAGUaDZVjef47S+AA166OKOL/YQaS1f4fRbgJ2TbSd7pO636OU5M
A+bsA6amHXFVkp9Rpq7dsbY4wxD3/tx3wGWTM95BPRCHbJlSWlQoOPGilGdSSYXaOOUh9qBFg/+s
ZieXhmhhK2fmD1zvZ5ll2DSgQgWmpuXN0cy7wsuKn30k8vWboSLNnUcQazMT9HBgdRDFavD0LRG0
5ksytNE6r5mmhpS5KySEl+Uob8QSHbOTRt5kRkSjxHjMoEF/VAAxpoiD/GXld/ca4QxLgKpUIFKj
tybo/vx3j9CLbIBGvMWsI0rGAf5ol2kKXH/ke2cZlXJEb5WCsFVgVmkam8VSP2qNOaEpUGhdrSxP
YtVZ4LxLPZC/0RTFtzE7cxqgdAEwFQUOAqb6dccixANWYmwvaeoa4669BpUalQ1+c0Yv306lQLR/
/4sfhvPRQRZVCdvaOotOl1ivdsJgYLygs/NNvd+PqSO3weJLTc/3aZA4ALmXsEJPshtNG2sCg42q
I8Ks/5ZHsU7w7li/RhJM82hU09eG1w/PGmt97pyKLpwD6Pyz9BCaow/65eUwF8kQm5nJtGv/nS+o
JbNEAFSGxVYVIPYrPVRDna1yuu7VI1WoSjhO2OU0h08FxhZJE50fRHD6ZrYeHK1HBj+GLOnZqq7N
4d36qgiuT9no2lxNKqN5Vj4CQ2yqEvhnUa+CWdJaNmRbR8sdqwEevbMylxNKr7MQRhfnWqQ148LA
58wqtg1myGvzgBk5vdMNVK702aeru2svlg6bCfwmro5ojhlWT4gzySHuEX2clF1QUDeL7k227p3X
H9MmktZ/Y+CUUpwHOCgGpg7CaO0hAJB1FFNUB5CrG0lut5eLQfPoqdRVrGeeYeRm+r+2JvoQQncF
Ri+o2iqsapU52/21EqPodb3wSFshjBgLsmO2wNue+aMTUbN09LhgYV2wCJyNr+UAscp6P2lvixcR
2cFwYhaG6oRlaMGCkw5WaGm9FD9A0/MLaPwayJki5ENitxmqKhW5ld3VSjkVYOkGyim0CCY6GT20
C+KbUSXt0sg9QnlK36vfSL+Rak5dPCjbPdZ87WkO3qznlju9szUWnXHZysPiex21t9o3ACBHC0HN
x1Xs4NIXEPjzkwJBE3+7/it5tZZzlkc3hSTLgquEjw2mh67blwr9KNIH2gBxGaMEG07btmp0hCnl
1oyhX37Dhoxpv4QcOFuvLFmg5bwYYJF5TkLFpoAM6on67SufrTpsyNtZwxvv7IXQ8D1ictjPYL/N
x/BEQcDOPHJ0SvIR999yc6WDASBou/4n82Vtngi/3fcVOGYpNiK7p00qAWEOGstM7C8dvHVKUOEC
j8iDBgucvDpx58D32/qDK6g/Fi0mVE/z3EZ8mtN/jO0RFFTswq19kGp3FC5lAQNdXJs1p6YKnL/I
dbUTFTPGo5/MHOIBkYjf1ZjSI53Z6wAAxIgfEia/lV9GQVFM0r4eJOfP2irKlcnAlTZzXksEQaFm
qbY39jUGN0+wtVhb8N3f486EbzIIqxY9oR2hDpiy+qijRDEan/TVstIL8IiVhnEAocKwNElvmHZn
sp3m6icny6hBb27aWF+tK0LBcsNOEnShf9hL8xM2rYJeY3v0gnSbQq3BY20J6d1VZZnmvNaJoXMe
u4JIJFYUn7LzwO367wCU5+XQEgMd8wZDpfdhPbeY0fuxclola6S7gphLlDgDPxrLpQKtIFXF17dC
eUnMLTsw/1UBToaIA+Gk2ndf5LkFU3pMKDW+fArkVUscHBTbgbgztxfMKhih5+QbJO5/ae+JdZvh
9j5uA5qheITY8fuMwVyvR9xhnBySfaHhIjRRsEfHAwEARc01ZUgKYCvirNHEGJkuRRReF7ZPVafx
ZEozXxrdrZ8w2ywCdZ/P2soHdL5Ua8V+stUHVnrlIAo29pg8vqJ8LGtmOIe0EC7558EiZ6Cl/zWw
4HxKvbQWIVkM0+DEkv78ukpRHHP3QFwjUFA6+1NIHOsSiJ2aVSZ/Yo9qyq/UZszJYjkgnqh5/Fr5
Lnt+rucjWsEwMJ/2HpGm/ejZfOYQ1WR/HjHClL5TarPmOq6c2XtjZ2WM18ogxb312lw47FRiP7sh
fEJ7xD5PruI42mJI+2xGl2xbMFQi0kD9GK+NN7lRiBbexfdzxX/+9mURMSQJEh9BfuuoJz2i/++H
7SQ2Ft0Zf586uyluTJYhaGkibhJkLTXG0jQqaIDhJVYdDcVTXoiF/kZZVtStmMpULPn6TrwZe/8s
3ilBMHp4aZycwWVDhqXAHhBZRVRQj5g/M5146QebSRVe/lA+z8VEj6Kj6BA6cu5elzFB8KQEgE21
NCvV6guG3QR0UvRC1SIDmO/D09fS/YEMoNaD/NiGPbT2eTuDncaW0d8aX2hTzGvGZAGtTVnjI8V3
zcdsLsnIaPOjFHp0nxX2uhHD+9nULS5q03u+GCgjYvvcEfljNLl1NTIQV0c0yYtO8jsuByzZc5bE
NN5HDW0FxD0Lyi3gC/FR5C0hNqhJG5lvTfcTZKX2bKoOn1pja9CBxKe8TbdhnCpXbqJMb1dxezET
y586WnpPsD783Wqqyc1Sx8NayYJW5iPj+CgqbobBhzSIsAEd7XmK3YVzBfnRzQTuKZJvirrRCMaV
MWCckI60Wh3S8cDcTV22u3/QKGOsM5gMih7Hq+UsV0B6YUfGjLRzzjIYyNyvDgoI3n5vRG6N0XdJ
KetaiBsDHYqNQiGBKuLNXqg0BvWyYA3AQRVI0UeSSS70frdpa447XBaXcLEsU3o/z19Wm7Ppjrby
PPPprg1JEEerSNEMyFmm5wRAG6z7vg2frxDdkV/whDXI7st3S8alPxRGpx2WWkuKSWLKx/wpAow6
YMxTWhM6JDvQbn9dzctv0c7agOryqC1ZzoLyvdJ0asusRiSYpT26RGQv9lvfDBycSDwYNVtA0u3j
pi8pO88KEdyapJslWpQ2QHdagJWQLisHZrDn7GGiyMXYJRgQl2CNOVcZsMlhD1z1LLDO8d9OMAIs
+rbwnbCVpk/VZrTPqlMV/hhWt3NRaFwRURRehy8/QAZC11aO3AlkY0wEmuwur3uXSdeLhXW/T58m
7daQlGNuqRP0hep7aJRu/OwQ/djpvmElfck6imekFwZWC/QRYPoYFzjGslfZ90bHFvWkpoNvAkZi
SzYur0jCsZ8O1kNgPF2g6PSHD9Yx3IBTdlFTllnFSluFu6RtUMBSIA+jBMNMkkV0Ogj/OJ4wsXXm
HVYm+EJNzTv6kNRGz+ihwDhUCve5WjLaOL4zD+Kf81aftrBtCkypnxGrA482O7H77iK5vfStP3Gz
II9SeXDuB2SoafPRjAXNEPsz3VwOxRFMv1QK69LFDhqP3lNVkYevuKWS58ODfl57SzatuIb+mLmx
jErhKi6VYAU+EvKZfvE7cKv4AxNlxJL0QoXQ36o12kpMgjxT7kdtoQ09Kau8sLO3vSL1+qeb9uaw
ZPH5meP4JmOG2NQ9MCQ16qnDOypP+S/CsuJQV1WawID6bRyhY61WnKnLEwt77xiOQ3pGOvf1/osG
I7Dn3eB95W/CDEhtBoySppZeFv04dIF98fVE4KHLOanbVnXFqkOAMqroMSjwJ4ugjoKhfWSxPnx4
lzyFL1oCDCi/HliJJIfmCwPHUwvHbXWE0GppaiPwTzgJXif4BKjF2GUyk/GGrxojNbz/Cnm2zawY
jtszJtI9FpsVzvfqGAENuDhMorBn/CD+FFZ2Ia9OSRwwPsDxN9/ciL24HkHYIP7F2yBhGHhSsY9j
/HXGe7UKcQIlJVlaaXlwF52jVJatAXJwdM2GcxRyF+TTyABA5U+m01i+rXdjOEzAcdduGwO6LBvv
Dn8MLgyD3heYwJNhPn0tx9mcByXhOyBuOHnPOlo06kICcsLabn9/cRxxnUeTqqJrRI8c+gEbbeAr
xHo5ykp6jhyIYNXwhmEQn+ol7jK5nM7pMTBK1XTJ0dK6sCDTfDqpDUCm3WURuRKDOz41vslPzSyJ
mu8TYCVXJ84M5/8NuG4407mjHlyoPHZTs/l2LW3ohG5O2QHOhFmXTWVsNnEOdGPiAyeDApR0bwf1
td2pYLP+H6WyXApgowXUtLZZtBMLWOpiqPsxeglx4yk4lWy0+eY/bOEANoL6PlrI8v6a9tqSjov8
2UCxmRjQoh/VwMG+RSlnHjeATh+GnCyEWzznZr1FCAe5lQA003i4cjl1oVo7yO8sugYTFViI4BSY
ZVc99egm/RgjTVO56vOIfkks1nJACnmseU3azFeZJ3UXzESA+lidNDW7uDoS31LYsQiD6LqmPWVS
01yuPPPVGp2ZGn48WGbogizggqvLdCUoPqrjzhD6Eh1hJzFIknTOSjRZQNHOTVSTKsLIK9I1TFYU
o/6+eJCqIlbwrdCTK3wOxbCNpkvgt7MFvdNclMlMLueUtRbA/JoOC166oc2nYJa+QAxWiLgseCMA
vbrDuH8rucO079yYxtgVxA2HPfiADzkMMTUj3SrGz8IVlEKHpioRGGcipTtrK3IJFLj8p4o4B94F
BNaGyXk4l6PtWuHFOMIjyEnRYktFzKvz+9KmNCVsmSYUUSA6K4dc9IEAM0Zb6uIq+lLyZxrFwCc0
DjqQsxwowHk8II4o244Dx3vcAwFlHGgIlnZijtikWtdDpIwDa5dZEzDixCuVGdVKCyzfhLwltJzx
yE76umarjQIofg+fJRX2C4ehlEvsGbAXumEdyYlqESyKrHHX+4BtmQagwabJxpyAqdjytn9FbMN+
AFXnu3TYyfF++22xbnX0mTPnTbwj8oCNYN32nUdUynrWZ7tu5MUn9yW3+VaQsjZi1x6Nma38DyuN
l+um4iJfOCBbUvXMMz91N87wilK38MyVYMx1a9WUxriIFRIsbqdRxEl5XbpRV5Hx+9E1voWn73bm
J44kXGA9VzFdij3LD1cshzbHnIos2Mr1pUQVqAfrmAtsz60xZmKSlhnVe5wnr3Ovcyy+xfABzSjw
YXDHEauscD3xaDFPX2YtIwU5Bbp/ik+eGHxVUBySa1eCwXm5k/5As9cksvlN2HdY0YyDxITP5U/U
7BrGrsUBxbPBBRa8sid2ovDtlxuEn85SzVyf/gWPQmhZqpiz1Ge16jINGdnWqEX6KaD8pCHtvoDY
XR+DGQhqMyMFadVf38Gpelnu/eALmXwlndpPK/tm1VQvRPQSgm0YdBAnVltW2gC63B0Dv3k+0oLD
COpTO9lMVWon7TrAp2oxJLhv+gb7OcTPPaU6Y/oYro0Jo+8bc5VHbKpuvW99ECr2x0CLA5/zyEpI
CzN4Bqz2gMu+3TTEhmflT5OadzTN5vdbXNWvIcJQnp8vB/YRSvOv8J4EZIuYQQNUARteG/V3293G
ksp83MvaBWu4pqd83m1Pipza5C5Eb52OIcLGbbO0E8d6j1Z+XVr0B5TkpNvwYgHTEzHc4Ia9+wBR
O3MRy3XqVceAMVxCnmu6shOf7cbDBaniJspH/icEtcraOy9tpcN0EHhiqcwqbN+xVNmaZmwrTZwx
v+ftg+CosO/ZoJ3f/wxMBru8HxYRX0QNStU0Xgup2pyAmvk/STJIfGTJrPgrAa1tHNPzosVpt/2Q
EWubIWlU9CiWXrUaDZ7fKS3RneVKKla4LnoRnolgczbAq9I4hpjiVQs7IjXJYH6in87Ocr2vFb+z
UH5LnD6xrLnOWbNhe9jEwewVsvqgHE32irwjraeg2mEXI4ui5bIpOKNHKLvCU1yygJTGmc2NHCLm
S6mALchCxBqJ1+FzJFifuJ+4PhRcPq+ajFmggU5yZaxpt/XbpNYHaS+ZPm0FWVKSqWVNt6SRTars
KzeNvTWYRee79shdRNyjQUIzRT+/DXlF5xoK/bzdV2xsmh6U89FpC4mNWvYW85IjIq83tzmbHx1n
j3/4ROlY06xyGfu66sRwV3BFZveXg8Cpq7XBTukvG0Fbk5lxJgLx9ROjMPWkxKa4bvV8P2uzaZxe
9YLx1CSV4W4vJDrUGwwSNSvs+cEKTzklS3XpBPbqLxndFR/M3w7JS/9rJX9iPHlGXLJQ73pE0BNQ
5YY+LFNK24mrxwL3BvxY1mWhoM0NkI62sBEgxme43CXrRjZ7w8GoJzXPR/buOP273jKMfDoPpcb6
CtW4RHCAjcovrt6jJ6qZez0xP7N6kLiyILlXAVbv/d3v5xtg3DmBzOtZmADEdbcyEhWjg+8PSrJv
G7JbTqBmxNjc4rBRoctw9f6H+4IJ/Bu2lRODgp7xpOSorhk0AItPboNa4yW6Al56xt354mgHqt0z
7PWSVThSBARdYy5lUNfB8iXeTQaiu6Sr6xKB2BS2H2q2abNE36Qy+G/4dDB5yrQXPs1BLHNEisHF
FvbkVBNuFYstvNlXBk+AjgbIJOsK5SFgfqFmvPXsnE6HsaqycgM/AgACNS/Cl3lpwbsWnjYqeSuE
MSCiD1336/AKD/CGlgCZTL9vB9gtD8VLcTuvXtH/M4y6/xC+PK+dYhxt8ZgURVEfYKifvoitCOMR
5yn+J4/UfTNyOCWdP74KycKcQtqcOLhsE6b3I50fqwXWifglLg0ApXOBWyRe3mehCJS5bj5LZ8QY
jk06n7srWQUPwFsrv3Qu0fgKiI4TDMgUADkWl3LuLrX+/33hc5w994sqn0Gnq8yBAOPh/5U9TdDA
dqwNGvST+gSu2c54WJQVOKqJL4gaat+H9/3e0T8rzsG2tYg507/ikSNhLgpob99Te9tPf0WQbRL6
MoylbhhbrOs2RZ7L63qVaI2VmzY9/Lzo36DCMu95/RPQVlq6srtYNkaTG3Uiiy/Nd/dG6vzw3CQP
x15uZaORbwKZLa2Pnele9kpl1SDeWodQ8S70W78IDPk8dYmv2xU5VAeHZjYPySEzFk6Yg72+kHZA
e/li/KM1WbDDihiyx8LUx+RAOlGPGc4ywzVXDlrIbJeWEdqEJehADItUUpqYp6q2pfGnBHi6Qsz3
sBH8xi22t0J0LpJDhnRveT5NNotnFHwthMqD6eFHhu1UQF9Q90Djfqight9BrquGZ03lYaMuDffN
gjuRZNxNuzzNdBpWRw4+00qDqpStlGH3lI8ddCuIouoAnPX+GHjU59Hqt39qFmS5WAM1cUPTIk7Q
v3emAWMwJURjMHLYcqSjm75n7NZxKT5kCk82k+X3ClOXyHgChQbOAGJ5SxzYlwbz/YN5AFTLm+F/
y0gL0i9ZIh9mT6Sl/M79W+GJjOJMfbxB1GzNph0mJo4C4mGvUAATF2zvNpGHm9QWm5mxaW2LTFWV
6qonbPiMgkWppxAyh6Jh3poISLqWFl2LRwzC7PHbPVci3pNpo5qiGAsTp2lZ0ucjbU4H9kRCgJNh
IV+UueYnrZuU2eQ+b3IX/v5CkXgAfn15GFMgDCdTGAV5r/oPYv6LKUvye+gEN+Et+I1ZBYylQDx8
2zVmffn/+kg5suMA+bOgTTKDty2gOoENOGH8zeciboolx1jVXqTYwzjy7/J332UsuBJ+cU/SfeWk
2sUQaq4cN1tGlGEAOjD3F7fbX7ukRGJ1U+8jKhuXFepbGrsr4YQRiTPLB7051Ntczu+9PIyq+S8M
6t1GFWHGRpFZXtdMctsSsWG1q+/Ve2nxj7m0VkjAeDEL4kqLKNqw3QXknt1+yh8sQS7CMHmBJIeh
1psi12M2n8Yv+PNSOrPPpNY8pMTIem7F7edJTAR2FtRrVShuyvsdO7NvizNNyOfa6+XLhWNGbLVT
todOoUI71g6eks36bIxhnKT3fdEgLSHprBB/nofjK09DNPzhsGLp3KnkWK/mhY6flbFMeLZJ/2wk
lea0FHPub5aRVzaECA8mubWbKKm1qbHalHOwoLiKtAa7OhK9aR2m4hYvM0MmPYzHLtDqOprKoBZ6
r67TNCgtASOQhN9zxDfk0dKUIHTq78gzzrMMGVLDjSWYRGPXe9B4+8LI2xgs//q0qrfV3BxrBpvl
zt2bfba0RhvuVqQpaJpFmIzIjRfst5OGIKgHIYq82APBTFbJAP1IUPF+4GKoSgQr786X30pIxjIP
eCCczuRENNHhXS9+EZD4RwAmeweHtrS+FOy3qeLK2KBP3df1zCzv8Kmlne33nOfM93dFXOY9HVTd
fthGku8cbBbeoJIpFxlg3kbAQBTkRowPMXsGkfOkfDOwET7rM8zTA4aZbNChL+zv5qdyJCA4mdN9
xVo7m0qCxq8PTprQrawGQc60WH4JTYl7cAEOwpHjoDHyJT4Hu2BZuIotrCnd7iE3LnmmZ6YR3nM2
OmAJXStQ8rB5ZZ1SyVYsZjUhzZFMfNc2gjeHEMMLge2Nzt2bjVVTUrK5AWFznw8YCr643xS8xO/M
mnCVTu2nliL38/sCTxXnhDTpNbTuRB1U0CcILY/Diu5TQ6Etib5taHDRBVqGnLJ3zwKFsHURRLb/
FOlD0Yf5JeRaJ2ir7Xg1S7EzHJb+0OJlORhp53hc0jv4nJBTy6zspQAfPqQapNwMrrEAjA2Z9D6E
G/ugBIC/FvJMVN+GgVfwut4oQMJTOvFUPYC1bSTeD5YrS+nZSluqT+70qVFuJ3r2nTtVQmaZC/Rv
N9gZTcdp7Ko1VaX5pfh9WcGsxs7d7RZ7r43ta913hOkcp8bv1r74rhoImLEjqWLVMVnpObxTxsjo
FR8xItPn/kOWocS6sGRtCRT8cDlrVF7UfuarnZCU8W5UWS5zNr82na2UOudwT8kCNEZfA20Io898
yF2/0/Z/WTd78X1gVXtRTqE0AbCrIW7/OqjvyJHTBLDHL/dmh48XSqhrokDsX7i65jqihxIZWbk5
1jWFgrzS8s0zRf5WHbqsYyvkn9ZNtGfmPouYd04mMqgEEe65gNHSvbvbjgsfixvwRQSfCCB+AmRm
ejc/wqB/XDf0p8ZJ3tAmGxNX8dOJ1AYpA6X3RD6by8ozolBj1pbavGjI0mK52iZN+t5pyR8CumgE
0hW8mffBC3lJ5a8i9wGjNv7PL/TvZjkVtbgAgEG0QLQbOWOiY/loWuxmzlzxrzMqRVvnVDfUN6Vj
2TWHRgFsH62CZ7gv9eZ/vSJ4VecVhQb2H3l66XdivL6ualxjkJPrrwv0nDEg5m3woqYNf2n/hYBx
uDAo82giL93etrOpJn4yNaKdngOvg0Rxae7fv2PvyesrH0zXwA3VePAKop2QIIUaWxMQ1r8sZMrs
qQdm8HC03NLV/YPkQJsj0Df0GCphU0r6wpwd3wr+W+Dqvy9KLiE21OyNm2G4AjMRKjG1MDYkGbH0
ksdi/jh+4v6m6Ne7GCqibRmQ8Fw4aDczfvTGNa2P3sZg3n5XCRTCs13cjH5hBLOZfQUrHZeoC02R
Q7qSpyW7Szfajt/3+9Iv9uGGumoA26pkfBfyBYu1Qu+75BvBYT/RWCHIumfMXbzDkHuvCAPk6NQC
BCNLm+hHfilia5WUJ7cFKfia/Y7GT8Ax4MTAEXwQIUnF7gMa8vQMSVl+23TOGvxmiPFFNfZ/F+tb
FSHUqRyyFlE6avYquiP9LsYzOxtFsK115hlMJfUjb7k20NkaFo20YCDd7IjIa61SA/erBTDQDrJx
R0qR5rxHDxeSu7CFj9yhiz4+6kiZw4TEtdu+mLLpWgEKtRXZzohz65V3jI+KEhCsf7aCBg9nY1Km
Wp4EO2DF2XaYHZmBNa59Sm+b4TIeWsH955H43xlEo3HKatNkEFyLeIC5cKPYol2AXyZTrhRrJwYq
UA1Ot8Q7TQnvW7cvVI2Lfrp17FNBYNtqAxCjfK9b9eXXnUpr0bXfQ59viH0PXrg3Hn6SfDsq7tmn
YptQb2KR/0+04/65W+lvJeolJ2tE5d6vZwDQmf8kADMVRkAAcjihgEo3LcgcT/TMaK0oNKjO3mmx
t2NCQSWXBVxvP95cNfHhbYVJIRc+yG+sKp3kVnfGPwnn0QTo8dDWvVaA3XCXQq1+tXZghfOE8c+i
2I1USSsGNnaXFxIOoEYd7UQa+Dg/xtmBkYUFTpwQCj5zaweNxEjfBh7PDtr5cGWJEWYM8riN/8ss
oh/BbWC9AfwZIdcDh5BJpFt7CP3FPtX2kNsT5HWGQ2VNa66igxVLvtAYSHgh1NLcOqcGyQv3VMb0
SeWsC0P0bGHmQTupMcntLzuFLa86FQbqCwuGq5Bh694klIedUOgUSoCnf3bBbjHk8rXDKEyHPZP6
3wg//cp6EFWIkyGLKekLowkcHaOgfwHGYMSl9gRULyg8d4yqd42W6TBFrnHqncX2AEgi6vDLUbCz
IA4QEzsFpo5M1Z6AmGlCSENFNZb3aMrdv1xZt9cNSKn/9g4J2WF0jM/IWysz9dlS0bfnJhn3KgIg
+UraP9vSxFHCnKzJ0djRhQwsIRJgdALENSqLbMgLdNNe1f+GIwUdxa8ceRWQsSedX5LuBKv/hKv7
NsSVm+RzkvGUSJA3/CaUYchSqHTJF+MVNyt2j0nlOl70aYzQ2l3YkSe2GCCeGk81QCB4Mct8cd0i
ekWMFDQiuFY6qIUuZsHwC9OSQL3t5svOSFMMqKV3IhDGF9z5kJZufNTq8JRd3axCs3f2aAhZoPJG
B21F+0Uy/OI5LYj3W2nZyqO+h8BMFAJUWl0y2NilJGgLoT5aUzbJoE9eDtJXmzFJ4UASVpOld04N
Hnol0SbSJpNuSbnsxvWYcx9mYth+i8wqvljZpCb30lAoy3N2ULniVTo57IETM9Rk8sSfTvpnd79i
P/Jcr9BzaMbJb6SBHHdqYCmiFD+s3M3HYcnaxkdmXTNfqdWfdtgGGuoi6qYYOndTP399yovUUnMz
64BtRGulbwIB14+7hjAXghjQL+4wPDSQv4OOl8LOQUuTG6H3rNGjCaXdN1F7+nMK0j28rjUqOiQa
jwcN5EUvahE96a4nP76M+7X9QFxEUIxBIXpq704yEaJGyI0KxE5sRke6C+6sNKeL7fO30AOlTFTm
PrSN0MD9KsYndWRN6qwuJdzwRorEXb0ZP6fFwNYmd0Ac49XSJ+WBfvVBQ2kwj/Mxfbp0edgohacF
0Z0/vQq1DLF54EuTVFkvhcJ1jNsklWlfT0S/8iQ/rYZiXcu+Zzko++SwDS6UA/zVwspSjgFn50aT
149SrM6Wpuju6ISuKH2c32xTa3eYDynKVAflVYCl+qKsy25yHJlAP0ScnMyIrTRmTK6Jz/UtsyqQ
gmg5fgTS0gwpoId2rOk/zEmIOJsp6BtWs3EHH+ZPSg3Hos/bXLozTP8gF1r4b6jyFl3wR3wfuPrP
r3+oceQDMzeVwDkyP2hSHA4oCmYn0M080mNuRRW78275UWfzN9I5Wpc0NmRDZFBGbLcSHyOrAJuD
I0VCCLfwI8Wu1foodYtkefF6Sdod/0r/n0AY66aPIDSDqUv7vauGLWy/Q5xLlA+GVUPFOx4nSOcK
3/C5hrL7V2LOFM4D+q2HuzK6edN/xxfaDnJYM5du8DM9DybepvhfijjwzTUWyH9sSqUPtYpz//lS
RwBIOiSzCZ+zCXc2DGN52qnpOdJUGIM9y9xxYLEnG8adzSAhLszi/FJCGtjCYDosPx/K+P5mQ0Jp
wGb8ZMXeYLEzWTWDF2DRVa9Q9NMtzojxfe1wjx8UKgDBk1PhHctUz4Xpxx03mjqRJDPLehivL75F
1Pw2T+JcE/guU5NQLPWIZH11w3HZGA0P6iBfxzdNWTwJbD9ocugNlkXbJ9C+LGJldlfrDk6yB8Iw
wiGCt/OfRqM0UVyKsnB6+Y9ZbcBsjyxLYfMZukHmk4TKxtlQnfogg8IBQTh25Sbmb1h1cc0LNwOI
YmdSEWJYa+ix9bYqhGuyLge+9zcNrN5cymcgfmTFPyGL/162KSghPKvmM1sp+pAyYB5NbVFLxY2E
wXb3WxaFsWfsPaCoZaSOkf8g/4mdm8vAM1CYX+N7QDvGksxZiSnheNA4ekOaU+E6dw84w9/ir8z5
bcwc0uh2LUFCkGjZuF7bYO7Xgf/pKNmOrFzJggvqGWVyTQkO1sVNFIN/yatwG/0uESYHfNtJ6+Wn
VgRIFQ/w5I+W2Z+WBMBGC7h8SdKwn3kmKIa1gZ4VuGrHeepzHbU4yXZGnDKp4l3ol7qf6Chtr3jO
ch3MchWAGcQFRsVFb7nMG9u2Vj2/VWEMTNjKZMZBcnvnpNWViVCqkES9inVPvBLis+Bv9EGl2LMc
bCnT7xD46Rgrs2l2spKuxoSQURwwEEpRl61ZyuvnaRz2z/IwrN65e3CpiE5QWduyRfATSnvkr5+A
6PctiXtCFqXx79emI2586jb/wdRZe96c9OQ/Laf/AmWsrYP1Jk7Ok1E5l3WCzXpvrqMu5zvLReBK
Bg+Lsu3S+SI4KfhUTX6j6pGvVJnKMswseeK9inS4Jcbw/VamQ0ckGsoUfKC72Z+ixcj2zqazjnVA
H486e7aE/Nbv+2bGjh5+fQkBPGNjv80YdGlw7OinJqVqtB82mhlkFNTPSikx9yf7Yt5XwsW3mrzc
CkTbe0IVP/HjHE+IAm/tU7gQRzKxLo/lyPcrKzp/T7A9WU6fdAEiLLleXFwp+eiHIBjNFvVe7znJ
kPcpS7Z1+klqp/rppYcnffUk6dyKJro8ef0FfrJvVZT0TFirMNbGlDYsZEZSqqKi+/tXfF2brA3l
hd5HjxARzwQy+E/16KzXbt5OKYK/Rp1C9qPB9j4zDLFGaQTum8jXACSLUrAUh0eKamAs4CtO1t4i
8Ly9DJ7jUoh6Fs7RcVPtxyMFRU6emKOS9OylS+d4pHiLU5hacCPqRtSSMtY/L4dy0n1W2Q4LovcA
y0EtBuu/599tO8qKE0H/ckwxMrwgmJq2TkzeQw5Ol2tGMQsbUN82GpU6IFHvrPrVzwmsX+JR6xFZ
p+z256ZEz4wlNPNtgTbm4bINIcO8kPL4TN5XRSNhla0PfModVfuMsbXk1TKSFz6EDMUujCLnDk5A
A+GBKxbOi5JV8H+snioc8Zb4ygGmShrn58sMRgDWsmNk+wh4l22i2zpPil3TICTMZV2geg3hB1O1
9mFzpZuDt9C2N7MQwflHr7PuSA70Zt+jXXjzoV5W3pFRUDUeG2ypyg5F6ybeY7oxUDIZqELL/1UK
BojaSXA/pZuQk6HwQ4pPD8iw/NOTlOZh4abR4/PQ7dW2oHIpgDWx64fMvSWOs4mqSFzQ9fIDspmw
2HVAfVi8PFy8uXC0tVKCeJSiBC/745lsjMCo2wm+GhcnLBF0bb1jmllEvJNWIPjJ8BVY39xHwrPT
LCkJgReXXSuqBe6gRKu5dx8C9EXrpuGuwBNMEdMuvf0LcwPbk5CiaMJ+/lQVlo2BPP8Zny5Gub8+
O7c3GhMmeMatawCZaMZPHEZAtdaoR0u9ODRw6WjmecCyRWqCOHvTk62Lqq5z8BPT16oZZG0jxzsX
fsQHF4PfpwmOLKXR0ImZ/vx9rMziWWXIsMdx0VbwzzyM3lqrRaGxSygXFzCq+ZXpHoEAaZo0EUGX
cQVc/E918fsL4EojeH3MOPYHopkvXRpM2HL+PlQgJktjNbazPfWLI9zXHjHKboBPLPgHucdsdHey
g5/xcCqWiOBRvOF5r6UVddfWpRhde4WBNF8Ndxkq8Vd3RePpTBF6Y/Gk2WnLj3MaFKxrNvM31eFP
FM3FmYT8H48QaTMdvZpt5w9bc1T+R5cPAjUoETCECWE2FX0zAL607+Rb7xj5c1qEWV5AS6YTnUpG
zle7B0WeYeaad2gABDSNZ7X13ryM/ddpJ+qFsmvLvrah9d8itr9naYrSxyOA6DVUlxMXMHkumYVv
hbE6vIn18Mg7U3DhBJ9u4DiNQV2OKNg8XCsHYmYI30xH0hF4pPLsPjSMwbBkujV19sWuSRG36LC3
jAJXkJbYOXCikbPU12cfK53tfpyDQq+MKhDE9LUYLMWZcmQXUS5m/kVk5J+jjr7nWq+j5/zF1Tob
tOwBdjD9Ttv2kg1j3IhWXzpBrrIwgJHSHr2S95IoSAD5ncY6xkl1abypfdwOlhW+w1i9Jz3PPTkU
jCM/oXtG7o7TCxYiOLhAwa28StfuRydQdobmqxfD+wasvBJo2v5tKjRxhjPaTgW2yErqeBV9Uejl
kJC1BAq/nMeCrEtAdaNbPtdm3Hf8/eMN3VTC/FoqoUIgy+pbBwBuLT3UNPJjFJbEVZnJHbdUPSU1
mpur/ff0S2rHC1cB8wHxLwCezpygagYavyq3fWUCSxGfn0NMAZjZN5Ry1mu+p7iHAKeoAPOC3nIA
pzNgkLBMpw+dumeXOgP7qur3Dk8qUoUld3XcBQcIInj76gwC1vUsbPCRnb+b+Jk+nEDxgU6vc3NC
H/zxM+dF8okEB6U727+gZj911SJy/AogtDfq3fZUETOXBCmO1qz+qvr4S+6/qldiVRScONOQix8+
FZCF6ApGXdPywUOlTJuatsQfVoGIbmir0/xXgC+KBompmA212x+Wo/ThhUO9Ea8LWfBzO7PKrz+M
gteCkXL/HFJhpJNM2Ftxlw6WwOGEljawB9lvX0ajAR42nmis5b3bGBksaQbNjG5RgXoOV5QEzlk9
DggDJjPvM0A+dtKv3k4KcphMIhg/DhURq4JWrWjV/YaJqQmb9/q4bienekdXg0OONIjqGjJfWVG9
la/mkVrlwhirzPCM4ZGK4k1G4s1zl5nbS8zLVxuDBlkaAinQic2BoCVWN+ojSi0L0xLUHQC58E9r
Uolv8fN0DpgbN+FWvtN8ZUGanfWCS2EjjAYjJ7EtvJS1VSj6tvSKu153AsLpbMkL2yA/Ts6B+X6H
lFxJ3WVJxuArXJWLTeaxMXx0gnevXdq3cIclwm+OfaVDE+PXhtjzVfpJbZrEjdQhKk/QlwSoBida
WmA7UoRSpEZxYQyJDTLMr7OBx5BGXkEu9WnswSSYax2j0CqG02K82i+2k4UmzOm1hZ5F02oczAnx
qTKCGPJp7XBi4bhYOi06wR9RDxiw82m4nmISsFPC1TI/ffOyu0QCmOFlFyNRtGbvCrUjs4Ae3WYl
8h6jwKlS4kxQcXK/a0LhKQ5Nkc6cvBxca1zjvRq3UCJ3i6j2KxQxF6BrFmwO/eyHY3TZM+Acm9yz
Q7meGtpl93F2YNt/QhYoXUdhnX1t5DZbDzVYPmkMrEUUFt9g5Icoxgc2MgoxygSvdVCgfv3iQweY
wLU5sFuxpGKMd2EJxY6Zh19GHs14lwRq9xMXY++EMXBCIeiIJJFquNSZmYUq4PZU+KgWZ0o72Re6
nRN4G/WoVBFBIlNRdMhXlf8Sov1QH2rFzHAIJWULUS3hCpctE+1JFYjyIFttcUdbj3IbSEEvFdkN
ISQkNJsb1ZQA2UxoXUV5bmkucyZOPnF6DbUHgve0BxfiYJf4o7bw7nNCTLcLbIl8whkgsPKj5MYl
tO31yoSPWPDOdaUgS3YjozpHqGpWXmIz2YbxF+FN4sBvNAW0vvLyHzyxtI9Ek2fIcwqCGdExgFON
5QEt0al5Fmr21j2VSB04USRfYBrmpaBwpJGrz9qqP4Ec5PO0T5gqQzlSYJ0/ZwxTZ5faT7Lai7e9
8xipTOvsPDXMKzjVmtnRQGVrEBxnlKevLE15YTOby1H7mWlV0H2II4eVYkEdaxN0VJByqytGqJKY
asQaWPDYaY0saMSqktkqD90uzPONNyaTCfQ/N2tAfDsJ84KkFt37ote2Fzai+3gtE7KD3xyvPYA+
YbaiIkCs8wru9E3BM2QD6ZbUpIkVAprhGHcmciwxZEzwBmD4dBmMWQuCoQaHFIRUlmbSakRA2A3L
YtTDdyb2Psro60zxWtjdTONbhWqSHc1wmC0eaEZo18DVhGH6y4OU5rGc6AgSakF7XpP4N4DrFKCI
L0MaWqEn9mzQFX/ZezWZVXXTh4ydE9j2SH+4I6gp8rJlkrDam0/uoqUwlMVl4gmSneChMx/X5QwN
0Sjfx6qhA9G2SZhreSQ6TkwQ7Isbmv6YXdT0ZaGYc67lCiprJYzTrQAWWqThCqQ2W2FTw6zRHYUm
BkQh5s3/p8RcKrnTn8prulamV50xJOnEJOnjWuRlLDkcUzffwqk+GfrASo/ixCRFgDtZ9C+Z9C8r
BoivjO7dm0M+6BNUpn8gIUB1e6T7FmrQvKdM4QwioM/7HmRHJDcxVklVzPRa9JYqAc3A4ks4GvjD
YD8rFemhIBYqBygdbw4Akxju+NdwLP4VOujQT7F+dc8FAZwR/he+443aIx1B3SqHDa4T/Jm2zUG4
/u6LTumArljEbE0kF3OqqPSy3exdBYZTO+kcCxx/IXCmYQnQC0IRR/Yz4TuXeQ2QaZB+Q4geAsHE
wpyutJBcxOtF2Cbmi96t0R3FU5J6MSs4wQ1HCzvmBGNXavPINQDLVoZkqcRVZBTWUWadefV1u/mD
0BB1TfGSD5bJ9LGMkbkg+WknWlILICwyAVkHPfgNF1i5YsrlrTvHvp4QrsVzouhaefREUQxu/oNl
MDVyborlFaPJo1EgRdW7qQBMPJNgm7YhhD89XdRwn1XonrgfcltE8h3FIMmebJzDGuP4VzWNfWEd
yDWRuhLoXbbwLUZap7g6pZksFXtNlERM7ScoKwdbfcy+EHBMkBvahLPaU/jUhUPoNkwgzMhflB1U
amz0QUdEK4ZUUpcitqkIMcHhUjq6gCMaSMkLQdBNOB2HwgVUkk0NcNCdfa05S5qokr/MrTYTt1uo
B77tZeVQcMXPFf4Iqn0Dzu2uWHomFSwaVKBClsMccV5yuzUHBKkffgU6vQHIGHfmPzuMxMfTMG/w
cST/XsRsTuZWV0exwC4rRGTzUXIYPpml0+zo6/TPmMA10PKBMcHVXLDk7PgBoPBroI7iY6PXVoyC
0W9EFPRnVkxiNh4MApAgGq7m8uKdT1uFTw4/KNhIcz5PlYQ4tpGYAOhL8gGkq8AnyJEjOlU1neuI
QqzwHJBM8ZXOujf+bB6S8TbbV+2+x7mZHpecvEXjBKslfBdcw8iLHFoIANpPi9p8pVEvwq4+LSyv
EEjjfkpxVSPH7k4zKIn2+YWws74ZYgmUbuwsvjwLNzhBOMuh327gM1OeRyABzhIU9O6xU5C5ixzu
iFqsuyGy4de7OoEYnogtS1eIdXQT+fdf6d+4Cqw+OsyKen6YDXPti1HiG0Vv88dMtm/YGCoCuQgf
/gFGWK9kL+RnwzVDiQwsvWmvSlJAxjOFW5NdT6nRpvnOcIhRQL+K2WjMasPULYuTBS+CD1Cc/P0L
YmMoKsytkGIaBNDWdUYB+/KkOy2kA9CyugLtKNEyCKXu7yFwYCE3oTymg+yvKyLjBzXdiBYAU6zq
aytkMa1eJteyDRSudv36cD5Ld+Kyl5MaRibgI0XxNWTzw4zAMkP0ZeEWtGvpKXsjojk5U9FoVoRA
7Ta/T5nfP6LkdyroKU5hML5vkvdMthm1SZOoBcOQzIKr/prdHX/IPVNe7X84iFHYbO26IkLYEKZQ
K0aIYXCwgsXv+9qCRt8YwEftQUx8Oa/Yj4g7s0201w/e7ZQxv8roPmh6yBUV8B7XznLQHoaQ2xW4
5b4KyMz+9V8W6gKY8N44eCmmFYhvzXdPiOPJjVXvLFbf1Sa9iDshzHF0shn8XTDuME/KrVat+htn
/79ghIG1HAwAqnZcdDckQvjlYXB8FwCJhSBdVjAwtroKmr2sCujuntDslMCjZ4iU7Rdn+m1Z94HT
JILrevs8XCmd8GRDtZ55DND2uk7MpxliFrQ+j9/SCY2MAq63J0GZew8G4e1ME1/V2A0swh/t8sY6
UUGZwJw7aX0u50poHn7mDYtCM+0CcxKKxR941YA6Xb/q59KtENZDYg7wz6SgbwnNCRLxjhHsZhN7
1XfgGe0iRgnF5fb+jabFuaJ69iBHnpKSVuJkKeZbIhDEV6vNpZGJD0dclYM9TyBMOI9m1QBR4Rkx
Bao7LJnljITBaLhAtbTYPXHBgD6LQ5ChLyST0Bi6xneEMQ1fp7E6a5B+onqaCc4RA783vd5SfLdy
OXs/evpqoNUWFOR401YeFAbL1pIZXEjSg9YfC2W3OrqghZUz5S/B7v94k69B17zJeJ74bl1AqOUR
i8GjU7SPWZFvef1t4KXpAQdY+7PhhYregOvZezLpcQkaFIDrt/FwZ+b7kfxjXXa36Ta5a1ljx/l9
xyW8ZTCYp+FQTol47muvkeiZlN8uQ0KbAOAq2mEWYOzmKlPaZfAZpJLxpEf22XWovrWwVMAGHRg5
5x/n9sak8aMDdQQ6naysq6nNhsUJqjITAoW41kl2RQtOr0jlrAEJwpeVbsDi39995oBfoHORDN63
ZvQwGJjJxsnyKxosqVD2R0BJnhNvAevIIbLf5GHiwBhycQ/DTDXpaC3ZElxLwl0RU0dKkKQUuTdy
JC987STWGmBipI7z5tkdlJdw+yAZPNiFB65ZEfBribFM4J/o5RnBt0tmorw+CuuTNyHqR20Bsdaj
jy8//1mfGc6lC/vplf3pm56sMuArkbhwYEHBX/0JqjeP8TK3lpDVADp0/ux55Eud3X2enFBOIgz7
KYnKmaMFJNAjtnfihWlxX2ayOANEgCWJhMZs37agHRuMJMAv3T2HwdV9KoLnceag47CYEIMxyp4b
J1WVVmIjmr5mcw9TBkK2pq5BoFOwxaJtmwuorUY3sSeMfACHfvxQTa+s41T37spxleqaTRPIzAdO
LxaCmDWOa/Omls/pSWCASVGjvJtWRrwjRHeD0DH/9fwoFJCoQ9r6lUheFkKA8VyTKWh9GWYcsN9Z
2VDzmAnBEydN5IPjGh7vtgh0kKx1FWaoBBeC6uxcsn7FU2kHsgtvSjC1eoXybmKc1ejtxvAuo5Es
DjyOkhR6skpr7C2fYt4ZxCIYu7avqqPvdWwx54qRNR3ir67Y3gDgWGTr96IbyfSv7fC1RaW4NBpU
3qFrhXaRmMK/69hT1O1BFXPUT2db7X8NkJbaxhESXKRW5I3t/yJl2gMaFHjfK5/Aur3Wao9KWDKb
ZsBFilUt6PUNMDEd0h6mbMgHdCO1L8JfklSgWnOammr1RzZDyft+ibQjRkrzRHebwqvT94t7yfBJ
fIdcaMOmkvpTZ456Zot+n59bxGx92vga+Mi9KbmgR5zclaayGeisrnW0yyg2l+5lsePfsxm54Q9+
Oq/keKDp3ANJHqJfYpzCvG3unaP/CuHO4v7SOwn1DMGWSYFWx9mPAnQ2wwJpz/gs4fxuunowjjXx
loGFIBhjf9+reXeYBo676DNKbNaEMMJPlASLqEQn4OYQZphF6KvfdAq2Vpbm1au/6Ge0eLa7kcPQ
wayy1bTuCLrXZQ9C68evpfdAvcvpgVcCFb/wizdVQbRDVjZNuYQY5Vf1CzNsxu/N+GtpWFFKEqQB
epKWMTdriJ63LMrVNbI6gjMjyF+ceQmt7xrnof61VnEZXq2gULolLmvBNkX1tN3Ou7uYKij8cQ8r
SS0Zcj6ah+lwlAh3sx/5sCIHRTpvOcCTZJtM6p7NUH/QgjheZNEI8LKBxli8hWm8IYR1uWhkb+cK
OwYc1QKOJeQm3K+Qdo9dUyaRpGLAVhqbX6kYwPyldMv4dBAaRw+0WkgDq88XlKV3lECE3lLmYXF9
EPeVJ3oA+GtoRvnMpU6Xgij1CxlVI2clhRlqEPNoXoZuYJbkHVABDActvLGy5Po5eNh5ac2M0GkL
vDjuH3yycGvNSHv1zu1t8E0aNChsB3S6YFrcSeolfEIy/Ni3cnKN93mZhDAb7Bz/L+qeaf/GzL0s
EsetMTle/DO99IPYHTpAD/D2u01aP2uLr9ls3uHNTD0h9gIrv1IwiQ6mti/8mdVQ6YtKGT+wvRyq
1CfyTO/RB74ITtkMcEkWltn7YjtlgjyF04lAROKhgT7JZ7TqRc+KuzbZFynhDILfu9ZOJR4pOSFx
BTp93aSq0eMiGZ9hiRZPgmfy5WBpz8g1kOqaTDUEroeYIPVNKA7WjSopigd7MUVwldJKkKSrLpdY
jTbGJSSo3ayJqM2Hsari9889M0ne/Ca8My32qLGIuYdmZAJleuuEDp4vFr0kY5gjKEkV8zct8RMe
w6YyrjxLYBH8GP7OUJ4wBy9lpNy6wcneenNVQsZ/h44PtJPVQ5ZlIR8WcA0sqNgkQBQpglFR4Rju
OR6fGiMKpXTCmsCA/0DjUB8ne/YeDQuasz6l6Q5YGdqeT3S2HgGAZDYtToY6nLP1Z1MbY818nFiI
wIo83bYMnEWjrFA4MgB2qMKL+b15okHokXHf40++eAq2Iwhmt+/BM4kRVEi6I5g5r8zoAnvekml2
fRGu6tabM5t10g8oXfJxdq87kJzYkBvIwi//EuV7PO62FZf6vY2pgbg3dclr0OTXV1Hp6Ae07RGM
/oXHXZBS3ZySiy3Kc2vw1xtO2TvLruaYzbujwzBlT9rpi0fCi9bT2VaH0hwhBRyB+TZ80E/72AX4
zgdjWQCVO8Z/l6c4nzpH/guf+d0JMXSlxO2gv0bdAemR7alszepZZ0o4ySj/P74TLZVBc9IdGywM
D/c8id26r12uBnoGI0o2/JvM+uIXj/1muMn+7IsEaDyU0d09KHppzcwXikcUBfbUfzb2x1geauz4
CAvtbKBsToPxde9CKAK3nD8nhpO4kTNaoK9Uc50G3YT4dvDVYJAzWSqThrc4s+bOdjJkWVFF5l2A
IEEzF0+QU9NSkYtb6w+fAaPMfLmTcbegbqJHUAtRvnnB7IB6e3uvJYhVsd88sYCp7n7rb4vg67kY
V1xLHCpU8K5j+jo7hjs0wJTq8A29dvLsmF6hrtuKO92pFjN+8SlwqbGtMvpMYd1KImIvMHyNZ6pE
OJqXE5Fp87OeYJzBMiO6I+Z5mdVmgZeRyI/QiMA6rvhBqmNrH7GiEqj5v8Oz9IlKzb5slR+yI0z3
cuQzZ1+ZdDsUip92zRKTonFZCB5Hc9cj6f2ewmY+rYYdeFh1yLPcu1mg3FT6g2PR3CoDFJH72f7G
MHuWwy3qX1kX3mZ3UwnpCx8fpHQ3Co5V/y1VasRut9G+ErT9Iowa5veA0cyeAgfPxMoEVLygRUGk
eUdP2VRj7Ga5gAuPjjPr+koJNzBSa7mrUy3JR9ST381eOjIU9nRUtyhNmedmzBY/DDpybn3t4bB5
6W0U7C0YN6E4jpF/UEPL32y9I0fBlPiW9MGw4SYgYOgCl9g1RpuElcOhFeKyMdzf5NMl/s7Awo7C
oRZbLjhiNhrJInG5mIcjhZ4UbGGYJpvJNPVPsDuSlt+hFrqnEZFKWgSFOU93P4VwCJIxvC/0MVks
XpM4UvrgEa42/43d5rPRX5qeXA7GgEuYIIhNjWjFs/9bNQv/1grq7daJpAeKcrLHDPe+W4bzKN5M
lDXJY8NCizX05Q0SB8mRiy5/mGhUDUce7/cxqelOYssT8nb+WtlegfaELU38DXRTxGLE7+7jN3UR
f8gVizwjkf81n+5rToBuwCxoxuj71P2pFArShU9OHdhDF2X7gCsP39VEYNvLaw1/9mBWnfB+j5lj
D5mqunA+McHWml8b+fEk34pG/UFslWyI2z1RHi1mYQuPk2M+XY1/5WrX82Z68/dNme2nLR1CoFS4
hY1HWToOTZIWjDDBPZVMqRORdUjE7V6U6mwU/+ltvvnqNwTphGc0rRR5WnDgjjorUF02WDvgZ9xW
6y4L/i3MZrxdUmS8r36O8VYCfmyh1ekrIFnbfGUbgFMhL3RjHE+j2gTK4Ga67dbZlqJBKTF6Ksg2
FhR1URp6N9HEg1vjRkPq07/SyFospUjt6xSKkbcU3xjc1I1zA/o5OrKo28KNKKI4pkgnshu4MqbA
FkCzNoX5g3Vv07gdQ9zXOdaqtXcmtk8p0hQHZO1XdCkA7vJyZBzXxQjxLgXEv8WZKw5DNkKl5eLR
dtiIbB0HWBolhyu/s6nFByesIJN5XLHN0IboEG+D1t2fPvpFRIfUL3deZRZ4lsiGI4EwAKdkhIgI
5Oke9GRbKTqgLLanoHzBuHtbasAx+fBFRovzkgamjKquppTOGWNsz+QWodK3WD6Gsr80ZR6cxmJF
SLa5ZNYc8mF1HsjCkEgRlrLyz3e+fo7mLxImitXkJH3yfwmWL/vdqMSYGjVDRU/M9kMw6S9p6LPP
WxCSrGN+VaGFIkeHkg3k+P48sEUrv33PB4O8gaRqTGKibZYz+tfH+IYg1jtuaFhWmijdC4L6pFDb
SY+4C2InWqeO0EgeXLv36C3IO5V98WXwfjru1wUN6aVEJPQijTXNYnM3+VSgy9yfJkrcM65CDOkR
QqvDL+eptP+rcer0KKjmZfPvNf1LSLdK7h6sOqX93tV9Uw67AtspzyR1uM5rks/uxeavKjJ5yffZ
MXRlbiv1m7TjND1CuwtTeRjdr7ii3reU4OFfsMWuigDCAglb6k6cB6ZjvUmAmmGMBiW2+72ZLVmH
zWn8bLx4XdBv6rcGspi4bP7EQlW1EoXdc4BkDVJGlkLhs7yzoEOmdGwyMxv7KlA613gM5zQCpujE
lZHTkDYzzxU6SL3Gez5xRx8gYZT6B3x/6E+zln5EACncr3gQe1zW3CGAQ8eJoZUGLj7Y4WyBYWpa
/se8VuWqEkQcmANJBthLlzVstrEtS9DjK+sll6uclH1ciZAhOQIZw3aO9K/hC9ezMY7ElHa/7/cL
Xqcz6eIVCADgAEifC0pvmbm+1cGV9R1M3Mtk0xQSOmBmKr4qStZFHHaOl9Ew7WUOe7Q955oIW4aE
aDQsM6+1VbQAteLdpibvYb3CC/SFMo5jrKQQa4JwDlU7wNm0Qvk4enZxPbEOv1YrsTCcgVl5x+7c
b6Wx5Y02iaLo2uA03F5XQARKZD3xOP+9Z2ksz+vrSU3/2tu100m3dKYbTb6ohiNapLDfCNQ7szKo
E7jLkRVRLcJg7avm2Rr1rJvAe9oDxgCs/pTG9LXCt2OyIdWqoxS8DzH+ZfSsCYNQrBSAZSa5gbTM
8TcfKnnWY/HeC0wM4uMw7RASV6XQJKW8DkcpwcKu6wII7bcCejR78oekV1HNdGVo1C5BhnaklI8U
NYWUP7TK2kvT8Hv+ZW2NyKa6CUvCo5cTKuqTrYVqqtibhqscfaiEbYCU9z1P7TVQX1vDlD1uS4Em
AR+x5NqhzmXCCRTEMxotkQJgf+ELMrzIACvvOYpOug4UsxWN+lQO7fVZFXEr4xRr5v5LFGmHReKw
ndo/Jaf2Z/sFGdlIHW4DJbU3nomkaPe0WZ1noZu3SZ0LnixAQSGqjrThq26gzTfP5zTigc4ytS7W
nNBvtMeVbd7cq3fz9/CvNApIoegeLEwp9ZtN4H5KeT+0ycoY4gQsYjxonr9MgIqFdfVhJj3a4Bw7
vQcqrpp7noKooNk6C8qvSDDuV3ZgNnkS3KX4ipOZ6hksjWA41lFloEmc2dq75lV/55tyoHL+xAI6
h5hDOgaLl+qXR94F/DZjjVB4mV+1ZTxJdeyGopF3cJWkqCAdUeUSa7TXBG1jwmh7OV8Avzzp/Di1
IfAxHOjPgTb0n8t++kDEXsR1J87frsBwWWpIkqJF1Vij7+1ssPVE9+vGcZo+J7eprUuz/3+qclO3
qT1L9pgEfJHG9mIs5pk3dPntfMbuWPmhDXuyw2L3FGmsSa0rkvsMTYZbQgNEy5KB806EpVhYYs/O
BT9IyE4R5ydPAOQmI4WTvDvm8bx+NnSisLDuq40U+Nj1X9+ps3NMhwly+oiQaWuCNMF1+rbSI9of
gmSUDbfhbA7NO/vzGOm+ITsNjftl0kHhtRYYI/vcP3EvioSbtAhRGg6bj3XzswzFYBJKM+EaLhD2
5J0/vLTzrhxsbEIHxYLQzFM2s8MxPMehMViD618dWrQNIdSd/VwCUSXb4nDSbfmIhU5tOdL8sQDc
utkzuvOUGhQaB4wWeXRab9zQmECeDN00zkVsAdpzs7vnRaI6pTQsbexRY49smKoma5IEX3nveiDl
940GonNoeXEMVzy8euc5laap1OoZm1V/rHf1I7xuOtpA9zfRcHWActQ3riceLx3yWBZEUHVXqTRF
gZD8DniMQlSxJvIzVVF6QIagiWFKOzBaKaeIEUNV+3Hp3ghCpMcNzO2/nSLCHZ+DXmw6pBJVeAs0
qHvva6iBpI6LTedtJVn+CH5GoSbTNe29x6DvKuof0uQeNgJkzyrR6O4vrs6go3uppGB7CdP2j1K4
jBcf8+sfB5A+rrdkIT/BEfh4/MkUYESqskex24bo0gsCg6IwRADrHi5GO85p2Z32mySvhCKzh+fy
/l9lHSCrcu/Wh6DxpVwzh+I0qhiM4AiyR6MrMQA5MGgjXRllfJDTodhOpLVI8yIpYSwBrkSBhUPR
EuZkzIcD7Z/qugiJc7tCu5Z8xy2IMY+CfTOcvMmE5p2Z/Uuy+l7pAsnTUoLeywrIRgUlWlXRxxmZ
8lUtWe9F4QhSvE3AYAjP+PA0dIOnEdnNwOpciZbbXgbrRBLEc38vP1KT4HbshwkyvjptQyDFLpPh
dToUi8AiE4GOssKX+0W6Lo9o65vdD0T/CKNEFHQ7B57nW6uNNGRvij6QTEgln7GCk+LrPES8QSM8
qIMN0js0z5D0bUcjNC5Mu/X6/4DmH1BALfC3kXZIUaSF2362+Z/qsgJt0vGlJvMGH/nXaMbyKyA/
E6A1oeOZYq/chy7jF7uUT2m14t5sdpe8J2N9JehdrCDHL1UdlAibOaTP4F8QdZeo+qPoOjqcFcUW
IGeC0v3Qdp3pf3dn0CZnns9dcEEq4D+DdumzqFhVAbsUtEgwKRhDonKWocLGxOsQe9izpYAuNXsy
7pu6H6HjSZtQwIFcj1BC4aAdpCVUNGG1UoU8Dljz627xSfgvDWVaSnQg6QNqtLMUl7Zo67GD9jSC
/w04EZGzHzNIqp5E83UKqLdsbZ3JJ0HPfRzrPewn/nPlRowC22fFmukMzG/yeEwvQ1bgdWynXPSa
DllM51Jzr9gGCFUF9KScI2EmqAw9jZoV9BsVHC4rqw5SVMtwO5PNU5Fzj+2hbmB3/ajGmWtmCZPH
eKEGgMR2f4MaByoRNolswCdSNv2UsiCpGHu286lq0QLdYjNZpr0ZzTs3bf7Y6vZ+MeDGlBocM2oH
V/Exs1Y7tOX4tg4tKO+TLOyAkVK3yFGX2Kbxa9odYcqbuFh2lG7NCxy6o+J1CPslSUuCZAqfbfwM
TDcXW4wE+pHC1HXZ2zJOoY6ljdNTercqwB891iwFQwmoESv8jqqFeqePmxOWFSnTT3SAoOQQeUxX
Vx304v2AxvOO89c1yXfTK/lQxziysN7qcfkWh8Qj+BEvi+DMrpYsMkMJhDISwuXPxKMDwkkjWAD3
seibRseERJVqC5gZM9iNjHtC1qvvNbPEi7sH2AktFQxylz5qkRroud4o1LzBSBatpFaKhW4W7Tjc
mFDmyaw7M+EC+5C9HxUdIDc3GPO7oEXw2thmIRaXyzDMfexvyGXLyeXEfk5+2xz4n/TzB98UZQyr
iYBbz8/FTVWo1CYbX2tC5QIfdDBVtgh9YAo+RajtsjecPLT2Qfta1K8hdEEtY4wmkaMH+A2y4M4c
K2q8PcIV0FpKqrKH8rNWUq55UZeUNltBN1lKRRsLjjAPzcs4jE2K7A7em035osOOuP0wrkedPfuv
ET4+zQBvDCaH5gxjgFzqudjV2tHz/S/1T1bgxKUBqV6JjhO+jUk6s7mP/UgzAxdF1K2TEFo9YbfJ
KZhHr2Zq+OoBYwmJ8eiqCkIuxgmUECpMSTK61yOx8NyBvYnHz3V94jgc/eQLaDQEMcxiM7HTg35A
YiK6sKswSdViWY8ZZR3lVlYtIOpECuDNk95MPRsexRwZ2wxO07MBYuO+5PCtZxYjWblXKrUbmCsr
w2d232+BMoRgHDOm0ZM4N7HLXjO7vqVCJmpSuWYnOJYtgExId/oZndRmVuxjm1OJQ7ueP9aMjavt
3RV92gVKP9JPlvHmpfmJ0c0y7ELiwK9jEG7Ng9D6pDKqUEU2+98E91Z3T0hoTYviO/obECL8cSa7
jS2tBUvvOqlp6NVRpTTvLob5mjLTVhfR85Eqm9tYaUVh+e9ppBs58k5mahUjtPXGBlT9snCqV93v
nkoOxqOfBGe+8g69rLUnJwDiBKBj8wECliArwkDuwQmCgFxzTOIwKrND6NBh/Vj1BSCNTKFxXC96
gpGGIfZurLFCCkS9Ji2eb4XTw53iabFe50qHw35LHjIdmLv8geM7y5V4Zuh/rsKHrx5w3NOu5GpV
uMS/EHf9RW5VL8vxo9tE3ju/ya59mdhmFSsRXy9P6R99ZAipsDTlhMsWmwuC2xxiMCfxZbNwAzl7
BYZbJsCbIiiGaJXow/f43YWEvY8Gbma4H/tOFRPr4qF+E6MN6PuV1ET23Z9BRFnQOqAjNd0GVSwx
VbsfpH050OIf3DBbMQ165aDSLWK6PQlreo1wffNB9gBzfGC3h8GX4DrjL6oUq2LRtw9ltvMzOFzw
HE+4tGFAFk0YGxnKgmqYTU99Fu2zj0Q7wCdeaBb3ThoO4fe/EcZ/EFuDIBD3z8raCLYRcd49f1gx
BtC+WHI9V67ecrX1qUBYPlZcg3MrRsVkykkaT99yrzNkCd1eTByB4h4Kvem+5AVPMRiLwU6KRC/n
0EDW0yOxK8VbSqshuDh27RpCJxDO2YNEl7mvXDiJftqjQXbgNmjYwbKKd9B5QBqUubuYQlbdpJ7W
JQywWmxzjbOwMhPDFJd257hDI4+nje61/5wsoZrz3ZeNypFLdzziLpxjCc5xe2ZAILD+nMmT1vNu
GoUMSZEblf9V+RCeMwf49B/NE8wx9MyLwPkdE6ws8ATW9I8zXsnpS4KzNAEThUBUlezbEaxw2JnP
6n1O7alIXPF2LGbEcOi9bNAa9lYL1h+MTMbuDD5xKIJzdnAqa0UtewlvP5xniYxluzFI9GXTKGpX
QxlDO3geSbbkzhLLCsb7t1hOcsEbGp6INLbaPqWAFLzKvWW4gkbnsIjj0a6bt2Bf78/crdl0Ta0O
TDUxo/SGS+m11FCK04H8ja6MaSHfnxFRZiQnUKzDPQ5FpYHkVh22MIT3uG8lSktvVqDnEjQ3fvao
f605lBg1VRUrmnTOBfLogOtSoMe9HNVBM1wqsaXEJ8Gf8mRYJobW4WH0PvY12NQp1Bt1BvPHj0ip
LqEVGqWvvf5vPr0COpO/UPa3T315d17dchADLYElubBwZUGFWC55/qEV/VjJPqO/OLw5Xq6jitX6
Im8MA7H5dJ8teJhOUTnIYRchlfkGRS2iR54cfVnDRqxE/8V8jt3bZbHdM6i98JXpoaQYTJKjAZ8c
biTf4NVScW3sgQW/ODetTi1Fq+QBx/Dl1WsuMPkCPi2ZVUwDVmweBNvMet9QcZGkHVWR8jGWRVGF
EVmGp7QhtFdhKDaCHp4KofxbfrA3KTX4xdhKMA3PYj8XDwODJCUo3YXy8O5Z0gUkkiKtrdaFuaHC
ZzNQs4RSVsYxaf8D43sbwKWkBw87NH4xxIyrv9e3qpapydadYZph0TRG2D0qckVUX8JO8BHVRhff
/kV4UttDmyYs5cqP68rXhj0SslaihfntGrKwvCEhEHu0nskYZupYAkNwXmZbWioGfPtjjc5Rvwm2
auma8v182+hahsNwQocEuckv5tWVbg6aIsUtA/OoUt7s9cEOqwrJrm4AJBy14cm5EliJfEzDL531
wc+Voq6PQOhVqMMWgTcdja5UIabvVipmGhlgUTw4rkUogb4G0618GuYtBKZA29xt1/j5OCme+t0g
NzcKl36aN1EJ3XtJ9XddZ0ruIL/rYoXxSlylXr5pdKEiJmVRA7MtuyOynlKH9RSPFNVHPrt5Uww0
J5NiyhltNXryfyyI7LP4T5h9qMdFtFmRRBB5VnqqVbwVNX8+EcE0KUtZASZ49pqIg2+h0cRacIZG
9V2WzbZFlwb80QY/8UcrISX+3IKLy+VnkVmH9S/9BRQ/hUUgh05I/DmHUVYFGWhaxeGiUtiK7j3s
8bTg46vtz3C4jrClqjdgmvr4BNaJJAP6aPQEpWkNdza8RErEM09kZ/Yyz5hLxJNos3saM94AJ4tF
c3UXxM6DrHJ0HViI4Mp4PVjBOpAYdXMNoYpGsDvV1cFxxeh5u9v4YoI4e7FVEgZyih67BabRZATa
MbwLk95dYRXe2X+yZ59gStt1wDWn7Ah6G+WdGZUi1ApJlGjaYo3jbzqLayWmnZpZpEBfjJU4pepe
mDcz1RnzvSwl7XDhu4drew2M3OR6+oUsmkpKh9/Bh2zMMNHHyRU+L2ePdJ6jTYrB0Ads0gLXArhs
CPzk/wV2A2C++pSy5s9A9GQ+lsVaOzUtOI8wj8FgxtHY8F/bVFuwukOLQFDOsDI4Kq6ZlC4F3Wi+
tBvZu21CpS3MDdzCPIl7pmRy86gKq0ZIOdQwG+YA7SAEcmyHnBDIfvJ6Ap7uCf2h75rzfr/2/sZ1
7LZfqiERvql9JaVi8JPMrKglz3KHwFaa3Fb3a8wcy0cmk3TNAx7i6UZexy554BqGVe5vsBPezKPe
IH9f93+QI8QyiipLVLxfAt6Lhyd5zq63AhbCL+fTTURBioaD8nxk1ReOXsMjLLT8t8jrb1WXpKfV
84OZrPy2ifQaP+8XeKDmDPXC5dZe1abqnAjc7yeLOwpgWCwVSUdmFjR+Zykw6wdn7wLZezCygDQb
+Q/hxNH13b7QRw7S/WbtzFgEPz9CjSTXbOlriLhA1ifCVZUDxtksQjw0R34zyF0V9OTcgusbVV+t
f8H5yFYAWKSZwLF58JCiUMTV6IzqLaK2/sEg4QfFuUfh4/9xGrcjKr3tXHKI0cDW7YTOSlDmfJ3s
dOK7NBSv4Idr7km13vZ7w9TAl3yTW5jeupUP/ct2+vPrO6CKlEpqTN0SwFJPWTJYz1NaRiox5nF/
L4PLDvs+keHs7o1iUWeDJtCQQSxB17tYhMkZGnS5cPkLWUeVuzolMzNH81xW89masinpSgHJ7un4
deytUC48SHcJS0yCKS8c2lIWNCKMg/8FcbiV30BN9Z/ZHHrXkaQAZXLMhfOWbDex94hiGpBmYeRA
M3GNqVK4hh0VvMYzt2M9QsRscs5fhk6cpSunQRvpwUDqYMJPZHZzjfdw9mwhQ9jc6OlBFmezE/XK
sdoj7ja21BwLcMUcq6PdAXCIu9JxG7CQjKoECm35WlEkJggjHM0+1lSaXWvpxvcPZk7yiB32IW/G
kHE0Y3jC+oR2ettZXBBh8TNsM7sX1bGWPcqqv1KTDkP702hVRsKvAJSguGcs06gXeJF7LABjZjCL
odiAVLmdwvhEwQ1/IG0PDR8O5VejlVQ0URSLS+qLvCd2r3TTgkr3Dem1xxR5TUspv59gqAXuAQH1
NCsp+IPBv0YkL4hURBjUxClnGHVP1NPHRVk71vKoIWeLMrMPYFTqkerEzLX37ip7bSbNO6wOMkLp
GpomLyexE2WTYu/6CtLrJ5oWqvuDEy7QafwRCD5iDl3XYDqflQ1exX/W0RRcA1irlaIGkxzg2oDF
CI08Fx7Y0TGH4ZcYQev8EMb2MArfYRlpV9IgMXFmwz00Ce8l0tQNGM75YhSrkmJpCYA27vZ5GI8O
5qVtUVqDFhCpsJOKDjvl8UwMvdj+W95V3a31WXYF/sAjRW+YcoUepU+bloPIZMGRJtbveS5ytnMM
UEk+7+kquMUB5r+y56YmF1WXseiYFJ2erXFhhZEwoIGJN4PcfSF4Oj2j9d8aSLbVRBF19PNZN5dZ
SnFKrIH5E17Nc9EiU/RyRenjtvvF+Y5iL9I4FLOrBzhU45oSC03LdVHGe87d+3O7XsYH0ELtyaux
e4FDOmLGUTbzQMC0GrKa0ykWugrsC0cXnz96PlkalMKqO7XQYvpdk8h7je+1KqImrmuss0DZCd5u
ZCpmaX8sUIrsAEuFXR30DZaXJ5sapIHZ2CzJP9BIuaCr3YH0xVuecord/jankHt97wholRKdQmzZ
FFbJ8h+eVGxox9a/N08Ewe6qNb7ZMHaD29OMgvlGRYdmHfkBgFQDZ8CF1zEiaZVpzZu0fXSzJABf
K6//jqq7e+2Y4bcbzkMpPZoOl2Fe000UvY37iF+BAfeN2Za7H2dfwIfVb7VKhjb12hi5SSHM8hO4
BtCzFLS0/+b+8ZvxK4SG35agFHgVmWoICDzT35QReHzniz2TbM8ILEQkZQOEThLBpMYzOK9KN9n3
zzn7kZqCNsDqVSl4EsE1/PO/TZ2I4a5e5MNaeqgx6Is1FjM5R4IdBGUXvXoXBFOKF8EtLkP1IfuK
2Rce7TBVZOCcAR/Kbnagn7hUH6mOep2aQtNRBoeG9P4W/VQhLqOF70cbWN5y+JdDgcX688VaDKNZ
pBXuSngsURjmAoQPzbrts9qqiSO+J3P7BMzTjmG7H+nC+xGpTfJzSeBWWJau2ymnjoXShxxlrVfe
dL5ir3hC7uqUuNN8lLxX7tSYNFjrnZxvC3Uv2k3gE+RhwtxiCXj/irAwv94APScznWDF7e8mSe9k
HcQ4F+55QXeBi0DnEpwqvlhuOZ57qdCH0hJgDh1fMDKgvBAN6uQ/INVQ5d63zSeDS+b3Dmv0OC7N
ljkYMS7Bz3kjamiKDxm4SBCMYhCbBDKIfH064rVxK9YqBI4fYshgadQRajmFzuBZv0J2NSV/4lkq
CeZ+9r2MGwcwg+hBLAdIO+tMB9Gm5yLk+yZDgdPRgb7C4FAda2hnbax8hieNrOI97shHky/mmhlc
RyFaUWAz2I+svXLiwY1a4w+++ccQQbBoIwGI5I8kwqzZUU2uFrG7zwEMrQeiXfsXQd3TWlXPytXx
z82EpfI+zKYP59dVwAb/puOmBGXOwzyNikSFDDgKgphMqHtvZfYk8iIj4z0ofPrE9YniG/lmPQnh
sqke7ZOZZc5kizQZ8FAL3793lIvqdeJK5m1hOZzZpiEzsy89CLIEyNwlmhexSvqfI2XvJG5DZhJU
oDRblEjM4ZHezeR2x+meK8L+Qhh/y1FBK5OwpvzDN5iMT3k+oUxSJEyV3n9j24kqdpbEDU4SRRSi
nmxzqCwQf6IfuusLzqXgXjjaaaz+saijFtyLcuCmbTiPuz6j963dlqrBPsLrwdDs/eGEb9MInR3T
40C9/NHJRr4bHGnQCTsMTYtyx9pRMeF5PKEUVCwikrGL6gypmSNC3YyfIQc6vNDiiiwLZQ8+0Mtv
BZ708GVO2ltD6EykIUTL4uViN0w/uOkfqz/X2LwnXxBqBJQXm1uuZvHl6vC6fL/On2Ag1bG3HA0s
7+ffteQzdeHo0Rfq28ybKkfPBAUokkfaIQ5kcW6QQzOUBlXunkeu6Zg6nH00OFQvMQRagN97b1sn
SWg87jvPSIaPoo8KQFgGH7NMFwkg8RG7nbNppNZ3BKNVQUIv2N4ODmEcAxp+uIwDYKS4Jh1B4Atv
TpID+qTFv/kOYD6IxM9plNTOgFZd1I9dHu7TSjiL6bKUrELot52svmYqxT3HNK8Q6kmx37ACA4UL
F1t1/cXefTqDb68Nm3pclX6P5c6xKUHQRlNfW+fcUJBc06Dv/G0kUGwPYadH/E0KCvjnD8VWrw2D
XBsLlItBQRM35efhGESA4faW+z3c95fYS/yBd859iwC+9VQZ+ypvD5YzAAuKEDNMEWUl9dtqEdMj
V2lPT7Oa/NwOVDhkNYv819ykIiMqSqgsOaFkATMaA33vcYE1E5TycNQdtFP6kTxAI3J6rq8F4UsP
rvlfDOtqgOawJDqo8q2eZk0GX1B1EJ8vLl5ndu+Gf4g++lm/EyYhK7sh/7ad7CxNmtd7jOzzKkcM
4+7jxDwOclGLlti8cfttp/ApTfo2o/+ICqIOUQytxxI3WwSESFfkLxhVev+XghwXFUXF9pgPV0Xi
beiXwjDWh4MgvknrYceSDKHDfmigp30zUdNJiZUd5N/BuKg8Ri4rTezl7ERfc086TAJZCQqg6OUm
yG2z+jc58k576Z9HZP3EIBgy7qNUNGhsTXeWQbrrNgd2U01CC0rYa/8WuOLTycfyy7qGysrKWLWL
mF3tlmm1l48xB00EQdI8HEQv5TxXdN8D79Wq2HZrOz3+ZBcJSZVNJsmBangcThBTKiYaxnRg+JG5
/u1IUh9Zm9lKb82wpslhVGCX+ml9tVVPxwYkJlN+n4jI+NLGtWZluuqoyhOCrElU2yy/t7pYXq79
Qgk3alXFfu94O9lxeLIH4PSgtfPsVpk6Ef6/pp60x+6SyY6R/cPuGG8ZnsAsu3oxltzfrqBtguVc
k+UQuR1t0Iy7ght5Nyahiu+rjcrO9hY0fs9+ljmj0d2/k4kB566LWvyE1jzkcQF543OLPEbKbYdg
kgBvuukH6Q0HhIsw5NMCAuya4ETTeMa6s50iNt2ewe8VSW+o9DdJ8GQ6vLTCKXPZiw5MYpxbHaj2
4YZCZRaJ0JsLv2S4ocvwgqWR0MwncjjPeogCbzgMuAN/MbFaUKu5ciuATZC0+xMNfdsEzWQM5QBV
ZKL57k9vY0cOARU7Rp6HWuQcJ/NdOTJCasb3pIEYiEceW36KUY+a0VqTZZ2fhY/6Fhc1lfUVrx9+
R0QDCfVWVS5Xw2/NuhIafYjTQECBL9Z5JIM5O8e98bkHbTMBlH7wIDY7ewbXBCPNeLheQc+KrEWp
n5SLGCLUGdcp+CyswyDkv6rQO08NcOXe+BtH2xvLV0dSwFz0TZVj2h3h+dfWYsnWAbxz/wfQf/8m
IssxK6ypsrIkpqW7Nqe1SUmX+hFdh65+CRuOWQ7arabZI/A/GAjiLQJgylQ6FDUjk4sFRFrKBGol
8QdmPYkg+GuJ1H4iHmbwwB9SWk24XCCpSdMAzyv4GM/4Q4tbSybXXh6UfEKDhi0THpSgJGUJD/yB
x8xzi3DOTD52SjF/cyHNMpTZ5dSY5PaA9bVzlvIYg2d6YeeSlQLbm8WjiTH/Cq0mqjySBQ4Tt+Sh
SHcvVWAXB02xH9yD9wCKlJs8aIUvyjPc7K+seEkJGw/lApZpTU2MBVKB9D/zNTla3IRIaQ6b9pD8
gwSFq6SOjmV5eZ8842UCSTYk0tebM+IvCEvdAwDeghJtfEgrqG3X7YoKF7gteW3AFpPonP2FUOew
Diugyl6GkAwgRlCLCChIvFgdrx1ze8IQx2hRR1rm2iVWjUmBIQ/SQmG3/VXGuSBz0irVPFGpolYR
VwQbeiCOQgJyEgJiT5z2Yu4v8nYFe2qqThTGVVxwJOiyo/2mbabAGJ0osqnaB7cSKqB7U8mbYiXW
mNrCL98Hp3C5XXNwwSefTcTKDl+U8vd718GhkFd3fn2AsbDNKscw7Ue3+lXvtHA1dvBERJlM+A6o
z841O2fq165ZSstQs+8aSTqIU2bh+ftKy71xX5CHugTgGWfEhB4S0mtbo+GaQQqXIKJTBVF7R8Yw
jWU5sFovlhO2FDjaosg+vgozVoS9aPx86hYsDAA7HheEt/vJGKRqyxh7bwC/jJ4DiuQr1TBGmOs4
bPjH2kYyNJI/Emv1GudIPyR5uSOf+WB1dtl5WkSzrxfyfMAzO9BZmQ6UqpyXh1fmZwKZuwf/y3fP
IdCD/4IQQGQyDAqvByiBrf9VEJYyaXNDp6RCi2O1TEdP3uBuWLnSZzscXz8Ria3vto81Sj0Q9oQG
zC2FR6u+BiJSXlCMFZwRtseOPZ9QN0B2e+wOra2qYxoeUozyQ0K3YoPKgAiU6/aZ2gKj08WvAgZV
UYufgaiJ23kvD8w/xVHZphweoiV+R5GqyWL2zQz75u71qGY1xWWm0aX7KBojLNsS8iP3kbNTJNXt
yaeTgj9DUOaxLPBchoMV4GSdW0PPsyzjRTLBxGYtnl7MEMEdUq+EAx5PkAtMdH2z2AvBcnJ6UkYb
68nE9wyyTpZ4wkubn6FIgjN6sOQvIAvgkj9YM0RcaOinnvonc7hD/omVnY7Yo7EFhtrjxK50dVpZ
NXQCrx5p2Z3+gExx1VsSjc8oH/hg2zZ3yloE+XYsLg9UCm09L/yju1v4aVUzsIovttvwBoV6JZdx
uaCJkzQsCqb+axm9i2sIbpk5bVuSoGCGlBUmWMpz0/ZKt1QYSWDqVK/8LQ4MXy2cdsgi25ibPmD0
8cVPkSoODZ6phJT+VCKMWmWI6PkwURrLDWTchvlkmavUBBtA7L2imIDBo2ZDXPrhxJXs46F4SbSP
Ho8PlEREIT3pBcCE6TRnDrq8qd+R886S+wlQ5AMutvrOkCdrIzQLsAR4CbiBPdK5wtivBpu7MGJ/
YFZBRoDanJWSH4TDiw8itV/QlZeTUE6kCGIL/pa1kb1Wn/tnhRpteJnbNqKnDNjfZpw2nU4agY5R
coM0jQAbVuIEfmA0Rm+jLQ7635KTzkqe+jgR3zUFyOHPXGT0uDdeimIHw7D1lQREDXxU4MWU0q/i
fqP4A+34y9TQoBH7c3ZMKF/3myoajPOszGQjDcGe3LEWiuV2EWNusS28eefNA7yfuK/i/80edBKa
va4kgbe8TIsF0NXdYSlUWnJVdmaGoMwk+YBffWr/3FzyerfAGNCQtpkdGDkTZGiXmr0bVJDr7j/P
fflmbtwcJlP15e2wcYEFGTpwNMEBo8+HpEVtrYB98RDcbf/BvmjGnSHLFw7L1k1u7S14EPvT592M
P/rGEaZl0SgiSuc8JHcPIoIFz+o4wOuYKXtRZvGh1PEwf3BU73bEcP9iREEVUjuu536zlg81T+S3
vdgIBcF6lrdrW6SIiCSHKji+S9MoJwgAQP/+j8Cr5vGSEnATiG3AfJl08Fk+3dYaOK61AjWoWvkM
kRj6utSBDYPb9HWGoQCymDhkJQhin4WCULwpmlglez5QQMmr/WS29uIL+k0szGaj4q9STnSQvMbh
hgri+aXxUcg9eRW+pgcqDC0fX0hNr2isQxZCAiwl+rAEb24Ztg8RpwMiwAUxsJq5qryZRy0gzwZu
tz5gCn5g/lGi8DsamsS1b8UGoclw4BAXuRLYfwrpCEPpMMBNQ2K8dGU3VCl+oJf1LJCNQzgzD+aW
oT1r8HAybc7ik/G+P/Bm5pJ5ekJMBEctvuoKhW9OjDdSrf/0vfePv2/qBa/Ujzluf1G4GyXdBK9f
Cd4FD5PsVEo4ZFuRjswQMf/iEBSxEZ0x8bqOJmaSm1SDtAGcCE4o5i3ohR1EC51WXJGpd2OZQHGS
XetUwU7ZAaXlA5HY6LP8vu0iralzo6QSmVLWbVGNHCoqTYlDbVvoFS6bnCURQa0WBghaRezXH8hd
bXAbTRssSkDjguaUrnAwr5bHBkkA/jTYdO5HJA/QG77iPXirWvUCepNHf4VqeQLuFHhd8WPxnaCp
NbftHD599KLM6Vm6oTL++xqW5nIjDGCw/MfvhlnP3XweD9nnEutfjQ/8MfTdbmEKOOV29aajadyB
c8kEWh8qfQw/n+xJ6HSclYpuLZ97QoBkR/LBliZctwYnJ/QWX7PG3kchWqiWT90HUySoi8FWQzyC
jRAvqNlud1s3KC46iTuEpWhMXtcnkGPE0pubjiyrJZUCiIX+2uLC4xeu1GC6nW174/RfimYWS27w
zzy+C6kQ/1It+Pv84OXJzywbypC/qkBaSK2Ce3auLZ3BueGPXlnG6XtckXgEUvX4phpDobBC857q
OWTH+7jHzgw7SHb3iK20MUsn5mJhlCqCzwNRB2GNNNWTWZfjrYyp602nVJSXi0qZ1hKm5YSKRsLx
yEAi25EDJ9XddoiG3bFBV1Wym6oxByyWBRHbf9ILRfiWUSXZYveTUordB5QKQywYyoZwFMFhqGap
qsdSMHmX5lZYZB8hWZsr5WRpM2TrRZmaWNh+FSjlihG0K93oN4yIx9Tu7oqVC/WF3AGsW2V74KwU
R8/7jcPYQVo61I6NqPcLGWqpv9tbT/hKLfBHSZv+BYfk/2I621HwWlkDKbLPoN/kwUuKGLIKxvlG
6kQ3DRRNibZn/Z2woa1qCxZf64duCzyyHE+6sIpeutdsTXfWKcKNaNnXlXtMzSSjT8RfYIqg3oCl
2uQQ/DO9d55WzQVAKefjZskN0l7lfLshC+ucNpZy9XdiKEOw7JTDzCPk2ZM5ZRzeDeOFiCoe0v9L
o8fSIVckJAkOOoUNoyBOiGeZ5chkMigde+RU0Uu8ECgssuQziEbGm7j6Jh/Kn/fQOyrqzKn1/1BY
pDlf76gAEVpLE+2MXDmFjVFXnB2vB5iL/+nB05UgKrYPbvun5TeaaPi3MCiq5KtVZvfj5D5JmM3r
kNIvBrBVWfJDvGl9xw+B0duARm9We1+V+IQBznsKlCWkD2z4HDaX/BmSwx6jkPaFMY0aIJV3yOH+
FlDshUPwATlO6q/RtKLAaSUPcgncrEiFyLJMlwpj18rs17MclqjsIrOnbMC/NleRWqkKaEGN1ARU
bkFJ18eR2DGeVQPzTDtBGF2DiPCdygZQ1P72CWf/AkB6cz0cpocIt8jeCIKk1/NmlBsWZ1/UejYC
LBAHjDTTP4YxKj1sNWEK++XsaGLp/YtQBtzrlYtgTg3DBy8O3JpwHvcxO5NXK6mgvp3rhwj3Rw0N
qGkeGT2+BPi74PxApIkEFvqeJkjbWV5+adqvtOOvYiQBT+LhCOK34qjLc3KQ6dkqUa/Xbv3tDISb
8TjCFsWRr5A1PddSfNfMNBaG8w3BZLJOcacy/6reKZuy2sc+YPNKEcSrz/aqgUtXhTL/yn1QDR0e
bUvpjh38h5OFL5XSnLfsIaoVkAeZNBhFq2WQI7hKijQVbk/Wneyn09Vb2nn/qx1IAmSQDc0j3731
3NVaPeiT9WVVXAxD86W5+d9uZDPW89OceUEEHcxsKNBWym89+ZxxVfjguSsVh2lNLusthc2TzETo
xCg798QTyhdfZiBNHzYKirnByDqzrxpt9BkP70gnfMT+uZG1nIKMTaTe34+3TOAFwlgiOBaknblX
0Bxdwmz40+ziXl5oo2cb3eZm5lgrFsOa2bp86J5CFXQpyE0mwtBnpPmlBPcWpIyIMQDhl+myYgN4
J7Krdq/kY2A9KQTJuvXxg2QcXAd9scMv1143wIEiyreISYxdZENknIwWtMizTTh5Xt/a5GJbZK+y
2eWuGrrwBIKzDKqOA387nJblcXF5qQXNc6LccT2VZ9xHB5FL0tJHIIXua3qcdXxteU6uBbz9H70o
AN1ZKzKGqMT29hNnCn5zs9Jle93tMNqn1EcDFJdYydgZU8CqUXsoPDNjGywt6SD1ndCGLa6X1Ycc
bL1AoHt3PsW3k865ufnAYzc8kJV1rzB7K2506R31hXoO0TpfJJJ8lutHqMb+QwRZwU5xEoKKJG6G
tTlCIC3Tp2ZQQrkJWRB0qirpHG4J235bi1PLa+izT/iB13LOGW5GdsAXryVl338DXh1Dg0+KxGFl
ATm9hAxEE/5mJUo7/hKd0rbuFOV4U4RjwFAmWgVzy4uUZ6q5pSsJ9q9TttykMMjaLPQjY4fvg8Fu
NIC6kMHDObu2UxpjiEe3OTR0jGk6hJgD+zjxgCPGBRh9fLagsMhnTQ4wFZiCvX7bJP6pAGqV54jm
MIrVzzOHysiVzgHoqXAR+qr0It3qdOwibrx3FILH3THYLLNDRcntrQpcYV6XfCdEHbsfLucx/6S+
5xaCofbPa1EtVMbMf2tQpyGRq7BNrTHjnLwJzt5NTlmnII+rU4P1OG/j7iQWfmLI6pkCTjx0OCPT
dj3YpWnrFb7H1Y4EGGb8rAakaH0Vyyog6o/0k6OmYCLf2IBTu0CisGnf+D17MJdi7B9tGzbyifMl
e0E7HVMkL+JNqQVR0QzK27IhI/tc8yVlOG/MiwmOSIMKYqBi3Ap3xR08XSy1xL3XSQbombkaLJQZ
oFIpKXJOysy7qMkZL1UrvZ4exR9MY/lPKk6OELduHelJZIcfbjN2WgEgC0ImgvNGQHEn+f9KHzhT
4bkJjeLlk7ND+SD2rWCUadrKXrtXpcs/WTZ0TdmjNNcbPzjLxDGaXN9Elfc5TV1vU3E8yd6L5EUh
vcMDFfP7b1W4zkLX93IWboMlpThUUHrW2xYkJ9AR0G2+h0B/OesLQJ3mat67ZmdGNnxo/Psl5OzC
d7JLXSST8bzI56ooDdXRKWnSBlGGsgljCwmgOt0CedOu1jS8nwzrQ2SXsaa5ia+1cfWQ8nQ5geRI
90YPU8sYscPSv5HOwXAty6f7vcPob0zVyc+9PBUxaCFtjew/iDkJFSCYp1Xe/UAggBkgTtWO5hMQ
9Uvyz0ei9nSmLAXADUuwrjTxQXGm3PnZC7fVFGs3KCs0f9gua/tEG+YRgGGHU4Cza5UddrkEnGx5
ajYosAcPMnkD53aMzbV9OUbBtJp+jZqKvfQbkz3hPbt2aJWc4gFemEhXmLIYCLM/TpRWF5J2ywhN
aRgoteUsnZzNW8X+Fg6GcQN3o39Rg8bDXDVIAJOP4uBVNMvf68AwjLM7goJh4/pQxbc/AHWfKnnv
QfUoA4h6EX0cvHVzkIUzvvCe5lSYBPM84cr0bgy4tNMrJT78UBrBp4sqp84ghFWiAD8HqFtTCEQD
X7QCe5Cb3Rug6BzaRl1gdFU5rYEIcy+wrLyzt9c/huqiLN5c6xmnL94o09Czvc7b7tR46PJmm5fM
0RIoMiRRZsMJ3iydZqjjMFCiIyqhP/OCxAgpIwBrDW9GhCESbgT4c2G6s10I+qZMQq9j1G9ilRMK
jmGTly5OGmk0dhpyoSPxMrDySMqb4c9oN6PvfAcF2Xmq8xY00OsleNInfwkxVnwZ41PNkS5gYQ8w
SU5WmjexdGG9yFuBhhYVLcj5c8heVY7pLwfAMHhC3JxQTzPfyIiI/dlS78Nu3Mz7m9P3Uc8hXO0P
uDyKP/X4efkkikhpXbof/1xNeosB4HtUkul0ShhkI8xg1ws6ObZ8jkzMsG/4Z7YyIdFk60YneD7H
liXDQypjAHPfmIBAPWoOprq3XaZlswA9Rx3PQlzUniN5FM/MPMzAiuHJAOGnIlMN/paoGqObjrkB
wMq8UV1rrAUrOlFgwut5mNUcjnNyXcZNRY9rpllYs1k8AULLW5gZqnRcQdaTP/0jERRlbr7igfh0
PPiPWkfDJz3QrkLwtS9C0o4rEgAkwAzj3ZRFmq+yRLDwj+cp/VEzMPcgQCN1b+ab8SFJCqqD/k1d
hoEFOcx6eSPNIyTgTIh+S4goHl/S8AKRb7e6oe9IpMe8P+6/jlKLQFwCXfzaCZ93sz4By7ESSX/Y
0D1euODaY6/Ig0AR57sCjhtcp1aI3jFU06xbYBueCT+RqtTSXCs4J1kT1IVpME4DaUUvDYzM0ygR
o+Nj35QSs9hML2y/YaekfB1XcAE2tiP06wQE0WNzAlZ0fhKDlCWS9sQnzvyPn3yTCZw+EnRKote8
7n+QTvOOQuVQh+LvnIbMFmmJjxePJrQ1NBb9iV0B3QcyW5tTcdDNGjfkZsWNtBnSS+gOiibt6Q7+
39xW6eVApSrRlo4KPj4uYkXud8LDZ5szN3t5IHuBd+MEB1Hv6jJUTOhAB+zS+1zSua3ZzEN8424Z
EshBkpLI7zMoOeLbm7hCfZKaYiUw7rFUI7EfXn0n7ipYY4q15Sg7UOnMsSBCwLjBn7lXViO5dG6l
Oyjanw3MQsSCVeVBVBWwlerGpsoflxLr0ZBW/tsFz73wgqmKwpvSfRC9qBI1C3jf40Aewt6DR5b6
Q/1ElBIhVnhHE80j9O575dhhQdXZ5j+1L+MZ933ZsWNOlO6nx45dNPCFGNmGv2IwZi9vXQLfUU1I
bSexPRq1hQIO5jMI3+rvpHhpYxfD+vD8MzfvUGy1OtcgA4OAqWRpCiawBF/srSTuxOVhTsQyZ4UY
sZFS7iJ1YIg16CK5i6ak3e4ZAWCLLUS5Q4tIUDRFwgSbDjApU+QfcN0wIwtq67Q3+mO5ybwG0Hzz
SxaDvSjuWZQ6yHeMv4nHsackp8Dgw59JIO38393R9q2q5nk9YamofJ7zGblnb9OGqBtXFycWRq3w
wLE1w7yPKqYnk3GBj6AXf1Lm2kS0gYPrCOjc6GEC8gLM2fd+usHiDyN5EU2n+FQs9UNwCg0EVPP2
+9NsgGlFqfGXlAmcFXYAUtw0O57W1k5NSNlJ6IbawoHhOWCW/O6Ev220t9OFP8pEsr2e0njn2wxn
1HT7PeSrJH47UXXkH66b+UHUctRbPFg7xvSHF5RHP94ePlfdcs7fKT8eowxBYEIJblXApjTp5jj7
GnpzV3h1hZADKA4+k91GczImfDaJV+cSUZXwlA9jAVxSwo9XbhOyqdGo4efKo17jROm9GuXku195
0uBq2qOcyWq9n0krdlymiD3RkpOy9PQXCDOgrv/yT9Fdt1XHvuGi1HZRmYrKkpHBtB9izksvK3+e
rIwNWcufcnLwJ/hiUBOnLTrsXbrLH9i5bDxdc7uWV9T+3JRmiM9tqvKoshXVuh0deDJCL7xqxU8Z
WEivjtzGbiuL5feuUFfpu77HXQ5IeAqo8saiM81pDZWsNyYlkew5S+kRMG0rHIrA+oOXeXLTIQzQ
0yq0RBS3dMdlUHpUXcKjG76LBbGON7DHpWNeL6eUq2PAO+8D07tr6ep5YwhWUk07vfr+65DkIpRO
GbmyAfSK2LiVvVGzuFN5CUo3ud268EfX87A2WtOpyMLmcdEJ9LLeIKaQbyZ8/LdQLjCFZuPomOyS
XeQP8Ew2WRYWwBw5M09uJilUrd6EEqrINN+LlFUj3Myrt1Pcf/1Rd/gwg18k5XYNdGQI3iQRWt2n
V8vUqrWLSCtHZmzBKeMMmLY5LlLWKpkKeGrxChSnvfzPFnSjRMXSH8xwmBGL9o5sHR3xqojOK++O
No024TKh0iM6NxCGgOLuAGC91A7k8b5nxLqlzFFYNbqcUfI1UEwh68NFtgNPzQEPbdRCXJ3rMWQg
/6oqa6bJHkUg6BccAMB6I8yk6M+BxilaWDQFtGxjKzGaB/EeN8yr8Y8H3J8acaKf8TX75SNIvmLA
qpmUhdSmJpDhNPXLxRksUeqdoSbcCnn8KlJDlHdb3E1vh+9QqoN4Opx1i51ivecRN7VnGdGGNyeA
yf5OO4Z8fxgXrjjLaNLY5FAvV3AAZIcyu4+EuSat3ASMYqWLT1kNJZkG5yhHEo3M8wWoOMrqBaSP
q83cBtIRsKJifcHavp0ExALs/SOtwjUNwtl/lA7CfWWSSm65vNkHuXPwOfukTVPUVIy0bBpas0HN
NVkkckn3aRp80vQfCON+/iKHb/7ch4vDaPAdYHvNGTDweDSUYSJoQuJ3QH65+r2GPeb0Qih2b0dZ
1Lk19MxZeUZFG4c6CvPDOaa1NixBF8nfAIEAjn565V9/6C8C6NlM3vKhwENsMy0aVMm7AP/Fs+ed
lIWCAcqFIuVSJM8oHAO71whu2R87x6ABX6o1SNV1qKRNRy/x1FL0m+CrpIq8/NVAaTsFlexEq67d
dzYKWVg0jdL5Xlf2msReME3Qbl5R1MyxuPJlORARdMbYj8mtsbYnbZ5KSJE0CgsaDh8WHWdrS+zL
pYRB2nGBuK3YPEwIJYcHTZEjvgaJtvASO+hkurlmq5J8ObCeLaIn6CyIFgr6V5kWz3JFwIrHpkoF
SBQafvhf7Eb2uHfhe0gcdyaHlVXK6UXyjm7djkDchOGLLZ2UeU9KgqTDDSzFjn7HuQeQzvBY+Z3R
xOTjrsphcshbpJ4U2vWV0y002sjf3yodhZf2Y3pKQunpP8DZ9PgUTsE+jv/zylKPZCXnPQOn15YU
izf6z1IphJNFccaw6cauaLDIh8F5e7pM1Qx9ksWeSrp9OZyX7W/p2s1zQCpkd74CNN7qSoZN5ywP
F6UtRFkqlN4RCbqmKTL3FjLax8vGiAA+EK6HgFkCMRN78NofznqeUrL/8C/HLQYkGuFpgVdcno70
zi5O1X3dKAjLn5uw5WiKY7UKYRprbvMwCk7gWM9QahHs60QeMlKc2ON75af1FtxamyVqKF2vv80N
phpzogSm9sAc2Op8aYIX9vnUVF2NTBzSdHzLcrG/5pCkRcKROTuEpDPx61+/0M4XNcWOUchLc0KV
Zg6o873/Lk/yQQe0a8Bt316cZVm/U6Npc4lxJMES3Zs08ydE6sgawNBk1Zd2JawgKt0FVf8QeB1F
8+1oVJVrvCKIMcgg5V9+45I5eh+xxSGpfnZGXsEMZtZchjy5h5lKdFqF5QUDE/eTN4JY6RGBQQps
nf828cuYpG/pFJTQbMT5e+28l8RM7V2DCBHcwZJedIwq7trIG0LWk9fIx5XuhEYNC2NbItx5GbUT
6iUhn+lxm7EnYoQ9o3PYQmvmMNYUrF4Keg0LTyIoEuM6B/TNw6HJ0TX4HAF7sK72BNDx+QNFV2ZG
L2OdKolvpQKkIGYhcW+McNHv0Si+9nZcFIOt7fB8Xs1OXPWWicG9zOFwH8fktLHv/ENJRQG8mcn/
JEUtz/aX2Q4HRay7+TyYLMGYQTFOuHGQDBnSbfUsNjCMQ2b9M+2Oq6d5tzrBPSNQOgnxLr2R217g
9IVcPml5LnbNXFqhQYn2dl8k534WK2KV6hUCgPAB1yytikGNKwE+jAkVZSyfhB7viSWpiZ2gGlN9
ZmMHBGdBuBnOF+HpPwFrXJ+dC/OEHIPztoibQJ3P1x5bTz6tKtmBAbpUeiFkaCYxZj05zMDIPXWc
oG/bgOBDxcHENd5lzy09+UB+nYxSXbhulnbBjq4/xC/jYA1Sb1MZJSkL7TnYip2xJ59vOsJDqtUv
ZnE7ipoRZYCXM0hP45DYRsnCLTMVwZU+eCkoB8OB0Bh2mqwBt6nqE37YT1P3P2JxXMCe4cgD4kmF
R6BSuM24VryYyEb+/orKU7TPhkxnb7fvYE22m6Na17lSv83be2DDUnVv51y0JPswTUZoEPEkyu2I
qH7iyFBO1p9+CREexFjtMXtQoV15PlNCy3H0o30UgKySLpT9KyGpzmaCZPbjZpZCTT8tbNUxvAqr
FOPaetqrsNc9x6cfURmF4TS93jiL0nYfjNtPlpVEfAXO02HFHfTu2FBTRRKbKYg/jbigZoxf/rSC
zlhoeLQejIHdGvr4j6xTnES3FU8nuJdOs57MFW3qBntsh/2TuPFgpzLDM/hJekLe7TIrzi1usuxz
0fQojumuxpGZ8ijA4Y62/07LUaCg62FBwpCpjgpEXaVpULDPO45V8KT+SKRb3CR/JozdjG4EsRqJ
MQiA1WumaMDxtlvruf8hTIsZyq/+bzjq1AZWMaFqxWZebx6Gto2HrmEY1gsIoqknDMSUZgvVIxgS
xvDly9kSZ8bAYxW8kgzpap3CI/a03bTo3uqNx0+K1vrDraaQZR1xnFokep8Er2ceygjalp8rmmNE
JisoMI7ZUeo014NuNWkTmByavARjVxONi5iL8mgVrT3174Ak3WrQS4LspJaoE+8l5t6LuC2dUbqA
5G8aeSliDtdOl4GJtufJhKbRKJ8tycxVrV7VFFBvsdqlzOo6u3fRksBYBo7YgVvmuLYIcgQvQrtM
lVJdiN29IgDRj6rAT2mOcnt/WLRp7w5yuxZQ1TSkd/OgTlBrP/VGy9zFgJZUGHGGKCbzAdMMgmnK
e0t9Kp8ZK1hAbXqm3xzifnXWUTZGYRS7uexG50lfpJDDUe9poqyxqDJcHmVmLbGo4S60zIyHBlDI
rtL7dgp6oL0eE0JD30iz5fO3RWeolF+da4tQG0w7SFkAtqSqyqQyEP/Q4qw5RCd0Iffbiw9f1yrh
27TdTsQi0PNeCRI0GSkqpFsEDw6aHkeJseqpoytsV7hHxbsDOdyAkHEf543aeTuF12crvYP1rDcO
uQO2TkMXouN4ErA0dvwNfow9uZZ6weVUfXSeyokLczZ5GwTw1XrhR+BgzbMy6KeL0TksC4VbhuKK
jt3i9Vu1hMEFhvaxDGZOpzqTmfy9j49V2v2g8fx1+2qvD7zcg4t0iOnFw9/cZkNJTLQiauKJKnSt
n56pq9hkTTjyOPQVx3q0Un+ZorhMG2SoqKUKp+wtHUs5taV8WCChkyy+D0BptElBDhPLJy184zrC
SiMKGvUp7IIg8/zqSqfFZdFngnJA74BC+BOXAxJD2o0StoyUxHM5F6rMoW2+lM4NpaNpg1u+wFDZ
j75JVIHZomA5nqeB8KZgymFOe9iUh/eNFnQWfoQmEy1fXYqmZwxif/3hQVyHenFGpE7qy0lEeKg1
IbqLw50Kq0k5/79Xwz7GzIWwUiKB+1Kr+p/A2/CwhyX6urD5gszX6DegG8pKW/KkgzY3yF9rEdYO
CCYCIfrJ/stUYKLNvYqFsPMXDPRurfJlgiLrdCtkav9227CWjs7CD/WgUfcCuPblrgpG18Q304Rz
zpPGMQYCxAK1/92YVVI5KW23pIJQaYG8clrLH3Slruhcstaifw9t65F4CbU0SRDPM7ZSbXNj+wKg
p6Gb5uR+wFqFzelhb7HRVPLK1Rq9eXbC/oNeK63Soe2Um/JHF+Ukz6b+x53u37bNZAiSJ982LfWg
d2TxxFJqwlchSZ2ea+HAJVzOYSmuS90tuOMCTZtRXbdZENarz9qiv4dDvHePMm1FthJKTOPbcsl1
5fyQDMIIMc2my400cv+LBsQuME1bM14OlJWnqqsotnSWgrgj9DmlQV24LdBEaahz5afQ1aL2Y6BF
eKnLvSDP4rs/dETOUtDCmoGAg/9ztbgnsFXdq/vv8SPg/9GW2PrR2+m/1uK/yAJt4vXdjhFUFO+s
Drzogx+KiYiN3GHWWTISM9yl3ZPhD8o1h5OKoLpF2ZqYixCnUuHusJ++kg0dLU6TAkcJ6Zen4crm
vyYrnYWbqk1G9ULV/0hVlqToaAPTjxKnhtlafR/0+hoGzrWrxZcoCRgP8iLJ6AGtWhvu/2+5XrHo
RZh8LvnBYVJWNc5+K8uqswjQsebUW9SJ0oVgd6Xam6P+/GWp7Hvvyb4KejEpvX8iZLl9U9r+aikp
xaOeb4VHomXbmtvWB3iX50z9tSucFhsd8JQBrYf6AYZVj9yWrHnqYgahapoZCYRSzTVokkGSmCbl
0c8HF9VZAXnrt+ULr5TeZA6/a7KDDcM8pF00okoSUWqNPEx0Ak53CABoeZdI0BKQ80FYr+QYa3/7
X2Ai0lb5dpxJFC6FVDKEIVVgkDgvShRiimAYCgNqTIfWZpIuntMC5qaaZg4HzSdBIbK0zFZNOhun
XmYVOyXqitix3DKYK3kYTa0gFNmmRRsxeoaRZUqbUZaRbtQx96VU6TsNIjMoZGcAC9i/dlu/Kypg
x+ok9rC6CFAIh2/M8AA3zRh96nKbVUw2v92FQIqbSeUH4eqD25w5zPQpn0aXWvh7fWRdIuug/6zk
rNl81jKDzJ0ebq6hXT+oAfQZ84dfKjzl/L2FVet1h9wCaZ0XZu75AgJI9lyYwUhYw8GBqutz6YjA
oTYa0azx2gJ0pNo8eZy8Z1jyVSPfKiVWoT8DVPHPa9ZdXq/A8RNlgzmP0xZcdzmnsVPQdxJtM5z1
j27zlsfytAR6gDpNXTb5n7HGaisHZz6YdsPvmQ29LcQFRCM3YrrCzd/llE1Ac81pt4GHxqwMdMrk
U85zQFxKUJzP6GE+++LKf3ZUCxur6eyYhsNU/z2lIcna+0jBm+J7Ic84TBYZSNnJn8f9zS5Z4G6w
MIs+ZWcmiDJm/V9m9NHjeyaUjLKZUgXi2sZ+NqvqUIrzuBXeMEE+N219Tv8uOXfPYt+v9GhhpuRo
Ulfe/W5/Wo2fw+kfRGfxP/vzjscrniRvuGOTvGXewvNCDUKSgUGaHswqC2hHORCRK84x9fqhezjO
MoRqNsN0ca8DZmrELuDO8xeCy/RwQ5LExkSL/qO8p5bH56ek/xxbvXuIeu7pyLwzxXqv7NuyCavv
KhUuBIM/p6ORPukSLaNKBdFXC/JfUYsie+RUDZu9fhq4kX8pK+Wgg2mTOF5iREC4axA12r6ju3E5
SfMgsO86j6rKIOKqby1/QPj1dAiyBqJFtzWGLy+xIqlEhg6qWRzg18EyPdsUofAfUwhZbcGzOp2F
gNr/MzE4kQfjW0HGU4LwyEmGSPi/l4+IvheOnpBnLST3IWoALFUHa0INeCKzwuTk4Mc7qfnYOFVj
FcV09v8ze5aGnYANHloPxJDjER0HwopLi8SL2zjraAlC0xKYNWBtsqNhYv35uL/I0Mv9WPfr4r05
HNg7XlfOZdCt2/Ogvnbqw1kh0aaVD91Aab0SjKnxW0TK9unAZmcI1/L3yA64i0kUUKFKB66TLYAu
AtOWQtfM0WhzScBHETQLMKIGCXyHlH9iNz8Z7Uf6yHHMunuxStUrscSiA2aT9w0qqADPO4zSNSyt
1HA4tPGGXxruiaaVqLWWJsmghcASkK7byAYSaTFY2F5MZ1cv9hBeOJsWqvAxbX+04p4KdFxf0qVD
40HN+03+dPSI9VqEe0HJtlYY/JOIdmnahxVc1qVtDIJ9wKX7HmHcboTisllGQnnfJo5/6SbrymV9
lVkbq5AjntrNON6LQRvpMejwnCGWe0e6fkaLqC7yCcqVV47lWRA0e7Wpe8BWvM29OgFRlCD9Wk0B
ztyMwu9e36/1uQ5VfTqvjGDwnPpJlrSwjnDXL4Cmob604VJ7kd/0UaN4bq+CKCs+nP9oiUQGpc3k
qAqCWlTdKY82FTGChkwuFVCxzlABmKC4vANhBjqt+CiYm4iOxriMHkGNyuFUkJfXdjOFkiWlpIXX
LxFeLvXKnriYLc60+I9BPlj8ox8r03qCrumEFcy4jl9YYDjZVYtWES3y/Sqx9CB9AaNifcxFCw4A
KM4n2oZGq8SRxIjVKR7h5M3W07k9AShUo9oevC75eZoIEx5vSB/oDJOzf57/y6j952FL/I47C/Vn
tAqMhzYnt5ECyG1aYwpstk7zEEIQclQF34EQwRJWaFz+7rrS9QSAV0pRoFxrUFii4G3hgyKDxRzi
bqp8LGC8qM1D1/ZhWMAqOSrbR6YKFxYZ8alyovYqE6EXBjfNzS38FWsj0TA4TO9ggTI1SS6yuhoe
3X7ylUYduva9aXijBXXjb3qTrd95HodI6yp/5kQLlABvXZp8Iq+w0/8KqqaKHzPtmwTyXYV2I5d1
JPL5HLhFLb5oLpUXEQo0Z3t3WBywUqg+bvP1FvknbaHa4II4pUg+q0bY4EMjF/lHIKOjUs+x83y1
Sac0k0rZ7/yWG/6fONUgNZFYexg/aCsP9zJvk1Cs3p/oudnvM3c0sf8hYYxCI/AY3LywG8H9qVaF
CDiDhOXIr+SzWv6tpa6LCW2pyrtCW3I+iXBv7HDs1txWQRC0wFAMvLBE/9atfv6y2zgSkCgxF1g/
MhonMuak26D2bCjFxJAUX6gtDTB6HJJ8Jm7Xczyh/wOIZvD9TtT7hnfO20qWxnUmInULGLqiuqEf
csQJIqCBeozspBoSXnZ9N5OcKRIQ5fq+ZdU0U4yeEgyZpXQwcO0+QusBtg7F9QZgdciHv8iGnyvp
XvDxPr1Nwf3oEK/JomR+0hvTjMQMY8vrNbaFOwbGboI+SHwcrbGJ2+aD00HB5cVKlcuwvrOBsx2a
aTJebYYDUF4rffOSVwPPQ07GcLFHMoF7ncvEucK43mXM8rGJHqJNDGbwuVNl7WDzj7XeIc8/1TGg
UF+11/6Biupn4MrIHms6evgQfi+kRTWJH07G9OlIEGAR3xOH4tIFKIqyG7SoDxKEoYVe8YQ125Vu
IxtelgV5r55EGx2LOUKUNflTw7IEUYI3OmHBXoFPMum6GAN1Mn+nWE+NTekAeWm6nH/mWI6zZ3Gu
4udyTFrT6p+Bp6sx4c4J2QQusI9tjrROWyZea4H9Zxu1uZ1C+A8fOeUJQFPEn8jzq8ulTkaFY3u6
NaHB3e8o1hWmEL8JpJM/72tX/IFG3aKR9RmJ42XXhe7xr8OGprSJ6DQlRz7lvPR/uEzFIp0LJzGQ
3DipXaUkpHIkI5iW8JVUzfvLmV8z/ttsEBI28wAcLRn2gLeYPwjgD1oypUhi+RwlEUByRpYKqKFG
aYXBh6l9/T0un33c5kqKTKudM+XBgZLq8NSyi1g08gYjWLu7M7v3FOUYHa3C/T/6cts2I4TbucUq
52DYGBN4ai8iw7Z8/QGLkoDEIgXN7Um9lcrqwJIQWVjgAxLBqjbpRgD6ZpTKTQk8je0kOWLkp2Tx
vOe0YN0htUQiyMCbHW1UTjNUG7h+pdNmsstPWQI4tHdBe20Cwtb7MyNcBIhPQp+tDg5WwjG4m5N1
VACR0xwx2p5kKdhXcbNE2IeJNpcgew9F4Dbi3jStHMBTLIarBgTUro6o5YNRkm0nln+V3EdG0AHW
FjDTI1FbcQOnepkEBavdSOgnr7AChRriPXzddFJgBVTACiLf7rbtYa68OJli9Qrhk8Abor9r7J5o
9OhgXeuoqUP9+jGGgkCPKsKAirMj27MRb0YGH3hO2v8gwhATfK9HYn7/kAkJDGkXHKr20PmsFLVx
CxVNW2l6ENLgM1zmZoxXHBzA2xng3qbZ6Y4Q70DMqgwW6gM0QM6Cu5UueWk4TWk/VL8NIRDmz79K
wVhQmN/yt0SBfvRqBcKi3uV/neoT4yzIc9UkGeqFgu0wfL14ZqOQ1/YM05UUhiH3ypbvYIYxzwWC
2NGABzmr3k5fp7yxSfq4eASyDL1PePjxRQuNs6QAguZ2rCSybmIygevUOSz/ZkoxUmZ2M2imrcLa
pwDOXdhOr+u24GhUE7D1FBGCqAVvAZqVX5Mhf1+Hdm4NtqLD18eSIiLgYJXo65MvQxRvhY182D73
Smyx58FcFy4hegiYxOIl+9z/UrveScSNLYtGcUtTpkJj/yiyxCO76wMPDTQDwBaVMUtGQsQPdoQ2
GgVNI5mZZvPKV4P6HZuLc+geklFs3cgOJGhOtPugpuadVaFten43ySZJYXUL+lEq9cfF7Igv3aWT
vPPffau1LM515xB8l1+QxwuafqmwUj93jB+wjpT1GwyrkBTSTD6ZIAHG5nvEG45rgCvthDt71+Q/
bZWn4z/5O6xczeX9rg9H5FwpCgd9v6Tm+YtHBqgcUTN4a5gXEn8D0i9qQ2swwbtkuD/9Dh0jiHZ4
hcesPDLVlhtXKNthblf+Ino3tpxNukGJSXvtToqfYzjkh2h/x/5Woff5vhBDlqqw8cGeBT+RFurY
DW/sQMbkNwMMEAfc+16oBu2J4Pb6nL3NAct3ARWvPNoH8y1NYGYqdvwZQrqpB+aY6Ts5Kr2mEtmT
SNuL0WWcpZcWUWFLIjaBQiCB/tJKlwUidOyCB6tRkLuLwkKtEK//6bgw2P/hWjPS0Cj27Vfhmm4W
q4Kt6rWLJcRNkCiDgx9SqerJHkKUqafO/U6xgHG3uKBCWh5wjiWc7HmwgVUAKHE65OSrywWzzbz+
55Z7SIfE7DxmtZfVDsImSaXC/IKInQaKR8Mril6KVM6SLk2t1wtfoqUCEN8R4NRKNdTNHQLRbTkt
nkrjzXX6IPTPvovGIrqxfXhKUXX2Ci7ytq6252tqA7WHe3ywmD1RivCmfqPlmLeKmnpftVWZeqRh
eou0VpUbjvUAnkxpya0BskM06kkItJPSLMnAMMCXd4Eemw29Qoy2SwrnApH27B/HIwQknm9f8zR8
Sgls9/eu2oJYPwa5p3eqDeBEAAfnlTumvL3ut1+4hDRxvkoUZctw4lmbOuG83FE5Id6Prqv9hOJZ
+J4wWwBRLCoqUle84GmKNy8cFhZhTRI9pD3qG0vswJyDMfi+o6yhNLUVXQApyGGROiIGqJJOed/W
dXXKB+LN3j6mXgw11MVDCIwVREli9fJtPqK2O1rAM/aa5XvqHH25Ue8+iJBsTQGFnDecUF7qZGv1
lJHa5NjpfclIij3h30aK+L+jU/ByAQuBfoDn8kDIM6ZKviqOmE2feGAiY+TnK6pbZLgKGHcP+Nh3
j2B2utTqxTZ3YRu1c1s9wp1vCpt1L4DXw7P6PipSPARUoIHek3hU+/vig2ajS5HzR36mbGQKi/KE
i+ThViFFYr4e+n3OleuPh5zsGZTUDUk/+XFoNdt7aAvnu3gX0+PL6KG0KmNpxcMeZphJHOYsI8wV
MVhAo3Ytqvr+4K1SABPvEyB47GXIibMwKLTof0VxC9UxGphJw8k3Kzg6v67h4die1+mV9SOo/CNl
97Aff3aXKmR1yQHwcQtnnExfObxu+8fmSe6CKUlwy8t9hxa4pw8S8LsxmrC8GimXvDO3Jl2Wise/
4AJ+spVQ99HghnfLYqE9RrwT6kx1SQejJx9XHGvEVCXhHm+c5Fk+mZudXpSfRlkzxbko+Ga2DZzP
7IIFKNfLPpBzQ/TDDCZYvP1uFlRGVBPKm4DJw2KcO3kD8RFGevEajXVPDsfjJV2Mgq+f+hQnA2yw
sfunqmX+epE9+b7ekmJJEKAOR9SVfogBIc0XTiLdVRah+hYPDpKccd8RWPzOLLVpYca2f/ZTFDAz
VKqZ6upCGWMfoqF+Se1ZlvQuL1QLwHdbSYeKtcy3zSiUzTu0g1KUnLE+WdEpyyCoRYMNsYPu09e1
cIejfPK7itiKudtBtiVcRwJdgmL0G8kRi1Qurpv2K4P20RU6RNknl3aXIRh5anGCWbXpYH1+mFGZ
G5gEEPByfopLHtplRXWdVrRxxI4/hV7Kd+qb1FcZOOKJi92DaWgVEWOUmktSZG/ueGJPNwZTlBpB
7R0eHxmn72rDs6UfcoJeqDLA81zompA3sX3KgYofWWxtoGDdy77+yDmkY0qwy8BYu/m2a6QREcYM
SUPScqmZ9wdmJHtkLf+4mbR1v6czD/3wP7SXe5YR1GCMtCsKKWlqrZMpaW6e/UHr5RerhXIW474j
266Hq3OaxRbt4Pe9019EUd+4UkvFeNvAVi2OXVUCoTXgiJqym7HofHrWg3npRE1ZLNqUjEuvsopB
J1zXWieSG5eiRT+KtTOViUE1o/sYrjQ52kiqIx3F84f1GIcmSccp10Hg2uwhvQvBrw7c6munmPXi
YcTw+hOM/F1dUWSd3yj8rvGsTPXdzISVjCkJDKI4EXLw8qghoFpdn2nNVlf//EetXXHpYgK//Fo/
+AoEf2VLV96hwb7KVb2HNoaseqKKnkUThvD4lUstW+K+WstT1HyypYsklukNT0Xsb+ZXGWf5ecId
bmp3bym1jPlOGah+R8lAKA+Ve5X3t9y46JxxqnUmnwnLEMwNUAuFs3w+sq/igdfCVfjK691eO4XL
nP/GY6MSE4wHYTmokCnfZMiKZM8IEdJoR4OK1WWr7HHXkuip+tUKeguKVoxMRnmjKsZudI6Vg5S4
0Si8jnMnz7Zf/bn0S/R6HYZhxnqnG/PfO/V2eoATLrOcNcASjpltUbjjGmGMTF4fxVbZgE87Fszd
sjmjebd83ojVQPOfozJDlSz7uFTK/vN2pq+GJeOA8Mov3FbXNY2I6rv3MR3euBR+x04XrdYKNrQS
tW01rKYRon1n3/lYJf890hK9ZQ01HTX/muFteetSq0Kq/M/bBNkSOUTZ3p8K7ZVa8g+vjAbECXk2
ZnyrVfCo/7VTrkwd/a6B99KoIIBiNdGHJdY34NWhpbzJ4nBiEHmXFLCjpP9XxWd/ZyPzw9iP2PD8
75JUJFrx91w/QpuzRMckhWHmGtmjjjwxs+hcKDPA5a5Gp5NBHIKXfyjmBU2OYXYuJiLFidaV/xAm
yCMZqmJ+OYtfNZPHOzyCCgcBXTgZtaX0ECWy6UJsmOSuGmIR5CAs5N3iU7CtyfXJgzVvvWUKUGmW
fo6R4fQXYROvhLJkjvEyepd1H1Lb/DHNXXCflblHGSwLUI89rc9Dg8rncPUoSP/Ab8n5o00z4XUn
yYJGJQvqlKOLC7abS7mGf79xjgsK99I2xsAgLMq6fQSgrZ6Up6iBwNvUWy0FaJrxa00qOD596mG8
0BrBhBZgA5+Kup5miVkGoWPfhQxfSzep17lfLzxbAIj4bFAPiJql4FhB14AlJCtGQNdkCGT9BU9F
2R0v/PfW/EAeMO+ugoTgC+LV0hDnACv4BdxQ6cF0SfVsh8GpeqJVMCSAaEi78BUahCQJtA2K2s8P
rLn3MBwpGJiFPlJ7TpQy70s7sBKDakKQsMNZJ5pcb7nrzu5T4vGJIGeeLEye77bL+rZIcn7stJaA
cyONrth+BzxYQEHlEFNnuBv8Q9hsXQELgLb4IXdnraX59M4g2YcIKYsSiGyiyoek5QOSN16KzXQF
rPb1vZU9jO2S2XQ+6wJalOyBQ5K5F7B7TToBDo1cNJ1Xrndfb6SeJHoge8bwXl6OeHwd0Dc2xB5x
jeZrqZlMxrlHZDygJtvGD/fddJBLs0IzmVAsO9Ej3MbOxPzfTVPfer0I+9ApyJRmJXzSVRe39l/R
3Ym9LjC5vvlLJJtvKjgcr+i6OQ4mI+N70oudFQm7vl9nAMpBdZo8jQ7TtV82WBpLUMOhxObK2raD
KOz9I2M4nM4Pm0hYRt66lR86Zl3SBr7DUv/t/IEMMyTwLeFfO/n0b7Bgv/2wwgKilqJBiHzUBEv+
UEulNbOz2hVTHE65EINVfbdY9xXREbRjc01F0aVPtytnAt39Rlrgb6vedC2Zay4JykPrSYySrP7M
SaEpjjHKgpqRYWmj/oFEKUGFiLxbxyBlEXaiqyda3JqCzfYCuYQT5H8j3R0J7PksIySW2RCcCIk8
GOKMcbGfaK2cePwcIwUMn55p3Ikggj8HUEf6vngT7b8k0wlPL4bpTRaSuqAo4z4fDUxQlLbzJAN1
F/Fbdh/0tSsZpRUMYqnzSWY22HxtIpKGhffoR91nCbXDtTChg/iazbRBEA0+TVBNv/Jv/NDkbMRT
J7oyxvIKpbc6k0HkEPpaFmgdzl4gnJJRJiMdXBufCdISplyLC54OnSV4SEmSrez1JSLIMaOgGgyX
b6/TlQR8lbrojmONNJW8uhu5bMTGGkauAijwzWcakZGAGjKPfL9XpxiptbejtcatvlIHPdj4LFMz
iwYOH+RVeMJsSTt5vzznjlRg1JdTvfamNHwm6KAC/FPF8FsD5fgs/z3nptAyO3PHFHGODwGUh3Xd
C/bCnqRgQj7kRbstkl+fFXNPPggsTc1Ze16c1bdcCJxgP3e9mRs2hLbpDM+tcejNUk4jByoMTyMF
M9yxzVXmqrxaS3t8PGsYG554FG6hqkEsTco0XgovRZYx7Vl2ZRmyCnuROFlTc6nVqIAfTkCgvC7H
JEO/NFrdqqLfcPNfByekbKCnKWl6fXwAdKQ7DOZLJnO3c7sGGiosooMMFCJ/fnM7Z09zzQwGtlnx
FRwVWWNcn5rphsU8VEecnvAEb4+c0c4Uf6hFOOGIRiYK31RK4hqb6NDOgy6zDogRdcKpHtr3GVtA
iYpE+MjMffsno0qvVqOUiKnqpwE//zoUGdbus3nSJaccYoUJA5J65QLt3EgyEicvMz7JAxNXoM12
x0OSVe3TROn3XiRX1VokkN13cFAeW6+m//zBXwo1Snpw/ALFkVD++bVj2ulqz4kcw0vitaWzApz9
AQnf7Wl4yGJd9vxXgozGzJJN+Bi3+1hBIcgf5Rvv0Cv1CzeajwpdtSMODnMNBvqbAf5MqQNI4dYK
edu2637Rp7B/YtRZp39c5Kelp48l2iuqD35i7PabP3JA7uWwxYCyTmospcAta40ATIflJHr0Cx6B
Nh5kBt9XUVDQA8HqewQIppbQ5gdJPcfGyj/85IRv80MvkhBVqQdNu4PRbOQt3dQAqG290fyWSox/
0Mk8CRpDRyi1SXDfHQbvAjy+xxtEO0VidsTZoTo/lcY6xn6K2jAFDy9ZvcI6ICEJyOBvAN3ONt80
2fVEii18SKPY73isQ0ZG+U92L2mrncf5TCI4cP5G9BPmYjUxeac3a635E9weSIIvObDr2qnmjVs+
Q1ApcGAHU8+SW2NZv/fYxZAL2h9Wv/JUhZhYXsGVjt6bZYIx5IEbuWWb7C28mUakBBm6DpBYNRDs
fzOylQQ/fcmMyui1JOL20Rl7kOCs0NAeEBLMxXYKMRDaf6cmJCPsQ+DF7m6hjhj47vsF3rFHbbzR
pxGhWf4uIK2VAwvquj0ii6wJPEx13iwQQoJ6FJw0w2n678AJgcb/2Si7nKAmreOWdo+UyCZLAV9u
3sfWXceTvy7HBe41Oy0wRnPOSgF0u6PbKVFZwpnYoftLbbi2iGy5VM+i9aO/Dehft4fKkFtvQBr5
Jna8MHp0ATEivHDJnjk16F3Q0AMstyrMX1nz3iW482OIiIfa+LAktqzJi7DAvwMK+jUDYCU0LSMf
pdzOcnaskrYypxtqxI72oDkI6weTDj3WT/9DWPoPjzUTkDYXowIcPexLtqDEHdrHfC5x7a1/0Z8S
cHbwMo7pkDf+QLdyCws4M1CKPLXyofmSaaasXiGWAFTKvHjpq/ZvTZRlw43Ww+M7pm1fB/XhANZ+
MjEmzN/75Zo5yZHHjwV+m0lKlP70EVreqHPWNt7PeC0bvL9fV4dywC068To7D1/BhkAyzJYyhWw/
WbO1qtXMt+HAx2i8Dkn6TA0iYYsibEyozjWyXKg/c8Nx75JXhMLj+Orbhpvnd81bezIWmtXdeMIQ
+vn4cEE6FAetHWHHtmtQOS57wOz031rk6S+wD7AyRRivOl17H53Zp1yU2PDzbcdJuojSKfin+Ia8
r1670crihGtIoUA6xu4OVbVrETQgKHcrUSLOAoxQJHv622kd+K2cAlOYAX3pYCleQcM1VqeLRzNB
25lAfyiIIcULRIxS1q2sWIL+Dpnz3jwKTOgJlpnyzh7nBTHMlIwXtyJSG66AiGu7nPPJhdWS3MnH
KGTz64RcUbPyrv9/MZMKsoHoK6ld92AOPAW7W80Vgdb2mrcjLB4jIXHs1CbBTB5lUptKQYaWJ7gE
o8AfKgA4oBq0miC0zSVfPTzXzqJ0Hgug+54D5h7KfffDaqdCC2/jUQ6EZWEjWxsaosyyjBsg3DIq
SMNlWv0eug6BvSUaiUL2kekXBW4kwQ9Pp2+5jXx6ZJvE5QFSfWRivKaUarciorCWSn/pbL8bfCz+
whu968lKfePwNINk1y6Ea+J6rrj0a94RbndhmZwL+xvvLma25K4/NlNrGGBHwu9eHhOl8ONcb5PI
VicfmxxjZNOGR7hCMmMHa5S0bB6BE94NX0/xnI9lAKttPIoRjBtqG5nrdya/cPTMkXkw1ZoDJLGS
zEPIt4JTJ85VPrLANAH07KKcymiLsMGcEkQTCHORTPWrK1Prmp2XSfFQOKqDosvXIECpKGrC+LWG
4eRTNbvVG4lvL+G2GgiHkpxtbOKT69QvrRJK8V2yKMaKHoki0Q2iK5MD9+hXOPBwyAwORRclYHEd
GCzxpoGp6wSSghGmc4fY5RSqmE5AMwx0WlXelr1SrPXRKphY5+G1X6ntz+Xakcw1wrGY6ng7xOGk
tgUM6l2oYsLPXB6RxfyfOGmcI26Uy79XMOraqlY5YbyloQMLMNitL33ALe4iIyiUEkimgCW2AwAD
twvEfm6G4YKsdvvByQ6gglJn5fclY2+3GRIG8fa5iJkIOJDhtGCikbrB+Ec8AR1P/fEQEt1qbcT0
KcDylH2EfG51rmKhHcpmdHXyca20DmMYwjf1mGx9F3NuOJmWMf50RGh+bFzJRklO1t3ieGTGRBLf
MGG5TOzbtZyDPM/2wFqOfTKGn5UNPvTOolW5ptTeHT1DYL4yagXfSAMpaEHm533aXMK7yFxImH5V
8om3QM/t255kK63X9w4LA8jD5sJr0aTG7awHEiW0J8DlvD730B7Xke1FCm5aaw4QXhXjVNCyrf6i
8g6/qTXIAln5PC2nNHEi5lnZvxBoa7FjVj3Yc/nt2cX6RehACUMebY8JA5S4dC+qtgKo1oEHWIX2
BZ+WQDDRuP+U0IaSe9VwZrXQ2XmFQR/w0ybYCbWIKhSVdhEWNqV5TxMdsFbnaTm0MNHna8S9IpF9
Z2aQHczsGg5M2QMrDc/5hQoyypZ1lYtJbBz7IxhLbrDaVWP+4GPAT18AHEm4NoBXHfmddEGUxEF2
l/J6DsA9HAlrSVpaoCT4tPt5tcYls2tJOIO567HaAVCTIuMcpJ1hOA+jZkw2uuiw7U+hU4SjuQUS
TFkyIY/RuuGXyaNu2JgLJ6crxKSSkxTuHksmJPSkBrAJWuK46i1usRvWOB3Qq9Mdl1inZh4srZgi
84SbrW4xh1EhP58d7L4Ea9mrHNtlk8gjFv38lrK253Jc8elaqPnTi2WTXhVfbiaqXjujhtn8KL0p
yV+BsyFe00VZ8NDGNqD0He6DrJrOMCkOvTJavm6+trMs10Bf6iODkfxoAlRTc5BiqqYAtuDdTDrt
nENcMWmoX9QKz/fSzlKYPLaZ5pYLDJFtXUAZQpOGec6u0SlYE9IuRGVf0NOBeAetwINQllFJpa97
JZyW86iKoQ8hj8HXHKhFyP2WsgeO3GpeFKRScT8FXyZaK18Ks02qsmWbkMmDmG3zvWpC0P0TqVKa
srx5u5660VauIEOme7m8e66rKg2lKceaLZiUlMw3+S6SgU6i6kqufOnQRFT0q/c4Q4jTj94y9syR
dM7Efcf9iu8bvOr3RgJZThcV0hhBrQemBACFXBUTJOdD9KK4I+VWPV5jcN5nbC7CQxiIn5vMaJql
wUM9+nzFDSCrSh/xk4wuqZriNKhJ+eDXvoBQFHisGE/sZwioiCz0PGRwh46QxHdwD9/wFiO9Gw+S
w9fcJXDU5moFoIPvdzw3xY6ZhIh8aKoEJkOdD5P0cri8W3dDkbEZ4/VILf0HACuhvkMVN6WHTkD+
iAn1hLBdg1bgJbSkWVfm3Xk5f+Bz+/31f4YQ/ibtgFc0VhpJNk7ohf5VxePbdMixSjPfPdaJlmf0
frCClyXfw74LL8lRrQ2CNbHoK5HzuJ7wyBKxBD8+PjhAv2jpjhFJ2+RrQgO6ITm/3J4YuNJJK0qN
o9WzNTF3hP9bwKXOZe5qX4vGYambE+X7ejDE43tSwDkgimczawuSPuip5LYjHzX/W4Fzx4Q1qyn2
g7OGH33RS+GGjHTLf5f+b3qGhnJSHHxKxmV2nhjl5xjwWpuVWpnMIGYcJ1pQ9X42WuhV36fajz9r
ciLcOEMIBTY+0qO0YB+jtL6Nfnyk/HmcU3yPgUIJK55AizFlgAFSj/hv6i0wnR8hx3OT53UG1AhJ
0v+m5Bhtr2OcvNzvfkxQ/ry2WrjuAAWcGSovYIa/uC5Wy/SoDq7Gfrb79xXs20CnDVzlvQlakXnq
yUt/K8kLpaeNxigeT+wHVppZnK6igSsszQBz1UDldnNybkpzvH+DHFW3QvIbEkMtBtAmZi/6Y5vz
Fdj1uLTV7wSGI+j9OCo7sJl/EdjM5TrSPe7xwuzUjAK0qZnmS5U1Tk1RR8Sdzy/s3f+JHvV96Qzp
voRH9Nw1Pn6O9nafNYSMGyFleW8l/CqZWruyTW4fSMIcAEbDhPI8e9pTpAGifnroDnlLS53VW+Ka
MOenVVrOphnW+IiA5QvMI6PX3GWOZe9W8xmIwqSmas+BbkFF/8KF1YU6PjY1yToVJEqOeP5E+Uzd
K0cWl/VpF2mkFinmc0d2HkJJxfdkvdHDahTohLwi+7Bs78BFo+TGIHx/bBjc+4fPkPUqMaK+K24d
VG+ip+nJLSLk7yEMH6w3CmkGmEFSpO8v2NESyYfvFynQZ5sjyOFt5hN7ZAvdsvAzdE2/itlFqlFc
otVBNJabS0PfVcJwY8wrAutVb3j0u88ABTq68jRp9BXxB617YWn1gWaTIW0rXIIfYdiyxZ/T/tO/
6xIienZ1PHXrNcBQoHGB6OcsmHo9oWP2ZAZiDVWA3fh5x/hUQbew4voOVz+EiVm55Uku6gADc+vx
2r3WA/5aEMMxIJjLO2iPchUYQNf94dv6BucUbuZCChMp2KKxuoYffX1pi/UHVmu0BuNhygSI72PX
XklokSN/mAAdbKuuE2qupy02WTOrB2+0YD6IIlCsu9E7Vv9hVOYNEMhmY0fDYgBaqR8ED5RPLMgS
pSzFQimsioRXTU567IltgKAOI0ZI8Z9JzMKPSBm5RQBXVcE6RH6wmZPTqbFK9O3UmpVl5YSLmKPN
AfjsTq/GDfC0HH//SQR4AuHuZ8pyP4qXOrqegxXGHWAhA61kZmi00FRWwjiMiZvkZ+gRwfT8T1wg
hSC+Jeaaa5B/9DxdTb2vCXuw2q5EyWwkY/unrrnHnF7jXoEELdS+HxAOXD+JvKMs17n55Od/Wj19
z8fry5uUR3f6XIcpH6eRNJzgSRpqZIYlbpHx/ItLu7h2gF1vGHai2r0YdRzZUQn4oNiHb7tHkyjL
Tbml5iyAm0XMnJf2rLBhpurzOn5SePwT2zCzu/UGOn9IIS3X2n7+DE5zrgUx0yaCPVeCiamgxyaU
t6qFE/m4m/KCEnwsRX4lhihtB8aVlvHRZ2cEjAO+K2DJeFBTX6bSXYM/JEReGSgC4zNcfc+5KcwE
6ZSUlsFhUOqVgsTeU6LNcofExn+VtNvdC8OvHhjAUasI2wY+CkhbmQkJHKNc1//YlQO5eY0726jt
JyGtHgc1KX5jzFFIOsWdZnuWCQOI4bNtdBU3JUK8m0X8F0TF82mOox41HA0d1C8loIYcahtMKqdR
3cdBz/A6X6E5hx5HrQ9M+G57YeJj/dYODjkleSAkhiAx/gBimJBKyuR9dsQxZ7BBqSbeR9K8lroI
2eTC2+oWT+9168vGXUf2mASp68lI2r4NJiGxbiio1VXWG5e+ntwxRto2bVXW76y0z0DacEvXq8ok
rlXH21mztuR8KhDCCOjn1x3U730u2NCXYyebJJYOrZ1SNI+CkE8n0o75VmtduuqDKMkHrE3SQh2b
PH5Egy4Rux/KviTs+p0rl2WwExH5LhO92vQO3E8dS74L9wdYvP1Jfhh6da2SHfVLoBG+MCeYaPXo
aPtq7xG3EBd/xqH3TlsenYn3WLfOJ+Xynn2dPUOVdehilWNa/VJaainY0X+IfOu/kHhwGnCF2xGW
malnUIv9R4RKNiVjPkgS27QgDTfFoxBNpv664IkN+1VOq7V6W2q9lZFz6OmDrMWd3fAouWCuJ7r8
8sSi94wcCT+n1yprOeMtFBEyrdu/UBKEXlGu1nUE8O1Aq9kmxeC4BNBNN/WHQ2cfFkENo0FpzGmW
ybFtnZlKOS8dEOrCbviXehz/B7wNnNe1WouRHU5sE7htkPjBq6sQbK5SEl8On3ao35jc3ZsyvWPM
9V2Gtv+1JqpdzW8RR/oOLWsJrf2x9Or6t0jvp+8/O9GFIIfPySpi+GLkvRoq21qwynCySw8DIpnB
T0rnvSzoaGzyA/t+MoaN5pdpuzAWG4JKlcKh45MiO7gatmUKJsxLwlFlMVcI5KKXSijZnbMgT2zC
B9NKSh5PQ9v1yUs7qpZdNZifyUI6OFxSHwibezroVHYjRZiuQsu7yQ8igYE9TZJZeDmB9kSdT8go
FgF0I3WUEYYvM6tgUuit44K5lrT85g40WCkfgOtriPdMnAQHEIsbT/lx0d0Yx4zHEsjnXvbNzHKU
43i9pkg+2Q6UC9GpvZAn6OV5D/qatnQcGLQbA5oao6bAI4O8wTuqXQ1/53CPxYe6FxvUo14ZeyzV
0joGeFPLmuTWVSdUhe3jxQtdCdRcs+R2TCzapkgCJTICx6+6eOZwZREiuJUgX75XXb3oiOPjLWwZ
qloLsNOEWtNE2G6wAq60I1o5G8qP9VApvl/uq0YpYbESZ30FmUQa/wFNQIz+meP0DvXuICiV9UMb
Pand1+sSf2GwnEnokANshEYb8ZLQBu3LmukmqmnXUW/nCH28tpOmdNpF42MMJT8r/kzUVeryBoYh
YiDc6xPqo1FN+FhsZ9vX/aBjROhjn5b6gdXA5YJ9+ivhWVITO6g/OODzKfArVNT4pnJ6z9MZDamy
72LVM9wT/g5ya2g9LOSXpulDV6uMVIcRzwI1EwLmefP9TZTauaKrYRc1zAtl84nkLBxG2FxfXlvO
cprHEgh9aaePPSm4qF2bhdPtlPRc9ShQK/jwsZbiXAn/u6ESHxL922Ro+AmYzKXtmX0o3Mf/p3+K
yfMUcsZitcIrfZ8pBe1iP9qKCu3IsHelYVz0DiSrFQMXpGA4ZxQoerzZj3DaSfY8ixWzHQAB9T54
oeXENXfxKm+L9FxVUrDm3BUjxOq7LkDSuNbRFhHGV0dpsPS8WPgKoUOrJa3m8yhxqltzQqUQOWoi
N/g4B6huXly6ptFpNEi+Nufzromb2XpIfBM2NMmT+j04hsj4xEnJMrcAdqQm9r5v5j7FlTk1zkdy
PQpenOwAoxWEhS+Tn1sNC7WtlrxamBKJW9Yv8I4ImnmcYWURGe+1lPuenzZ5Xj85VfJNloC8FS8m
ZcJrFzZKLZrPPXKfLNEOp3WRtggTENLf0BAUWOUvtob5MN3cQnZjvl2xLGeyE6E2Z7wWMh91Hqgm
yG3XbGdxw2Yx4I8iEUdZqQM5XRmALxDcUkiUcr6ohvZnZCPBBfwkXwLwfODiNrYiQWj8BHdmeMVl
dBw3ZqWWUrYYWEai/XHkiAUgu2YvmNXYjLv5Q9ErgV5eZfQm5h0dPNBo2HiK9lT0IcQwaswzoR4a
TASvko4BxAldzVe7JHT53b+gVqn1+gKWD6V1iIuevEXclKvvPK3rJ2ZRH3TqZrNYfM4BuvlmLkRW
6/fR7QXi6OIjE3OM+GxOV3ztaqi+ZvJfT+S4+E0/ecGr5eCSBQVuA8NTx9TblntHD8YI0dbWXcD2
qrBkrBXC6xT41ueP1jUoVdDs4g4PwKi+5MlvFrfEy2YywNugePcUHHJKD4WwjWzqOIin3dfwlFzE
dsP4Dznb5hFm9PKAzTFKQupukh436yZMQ9faQof1B3OYnA+aZR6EG4GHLMMGzI9bBCoKWApu9EbX
gtZ1eHh4dd3mM6yVS4FVzOB/GLZgyWZDWO1v3/btLaOennGVcUsDdN5jfWUMO4rwPyM9N2x3Bp9+
EbSJbCSXkrqp78Ei4aXuLc0+O+b2f5eMwCmQaWTygIWq/7GpXavxgpiMm/sim5+9mvvDhwXbnbA1
0+ymcd5ajpYEltenx10YlXOG9Al03Jv0GecdzdbbDGYoppqVpSaqI7ZdKoHhdtWtQCNB+23UFGjA
4fnH9PrEeLEXKp7EvAJGgVmvk7QzJXOBQkDlvjJ5/oh9J/Zvhji8tyWCxWg8h3AwaoMNukJcRkEO
xfPl+4TD9B6L0QI1p4AYtH6cJlFlB5UUf2uGpibCFD2MU99iNoJKleKkUc01bHqAN1Vh3Pn1EEvv
n6vtMlsVfD1vOL7R1gDerqsDzR8k5FlLYIZP7T8C8zMylloaoUPDgazY2Gc6sjlMKGRHAAEhhA+6
9DZPYDQOl1qlT+te5lO4YZ+G7Eiz6JgJAaqxnWG1ILzbtWOHMkcepErCkXzE7csJWGfFBFHxOL18
OtVyYMqPiYnJFy53kpfiFt0cBb+0Bsiwfre3ijJD6Va9b9ZllvnN9rLoyzDUfNpi2XRT3bHyv/q1
FHDPXtPeULamexDCQ865IPaIU/sW0wWyjCXgQxoomygJ2cFYE238B14sWVw48UYvkBBpfEa+fCDX
N8n7s9iPU1T5d35X0dc8+Uda9MG18Su0hv40aXUAvRS1j74spQyf7aDPv6I50auz0UTCx3c5WkKl
MkgG75p9u+XXxlOM/ia0xQ77aMQDpssVQFx9/kH1NE9h2+H82aV5ffOWJMVIYhK0rZ3m61u46jAy
F69LKh+X4KWdCF/CI9pgPUFtyWWDN26T3KjQnxMersE/PJgNDDamR9xipzvtm0KOauQ8so/aDkOk
PIHi4KMKWepxF80lIFrHEIjLmZiu68PLOdcoOaZfvjcJeAW0EL7BSp0MrNmSB+RQfBoRwU+5RRxE
h8wJh4CBLvgLkxBMskwIn4Yp1h5f2sf0zwZqudzar3JzsBOTigfoYr4PdUhEBBnCj/MQIqrHZMG6
sGnxKNOYWNIBYeJHpyX/n0i+5DR9M/u8cCthq82fVkENKysunqOIDd/PBa3PZ4oVBfa8eUTYR0T1
m0I1wk9fwkSRC2I6BWRjntakRHfihuHZbEs3s0lWmb75ovidfe5VsdFDRYpYB9/8g1FKQJlhjnXr
nEhNY0w1w2fxd4c9xWdSzb2Z5eKIpQFvI71Nu9LH+uxF17derkxNXVZd4TL3XIZ2JLmterVohAlo
ezI8rNU1iAo5Nd775s/JnVD1y3w1OyvKIcnKJQPx8+lx4T5doVdEOIxCV0kC1h3AbhbBxtCEN3nG
rZD/Sue5Hcz4qvvqsOCPFeunH6iyOedV6IgEg/puEfw8PRrtSA4NsRFiJnFyZEUvrUkwmuA2Khn5
ZLEg5KSp2HNeDw053+AZUxARuIJLKJo7L6L6iQorRVDKvUc3AWza7cAYxloJGADg/sbLp+jgqPLI
No1m92ULdsJ4VRtzhD8O6qdMARTEZI7UgvT5iDx3ozgEaPgMxxBpvtRpTf5j8DN+Pkh0GowPvtsm
wY8gs7JP/TyhfPNE4w7XahLhlIkZXala6hulApI5Eiuw15m1HydpVzWitDbr+K64RDtQg0fpl9d2
SEj7X0LJvIOs89nGBwC/Dp2G4dkmEIoIbKZX3o001FseNKKTTjm+Tlye1Zw9ZImi1F4sLGGYRDlf
/FqfFxcawOGzYPq0eNIMl4Rs/Xkhd122pX/6nl1AnssYFX6xZBaecEFlKtKHDaQPX36JFUCh6DI2
z/pRG6U07PidxjuXqtsb7LQfbKE15c551qFe7v0HdSgQp/E1yZ86jaqRi2jhaamRRhXUqFHaatxl
WH++zNdDweBgIEUX5qwyyPvtNS4Uth7cIqtJooluTwsnArR+qXkHe/w2RNG00wVbLvHj75pGjXXp
HOOt/0ia+qZcBXnXy5Iul/+hGbp8PHo6B4UqMIwulMbGAhFgSr73t/QdTh2EUDHQeAo4e5G37E7E
n+LFUlQEj/55UlDTbBQvnOy3w4l1YBSvwnB87uqioon1HG7qh2VMlPjoZbaxjhN3HYP7AINSbmf5
CUm4ZWj7Zqh0Gy13AqPB3/3fzDSbw0d6wplm9KVO2h/gBu9lgauwJ/z2o2MY4KHGXj0+ZU6dJHz6
k6bgoCisrgdEqqZyFMUnNuE+XeAMpuMHUA/1cjei/1yr9wUiDD720ZdeEjrA8Jwi6IfT2DT4GI4u
QiOHlDQHTTfUWYuxHYJeUpbG1B49ltLxu1gUExlXbSHjjzkwB0nl7EnxdVoCOIDw2w6daaZ+1g8S
msonJQK7DKAyWSEmlt2+vW9RVEOdoNVnhq9SyXxO/GV2ofSOClweVS+wChXeU/ef+54JPz9B+BCK
YDRN9qpgUi7g4+jtDOlNWkbETZIytk7/eLZLKbX4MymxsvO8D2dzc9KBOmE57R8MPDcdMLzBsHK9
HxGiaY45z22/0y8UOkyDI6KDiLBVjVA8fWwL3T47Haj1v1TrVN8Ut0JA8W0z99rSIugAqmXdQEWG
uyNeClEib+rY27lWgXygueYUKUFnw9wE/Kx5d1CE6oceOEWgIDEre+UQ3BKmVMR1x8LMFHR4XQPi
IDkrnFgFVb58PTXNZ95WSI64723/ZgMfVQXEXWKz3kCI5K7G/nsdKtpmCvVmmf8kGe3xZoyyZ/As
TNpUs5RimzQCVbBKgOHd79xHwG3mnpBEf1djN4V9J+Hv0pNfbTC6n+LYEShLhrGUMYr+fCwDRXOr
6LA1x/BCyqLlJNBsD1cwo86Ouy1hoaSdAWBuI+Q8KT69W/iUQEAjEPzpU40D1GdDyo7ar2yMBO7d
C/WwJaql2KdnpuNZ5Kja/6q2zHeNPgL/CjFyadkfVYNM/EtG2pqmmMcboCngTUkJ0GZ0nJvmfyxu
sule4Q/0kFPlhDE1sON586uxMGYqMcXCnIMzd3/z4A8OfBRn0izeVddG2ZqW0ivez1uaacRLqXcT
3drWxh+aiZFnVsKdit1PCKKa2M2XcDWh4gFwqcZHkviUP08PxJLEXcCh+knqDSqDNhWK/7vjiJKT
FZVvVbLkLB2StQn+W2VnJEhFy4IsNYJOTtGzOwdyY7AJtQj4YMfvqDj13y+Q6AALb/3+uOMfRIRP
Shzfb+lTtReEmk4NBVMvoirH/NQh+998AFO1IpjGcz2UrVxayrBe7KfYmNnF2h3nVzt8DYpBZHob
wDYt3qXKWeFL9fIfzY1E0PRl1GrV0kufC8mwVlCDjAo0uNpfMsE0tcMFQItppE32B6vcX4yBQqMt
jvB0mHsVn9uxWXSsZrLZC73gydwhvIbXkUOoy8P6oNBb9kCX3oJI8i/4ZVEWBguTOi/zvGHpHekO
UdvyGFqy1mYMl2jwfZbIPXsGj9nuHFWl2+r94zcPaYTWVrGUxMdEp3A+Cvti0KHsParX9/RbLjv4
FBOcGDuUK/6uxk/qr9E8+jFSYdRydGByf4t1jV1vZzmaTiqC7hF7aoPz2JnFzyIeB+OxwThZrxuW
mq8qLl+rdStP+wtXFKLe1MXe/xlD/CplJfOhDD58fGJJNNXETnJrVcTyp/7Wpei0fW4JraheOGmA
6Cp2PnspdQ1CoMntNiSoQLon9z/cGa6mqNYxfJIh3qvlrTmz3O2yykfvrIpTog/x2QqnKmqLvK/1
qAn+2D5rel2950BqAE5rVRj1RBhayBZ2Q2v6ZvKFfQB4y7cZKBYGODw6owKzn7gjypcGARm/WN94
rrKQ/XzKMHDX64RrZ9PWkEM/Tv6pD0HEp74RcHEg3bJUkTxVbkXTfh9FSO11a/BxpRIrGjYCLp5d
yiV1PF3nR4PEDEdF+VH9K275nhJtrOV6OceUK28bzrg8Dec+8+6+tWBy8d1ShVYCRwb/2dKpw0gZ
XKiJBNqBW6lfGOYi7fEh2Xz/ecVQIREsg+nyFp8tTwSr0fbDL5qyzNWRZkPeWbIpL7QoylcUkCkN
/N98TwhqC6vgWUDtD1JZ3abinpm7L4scu3SDpxLBS3FGkgU6PQmggk+npqcNTp//Sb07/GeBGpyh
vipG9nglbAwX+Tb5iJEInXe9IgRbfowsWQduCHB2PTpgz/INi/S9wwnWEvAJApefSLTyzSxhRUVK
gLz9iIswDmqj3Av2mGyJLzpcvG+98cEpowSCv7cJIc06/Fi7PdpKbOggbjHd0hmeSb9961MuRMsO
a/P1UUCF/aySpialL+xgdHns4u2TNmEGLCz0AvrU21TGRcFp4PbvzugimUAb+gBjlPDkZuHNb2OA
9sEYaoUcTHauciXFdJBzfuzGohi3mZc9NW1GLn73UX2dkuwPqYDl7UagQDcwluHCd4/FwDPGtRPD
OxcejyI448+6Y7sgZf/XSBMjj1bTpzgFMRf8HhbINA4rZAgwwDU1afpmuHaLYQ9/BA3qB/q4pfQi
ndI0NFfXoiU0eMvPKmcaYcE1GuWcF5KZR+Vr/TaWVPqJGq1HicS2yp+nahP4Pylo4gZn4X1RZ99E
2njAl9BcAPBJEjot4gHg2Awf1p+xm/5bxdUIj8kPab4uobFleTbYfPrj1LQO5sb8NkWHQ3R5YF3L
H4VKkOcS9tUQdbkalwZtDcT8euVRn+YJkX+D8zvfQH/XdK2yiCKenO2+qsmhMRSVv1BF/majO/Cu
vsa6TfDf5ltbbMhpL0U4Q370w2PfgvpyWIYB2rJnQJaxFZ0fAtkdWai/R5DfjlHxMMj93N8XEIp2
XSDHpI/3rlLVJNGtBTPcNgljJ7KsLm3L0Jv1K+MXrumdwAMiMOF4eYkqaNM2/KDRCsGIo6xApzUp
A3AXjxWpSZFZR0CRD75/YE5kGPBuSxjD/9WCMS/BR8xywWC3nnY71plJ2DykOzZMED8f6xMbpQxG
4FKi2gTCwompnl6IFE7JVRWKH9ASY3Qfttwj2rTs+8RoP3o3jn5AVFSNY0zrxNE+3VbMJUjl+Yst
74hn0DTaAtS/ZV2fibJDFNWrlAlckdQoejwrQeOzDAgvXCW90WGivCxtFj8u0JW1b/y0pQ9/iQrx
Dfn1vdcHlC6CCrPXHA6yJ96mip+Vl8isg3Taet2FhjwUdRoU5GqZt4aq86uchsW16tKpG7bkQQYt
HHK6IBj9xQjQfyCJm4ki2hK5YXVSM+RGP6dxrpThYv/I2msmfX5TM5PdO8VDTgOoVsYZZRtk2tPt
xqkqq+cE5CTHOFhTK+kvla2E96OY+WRxmmN51W8qKErJL0LawnhGHBBtEwHUfeFOKEtewJ5pw/Nr
Mi8iV8BelLB2jXNMgzVizNLWicCD1mcRJRO8K/lIh7RNSUchuxf7EF/sjNlLwX0s2nUWBZcvt1RW
R1z0V/UgEWjTJN6lRreNBWkW6hrTzbib27ihuqKundYra3WMsvGdiFzM0nb9yrvhfsCzkuSN+LTc
fiEq7wo9dBwpBznxK/ojR+PHXwFIpvg85WcswbN8qoFmi7eCN6Wv5BjQvexbfF09UcvU1nTCq03b
RFJWjHa0Og096iiL3qTEXVP2fKhDnuKuqnrfU2Y9SrdtgCgZrXvCBzl5ndgAuiKamwtQCWi/M/CG
KLQo1idQocMQ1caNRMo5lCb5Z7MzpoF4Ra3EkBcLWrZGWIxmTVAo5dGNDh7p2pmrLdedRf1qa+m6
HUddqolSV4jjQfM8I9uIxRINJsYLjeMW9p/Sx7HKGR0fsjHcWBHP+8xcHC6Zmw5GyKNFfW9xENqj
KwXpDuwlLvBwJRTIqO/pk6gECzqany3LTtmSTg/YKweID4DRNRmzt7++q8HlhasSW80XtYn1wk9N
EDamQgU/k6OyHgFfR6AZBmqm6ccGkvG89drtiKSDtcI4JDn6C9WfWRlALgns5gjY2g99cHJpn99H
G62u4KW605ti5R6ln7psdZokDnORbiefByNZntIXuPFRQaXfH/xtYAsXjF9i5tPbWXJTxzHUw3bI
dgS3Q/wlk8jswz/uGtBFveHEgF2CkeURwf0QyZAG7e+aZktLIEfN3VfkaEcDv2mOyMRsfBqxsUFf
pqH+fZXjPNz0K5/PC2oi3KyTQpcnsMZEhOEvRaQggI7BIqOd1z8cvKcugfYdyOs3dw/uqWWMsZK0
2kq4BFmk955Ei/y/zy5dJO32asHmyMgM9vumRqz/awWL/3lDMT+CekzJh0aGQmK4keETPposNWT5
tDCHmsO3keJChas9zZHzPFKvo2hUeMRVXpdWzAlJTxowFXCpu3rerh4ZIwQisfcbyy9ePCyn9SFI
2/e9o+Inwg2C4VvDwABSQML95fVYqGVT2nE2627bYZhrd1wd4yJ/Iz64espHxQmvxNz+1ex3B+ke
67Sgih5t0zeN6aXlYtvoK0pePNSSP54984aaT7xkiQv+lpjmcKuIvbSUqmUfDV/WE9i/4RaHu84a
58MNnTdanfOFAp4OWCU0/XHvGLVZw01Ck0XTZDh0Eb2vtgO96z34lQiStecq8/WMaijZFm1PjJ9b
QlMh1mKlMHF+9LUbVk2VKuARimSwZTDLWh3sMddLndDIC+8wrkzWGnZ6oW1U/6FAe14wJ9dhrHCa
ErRtXjMDlMhjqgp2uxrDwVFfMhQKNbd0jfu8oZ3wOljfodQ+RFaks9nj2VCfR12FlFHLBokVNqYb
lKu8xLCfs6oNDov28CwZmlnUVKGod+DSu6NjL/lH/k5uoLTLyMW4DUes6S5ZaItImoIjmOPxEzJ+
JaHjlk9Zqx51FbYCqT6xHyITmSfwRAkKLhk3M4unBwYUgWC1+QGsQXyZhJGAJzg7b0/99NiKNuvU
Qsq5Zs7UUKXDO5TYaRebFY1Ky+IrKbom9oib6pr4FxVFKrZhVAUmD42pQmcNtbLNb7GFRCTc45SS
VoQ1imXARyn3GBoE6qlLKG03+XL/9DqyFvNKjX6AYyj/LD+tYabrhao0yeRbCjFQapUtjuxD9nNU
Gotf3n3Tsf9rf3xI+/d8VZxK3uzInX871fS8pN8dz4bJef8B0gAPfLKuyOp6KV3IYhRkeSANpwyY
aVTnxfEbksCQCNTys1kA6ey3IHFgFanl9dlLvRzeeI5JPH6/ksNfVltnScJYXh4ejmoy0iWO6NRp
OP/EDUJw5ePgVxBhYEi41iXeRMPTUdfTfjXRkZlbzFvQqu2DoFBU9Gp2dsrpU3v1P80wkJcijMHO
kHbjF6HH+mFAvoxsQjbXSuSewJ3r23qyetQf0pH+Tiok9CLZNWZhBj9t/xrZweucXNZikK+unQGo
9wIHR+Lq4bxkvBN6KO+YBGeI0XyW9w8wk3BbAPq3z488qfGLVakocYyOnz8VD5gX0Jk5OPj8nrne
LWdZlMSXJGA7uA7GyTlm0ruw/g4XUTU+s4CwaaMHNG/b4VzI6lj6Rvrpp3RAEPP7g1fGDEG6+yr7
TkMjW9HTvBdqHm0a/BF4O4rCXvRIRkZZj1A5gUtxeme9ho4c1jJKhW64mrc6uyrn2a7MjmH1h3ti
QL/brnADLrBhd//HNOJr3XPJ06VvfLEZD3w+rgTz7ZlLosUCtm9Iz7xTixf0r+j6gXZjhBcAz1sD
UKElTCT5En1WYjDTRXlCbZiWGXfq27jgD4xDuICOeiMoR6zpyTfsnrvfUh0TFsNGeb17DXA1Qt+B
9j3OrZvUbC+sgHMQVE9QbBsYlEPUhNgtVZTUrvTYr2ehvhazm2kiqFjJtJqCK98MLA8oO7WrTx8G
SHohn8ZZ7ftWqvLAMMPTnqzmX7AaM2dvaosmSMuxLdrub4GDElFRdRrKjBPdO8tEIGCqCbr+qcuC
OlE8khadcRW2bf5PVr+aLYzITBc55yyey/EhfT+tRKg0oIZCirjozWZs50OwEHzjluAMxoP8NLoW
jIaHS4ocopYY5NeUDjuBrVMSaIOfyvPxazZ0YBatLKiPB8XFMGzASD0hLBJATp0/8TaFtPFd8Cds
gFtIKsuvYgSrorLMIMSzibJ766zLYFGLA65Nwudos9IGAT6PzTs1piXXsGGKH79WK+cbR3dgVd7S
k/6XwOyQsopms4x7TK7mLdXTImSqcwEn4nMhBL4aOyr/A7a8s3Fvn/ZrotD8feuaTv+Gm3vr+/K9
gwV+Pm0eG7qzykXkuKVTzm7WNCwDwEtZunRmMq6K0IWuTA3Y/loDkfcfPaUkgCF7bUbXOkaAgxVz
GjkXUVOPqdwe70Xv6VlgXmdKiitL7v8yOJAtT+vjgua0ffz3dR7ou+Kf7O6+IlkAx3VVCV66LcdH
fF4E+ivXnrzzb1S7URHcG0/Li89ljmjmM9YtoOJinY2lVFPPUsAog/DyRyTegm+sFYZD5tQBsvEb
apLWU3j8qGqNSb+RvUZfKIod9xVqQyqTjuxcAWG96rhGqIcwpk4l8gq+JR519P1uia2jIUHUQzQ2
oH4BYlT3KAr6qK6wqeAwGgEZMq7Q/s4q006sWHkbGs+fFfYgV/Ly7QOf2VVcIlnvRhALiuGzZr+X
36B5DW5OoWaBynYeAa2mqH4qlYJiyLg8GHYGOr1IUALnXW3MLvEOKrifciUXJVFwDfmaX3536zbg
RX7vOQWwi1hBDrlrEQ9Ovvgg8alM/9FVcWB0B0aS+vEDCBD+RG1hJvLJCTO15ZGZU5M9CMauoATA
6+E5E7E7OlrtMVBIv9sQP/Q4MzSn/v1JtAUbYnvblZHjZLvgfSej2yh3tKyXhIgk/C2OJM3+yPGW
kXtwZleNYmCL14O17r9ClJbYp01LHROcIfDN+T5EqK26ZJr9JGSJWfKzvRjbpqcpOi56s23+D9vr
va4QW2MRSFXz1mZRCNb1XK3hLZvQ4nWJND5ATrKTrGLNwHW+Ci0KJ6u54vL5hz7mhCFMzYiwQCEH
xbo3ECbg0H15hYK/a9XL9g67tlgheXMf34wRNgi8pPuQdHB14Y+rwIfdQipGYru11HZyRi6e2px+
SBGSXKNkxg2xgGKwIvwNwHiTBgFirhLXyACSk4uLzhNoUWnPet9RbqZctUL9xv6vl69NVlBsg6zI
rbuYoE5FMmtkzSxwrIfWTwgkRcr4clQVF0I+FIOupiKqbrY06DqrHjR8H1aeUUhctXMV6RXSvFYu
PudD2iuK68+38Vmfv+0EwOVombaonN2YgTsPt3jmeWdWDpWojtxrW5+uVRD3ZZDgfTcgjmn9248V
dEeJ2pFu6BEgw46lUsfVCDwssw8YVQlZZzMNyhxrZ/7k+7Drr4eOIc6uZI7EKa6JPty7UXi3OX15
D3tKPjhvXONBcbd6/xvak8QJLQ5cBdQU1aIkTPGUu3A7hV7yLOdOuT4suxO75U3j5swjmrYg61tM
ZYudNKJReSxfX/Jq+jtiUSIejiF+z13wSdvJSG7Xk6fusDVhoYkfoxW4chX5WXkvgmvVyMiJOCfs
9dg9gOtv5CNwNxWuVONzvedRHc1YZbVD2JTFNJK1/s5nVfBcmkviuFYveBdIZG0mLdZrJ9qR1/Pq
4DcS/P83iiy/Vm4UhsEoJgbtPDpUyslNY6R+mqYxCWFmvSA6BttJObQ64GRGTvJSbtPpxddH/uNe
7pcQutJsF73+j5e4BoHYLY+m6wAjRy+TBcPu8uh4gR+QbuNyu3hduM1sgaFnGkTXykmBL/t5gCCA
X+4yeuQZPLIirO6rQYPKZTPVARFEURDrRZ5miNpHNx+v6bqtkGeLk5CP7SfUalCPQ30lTjP6SC7C
1l7GJuHNEEdJXF3aveEddFJHshA6We8Mm7kQUjMSSbFuz2s1lI5Io7zoWgl4xo0SFRvzVRpBisq5
/EMciwvNn/6HAc6mO1XdA1KS9N/mO6fV49Sil1prcBdU/SBXl66gaAP68KoZBAaotY6Kg6VrtOct
ogkfyrqt+NhZlorfeZdBDlk4Ojipw2wQWWucTRxJwLJ5u8fuvM1s9+MQXJVkTzj4uQjaLo1WcJUg
bAIMtzXA2wWabApm+KZOiHmoKqOdY5Y3uhk90EPmiPEZOhmjTYYwMxZCUIhMT0Gte7ichgZCf5HI
p+nVkgZIUyfM3i0trjT0AVYVLmp/VFicvSKe2zleHWKNHXs0Ytpjk5bDne1uWU7Jamwa8sAJDdX4
owYIr/3hqyWLLFZwgcTvaBrTNBQCRVSS6KsAeKOEZpNJRDrEqK9GTT0wRSyFa5HCEAQdAphX4cAJ
avnQT7Jesqx92i4eqR4keS0N3atVAxDsiqP1fY9rJKK2fh3HS7NMQrETp20Z5W5EF4R21MqR2Kld
pvJHDhUJPgzXuxHnfopqsZOyFGijDjwWJ+qJLZDi6VpZJURHv7gEBSboZSPMu2W4Yxf2F7gtN1wn
CQioa1fDOFJlJtDoC20UfFH99kIhrdypv5M94za5x4q2Fps/OpsExkOORvMcK9+9vBHLz4vxuVNk
iA+oHrQszO4cBees5GIigf6qwiuPaSBV9izRrmYZYCjNL5hDLlDajXgYtjoGfeUzF3E9fk+sFU0Y
8fkmZFBeiZAdiDPFDTamwKOq92+uW8+uhdP1wZ5Qbv7126Q+gRYXIwErG1LlVzT9PnyPJgGbLfYk
dqr0GWFF9zopGaa4JZ/GioINqaYfbR9XBAsZhMtQXXeOXhIUO+aupvM9Za7M7LPLEbqdxtmXrTxT
DkEH3d7jVZPTyjUKki5nwJYVaPVNVdvSP+OccE3g1wKKuLL+vzpJVAtSm5JzQ93XT0DbCiFGpBy+
XvzZstu0tmCAXkIGhdLi48Pxy9+abzZwAu/UqeCo0aazD3+YhHm5rqAsBINnagesO/Pt49YnkleF
Akjy28iTbY2Dqzi5WhUr8pJvZQpT4H38aiVqLe8npvrSg/VGIcw8HaDLnspKLPPcEw43JXdNGtEy
aXQgXvDfhvo7oovk+Xn7p4uVmQ1MuV2VEyIC6E8/nzq1UWFbUxPFDlBsFoko7q/775ms/XUYAf75
/h1ic6dr2iL6xwgLkvoIQU790x6Pxe/lxor4Ae0z/w3TZveic6RGljQtgQQd7ga774Bt94oSPFPb
U1usdf3gIkOIg5OrHI0Yv8LpcySVveEWUpGur9AzWq+ziWz/aS1hnE1Vrlq49XJM9mLzk41U2M2W
aK4zezNS6WwW6JhWCtSEqG5Ld5WPLWv7wAAHYt/hzEmWNZ+2RfXJ03VLfeZjUehVAi0Geydb0+Kx
S8IIkJ5mu2kYe8CMb+NuOTL/PxsSzUbLHPAUbyNQfy9jgtJr+1o1QIHLSC04o6u9Lb+7UXKNSfRy
82Wdpa0Qw9J6P/OR+1dd/GN+4dLC8kNjqNibQynrboVllTEJajHM2SFKj0srB++5i2Ti2QyFBkmk
+yBqRGlvJ9SsJAmnQQL8txKUR5aAn8hqdy9imb0Q/fjAgtxmFMg8THmeNGg5fO0TtJ0dy1+eTJ6P
HxpkTp46LaCYIbG9Kjbk1nsoHkIp1hfIppqT/QjiHuHsD5m3yIiIaSCoyOnf77y9mZUN8U3AEL/4
PaWospBQU7KHf7KZSdE5hxQfG6/AgJhyA8vzHu41iF1deDMyaisXjfy/zTrT0uVTytF0+Dsr9/Vl
VJw30ylhfP0g5OPJ/sAe8HAp4YPhUqGniDZqsCdUdHKmPGWhjQBplW3Sb5PuZxkiZc3cbZNlRTwc
/Dl2qK0WXdPmcJBMNGT/2orlenAjwLqeoafr7Flu13QFqSrNstRn8DKzTZ82Y7JdlcJSvxqvArIV
5UPChQPXi3Gy3E3NNfF00IcDTo5kx6n3axGqvCiHdE6hp2a30koG+Ccs0a71m7xgJ5yVOn9AWlFK
KzwqhZG24mwQxxD4mUTjiwlbR96Ta9B3iGoKzapuz9NAzw+0MBtA98uIfFqnyzruLpTFVXNYJtFj
Gacpfvab1BNMHNSCrfSLbF9kgRPGIJkCVicP90j+ExjcIYyR1RvU+GBuKdNg2hUK4RVuUOQbSFS9
F8n1R1tNG2SbZy1zKAuMOpdAsy9vpmgG/iQluoyail8DefmemoPDsMTipQZ9Gu2q44Trp7Uo0X/A
PIbfIvkUieZEJrr1sdg3bZd3FdDwQJe1Ep8vpGbT10tmIhtT0Rk6nfJ9ZM1cbozpBAS/Gs4KWYRg
Ptys5XrCCgZI8TiLmQTsyYy4ikSCgm5/7i/100S2chrgInNm4IhJ1DEMcuX8gixGxwgaGpLr60fr
kOG9IfUILuyR936BUxD08E1Kvey4GJK8LsEExn4spBlxM0ZKg0KzyOuss68AXsM0/ngDsKYg7JMS
WPnRb+R/sNyHFKppN6Dw/SZ+OWyZHSaQl/QlA7tLxEp53YQaTvZ1aIgqoA86s1LVuAfkXFy5sdK8
143Pg6tUPC5oS7pY4S69GMzxZzdBbYO4baN54x6mabcHbZp6zi4u2cdD7I0+VwPU6x6+/3mso7TQ
PElVotBtMliASmMv8ivsTynly0AbKB/JAx1oeL8NctKHAYNv98mmO4t3zX2IijF0YffIrvFxWNM+
vF6IJbt5FaUJUdXaB5nUC1Oo9t0YYSThadrMZoR7FQJ5kcaVkALwCJVGJSg30QFS7Pa+UUP6CdFg
Vf84IHrVuJhNKoMSDcE8YuvJm4A8Iw2YfB1BpwbnobmH3aBSHUbigtqtQN7e5umlLDnsoO3bT9jF
5o0IDtZGgnlJ/bw3j3BnXHq07ES8oo2DqRITnMuxhTa51rsj/+FFRMruHFY1NClYdhsjG1+04HOu
6RXiVSNd1ZytIqQPYVyPAkvhNlvd7qDOW6WqZ0eZb2iGIc6B1TapTUpuq0oirfvFFlScdN1jtTe0
AMIf0CrlzLJpRtGObJWa2sNZtA7uBA9oscQw8QmiTxrjVP6f5jlULwOLIvngr3UZH6Zu8aX2BHrx
g8msipNXfpxugYzX4P+hEDGlB164xap8sSOt4oOjy5Q9Dc/yYOGgZo0lDxcjxmjLPsMYfON3CZoX
y4t5SRZHFyENa2Iq1spBeuk2K3jky80BeVg1f3f4/Saq8G2/OqCvwXDhJkagvgVsG5GQGLRbQ87p
VfIzJV1ngJjDq+KgWr6ZRaoaDw9jRi2cQa+SGxAovO9L2oVK+wAW+mdqwb9GtbVJdPzz5xBgV7Y+
f/hLMvvuBhXTEzHcjLSJIvZPrj0dStRfje4vEfKQr1ZZBOBzcUSovaS3XHSEKbfogkN+VJqBI5GH
pfs+O3z20gRyCrzPZgWOZS9nLy3LTRrWVTqm8X4OZ8LGkEHHcGPBGVjj1AdpPvJyyFTRH/RiwmdF
x9hrWYydTk7ynNWT1mPGUDbt6irx7aWvhaJfRbGNBl0wCMA3APbC7OenL1dRF7/4xM4cWxAdZWfp
moWlDLdwmJo+HwhLvu2tJzF4bUoXzbylW+lHcKbW8OVjGe+SSeLuk05lBHBCmHCr4u6weu2jyvEo
+WaYx5H0S8/nE88bIjxhkVWasu//sOWHTsDgSjn2WPGfy8nirWavqOA4xarrBs8BWnvBtdBL1Sdl
99rUM/LtakF6MF20x2HyVE2Lic9BSCQY5nuBfUbE9hYsOfKWzspEWKw3ICClatQDLfH0bFA2jqcK
uVeU0rgRwbMsr4OJd/y2YS0V0qp5JduGKrWBkb0rvbYwp0Q2zFHxBMtAiAESrWgkwMthdIK+cl0Z
t+G3G/aWR9YUvbRprAdOjPyrGMZytdae6663V4PjDUniXd+sq0i5tnusBhZ7Nj4f2mGsRMd0PkAf
lAkbJJwNbuc589ZJUsTRzPSlA7nTWvIxFUvJ6QTJWWv33OBUDl93k0TVQdZMQsbnYMvMkOsRINNg
x3TPBwjekHG339Ysc3AURjBnJMZOzBL4y4f6mbTIjP3S6rJbVzPEFp5wa6Xm4w6vvnhLICbHQmUl
ujtcXlqwHiTdDi2Iwa1QQov2Y1wFME8awu8487U0mE1dMFFnmjKC1p6dWuuok+aJ7G2uBYTcBcFV
wPMZvoKQj8fqPSyhEftl4na/V4F5mz24Vjd6sZDGluZ+zLOK1wPQ5LNxGMajZRLeObYbyNZonpIO
GXE1ZQqArKjeJSR5q34WivjrgaaopaxJSWk24h3jFgXjX/Qe1K+KOVmgnXm1lVCopF39cNjy6alg
wPNWc3oT7c8aHenWfnSWjpkSGUryztnKqfEalsk7GOl9RHahJR/RdcLa77phNnSt88E1YbuHwW6/
9OA/u9Ab2/cV3DB0hodMgQca/nPtwZ//Aka6p+SvMlnyN7GzrAmurFND9wmcwemrDzbqg6WZUVpo
kNSp6qB70yyvVnoprd9o5K4/SV1AL+srKJnb0Oj/bDF8kJqsu5JvZ9ppB1vtprsBwmmc0oewofXZ
RAv4GrwkbdjPmMNN8DPWyC+K0IM/IrRhOc+KZhOqlxkAxZJKYEZPluX86DvRqzePmQ1+iug6rm4j
iZErvl8MBRU/m7oQWRFPzb4HK5XMNJe2Q1SEZbUux3/L+Kit5nTPMwjdPUsvD/SuiBpU44KTiTP1
o0kZwPndpzzlKPJAQXlYCw45Wy0n9ZTABXxWvxW6rOV2LPePf4MAUOPtHCYqjgGlTFRAwYHM8f6j
kkvys6xkqMXb8aXFBg5sESt+RAbPeO4YORjgrm7bbW4+pcPSkRA3HVk/6KC821/hiAatlFwUfOGW
UKmXZ0KJyjh0Q6n7lJiGEranJh9G+cw7KCZh78G9aKTseEZKu1v1BjbpHa490AaEDEpuYQW+3ZPN
/XMlWyyA4K9gUeYvD3/w/cNJOFNJSIuFHWgM6JePbEtBcUqDrjTslR4j+VjrI4SUoUQUPrNZ/PpZ
eFhhq8esaxEIqefe1W3TQhDRxsCL20QVzS8/bl5YE6UMUQuQmu2zJ2bIlOXu9fyQ+nRxYR/b2X0X
m8Os+I53uCTQQCED2afZUmtmANCtBhAetVpSqXtk3Ens2X/dfxlBp1KdjRfp99EWxUhWXEj8iNg1
Pc1ixLNErYOFik7dryHsYr83TeO8gTXPUqRMc/NuuPd5XidQTtBmPuhWeiasGAbj7KndzBvxM3xv
1x7AjfZg1Xv7684af8mnm8Tm8AJrUZ/1N5c8jKA8AtU/s4DYf6u9slzEwmT0D8v1SQpHJq8P6AFa
fuetMjdRDOqDs27HVlUUufwZwZP9I7gUwN3J40cs4QmEX0FQiOXTjqzXDO67Et8DiBH9tZmw/ZrS
EW+7t64dprvf/GS4Iw1ogxAlEaJmKsWkhVep6Bel/WRUgvdonjGk0+rRaFM2rbJ0eMTyvB3aNhOK
Gsr3qGet85jQGKSCWSjlGJ09qgGBURUXjIbH9Gv+IMX6RyBNj4+Fs6A8dqVjYQmaHKPjUJ4hM0Eu
uI2nlUszqe0MoXiDAOO5QneMaY8pleVYgDCiPNl0PNvlxn/qC6QcSWu3dc0GmUbS2loYWtGC6Pv7
caKRtXVVKOw498dUKJ0d6ZyEPjPlISNjVMUoA+dVC1PKN2H3SJJ/juOCijOqi8Hi/dQP6idmsY0y
r2RHv+UdVqvYd9k1d9g8eu0YfNqIseUnT2YhAN7cGK3aILEKY1kbGS2UUWasl/1BDuMiL23qboqE
UBzewBN1XZxROreGV8VUukuAYzPgujZvLGZm5Ohpc4vIVnLoYtoEolF7wAEi7Pop6LMr8jyG+Esj
AuJpNq/DZ2pvXd47j6njO7BZOrqTtR9aww6cjkOV4DoZ4rGrRvkj6hOs7JGz5c1hQMniQXA7ivLg
0E5uDuVa9nCuXfLgimdsvPLYcArQWCbJ0FFR5zXCcCRtGInGSc1nuuPAq31nG82ynkfvNHN8QW4+
zWMD1qAMC9XXiY3bDsbQ50RABCwwW1pWt6dNGmB2tdhQ5WPxWPahigZBcxbcl8beBT7s6pw6JEC5
X8TC4QCoHUVn9i3kFW3gblHFmfs/bSqeHLHgm4hA3k4Nud9sgEsreTUdXYJdc3cQt/FEuK7Bwqx7
nrNkUdepe4JbSJ/woaKOjZ9k0o7/VESa0IUPR1Qp7DSVOd1LIxHy3a9YLTZt/e0O4J891ydO4Eeu
eOe74fq4AzDY4Xpdx1XVloo+hW/Lrzrew7lM+crsFScRBssRxMyCFq9t5RizvrhRlEgFSdLVI3iJ
HvxDHypK0HrHplDE9BhfgKOVuYyWaJoWvOYRdee1f7itKuNCjzBpamVq9GkF1pU1VVpKnipxgtLC
JQR47gS8Oz4yV4k2/JHjdOBX7MpVzbPqxiB5SLoepiXDMLo22l963eF3M+f4YSL4w9g3FvfILg2B
nI8AXrvxD/WJ9p8ikLB2EFaud1/UL8wLJdBT7mp6/zY/a9zrjbIxq2POQnjOkc8QwZ9ZIziHbTme
1YrJBAyBhNx5d7oJ0SbNQERsyURDGGX+CVEwFzptHmBfCNemOYYYwprRlYKlNl3XD5n5RlsGUE6v
qurUx4Xx1F7eP71m0y3u4lcj4eRgGRBGHFJcnjQzPRlZqemYmA8JwQ6JuyA4xhC21OKeDy+Nzi5a
pGk0DCA/in3unrNIY26iUKIePgQbyhe2P4g54JGtZXstNVxHXHs6vpBEu5dZsQ1uZw0ovhjXBOfj
Mo8HaZycz/QOsMBiE/S2oxfWC0PTNylrE0Eotj1AFvhv5UkAb4LuYRqzySkWChkfaEFomElvVGG5
fcU4vTUzEE8Ik4+GSkoIDOs4C4jklR5vzcUUkz3j4eH/q8bSHd8gZplMTQHF/QtZH+qQLPGCdOCB
QGGXxj+icRLpyZXL4o6QewSFKl4azUjQ2MTI1g8KVLHBmUqicaAtoX72dBoK6xcKNxnsnFp28TUL
acl4SYzFH9R5C1ivWOsanhOacfLtusC4ZjEgFvABweSm9X0+nMoyxPPlVOGtXBajxfenYONMYahm
Y9MCnHHYsODGCEJIlg7Y3MqL6S/u0MUVe/DU0pZ0hQQvk7vn/EU+eEjEaaywp0okMIt3yb5IrRzW
YWt266kTdyX9LSUYODSmnj2mcDYJxqjUZKzVAwD5KeUcNcTPzFaBqDzy06aTrjrpJd28wJpZLk4Y
+X3sfPmKrXYM7RVcDQ9JBLDLcSnOp5P5UwiY3wrB8sn7a7A/jUkZAUuoHQ8F17bGjldwQdUn6Arn
FERkQoV8aytTOT92yAuPURBPnqEZGb5gmCnxBbV9XN8Cs7krFkV6Q6cfbi3G2Kkq+Pv5lM/FjHfT
PL35mWGhnoLrxVEezyr7DZBZddTMnYz38WPy8O7//6KQ1ihN5Gml+RxpXE4tVqHwk0g/jUfDk104
5+HnBaAc59NVWuy+9kxv3xCC/mrVV+IXQvt6JUso+dM2hN1suLJZTYU9ccPrh0zMIzkFnLWIn8+T
nr9d8gn3/D92QKdvRDwM7ieoSmljF00n7+loC05pPXWglA3BWnYGzJGlA7yrU1Qs0PhBMRi7NZtK
Pw0Qy+pn7Xff/tHynoFaXGEi6QVSka3uRlEA+ZQiWb+GhnQqBljyj9dweNhjLiWX1v9w7DZw+l0A
AyIYjKfcCbrBA56rjS5HfOaQJE/FnAFNWnXAvrnjh9W/jCvyqfNRu7MhQ+Ok7Ru9pEPUw8V5+2dS
kPQx0BM2fSHSGjPsRZLmxuiG6eMWA1gopQINY8s2JMMybc9lZAY37lwcirz0fonvsdYdinhfaycF
TXCVBPFB1Ci41yqz2YYXj5GU1aKcljk1j5FQHnEHMCIA0D64x23B2UsihKr48OBGJZ/pI8lwgloB
aoojJsFCDM17w6PKfib8XzbEuv/MDn7QZ5/cGSGgxR8HTq2Xtz/pqX66yeqmIoyk3dZ3v10OiqW8
f6Bnf/B+wqa1nl1gSXURI22Tz7At+mxye4ZMS35lO2HxyOVQsL5cFzW954ns0GiYaHkKedJ4sTV5
3H0Z4FBygKox159TbGJ/CRbhTmBChAV3h8vmNKdMP+KjXLgpsQfkDegoSTF+XmWsbQy7juvhX0x8
btzU84rHDKLwocKAnZwZk8zMAh8w7GqU8fNmhwrxts2/K0RsLAUnKQg2OwP95HhA6fPzdgzxtwKE
cju/NkVxgFsHx1YHA/u6laUgDKv5aRzr80B8XhXHtiLmX1GzcMg7JyrItIits8nZmmBDUxX5UIHL
WU3HGWDFXMWLpGXcqrg/VJoaowVMVm2wvmFNxVsuV2XLHLuo1DUFGTapD+rYHlDCwf2vkiH6riSW
e6yTb5aA4VTU1W8iRNcccNFk7ZdUeXLXGnG/3XwQ0e2hjUV5jNhOWaduemZOEQRzgjJD0S+xCHxT
n6e5Ag4ORBuW0EcZLFP0Bu5W/W4b2yNfi753T+4rfUx75fTF+Y4w3fhhMo0iRU33FXstk+IEKr26
aZQkxaGAlTvKwcKhrYlLYKxagwE1aMbLzjaOcWZ/sIrZzRmJWvhjtalrLRF0l+p+4ecvnegeOeZz
ZyNAAdvOJjnfPx2xYYIxqooB49KqpZRfokyfZMvje25Mn5PXKmyIsAzQXaHDun1cjJ8dDva+6geI
3SXDL25gnwOUjMAAMtYuN6p0gEk1gNEgU2IYkbu8s5SIChOU83ecminXfI8rf9bzGswB8T1Qe788
UivR5hJ3wnQqyaflGe39OvVXcXqivckW6YeQR9ck/IsVLJPHMNZit+C8Io/DDrfRFuqdSyk3xNMf
RVfuxsEoZKzF7ONs7R5rMw4oBOVegJkRhf8Zgf2FhiMLLbaQqfNkntLy+TynFpBiiIP7FbYwEXOL
TH+AKt8EZ1Pf0bWDciD5GR9e0hgEqFb6YJPpt8jZc9pljpQX9sR+NaA1kw2kLu0BAUmYqM2++GrC
aCRsW8uaezoqREUMnuRQMUm5XNus8dfBiy6EH/YQZwBGD7KDq1qvm9nERU6//1GWs3dwdYrs48rA
cnIDJR4NjWIEbi5U9n9zWSHLPiPW6Js4wKMWzoTho2kUjVX3OLy//FWZFSRktTV+m1dNIHtMvN9I
Ev8uQeBPlz2rNMFg+VEh19iij0HBtgI6qC0AZStiFZFycQahmqtHx+FDBc9S7YjSboMj+c3v3dDi
xN2IEv0xQUmYcP3RQEu/1Uxa1b97+P164G/MZ4pxygEyOKet3LRkmvG/k4vf4yfk59Bdh86tpQuF
StDEX3QE42jMAnBzo4AwwdYfq2hdG8ZmgWGdyAqAb6cOjYnotahKpah1SNlxeqCv5G5As04OZp/E
HLsK7MWuqoJpxvi78Z5RBFk4qMEqcqGzeEpRRJLXI34/QuPpfTxt5SnWFfG97X6yArwg5nSiXTqP
Vw0adTKtMigr/1aIIRIlqpMo7KBJ8Nrk3AQ2u1SeQw0oVAItSjL1cjzfy2ajiycFmIu9jyzIVBlU
ney/jH/RmGsQ+BPG4flTcmGmWxvzO2djO8CbwPItb9GntnKmNz/5cQ4fpVDrQb6kJ3yEFAh+mxyu
APFF5ZMjjms768r2BopC3sbrKJNUGXSFloCgrciDoq/sFjb1u09Blu48BDCAukkxdIHVDtHw7381
ghZ0luYgMQVyndI21RCDcXqE7ysOjWeTToBTqHa64ZHl/R+rRHH3gQDz0oTfD5baDN+YiA0XHSgp
gxOr95NmR3RH48RQdryYgnuknPGWRt6NQQRpSTuTPjKIN3wKWRd5twJynrrXaOKa28gosc52qQXn
eYE7u8a9BLop5Az+AhSpxh8ZrGIfcucqCxXATfRyRBjAW9Vv/H0bnoEc37Dq1UEZCv4c0RRfxZ0o
oavuWi0qHsHLiar0QzlBNGHzmE4iGjjYL0CdCpg6TmddAd/JLbtea3a8lVSE6ykBFd5R9SeM+Y7I
gppjwTxBLaGPFNJdVVxHUvBKqaZdhEdbob7XAmxAP3+BYC3W4NBQkKXOuscrgLmU6Ex/vOE89KDe
34OiUH6IkU1si32+wPr5vmjjoo5HMkofO0Ysb9kHXV02P805WYhyoCapQnHuBbb5/aOEB0Upaja3
gQgvUnP++Cb3PcyPu+0UcRYqcjiCESi/7XMMh24S3sVzBTq+yy1OFlD9/WlEI2DczR5L+5JB/DPZ
Zwnsqyk1yqT43rvBaw56q0xLZJOg53AmlhgFrvOTmbVRCRnoFLeFdTkB34PMH0wc4s1GML2UKlgG
GtCyPRT7M3PEZrpCxleX4XL3hU9gW3c8XQcb8EC12Ei/To/5ugpCJwYxHk8i/PjtYsgoXb8eziZc
QgjecEyJ4jXinOCQtE1412fspj72aFSyFxg8sStxgr0JHV9NDrwiVcODbeCqhaAoJ6pjhl/Uq2TG
3MBjcsoDNlfvGG42yC991UQkoh4poTtuf1/114O7i7fGlfPMFGkt/dG1S8VisaWUNuq4nmJY1ZnX
XgsEtqmlMJwUpmoqAwQ2TuRUMaNOnle6IZTK7PnbDK1lNnJ5fNXe2qaPqlWInG5MiLn8LyDiH1Ah
ZojAa0J4KiUu4TNi/BE8yVjoguweEwdMZeLYS6+N6NrPY2DYk+VLZcgHko+AgGkz2g89jaFZ5o6B
Sj7rvccJPEMuBkfdFfcWswrkV+rQk5MvHWFkPxgUtsTjPcRfKf2osCZncKRCRdYZca2hajWvQqnJ
pbTdPHS6XAjWGrXhhZTLXe8F8kzQJ06FfYYhWFOlZzaEFkuyLMeD3Upgf4iGpz8MmyoTXpJKXhKV
p+2q/dhZ66diN6FXOMuspCIH7hlHAqmXOllNJF0XtpG1YaXhuVl10mDNtRzkyp70fnfjW5RAGQD8
i5txVs2bcgPQqSDFjmop8bjcRxMyQ2Ar0UDufkCXkarE6rkHycgnNj7WSZKkfyB1+FFff9qz4eVD
HkUimMuAmaRAz/F30ZYwlZf0UKO5bpuEnuwLYMnQk0WiF/0mgQXE2/1jZNvB/irA2bm4CO/sqyZr
MUhaRBIkmZsU+dsgqcq2XptIXaHCqwZUZ0jy98a1rcScEN6ME15xnokb8Cv4bl94C+vIYyJIKuPV
BrYLmbrvi4gtqhLc0qn3jQ6pJNhFTFFKvudVY3kPqKrhj9YICgPWl83+5LKEgTNm3GjhkmnP4Tz5
FqeGj1tAHWRu5Olz2hbpp7gFk+2SpXYCwXl7mCVQYvvDyuJGhrDLQPz25A2uD3L8jusRUPEArqb+
eGzplxP1YOVHG7GoLuSMkJAKOidQz8+RJgdSHE2LtlUIlc0GVrJ4T/PrCNA2kvSY3huwGdgJWX+N
5rfMoVVhM8HVg1QekUoS67tG4p+f0+abAn3P/dBlr2cATu+IHKfL/hnZImDzIMZkvZElJcDdGff0
vlbqwVsnkTiSAhyBq6jthLhpnsOlKOqQvI4YEIduqTi2eZR2gP2RFW7+Tl+OLfs14ir2/y4qY9Df
KrcaAbrnBsvdqUr5Pcz1xJjaMSVD9Zi7AtF4A/ckRpqAktfNjnr94ZyVPyTRnuKQQnMpXnel95//
9QZXgOglXAeR4KJYKJ6n/jqSaLYV7NzFkSganGYQ4V5LfCVMPhSjSfEwoWHGLHu+y83E/Fp3cMlR
0WfzY/tPQcLzYXrG3aPgrxtg+7170QRABCrnH17ok9pwROGW1jKd3yUDTjHOPpYwIjzj6jU/csc+
LHv3TKRx5rGgfEiYVqQhDCaN3y2jDSxw470Xbfnl7ntHfO63LGXm52BHMwizS1sawtwIe06WVEBV
3FAcfVXvETkhbPJnKPgvc7Ue4aAHtpqQLHkQ3VYjq3oBThn8wzmHrprgdPTOhzeyqqArXVEfjle2
fS90DClE5yxuv+Clz8ilMXBQfyP8TeCPFDG09IGeDC8rEm3o2ZZ+vigV1bqKJg6LNCuFcbA+6ymm
7LswkXzQ83rGXjn8yWS2uXXPKTgpNZYxmfny+hrjlnpFZqHDHic7tsX0Ih4ibmLw6jQkAC/VPM11
hgy3+Il9o+qUJ8XEh1KEHwvlbt3msMGVb4g44tkvZNEnolbDh3/LhU/ESC8eyeAV4QyQcmKJIwsR
HscaAuMfmu/w/SilMkj/g7XhrbHSynz1OeJ9A7M05CswIWClDiY6IzuM+e+sVn5Jct2hk+ot6Sxi
4zz+UlKZQQ/ynm38dogm+OjG9c1LB9gfCbzzaH7NH7T4RHZmD+/AA4or0Baal8IF0SqjyOkNR3dd
RqSQOriNknhJDb0uvr+eHJmSMjiwyS2IEvlWPmDq6SDZ1wvBDmEBF/WEG05Xrd3Yigah9E4iehLs
FL+v2+Sl+EoSXjoIraXK1RyhL1dcxPp/GUe9bX8QCOt0zT0bZrDfKf1WG8+fnpv9vttt+Wq6VUKa
rMJMBRgGvqYPoe3P2e49CDnAdrqNRjrl6vC3qBNAbeHIStGX4RMfv77PXNuxruxcV30fWPYVPwnr
hiqsK4YQzpyK8KWHiuzWMPRkMB+ngxKXZmmiIwi36m0dkxTGvT6jDmu8jeTJNj31iZHikxd2Z7mx
bJKbvmBsKShzHDLSGadK3wxCAZXpvAZcRYM/AvRHlDXcFtFvSmQJuQ5xsyldAmqMNeVYpiHIREVU
c0v6WUwoI2n8iXyQt3qsiarWSf6M30XjWDrftEXzCfrm4yQmSw9+gua/E210NNMGCs1DFDk6KWbm
WYl/jaSU7t0LRQC7wsd0FlpS0Yki/o5gzNsrB2TfQOI2gRygbavGI/r/K9+OQ7ELTyzmdMoG8jzo
/iYzzZ/4Nlh9ShfoZwYU18LFVT/Tq4nUOkRzoQRxUII3vG8xbNivyKqTR7cmSdJP4jQTdu304nn3
xC02lsineiovBIy3bSC60982zwJxzh0aX04G6Zyo9KxeOp6odgoala1bCJsg3jUcla7G9KW/AVKW
iv2WHuhvpcerN03AyJNxrUZyXhEXBOnGp7MBhCQuKycqoYIkhfBqmk3w/T3TkLuvaQnfQRvlo2j/
2IwOFG9zz8qizjM8iigzPuBUeSN7qOiaIDQAK44edIr2hp4HGSmrhZxnllLYrnUC/qwnrDCFlU6y
hTLZftM5O7DK6l5vQWubKvSZYgwgGaPNx+2iiL5A3R6G3QVc7OXkyafwCVyZc1KjjQoc7ANJDcs8
t30QcX83t2v5HhWkEL1UXD1TU6DaMvSMl4UWTQLJT3ta3lPKFGOUT4zhXooxizY2d3+T3SN+sjPV
eXSrJcKgOUPZ0ZiVhFDV+TOKDt2u6ICcBMJCJsRc4PEWCCp8mVBS6C3uC1Mc2DmjoFSiz0uLCRC5
uUr7uYBDqvZCq0TGmczeR9KM/upXbTakOq454oF8i5xBtX7FgOiF4xDyZcYPpOTJEshgCD4wbv03
vxvdzRiakLDX1cC9sN7CuOyexCGAFtkQth9a5/qp/XbIjDrmZA6feoZcghCKRcwcAqoVVh4drUDV
Z2hHe6oLi2MKSYCUiDG/nK8xY9glsDdvECA5c2DULmMRFYojxnkLMyGj8c9OYHhLIxqa27aI3yD5
9iP1pa/ASXVT3sVIPks+iZ9fED9CRx2+GnF76Z9v9QeTksIuNTvbHqyjqEb7uUeTedIJ27TR4gb6
AXAESbVdx7nK3YaGj22txXpbEbSlMHjW5iR9UrXSt2nMOn7/iMW9PsMctM/6ctpNy7mD+0aGBTso
07/zMsW+dD8fTUrrZz7qGyujA+HieajaMBic9dprG6eVOTrYlpW54mAW8j+3NqKsqzKmBrxhDCkP
41Vx7p707ZRD8x+RniWlcQ6AbYH07QXUviL5QqsfB3AqN6VASerHu7xdu3KMCKOtCeUEmd9uZoiZ
AnUNaG4WctFoMfs0E6Kd8F2Ar7UrvHM2uugbMwX+7m+vy/iLFFDTjEuxK7kqoquys6ZHztfL7wWC
HzDhwIp7HXckPiU9BH6miwjzFsF2Wo4byTaqt1zeKJmQzkNN/Dv9GzLA3EVBrctH8B7NRsa3DS1Y
q5F3pAMIsU4J7YyEvqRAjCMsMnDbTKFz1VcZ663TnecOiVG/dlpwFx5btALDUoDlfm6ex5WS963F
OUhhe+HVOHO8BRWmqmol5o8JKQvEo8yqYsoujxs6R/LdJYlCxPhbycnlNiM10jUICdvnRtonw9h5
+/WDEAAF4anGKVOJwGUMGQTAihvzLRhSlqsBWGeLOqL0s4r83vFG5NyCn6uDoUo/SD2EIi2LxSYc
pZGgHCkgQjU11nkxm8k2tgQMlJEPAabLR8bp/KUGliYyBDU6ePRyaHYgKIPez0uZxvfLIKZXjRhf
OSLpcBXoL/yQYMd42bYPKpqTw7mpa0/f9tx7k6W1rNr0c0uCKx4Q1byscCb+zJyp+FRJ4g9Ox9jR
iapnk9qHt7RiSS3AvaTDuIWPvH0ozB4tvuqshh5yFzn839pnyVaGy+7b+uwgxzphyduYGI7wvrs5
fGTPXFnX5x23B9YL5E+KUDCauAkBIdgLorMpIyOPdJmiG4oTzjJfcLdSu+Dhf79XzdsTgVjgLZaE
XuZ5YeN87ACJBnmX3i7APD9LuM7EQzIy/Cf1BBI/5p1oua+DY5V8dLnfjQ3Lf6nxpp1ZtbToZ68h
xP5CvirApocVz/ZM6dI4KyX9PPwT5jssk+h/SJw8qocuFPBdHpDnfqqyOGVCeODcWCZmoLKrEtqm
cBk8pBmHapouo6hAcrQRt+ocyvkcMsj1J15rwMxssBat05GdvX2DuJ32q6ucCg5iWTbfW7reBf1A
SRTxYktVpPyG4nQ8CXM46cOqyoxPEjQjsUKuI1ECwuVF6NV0rsn7ohSoqFWR12QscHtLq/P9hBah
SvDEhu+jv6YqO7Kng6LHQMNLbjA54aFrZ2NwdTV1cfOQ1ZWiF/WAi2PfOWWS3KcJgglYynDMspry
VTI67R2u/lOW5woPqxM8Cabr2V9Mmy/M1G/sAMrezA7O4R74NpM1/lE/cliuBcH/a23ACgCXskDa
LC6xV/b+pSWWGZqpzFbMBCeGrWo7FU6B4D21Ure7ScieeXzPM3DyYKdLjfodgDQFyn13SRnDfwSJ
wWaoPuoH1zHJTsmk2LimFrdZRqNwnKen6Cjr9TtfPkwSNEliI8Iv9+7EFMFWQweR0vqRjcRnNiKq
eRZmHViGDMgOUSxZ/HrmASjr+Zv0uQiHZ2i2LbmJm3IQdqajzHanvBLzCRFJSklba78yZCDdR8Yv
tSsmkJizGXjq3e0aNBYcO9mQpdPnLBWeTYt7g3vFrOdkGyhH1hc7fC0r83q295eexFvVBekop5Sp
oSCpd4u2I+VQJWNu285K62HugDVMXQSd87QK9Mf0lv5sw1cjtUZZx3yEWtLX1dJu1dGRojFXpXDG
WHEYBGksc+KoLpAfHLvXHF4Igc42g3Un5CIjTqauhGRf1NoxTx8axZNU5Plwceh4C4gCOUSS9IHU
3hrluwGoj8UKAXmkycpAf8ytGigr9lrZHpNbySiOmghqmlrUPYrCBS522GsYk4C80i6F7xggXwMJ
q0aSLWsnChVfmfzkOVrutq9qIKBJuaoITOud1AVd6n33DC4sRUrpMPjmbvfBohbpR283Pvfz72Js
aT4GAPribRO6qPBjn6gf8Ru2SzT4rSJOx7nEZBQEsCGMnT40q97NlwGKbfQm4HHTuXzhPVXY2J2R
oosaF6QdVLmr+QInQdcDdNMEv9wq85iNzRXyzM41VE4XvMfV1TcynSSDRaZoC3WvayYcojXd47wB
329Z3g5R9v4u08OYVrbNK4WtGfKET/O8DJH+RjnJwudNeLK0aKrogUGU3wCpxCQXBql9v/MuVnep
S+l2xJ1TGK1xhxeSpSXsaFFjlEe6YtUPRuMW4f/u2WLslEIg5WFZZrQPQIB6NE2jDPFIUK4UE6qn
unoC1lLocAXxArFz+QtQFP9VNrkcc6SBGZOJ3VjUKff5py42SvcmommHcnU/TLykqxO/TKVn32wN
USaSOZhTGuBgEksY+xdL5EeEXOg8XMAuGf4HpIExQ1ef8RxQdHgEMni8T2MH4/Kw2N95T6nT+e/4
ohOk3VIzLGhgNilJo70chRfKeqRLM1XuPkfwHHUspZ/Fs30Ig+kDLKnwVDgHUTJ/j21/UqULx7fQ
74Ze664CSfl4Y0ok99vSUGSXbXwxnJ5FAfRGLDPaQNW5s1ik0r6aJs/P1cifzmzmjRFlpTyJHwec
34iPrzhE6hGUXz6pPFmxtF8C1tXjgwDOJfsqPg7d7WNIdqNpMZCc/CqsXpws1QQZ7XsTG1yZWv5Y
bbcekamqUJvU8sWzFdWUN472jth/GSQGWpr0O9nLJeWVTFwhoJCutm6xEBbE/lYGjcixHNCk2Ep4
qSJfK4m2xEYF4BgViVNNuhe1J0YytazAnVy5cFfCd+XK/YA9btmCOodZ52gZBWxF3occc3LgkXu9
uIbnK+7QVGtyOgTh7iKgoIFCXX3kK7QWNn3BU/Dq2zrGKiS6z3b0Fr+17PuCHEwhoM0wwXIGahDM
8DeRYBVhgyIkQv6AVTSnyNBbviM3XnIrAFWUD/MaaM2Wm6tT1st+VUcb6p/a7/mtmzinNeyaYMe/
Z6FQjOzi7wVDFR+BniMKSsYuk6nfRgKcknOXL1x76CXLfzh91ixiaGR69rDTI73taS3jy2YzAqpi
zE3QtNpb+hAR8hvtbV2hmaSBmLF/KXjchGiqJiSdbJEvmhdBQgx1wh80vqM90a5s7cXtV2wWnIrH
X558SO7Qv3BbWnzVHrv+olEYKEPU5L584D8GteJhVqMgYyGqL1JHBWVLmiW0l5986eXKdKOCAPEa
50PGXc5uKQF5G4LiORHCIqsVTJKbgTPcqpQosEfNm6WbhB71svWA1NrjR1PgUENjV2Z4YnIScSH2
ZduOUNdIrrhlpqizoij79RheBCQy63asOtQ/uD9Yv90zRE2pJP0RNO5wqk0tvFxC3okK/LpOMzFs
fWuiEd3QTI9nRexGqa+FNHg2WCpwQvmE6jOKgPoNvvVdu+TvFYcO2sDcePZj+oHGj4YnmE7OfHIa
bVWj/jj+mGKtydD192J1OG5bZQG3r/Es0vJNc4pnbJBqciTRnq0tFkcGJDI0OpPfNeYBnMDBagmT
GVCCuUptwGW+xTBJniZq1EvYrlWn2AiHIA3drt7Vkol9hNdUZQbRvisdIo8w8g6QCWXlF0354ZjK
9nCyw/JIfQLw/o9uTJBglJg/PlOM9mI+9IaOT3rx874jcod/3Zhcqln1KeQZvodfcBvr+TAQEqmT
AZLjbPfreYk5wi/3fPXxzrwSRytOYwIJA3B155ioVn0pOB7kv3dnT312guUFNBjhTBTWDrOeLOq8
UumfPVSKeGCdyOJV7KsYb11MvOK2EpnqVgN8i7vPiNYn/KdNWV3sUFNog6lj3b73IYz2nCJK7eYo
bsQqnt/t2JDvKx/cu3JAQj/scCHZpPt3Mfnf+njSehl4NiO+nWmY4qmmWci2YxuAsjUNj8vVgMNe
y+dnYFfte09fBz/mUU8U8nXeptnMstEnXvIB/S42tFvuAFDojQ1wROJRHL82SYU0u+Vtw6jyy6nP
9eTUh03Yk9s/WwQDEd593+kGOriTkWruvrZibKsgwNUjhOJtCB79wu/GCJRVM07BcudxS5YL7u20
/6wfPtpX7bdjHhBAxvJaqippkNUhHHuUhcgStnCMyhICh5SzH90kMTl8qfDKvHRHje8g1z3OaQTz
pCRVTBB833vYEcBxeW9KJPBS84mLjHTNws6V3qdHLpKIGp8kPYHgo8xEacgOvPqjm5jDcEd7JffV
Gzyn4KDYj7aWw5nD5XZTkUJl0em8fxqNM/VBk4x1uBoxrY87yp1mQUZOizbEveXDuOJ1gXsNDx+z
Q+2KRihwjrIDR/F1FR+1SfJIMCR3QCMul2/FPH467uLWEh5MG7cKrLnlXmbJwdwPVE4NQgh4rMu0
1aKsZ1NRZJw1VDJe+tDa4m2B2+PdwrOjJADRgyZVvfyen4aWWv9hV3nM2xV5mFb2LGs+M89HM9pD
tiS16xh4BJ+ztdVczpIVW96oHkpY7eS0ZVsHdxnS/+Kd9hl9CTAY2Es0Znuq1cDp+BAawkXP8HIM
KneyifCKeNJP+JklES5LwZI1lVB21u0c/FMctzMbNejaE//ZThqMjaqYxKOuvCloJ3jt178RysDy
JRgRAcn7skRtVcbre7pQDQ07Vw/PXHXyeyin/MCMqTDiBgh/xdimE9igYM89+k33+eydz2jKYZ7y
GtxAP/u6vVT43syp8jaxhXY9G3wP3NYQBd7SX7SpTgFw+8HqpnWMrMwCWPBnD3EcOeZHr5DQyGT3
lpGZkqX66xlQNLgVYO7DiafWQTMf63cAkuP/65oiMuUjWgLI+FxVDt0IXX76siuJsQJ1COBBw/jN
Degv4zhqDGREEGPjGNp2vSAjIBO6J9GKS5NqzV60LpTrjkBcpMNqt2hctNE8qXyXH9XYDJcARl6l
sq5gPlSdZZMu3tKOHyyw6Z+L4mdW1+LeX9/oPsLQNO1DH/iyPWtml+4jhUxWwzPSgXjNF3ZkimaI
kRRBWU9/8X4sGGkDBYqbwtxm/u9SMQLtz9rIHWZMISTAwz8Xi2g5J872EbwFqty8RfWYUTHp1l3M
IZ/LtrRF9M/8ZfF3TTCYYMUbMNdt8PO2UA3Ujxnes+rBR4a+Q5LNcXGyJuyS2IB0Be3RQ1jzZY0Z
9pJ7cfrRASqF12NVHjgRN1ZJChfco+pH4awkS7zf6YcHDOCJV9sTI4ER9V73zoUBZn0E82iZXetu
wVfecoIoNFr/7iG5RTVkvPbSuzaResiDthK13nr/LzI/tTa9KNpIbz7sHZZreHOIa4OqC1g5TE5O
eL83WDwGMCqa9rix4Ohm5vTbsahFpxdN9WjexWGw509BDXFphFWxOs+Ro1Y1s3C3v+rGofrtJPoJ
W/d7WvoEcv1KlQm3H9w6GIm22HdzrPwRJBmxGjRjig41dRk/G8u6hNRjWkdkIDVGr8Z9uKpHgOwJ
jAIk9plaCrL0XKvktDbeZMPHvfqDQdJ6bxmDgh8pIrrEX1PGAqaqowym0HgcR/y+wyUFy4Mrx+sb
dyBm2sJKE8K7L8Y/JATn00qLHmMwY9H2RJD23aNOZqa9XVS2CgxiMm6N5nQnFgY6nPVUUM7Xja75
JUQHRynTstlTKlgKNN+OSzmgW6oiLlxvEFiOd0D4dARLdiAdprdeWzR8zYUGGXYcZZhyMTlROQca
blh4Xh8GYKaO4JLg94jmT02Fa0vWYUO5vcijSSF6KTnn8OtCChr0T8HHNz7LA8YnKQM6SzQFdI5V
S1pc6tcxunJbF88qZVsn1gaczU52t1TqSBNpLMJniC4Ot4LDcPaXIcKyi6i/iOT4RYMaQZ1ZEUYa
W/oGNWGSDzt72eBrJ6bwJOuaP173/vb5wquKzdL6c2RJLIA03jCEcU/dYfZw/oBI6O99WcDKr1rB
ia730Caxz0zTHL/IYbZ/d78UHlaz5BlvO4OUf/33qVE+WjtBakg/2OMqgyTSRu6lB9f9IivN0GDD
4zJ4TPYaOJMnqThgyLonnOhqewybcLdpF0N/LWKQhp5qr4F8cbxLy3bVSLrAo2H00BaLzYrIO0gd
745f33/xoVIYjw4YmRHVcg3nJovZ0yAVjFRvYqhTCEq4th0XGJCh4VGUqMnDl18GL564+kdejK5D
hd0g1LEOHZP0wI+dDqhN5ovuzFbTSdgcmSAENAbcNwlp4LieSCLNx8azKw4D52pDHrKh02YveJqi
aF9jA304R02CcaZcx7n1ZpeM9eymrTM1FO4jSNYHpS/H24hTA8QIy+7eyTZJAZSQtvlRWdevtJT9
J6rxpcD0D0+wq3xEhpq3/kRLtx8eBzuQjHgCX3vYacvlZn5pyLSIJSrrCmahq615HkvvDL/o8lvO
d/x2QCc0Ennagt5lY1SQrnlz0arXRT5nVfCZ2xiEMTEQIFaWnETLGu+F6g+7fosAoP3I0aVOjRPB
Ta2wwq9ec6tU/efysEVsWlZndEddZHYxwjgXlZ0mPqFPCYT8ZA5sTDBuwNYfL2qtDnJu2cO7dD+3
Jkggrt/rVJaZQLeLITd10KDXFi60bLcpL6kbsvKthBpn2U8SU6joymFJjarcClKS8wnkfdLOG1QC
ObpAYYKmxNujmHo6HqfQW7EiTRbvZXJcg4u95eXVlcv6v+UAG1UXItkDAnwhfUsEa6UKge0VkWhT
LSOUCv4V4Q5Qtj3rDj+EJDR19UZobilXCM6eBqevbE/noaopdxYjjDQJ/tS6HoCEAZDZw8nlJUuf
THoAf7NGyIf+Oxp5SeN0LTaxlwnKdG/GrxSWZxtHOhM1//iXPWjf74CuPLSN80ZfhqWMdqtcp5Lj
z+6/nCUcmWHUX4nkz84+abHyPpjQFfugI/TtW252Db4T+04KafoWpKMgW8WjmlNNC2bs2HQqMTuN
t9IxrvdcncX09dRr5Jg+np7lJ5bF4jqHL7vKIgtRiEGDfT4yzlgwVf2d/d2336iWtIc/pfOb36po
syOb/Vp9/vp+DQWcUbiKe53RLQpo0aDgvEdnvGP0LIMj4RG2El8manddb8L7iR9m7IQzlcj7NcEC
EX60uWWcS97jzQKcAgpcNRhlITPS4uYOIT88rZ3pN9l62SdquBPOoeTuW5j82P1j5d0yf1VTOs3V
tFpGTT6Ut2aPesJw+8yo40i08T2Db0BwuZiW86wyuz7eggY+OEZVx+Nrv4lvCALV2GLS8RsN44D9
ZgXbmGB4WvIgc7fgSkzeyTd7rTZOw1wErjOxtzfjhl3j/Xj3/G/dE6FMrl5dmQI6Kv5rBBZfPiOE
S8SadC+af8WSgRwxts2khfFImQtEGURwIFfBEfSkeTKTDikypX4BOzcAcIxdgGbHJyzX5UT6W7zP
8bVWDgYIf60vFpyOStWFBFzNIbTXv5WsZLHZ89m83PlrfVPiVWb0LMKlWZLxgA/5tpIDrKwyAFbF
bPlvJAj5ItftE42hv9I34q1nV0jhyJeMPu4/gy+sR7UxdT35UbRlfHGQcXbWtIfMteq3dkK096Qy
5UkaG7fYFSw06Vud30+XzVDjfM9aUHOzyoroTcGc2J3s6kauNPVkgoI9Ixc5Dk+CIhReAwgO4tRw
wsZol06pB0FMySMM3MvLl8+Ajc9/JtUviWLm0IPV9u/FGaKbv5nlVP5O52P6UoTYi2QpuhuMaXIF
YjC/7x9El0TTLgUvI43S6gmwQ+9ldKoRgidN4/eH5c5CqD79qfJiN6RfMPO6QIngW6c2ETPmAfBh
bI7q15NTj3yicenzcUbLpGgMNgW1t1NKmqPXaHp9WTwezAhn6hXaoVfDzFTnra022PTcH+lwExlQ
v2Ctbk7BHmEkkVzVN4tbAe2Y69aioKnCGmcMFfJtGh+jWgs9CC37f1XDuBXadaePpXDXThTJdVdc
coVryL8KSCmKnKCFsXw76FMQNQpT3UUo0+cIFjKMBcn9W3FoMszfuW4vLUoFOdbOT4JsF5UJlEpJ
Zcf25pGo/gdQuQTjzWjj/xBcIGkWAkcUR1IUXa2wrE0etiHLK2Iqp9U3nIfLNWg9FHhR7aqrBeLq
Zi9lch/gLmlAr1/yAJG4oYFxjKJkxj/UOT/FZJmxo9n97O8q6Tnc07aSkKPNj+YyMPOazJ1EazpM
kcKd37GQlPeKKncxq8Hpmt0+VF5oeVYZzbXjfRo2TAG/NnXREDP+9MyHbAYXYndE0/HihJbjObH8
OshTvdiXm1Mvpf775XYWU31O9T5NqeFkhKbiRj6tbwe3VvXr53cw/t9ByAqCGNM7I3R0/GBl7yOO
N7ere8rlHLl/JjV4g4VZe/3TvZ0o+i+8nGNmVGqIqTKvlUwCeWCs4l2dQelMunxscsqUZGE2TQKw
3ed6NX15sy6ITbAzOk1sHg4lH7fQpdDVoj3Iy0iVYpOzfkvwznfVfrAMEtEK/+enV7u9ot5QH+wt
xF8EDfgXDCvktaNESu9TD2lhi0XDrYHFWAP4LJws9Sh8axutyPBiLghvYA7vGdRmuhzWNSEzb+m/
m1r6L0DCXn50Bll47FAShT/Sqb9TCEbffy9MfsZD9AqWR6zJaGSwIR6g0ayzJ6MM+XSRfyDeal2z
iWiIqjqPK6aWNoiEowacx3rJOxE6JCYLngg8RgXg/blycx2pbmeMfy8+lQT3q3UPoukanGov/ZQl
SMcWrZNyuHmwHUxQsjKH0cMEbyg4kstnvfe7gpBB3DJuTkqFGtS5gaABHzZY8QxVl/OgEi2w4VRO
k+dutM+u8MW14o/21QuaiwEyx4QowEhzi6Fp9KkSHrZs0koVX6kCRpfJyMw/j7UgFXlFPpQH2nFt
esJYl1DglmnNXdjNf28wXoPXEqa9LJRxBSdXfXzxlzcBNgtSR99AW0oaQrt2DZR2b1qjGMXF1PsK
oReJFSkx6V/u5L4kSB1Zg35wwrXRWUOrpHloHyRDwtmkndZYxzEIJJ3GsvSbO+MzG+KpP/Gy3UO3
ZxwBfDrW06d4E3YHZ+yi5Cxe18RunyXGGdXxOWeNSSyJG75eIslvIZcFMWMbhXyxi6la10WbvQEL
I9HZRnUpHKXGOUjRyA+lsLS991qafsy1B9J/0Wf7EnBmIQlcxuuofi/yzNpxDkAIKsgUijWYhuIS
XJXOw18AS5oC+EpsSmFWYgl+BRArjhclIzIsuolgQfT2VBGaAjBSHArWDEMkh9EnencDvFp1iAD5
AZre8lEcbB9cKC90v0YpywDQFculLWvNCVoOCamCNJqMq82p+23IBwIRfGLbpT8L0NfaStkpCb7o
1VAhCxwCXvkZGYKrlbDQMWKrB6q6yu72iIp9L6A2PuJrCzJC4vg0pgjwU4QCass6KdxvnO8xa8U/
lrkhB8oR99YQqMjuNSOeK4B5OIHYCY7rj+/mLx0P7PqWZeQk6repMZEJmtMLaxGrRuUTeK5R9YtI
wfSvQwgosMdAZSAbnT2Yd3dYR++iZP3AFhF+Ma6MBjqoaZ+1+GKpYYm+Nmgow9v8j/Qpl0B+JDn6
g85FzzSQskcdmjij8qj/xw64Utw5PCnGcsHf5vCJmCbRfEfgIuD2jIzaR1+cZ3gN761PZsG8NKzK
4E14XKBa14ouoCN4luasLJEfeNoscM1zlMuWf7gdAcYTKJ0EMcya6wxVMhRkX6y6ZqoEJ8k26gl/
8BbbFGtoJCKVgMIGDhdeUxm9qKdQ6sgr21sbg+BrHe7ot+ktX/bUSNCllw60ts5RpArmBk77oYT/
ZlbrVlXI1H2eJ+8d5ySqiWrugyer5f5zwjJuzFsuluvCuAdv9A9AZBSTbUARIPR98bM6VyDCkyHY
boCs3femEE5sGPrKHlsmOGXQWoBzP79eiP+4SaWZbAwvDNwq6EM5ydXUAOEhURGbYnYdZid0Pkzt
z02POfIiIKMTMWoxmIcoodns03FUl1QRZiBfM0UIgtOqhxgEgy0M9eB2HrvN2PgEEutYbZymll+D
2ZgfQq+JYxve8HwLKWxbiZGjV3LGT2x80YW1C+B3orCepHAenJapMbfJfZGCU5MEud44Bddc3Pnr
0SKZYgKGT9NiBv53azMONhf4v3ci/cedoyxfeHDOnrGul/Z2e4GOLyMfZXch/nn1KX9yBspf7JSG
19OccV93RLnPHNXoOuuQsTPdWl47Pt7wQsxIjCxQGVIZbzUdCdAkdx6k7SUc4k2YgGr8uL49VJHY
XW+Qvxy4TZ3TCP6rHIt9oJlFXB+SZ9aszKJGxq6TQyf6+ip9dTRKzkGEOoNcdwJeba0OafH0aNQp
GjiOlqAIynP1uBjyqRfhO/5FmO/L2dtThovxDhSwlgYBR++NJuEAIuqtTkR70F3q2UCKth3wwstM
ti9MUoTtusAI51po3qcN+osxFjls/9cbTzqnSM+JOzkm0XUCFF/2x6pq43/70+IerYp7chqEP29e
WOquN9o93eBwHVMi6LKf8cH5LjMGplkk8gcGaajZwXcivfF0sOXFx0SWSwQrx6dl3fkv89HYMlaK
DvcvVkb0UedHzJHvDpAt3zY3N/RmyPt2GMQ16nplMCVSHwNoaQJwmUbLL4QA712SeCRgcK7MRuRA
3ESrxd34XTv7nmu86Lw6iDxjw2XAfOzNR9PPij82Um9NhtrOjOzwpAIbYeTsjZMZL1vJmfNfNYXA
daHmaE27j6dQnKjyK6K1sKxBStN3DAXBONwcD9okfzuEhB8K3HAG9dDjWAI5ltR2dqff2OIbVEM6
ml6Zov1DP7Q/j3ar+PQU/PwUu+NCgRWUs+YHPlM3uKtxTGC+kcUluHMbVKdGULwhLT2uprjLRBDV
Kqc3hmc05e9reVwDRR+Mhl6xOxL51pSVHZoyA14x2ds7MR01t0zIlGqdPg8z3m6InaDuuGC9aOOg
T+/fUFUdMWyTcWmHbibXZy7bKsRtpKBMSk2XMosUk9KcU5m25IPgGiHehByfZvF3aAJL/04gL3zp
3OjJqd+hcRqWPsVCInbNm73uiwQ+iDmlqiFJnP/uLqNS5xfIaS6x5ZIPe5A5/+DtO4UwHy44eye2
klqc0JhWix/TWWyL2Y7CJmPSbN3p5iWIZT9IfRElMIRjZTzbQdvyASWaobhoxSJbA/six/BmwJVQ
ZZlu2oy0A9pANE3qy66JIjIgxbSlPSprfT5UVPZ7NdJzltF3VtHIMzr5XoROoEI+S4iDIvtlfgKD
xkrH+QLsPKFtic0V1wag6wUbsF4DCSJzeApO+3QwjLMN52mx8NmL5mJtmoKT/AL4E43IasRTAROo
IJgebcKfVmxEaRCsa1QktSC17f9xyLfl518ixp/vwYvdDjIMmJXmH/e+3JzDCrJOyv6pVZbmayc+
ezK6dgy1pMvwooNHwPSjK6rPqLJ6/LjqgcRgNKZCo3EOeOCbysjslcmnJW2kkFxDFkXU8tcbSp4s
QA6w/KPJ0w3mcO5xjKndkxnXJfDEMwZjoLBlFhrowimhxCqAveoe020JI6KD2aNnsN+xYa+W6qHU
ya8oafQT3uKBDUJi72gXphUfcS+594ZxKgXHcLXPq4PNWjatepNtuwkqI0U2jN+jx//U2jve+sgS
ouriG2zSMeKJZbQJ6nzzReXrt+od7T37wVeJmWZZ9fEEae08Eh3+OmBDjoNdww3qIeK+faLGSa/V
v2fg9wdBSBCq0UaU3eOZYnY2IFXE+zf2Rqy22F+ifsDwFtSssCjKMnh3SpuPsy15o+tUMas03hxc
GTaaHEh8vImXftyduW80AAojb3HmTqhO/QNatgGAHd/Zwe/vopgz2S27MhBFNk8Eki4sKe7bo+zK
RBuO48qx5kkbH5LlHggbJA+xwDRVveq4I8E9gckQ4cZZS7lB+d/GDO4YxM44LlnUgLSgLKfQKGL4
g6gen/nZtKSUZkIsTfbkYBHvdqAcSdP2IE0/JZiRRpigLIisu4c/7g2vUCX+H0+wJp5+SDsSuxIE
ijKakQTDP22M8xxyiNxQc19YM5eshBquZOQHZCzPNxZLfs+X8jq1i58hQ7uEX+/VCtq+GJ648KWL
vNM7wPnu2eVcq59SPOjA7sYtoHj1/0Ot6HaPewrW2NKTQxxVOuP5r5F4xuebN6MT1YGFvMclDNQC
fAgJ+0zQ/VOcCU1IUz6YQKMpSQEPhHv7CrmnJabfAtQOUxIyIPqv6qk5Hd5W992otyro1TDwYvv0
ZptBvXjO0lip9Sv9wr5CDCXzFSgP/7REUuXT1udbNU6QrpUhshkaDalIHODsIgHK8p/rA3JgRp9Z
aWsxqjFMld1b20Y5Gzufl1puJmT0HQ6rBLpc1t//LIQ0gSWgXBrcLGNjfb2Zef7kkadq81x2YLZ5
cwe3p4/Od+VXGV6w/7zHRSSPZyvPbJvxa57R00nbYRsHTKV6uC6+qji1t6waOHUvE20Oewq2dGus
MgFjTwyNjG1CmLFPf6WdlWVJXvJJu7ZQcZudq1Ghsho1B/AP81uGPlGg/KTJ312OGbJFj5rBlbqm
8Fn29UIEnFicpWp5Fq6eXRy9JNPdwX5XJPKmHNNYaaO9gpkzLTmvC0zfe1ALlxaFLRcFZf0Vqa3Q
PIqFREGwd9P+ioT+I69zEFL5V1vmMWT3bf7VlQohuY1jNCwOpAZRBxa/YEO28an79Kaj8DYAPmgz
ZQm5bdqToR6+Y7v1QPgJztS1EjWlsXHE+RodZiagytB/joAfW5hC/WxeGDOw9FGnwa2zanT3tkOl
PWANqeR0l0gu6ThW0OBZa39tOFNKei2g+DbZN+STKAJiJEj+lYYcpHV0bqiI5W0KikwPBTk6Gn7i
V194U92HHc2ImG6rMQ8QQtEd3eR3W4ZkGLc7KgIJcnMDnkjBu7aAfDWeTa3Fgv9psX1KGjde4xtb
p3OuLc+rRGG2IzSfAamNj1rLQoPYzuWUEOv2aW4q3B+HsHm2IDlX5tFn2TN7dJzq3l1mo46eD7tO
LLol1hw+mvbAIvINFvAz1xws6QK0xm78WGpfTMpHhh7TlJlhUKsJa/CjdoGcmK+mQapcrauhKb0I
8FUdIUWsmTk/L0WdwDhbZuMNaRKyKpqTsPGttCRbkFK3YaPOK20vmwGp7m1MLj0yP8NH4zEssU6w
SiZOgJJBxYnYxhMsPNjxUGu2ata9T54gUsH599+6fk/Bdn2vKxxaYOLbTwKMNPcx+kf5JZ8bO6iT
mzy5+8DU4TCy20FvrYUbtHJYx1Szaobn0A7PzXj+Trq/YdA50pS/QP95cYH4tWvYAzHQLAfFjp+n
S8I37bZp+m5vU3T8FYDZ6Ldfrpv4BDp8kZmBf7jxlxgqlc0x4OLi8oWevBgMHazB38vqiBZ2fMOp
1NBD82c+O1lPbgh82D7fJ3mTEC8kv3U7HhxI0ShiB84BsBdAE+S0KhCfb6KkdaB0+N23i8TdWALT
xxUYaCpn0AWsywawSwxWWa62Asi/VX12ffez31zvtV69Ju3gKSFfAOSCbA+FOt2nK78mS7hwYtOC
jBT9M3r0eL3JWB3QVn+ewJOs3o4hkoZy3CXS0S9CedQNC1JjtgsvW0MBacgJ8JvW+kps4cwmyhiB
AxdNdEgE9ROVi2wrlz5AkMbbpN4cXPHDV2UMQO24mT5WrwDhhLJG714BU/1w/ChrbPXH7nV0TSJf
jk7kYNTAR7FOiPo9le8HuYs3ySugdGqLJ0cntbMRqI4agB545RBzrjHzCeo/AQJ8f57scaBg3nS4
5AhI22z4mkQsJboElXpIA4G5GW4P6Ohx6KPB0Ht4wbtQOXc7DFuAQuZ+8n/v4NbKdM1DQWYFXZQj
50zQzGG95a9vL5ngWW16ETlsyIuYWysmHBK6GpT9Mmb6Xd2hq/4iNgtAyBlFtaUzpM+11UUMLDzF
hbUsuTomMfwmg6m/jJ7r7vv2MIoqQAL2ekB8bQZIGzU6tEVv8Mp1pMd/BdqlnRmlmE7ZFPY6aRHp
niFE+eQgU/GTLP5Q+Rjv3KNb3KKJ6t5PE2vBY+WkAaTyltFO/4Vz361jZvVrStiZ45lDwtGrEdmv
Vn83aXcomqxyQdOErObz8vf5CMfyYWPJjiFlhtYg8YPPqre1L8kQ/8bSZ613IDVYqs4jeusm/1qF
unBi2NOEnmfMltQDoo58QJiyDrmEzv3e2NzOBeii1ebutNrmx1LI/dvM+gWKQaUafEGmiepOTaIV
QZQ/A7STlcguTZWCLcx0Nqdtn8MByBBE5u+HLC0/xwgA8x5n9J8dPecmr4DN0aIn/JK1FCyA9wHI
yPR8OKVfsGkU51d43xxGyrJPp0mIOQMZUhQ6MFL1o7bL7wbk6B5PYHL5yV/QeRXdWzDDSnnQevvH
0hwgjr7lKa/E0VAVNukx82LlXXqLK7lLU/KX3QoOy7Vp16zPuwiL9PUoWb1YPl+/1ygXZZbSj5nt
o4sbegp62Nb57WSL2fQsDkKABgNvHIeQjkRmNE7KGIeXi9YQ3df4F6WLCRTtZtwu0GOzSS25uSlZ
9OiNEYclSLdsnrS1I5hef0rghfoWULirobFJQYXu7/5456I8ysC7YG+oln9iuPZoPd3NMu3Lf/L2
QaNsI7ssWt/9/EhbZUfHD+TId0AHykh+wiYByK+7pw4etRq7YR45PNtcts83dYdMfaKknRDIDBlu
bxnxVo2biAduzOCIRysQtsIGONCrxga6gXOfp/BCDYURkFzLFUuNioI/hP3Zux7bNkWdWRp/l2iF
WAnjlvmZeIDhJBiflwxQldCwBjiFCMpweRp26w0k43AU6qnP7y+yH3/zRp4Wsw4lUTnuM+uO1FI8
GvA8Z8L3GzikWSo8KHzE29m7L0qT6WIIySzEQ/w//SObm3LOKW/hW2RpXbm5ryuKP2BrhOj+ndZX
vdIwlZwST6g4Y8oMn4sb2csGRJNIzGlxjDZQP7kZvl5iAY/RKtsVhyC8XrZWkojTuARanKSBA+Ds
npIoejHem+O2rRJLOUwW2ia8FM9H7yiE9xdrQs2qwIjYhU1wBAnfqv8gl3LFNtclF7B4GLF7G5PP
kf5CnNlB2Q2qi+wrvgmzGpiZ6NUQNndCGfpd4cB0J7I4pgWIxE5IYWZoln37CTubUzAsMZZb1bkN
md5F9s/+jJMY0SWqP5BTbXMpLgTKKu7+jjYHtk0XWz0c8wqOFEEv5i+JZ210O4/vVwO+y+i383Jy
NMKxXyCmemBemQfjot2uKXAbQI1C3cdW9ZoExCwlLkgLm7Nu59Zqp6Vhz13nCwxnH2qWqoy14i/6
gGkTBzf16UXa8+9//SPaAnc4aJKEWKppFGcTWtO6IwAL13Mum6Lx7qe7fRGAqh6lLAiwzeu32RoM
AZSsQneyAQRHfY42rAg09I+fFDYoEdCPXRJ9xe7SCO9qYgAV4QCwvHn0xXT73cvYTul8MtIkmurT
DHa8OFfFYFiN72zoYwpMHvSpi1RQEvsl+n7cDTHi/gUF5mr5Y2RwshdL0vfBCJqTqHGbCu4FSaQN
rTa/ezdazCnK1khLD+Qf3UbMiBxBwfOnQAAIwk6GQaLgowTnHWosICwE1zH2GO1jlVOW1ORZzbFh
X9E4BLZwPPi/bH9XPHlM07NiFrC0jnyVyjZBtAY60aSoQ11+tUKdx0KSHq6moWb9cd6JCL5/paaK
rAmIBlMXJUtngIpxq3KseBZZQAe9voPlRn2Vv6OW6SDbjj/rIS/PgYzgLFESfPwryvs/BPXrxN5o
pQpe3Drxd7njPxjFAPakoQY6qRGZK6LJLmYBMSBWgRISESAOga+U0xJKI3A+2RcUAO2DVG69DWpt
LNMrf7C+qLV3hKSLo8OnCAS6Gem/n/Rz+gWNs7afOJjfz6j2hiX7z5tNrLTzw3sJ7ncgGAFtYqh3
JOB4SeFGLPzLC+Q5yipl3yVY8vV9RkCdndE6fYR6Lf0ejsXzYtfqTS3LtM6nRIoEqh8FZv0qokq3
Rn36AHf9DwBDYMgju2HTYB2Yf+6B08sduvBRdxenqMsoioUyOEKYE/TZ5n3Azyv4zabiI4JxIsuh
ac9HN03lK0va8sVUOiOFef1C5JHNcSPGvzQkjvXsqsOxSfD1CPh1msJzT8D4IBvi92RonCks1pEX
QhOTnO6XA/VhPHImXoK/8w9jVnGD9MuCYwGKW7qdGqsPYpx4Vb+JYpdWyQjRigfvHZG+QJ52twp4
RiL2jxAtJZFwA/8QZhOeM9E0T3mJ0a4R4GbEBkLCBIPspkBOTgRl4rYTEGy5JbHAgIQXllTs/N0Y
QNMoVWk/RfLzv6RFkTHnQOXisv4WTAtXH3Xt/fXPyb6M7Lf/4CAK9xvNd3uAY0Lcj+u3thsA1HvX
YafvRs1iCLwgMWuJn8WQ+pDho4LDadql083xqv+nA2p6DU/9IhU/DgCU6HjDEBkYP1ByAJuzTOJm
y/DKCuHOgqAlMtZZuhM2e2R0jbwot56DrPwcLGiBnBUwVbk43r/DRcHoz/U9g6yr9sf+9+v12btR
ksxfrAyrn6ghHETGNe0mL/v3B9t2/dszKSP72+if37QPp/wkvdhuMfPz1uVCy3cwE0lNrqL0qIg8
7j2b1byWa0DAa+2y2v6eRXzkpbnWXngiwZVN8o5iWpHnn6XDn7da/eOVXyPmppgdWabdv6ZzfASa
JBkv7FNu6+BDEEfADN9uUjRk/xqFw5oS1kk7M1OWD2nHqmJB2K3hDIxTFaFTH0ecFmwitsp57dJ8
zpdPS4tvuVQeurp0FRskLuv3ErgVdBNlg7zQJNDuaKYFb45/rBadYYPAXMUb3rN9l9oc9AdnES6y
RdBqbtvIQB2ynf4dXqfNOVd2WmrFQt14KRiQ+VIsiH28b6Ow4fU3AzujeIgxcXziednRzthkoDek
w6INqljJOgYJJ5SWkquaUPA8iOW6Dx2yuqc8Rr6MvFIDLEhiZc9d6qnOmhsA3GuEU2lC6d2QIc58
J7yEHJlYSPY5MrtSw6WeRt1Rq24Q7CGcpjel64BRECTOAG73B7vozV1/LOL3puyO1oahg0Wn2O75
BK6sfn+JT+f7HE/hACT4TckWA6cGozfnHkfY7YtojfBPMsV/6JRls7wMlWQj+2s5CsgFxrXgv+BM
grvEciRApuuvLjFVyShqdB6UC0VAvERwb6LT+0pivaBqDwfRNa13lhtE9IXVwb4Y1W8BlMD7p0fn
J39hjcCrg0cdz0xqBKyEhWM0w+lphDuK89LrFFRb63HUkYH9MY4af563nigbtUadmII6qdLsIaHa
kUIRLHScwqgHIWrPJ/NnlXUi/GF0JGVz6wEBTgmtSDINlxGawKNKcj2e5NcS6gQa71aelU35mqL1
W2MuTI5bIfH9pS0j4vb30NG1ohj041TGbOdNivZwmgBBnJLyQ4tuizsyb1ZTQ4C53r9QBISBdJRT
LluuXOu7D22VhxH+BNXfDvLhiPFT/c2wMH6y9AkMuJnIgiLpqj+9SNU9rkSO1Pk3luheFz/+6VNN
cuWI2/rmIUZmQR5sCOiSXsBdil5rlxJvGSzCSyyWIB/CdXXtRfS4UzfNdKsW+1gBkAico3Xb4nth
vOipbGKxtVCyHGcLZxo9yXzBwjCHNkehe6TWypPIitUuu9rwZUiOini0dHKVidXk1Ol/07j5SLJ5
IcG3ji88i7Lib6ZG2lJ5SNcp9l8+IZ/hgeWde9j/09OvKVmkuyVm6dwh2kM2O3ARo9NwG+1udmRK
NRhsPpRVHl+ZsKMFb9H5+8WS8u1R+z2rUmfRLGq/s4pXeAnpupHibtr1+mzy+i+SnldE9Gze0cqA
Ot7EeesYric1LNZEueNxpTo3NiIDqrOGOpHh8kj23IfW54zi5WBxwlltd9uh7qtFZQB9BtkTSbmI
cI33tysYb2mIbKgRfpupEGD7Kk6qEg1wfXOdHQOuEQW9IZMCAWGn0Fqi9wuPJJgv/TfEngcW4/+J
8dXfW4Fy1bEfags8zUiyXbZ/xhLEO34BlbV/ENbJIFfPdFWxSn79OgIj2lcFB0U0Z2IUudxLByAW
Jv1eHIIkDUwto0766gCKRVWQ6mq6vy1JM7cxwBZyLsLGIHx4nrKwMxULHXkiVHJy43gk1lo3evdX
+BRZvW8+HaRqZ/LAMdYxHOPTc84GfAKqYN8O5IaGPT2p5UFL9kNNLvoJi3E8jssOT1AVecZ6zNcK
w5l0Jk4OMf/eLrt5OdOzvRL3AoAIkMSLy4bJzCG6ZV4u0tSYfV9jUo1w93Pg1NSbs5WNmNalpA4K
ykLPHqXcizSquYDjCQpAoKG7PhXiDcudHaOZgKv/QPclYl/B2sO6wDAbD+CU1aXoyOfi/FPSSBzX
tVd8bHz1/YSfiD1biKoebvkfLwdD/v2i/dIyd5udRnZEp4KPe5E9aWZRBM+i7B1YGe/+4AwRm+kc
4sf67/PK2xarUkT6u8TyRCPK4Pzqn0PLkubq/RzWrDJgBvwzlSfy/er1p45vXfgIlC5gq9X0cYAq
pRccTGG44pbFLzj85jc56qkFbybdrl1K137IptPg5/PlvFSkWV01Vc1pTyrA8ApvW20T/OyqreaD
LePBBrodJIxX1vw6dV5x6OpVB1w0Tg9/flIpLr0bd6EXb4wHSr67iANyUbx8kx7IVwX/XvC91R7m
GpuHMEVIJEt+lIlxGlkH11lTlMY4CqC35Mam1JfHfrKGPY7wCGDzIe3jZhHqjSXEa2gXT4zDR7JE
4yasAbXXK6nv5c7y7Jemma0GEUkV5895/N/oY2EEJtXEjWU/1eZm41rhHPRZ2l1sCoxgAYzKpK6I
/i6AjFb0bqUU/Zt1wbEZm9tbQYHFB4ILyytGFOtUL4jfJ4+0ZRUO8tXJjFEb85hFGli7VNfE3lEM
YNlRpyE+gMWnrEiLlT3I+9diLDUgDLiLWV3wC1QndXEUwZCyzg2H2JfvQ4uQI80v02YO45abiJbo
8QX27OSm5Kq1Sp4dRHSLxEqSjvSMYYmB79wzMGElZy9R6tz6dpXGtwO8q+KzimBJceUx2RO1nIv1
LmpytW43Ydjf7qzgAiXAobQCvQeWCKikyv1TaGlAHJ8ugrRALLKXG2cUh4u/bihAUWWtT7eauf0O
SOTlAcFHvyYRqj7XT9oVuKqPdmGfkRwLVnCKrFPVcsbKUdN7VJDbml2PQpGMG/d6NRUWaM94cAE9
dxwzAwcUZuHwZ25smakZSBpWGDQXxiWJ0eVqJdwTvjWHS5vah499QBZ+2qWljpriWMc2sHDBAiKZ
ZWeLNlFBwDSJqExRfgAW/5vbhPd4WgE8Az4EfF9BkKpsUHAsjQVLXXjsZjCb06mLR1mbjhPHdwGd
/flb2ucjnPKP3FyPxR4xEYNCRoYdND/7clJbt0n9iWZHRDftwGKK3Fo6Up/I1RrcIi5wT/AKRIIH
OUj5ibVUc/pxji6y2qq5QupUt2M03TwCP++aW9p2eiwcLxTRJpx31lCw7qQuEgXtiAPX1+dfYa/o
f3akhH3yxSl03H6inq6KeAPRurHVhKSi6xMZmyEe6c7aorUYk/LIUCimh3MzDCSC31NVNdeo+qsq
Zgv43iKxFvKy/EVgzsWAlcd24oR5mesxxNxrwMV/pZ/hRfotXS4wFrdl4X9CTngsOKEj6PRt8iBr
nLg7L0bs/WuiWSofnCJ65APqI9FBvBG3/ZzvNf7yXL1SrmJameESYGmFgIQe/tUjVmNrWcHyr4tC
DhEWs8RHSugJDZ+WfFSIgqcs/IF5rwsSkXCTNYfjqSYW/jK1DdRJofEi8bZya4ghnJQ78ryTb4iv
4M7YnwsgkExNsg4kH1Z9FY96cY4h60qXJFwSpm9kL6jjTUYYqYvu6DpGZKw4oDZMmZBEupE93Zpu
S0VA6YQtl5a98rXElI7lNMpNCKEW5HULdXIN8iKgURHL5S4qaIxYPgd00HXRZS4lZybJAPeq6VFb
tTt/URpAIOlbrhu7v/IMP22vGQ6Jc6MplW3zglMI+6qDJPnhDgUvaw0a7MqbahnNkxJeEVUBomku
eRlPC72lfnvJKDN5d/S+FtZ6MOWQ8a1bC0GUBB0vq3ZBUMAFbnTtqUtkjKDPLOKDQzQGFgJKhRyM
ITh+0mFPQxPRrTscWRkX+iI0tEgBk9IPgng5JkkM/OZHsQo5LjQsCy+BXvJB8x9JRb2zHCRQHQ63
o0SFcZOR1cZH//GsmroAngqUCj/jC/ifXD+7WS7GtUo3Zky80cj/GyIcDq8qEfDTQaHJTlkqcrp8
qyvhV46LKF3rRMRvuhyyOLb3vEgGSiB6rtlmBUMYlid788uEUonNyN0+VTZWNoN2GUmOpxBhPU3a
ULqB1Xwr5vIlYxgVysi+ztBeaN/appsKMsbWWNMjC+IALPrroFLcoV7cnaRb9mZTRL20CpuaJNqQ
02pWf8XZfoTC1AGH3o6VwLx1R1CrTtATSe+k8kqDNVAE9uKqqFyfuDk9IRgLRZxUmy7/Tyk0sk4O
AodeVHhA8QGrIWy91/REEYvTMdiggYVO2zOqwooJqrkf1HcYHwNm+K4s9MwJSsLa9VQMV/AMULHp
82qNK8UXZlRXPGoTmx0WxG0AT3wWYhUkpwUGfwFNrKynr7ZpkmVu3Uf3h9wA3i6R+s7aMXfSNw39
dIrAE99BIpydkeMvwL7LY4aGKM/K82bSkH4hXwU0Ayo08ITj0Jyq4h2fh+/V4QbPKFZKJWmxomK3
ONwXOyHJSzEe/jiExMYr1ulbDOwhtliO0fSS69QKO52FQof3nhoTaovaFqgjusdcPxHSq3iKuahY
RdfIDFE0Nxqb/sRnAfckxCeX2m3llJDupOu5kAjxhLsQgCr1Gm1+Xw9svjsf7pQB8e8EUImxUMOM
MVY77BmvEUcQ09D6scPFPfI2AOunjPtnhm8lcsN58U70lWnlJs+nFnZlncXeURVe044p74o3fHo/
Jfjiq6wTtt122DQ2sP01ovy8/qKY6yRT1F6/sImLSfbDrQtGtvab8ICFQ8o+AqcO+uYgNc772ap5
cIXcm8JwvfqwdX0gq14QZ6vtRpG+bIN5AVDOy/YeSE5r+VoNYpqCaI+hNv3ApGN+jddfzQO4J/e5
0z88ZFiHWB9B19e4mnuFrLVZWp5qW5HvinbkmqUH8VIEP3RtU2Vu4nZ5HDutE64enyfsbKBulkL9
T8g2pAXlQWK6Ws+qJX6HJCtUW05Dj3AiiS5Dx1MJAzNOPpH+mV2I/++TwDhHi2yI/9Zl/xOZNP9D
MrYYk0LQ8kkMczpvChmwGgDRNHcVX0r1O/X0xF8i6NxxHCYA8KOh32XtzjgbC5pyIhttBaJdVCOm
dEosA9Z8NG5EhJTHehgCYrd2HeWuSm4koyKs6jNDddsFdGGTKsPoFR8u5X1JPHXzPGE1S2aEz39t
kAOoikl1mikGYcT8qv4lB/j2hlDzz0oehjDNCurdAT+ok4Lw9YyH8xpdUBhQufBdaCuH4obZlnWh
PnYKgYjnDQU+qP69khDMmHW6tsPnCMwjWG2UJNg2SgKkVuEKKOVa06ndKLdBMrcZX/omRmQs7OF2
SLHcbT1m84YS8QNhBWcrTs3QXqYAU5mNNh+JoKFOpMd+qbyVWYOCv+1HE1/KGnNXDtDzlYGwNakt
R+VjjN1wYa4VgWjGrEqFJp+blTNGMvhHixnMIyMorFiDjHbPR9KQoGUCrqXGoKHRUVZUORkGvqbY
HEOhXqoGQc/643vkfrvD/V8re4Tg15NSpDU7HMXYsucFsls9LR4epeG75ChjkgiFFIekRYnuzfC6
TINE8hfuXw/KJvaGiWW5tA/EMsDMailP0GrjpUiax0ZlcLSE/AoDgOUdHtpdzhWXFlzkFx+g8/8g
vrvcfsJEVRKQvu/NXyoKMeAnW26KaPfFvCBRA1/3TkVahwzbefsBY7K+jFFlWP4xSutSZDeroKix
4xMiA5pu8ZEg/V8zn2L30oKubMwpaiim8Ad5bW1tXN8j0AgC1XfbnXCGLaiRCxlIm9ZhiECBY7M5
asWVTBxo+5irAjngUjPeG7A48g606AJm1hg6zy9XkByJdLVAcrR/MXLRp7p/HTt6woIoyJsNNBNs
f4Z5o6yjfDlE20BJdP3B7UHDZd/oboCj94FUdidEzotSFw7QuTT5yWQQpYi6Pkpf3/s8eVOBpoiO
YI4hQO46TppSdktsTEvAFAo84qJdqcfPwo7wf6frm7rsGOyHUPVObzWH4tmE7hRKiU3/DcCpxz1J
J4RfzGjeU6APEx5xlz4GmleaWvRDPgMwh+NnvpS6KMrI3AoQh42KBXV3H9V5/aorAQQ6g/5/gSJ/
kZsRzui/FyZ/UdD+/wjek/iISLUiobGJT7eq7BpXDCozMJeqxt9Hyo2Znwb6h3fxqIINXKmN+nho
Tnxcg61lXWQHpfATip/peauxhov78nu8hXPZQjs6KBLY6J/Zieh9ZkQa6ceDO1LZTcXDylBFnS6q
t8VkCzjH3FIGyIbJc4eiZxOgj8JP8IdgU2NclN0dG0JQiHrR0sWKOS05vyEFHeGMk8+m5rIzdYf0
F+xRrOqNM7S1TUDIuaNXmV145t9Uww6b67W93HUuLdjyiwr/tkwNRIeGLX/FHfuwX6kzcNRAhseF
z7Ht+dC513OsXYitbhei+5o/raPHyef3HwKB0H6H+EXfljJ/6CsupFwS3DLzZAzE55pYrFyaA6UE
hbEaMOF3aW6XfCXyx59uF2FwAC4KZkiE0QJoqadCw6GB+6zxGuvvG/Jcspe8OtPcqlkXzD3cvLqW
OadKT0PRVHU9PPxQts8MBkBmfRamV1hti+7br0iDZiPR1IUXDYPmCCwkRmBgbnI98SMLWl9Ru80W
cDzDevAQuecPh4LJrsIH//jKEuZI52C/IS4CdkFZJRAjzqT3Zm+VdTOXzhRGADfZKr7ohdtopNmP
dZTDIMbk6WtF8JpIBxZU9n+sTQ6ZGz9zSFj03QmpGjmnwN50Z475+kS1TsrFxWtwPqvwaJTWsTtY
QqR3+qe1g4w75KrTJHmqWQUh3o1SdlILtIkhIfGT5Qy/UlrhpwyTxNsqILJfrq2SEoVPaUjhYLtD
OeLfHqWBUdwk+Cb2C2gw3FXvJ6uEtqMSGniJ21cDSwplbq4T/YYBpWGYdVDq2YepXSI09qRSFqUs
+5ys7Y3qcD913C1kzbmeUxmfvZLYlzlvNdEgkQk26GyiiUMrfM+cBqKw7sbuFimmDBfM1kDhRcWa
Gu0kh8on91IbVE7tsYtgY8FGdiCxLr7D6W8+r3hBj98MbkM9AAk1G0xpseKNVR5MAJxDHfEi4YuJ
nvl2c4ZMpnUJvPU/yvnCtY3AwsqaHKMxXoKdaBq4cyCgbenWF2cKzVR76gwcRHh8pYj1p/fr+/Cv
EFGjC+VE50WikSa3MflHEMopoq1XQ2PbzcHt4rMvkH2DuodkwNrjxqHiIf0iX5+bkrEzYmePFOY+
DFLs5scyNgPh97fmU7jwXoB9TKpItDtbSsleKpx6x7XcenA8yUw7L45WDxeI4TW3xGQbt7xYYSi1
5ComQt4jgx6tnA7tH8xC/eLUuRvkMD1l4wT38dj/5zJJ9qy3s7FjYhIfc5QOThy/w0iO0THz7cWN
VvdvokdRBTPAsTCJE2UkWPrVVPYtuxGXrivtd/yB4DndPNOUHx2GrJDX3ZNYIt+uFjkjl14TR+Sx
qqxula8Td0vj55vNy5ZnR3hzpDhrcw6Ib30h+lLQ7yujDB2IdRrs/NQ7iYvnjNa5SrPqApHtTm5o
d3AqIUr59k+v/PaAjIjU1R1yJEFAildhgpl8KoFnjaaq4VNPY8tGJHf7EA5/FaTBRbj5Ich1VVKT
aL6XYnPQca0vBUZWIF62+5LoTbx9zUb9CYWeLuArn8w03DidWGrnKSQkTP894amYZiTbgh1ad+Le
2DNw6u3FqH+8z3h0rP2QHhA5qonWNvxQq+phJ/E4AQ+lEAqWhID2/GY0B9whewjMxkQu0shtCywk
cyvUGxeWT1WS1PTLX5XFYcFRoIjfcCIDdgnnhRjiRefsWu0j31OQpTA88zZ3h1ic+XkN5LaWKZoP
q6Shbb+KJzjoKgS6vyh4cLc2LLP9/z8KCb62SP0jSjfTcxjmRg57q1IvXwOv4QbnFMm5JI3Aoj7x
cKJ6T/8eEL5gKY4D93BSNQcyrpPzu/JsMFuvO7Ny5PJ0/pifAIiqzUU5UwoPukW3foR5wQmMk0Ux
/HG3nEKRJWud0kKC7IZlKgnJYfupodD9oZei67W78F0Fcg4TjMybMXsVP/tRFizZbmLi+glt9f4S
eJun/oGgfo506ngURGXhRdHNZbx51oFPFVpWyIfPNpUdgi9ghDgsEIJZhYDuNKT41lZ5MB99Bved
cF3i64uBHnXn9qWrstbOTmA9odne6LgNIMuBNOtoVEK9xdLOC+SlD1E8VhlU0KfwZzybQlbUpf6o
vY4Kd4j41t9c7R7fc0S0OaDc8zOtyh3Aaf1y5aD4a6pAwWk7+oLNurGRJQ3gzsknyks1XaxIcuXs
X7XL6b0yiNqp5sY1PAS77sbJ9K7eRFYxfNPnpyqMayW8OdOgj5E5ZZLLLXDup0Tkidy3B0BdlTDT
GoqE032+i1BPaXikyWYIqVZpvJVPLRiulsldr+j/j939GdE0pfk08MZCkQABWN5Qqkd7X8tcQLuK
m994fD8dwQz66vnpsrl1XmDL7vW0dB0mbPTaNY+zIKjhXU5eBSIoJgeZwfaCKhb/8+L+5FJYUhQ+
2tY03yhFr1YvJ+hEX90IGRh5xuBH8d9657JNliAE0y4GAyUoSW2n687RDRAELBLUcZQfRgjwJiSQ
zIernEl3KQxd3M98CWOj+zQAtkc+BkIkpHc37UyuoMtHD7Jn3A2eU+wmQsBi/JRf/PBe1EVOUrof
yQl92dTxSIxPZe8tvq+3kdzH4B9mWrjHwj4C5XdKN9IGsajNVWAJXitELrXvnkgBvYEwePod5pqt
Eyz+v9JnxqHEmgTHhl2DumAdyiN+fDb06vb77KqRqKdLoqR6aW6rSbqyikwk2Bs21noh/a8ylriB
gB6V/LMkeErzNjugjf1voKqTEfq4ZfPQ1oG0X/2pkNtLbKIfuV3E+e36be9TCQR2i1GCT3zkyeCG
wpfYpSqDwCCH1cA1rV2DCiaYPKKae8ZSkib6QxJHDxt65F9LEt2bxzcprikwtyPbJXD9jxGG6ksz
kVpxvOCAX4FduP0SUVKZbOOCj/K/Ax9/H374ZByMteB2TZ9qvfNvSW73qxDkyl9n3nT6qmeNFXiN
Pxmym4yF+TTRQfLMwbOoTcCgHBQ5GKDca/ZbUb9BW4O4P5nmf7nDhEx7+q99tDAaFeiISmTOrH7o
Z2O3AaxzO2PaR+fwzMqBVshlgJYt8BjKVwCim6q7f8Ijto1WVtreCIpK3CWwea5RwKRMywndAGIn
yTWYMmAegkU7h4BZEDIuKcPDa3H1SvkcajL/eUKHP2WnYVSyELnu3OdxvXfh9dCZp+uL/uej2nkg
KBs/Qw9btvB3Dh5xtGPTsCHn8Geiv723/bhCpmU1Vk28GAl5lBP+nP+3AScqDdkDcWULGW/QtFxL
yKeaa0jz1lH1rj9Nrw2Tc6GVuyZ7WPAGJ6nIl9S9m2hm1Iug2t5wC2i8Tu98lUzWBcMm1oU8glTX
RCnHi+dV6cVe7w4O4f+++CEQbbP2MD8aNme9i9f6aWW8YK/BPxj/dYOEQv0Lfo1unffDPyZ/3pal
0Bdur0PIl8x47HdAzD2dAf2JR3gqQYTmXC91yMBuD43HEEugwVj2cpHQWYpm/T3+y8HwKM4dnJVw
GhDyXBB7tvbeX6yTWwn7b1/Wq08k70DPx5MzmxMM369ESIG2Jqbw+AWjL+bxKZ9ru55fhLLR1dqs
+H7IswP4EtiCfIMasRlrdgiQqpBHNbrxB01wnF+ayMzOdU6D4VDuPiN/T7m21twAwtpwtnDCGGfU
imhx03gA2H2zAeGEKekbokc38cXuVbVIYmms/Usk+aCFEKHxnR6EMGL1tnFQXnYJMmvy48nhVD76
+OKs6mM0YuPqTWAqzy6uCrJ4R1Aao5Zkyh9oo8vkP9/m5VxJe/vT0ocGUgjWGd0sPPTqCLtKVLfI
n9TNOCE9+zPDhddfwlLwCCtvdHetgjy8u/Hj2TovAXUh7bTxGfwipFM5lkIqwHassCxLZBqwiH3j
FyeOJXEUkhpkOtyROwRXK/KR9vgBI2mY1ysYX+de8Pm0Ck50H9rCZVPxkarKFJfn4aGtCXxUDYoW
adyGmCZU/Gj7E9Nw+MS3VuvyJeYtlEPIahJ70VJouM3K9Rfxhbyn4Qc6Q3PtZ1DPJgwkBgiXdOuI
51vQMdEuWXO2ycehs4mS9JwP1va05tZdBacggWB7TB4ZkhBRAwxE8+TZP4XxCERnkTrEdJcj+06H
OeC+nZRVEEjlAk5+T3s/gJfYhjziWS8b1BQsIKz6oOLyo8tyYxdXYwsf/aXAS2CdQ5NX+16scHhz
6qXh3MxcdMidMIU0PCQDVGB1SYGa0TJinY4Fo71f7QuqsoaSt/riRcMRqdVqsXiLptxlFhlFRNoJ
HSMP7EbxWhy08rQ2VOT6gDKSfN+zZn8IsY+6Y3iCweradv4lsokvFNWUltjoeekzDvj/Eu4ZtL3C
kWc5x08Fex/smnw0Q7lCX12khSn8efPABC0ol/xDEK+3y7M/jKSTvZOoKIk9xhGsZuQrJgt1qLsb
mrpyaGtVgtIwrZHbohQ6J+wHfPt7ipX7GdvstLiCRA1PQ4MyrAT4/uTnt1u5mIC1WdcuxfrVOUZA
Ot6dVgGHAHo8ovPbzEtK0vHXcp4o1ARyHOkmW7LtTjijblnmmDLd/EUsj+o0MqezWCNlzySTzDip
cRzhnjFw8XhmtGvsG17OHolCiutghG8WHYrqLbbcTGm48cX4ZAGSgLPB2TEqUoIJ8endistH3Ckb
f5cWAMEAeOKwjYx/exg9Q9VgVNoC96K2gcqLgebceMuM53ePYF6Yo1jgQ9naHc1BhwZILAucAgal
1huN/dTVcKtaX4x9N83w8Vo0UTIQEQvRSZAKth+uUPQLGovGZGzcLXWljva/tr8Vgj7DNP43HNNg
E2ygjBZ9qGJArGo0f0bEBxRnGFOQzDwVucGrdPb+kSvlNIchbyVQhDtRLIxLtMM0JqRHztgYaJEA
9JfHPqMxt8L1uo5Rv13EnbcoePgxl2fgYIKmQpDrrX6gRPAmkn2yLFQIWJqJx94N5r0y1KlG7McM
SdTeu7bf02MJ5+YSQaZhIuJ1tVNVtroyrlWcMWbvx+jMP+f36HSRGO4Np0/6qZyxpv/ASqtp3c5J
Z32huvI1pPXohcy1PYriFqxvH6xMpq94iprvcwssZn7TiDokHXWDBJWRFs5S5EvS8vBdQKyNnDcO
HXcDd+Aany3A/5IYR2d3Hr90/PrQtbig/lU9JVzK871tAgX/YN6nEiPIkU2iFHtSMc0ONdThxGCq
u5HSzH7GBzx7023ny7yPS3TEGGiozu8YK9AzuugPu/0LDf7mfCx/Z0MRxyUnV/+RFvDl+/Phfy3/
kBUyGOtV5EejDJCC7P6XVNEZGpeX8YviIj7HYMEFTJAyi5yF1w8dJedIvtW6cMq/62d0js/7E9Rk
ZTV6fiTw/aoj72fTaoN973TZEiE4UJXR/GHgEMDCpVNqFJ0oTl+ZUFWx3uzA/kXcM/cpAWe89hx8
x0UOGGcxsOezwD7Eb7mSUxusBQrkL86AriPfDU4JFE1jentIaJuOQkHAWENSSda/Ddzpiblz2/rT
3shFjgznpu0r1o0KDQIFhQILVS8BXk10lMACpnW0Fh+TMhARtnSYme4CRm3RlP+8E6ZRWXrKaSye
GOMI1Hx92htGUpIOOOBlkHMpLqqI4VDRkeXdoBnaYPzfMvrhxTLKfEb6x2zrOWr/8ua+5H1TO9U6
zqTlfDWgsl6QOuy8Aj7IAGU8eomZzOr1wQE/e6qoy53oViUUeCgtZnWTDzWO4dRq7mB68tyeoCIf
8cqQTuQN8eP3JUGYQJfAVGCM/zXUhBQDLAS35IQrIQtFQtaa0XkDtrW+SG7CRUafBSO7FPzMZJzI
9in/gtIsHweAzPbPXg15/ebWUh0eMMjwZt0A5Mh4YYu9p2Qq7ZwPnrR3SO/eJhT+7sNY5kb9+Yls
tRLf3wQxKj3IAuBEkujPbBf7vgRPqabTc98U9s+xAgD9jqZO8GHT4D9u76f4DTtcCdxPpuRC2LVg
gME4rP7t2KG9xWMNbgwF6hwz63G/Fw+OZAzqj5+UV35cYliVeMSrpaEQz75cFHQ43N/H/VqSYwyn
X+LAcVhWWNCdNMuAX1LE+xuKg5hR35O8q+tksCGObIFKgTGatCTee9GVjs9wkGIjE5lmYccIHxt1
JcS4j/MZ8i2t9OS5Oz2n3fAKe6VGEhNGythgjK9PD+aKyA7QvEXhseVYby2oS8jlZnCFgJNhikpl
P8+YCMw1t/eVLLnp8sEI8kQR6Ib+OZKh7EBoczp/gbP5xWedxZSJdFdgx5BWmtObUPE7oaXVlY6s
+s+S9PvnqxEViSLMdS+Qi1GDxBfT0OmWCOr9OJCoyHnXqPbjgfsN65pnc+n5u5DE8FRWNhfVEHRp
6LmyPCtdogj6tjvAZ62Q3nION+X6jKlJ6ALKEo/MoizckhgF6+4a5TfsJo2TTxh7PCOSehaoAKE9
vrFT7HulQLosLzVlh8ouf57NxB14VdBDK34GahTLrdxmosMB0nEF6tYUOduChuzFsBUu4/i126wa
ZxBlzFbHzYKQsvfpdkCJ2wLBsO05/CyGCYxu2b85Kg3QwRTLfiInSUrVs0M6Yz9vW05YMTy+Zn8M
qGlU8n4Zj1UoHyVOvs+OIB0VUJ/fvyE5NTbu1rD/OoqQV6wzCAFT3qnTHq/6C1QjGa8P/BZqZ6PZ
KMyw4lmmjyuf+kLPIgNJ8Vrs1f5PSTR25OdO0AflUnj4j4REhV5WLY2mJE5iTKRmFEIZnnkNjSNt
fRCgbq//AL9OnidoElR0ouNPy9moImwHTjkJ4GmqTSyBN0+KgfWRwlE6TwAoOkA8Gn8txPbyjYZn
uXm9tYhXUBthV868J5ZoqDUGMjwvBx8L+uETb8wyQ0YCZXUQsKm0G+5VchyE5HAYN6gdsf3JwiFy
o6Nu2dBt6x3SPaTTAXa8mnlBdiLe5JZxykpJ0dtj0rZ323SU64C/0tmUd5GdtRbNFGGPfcmq6r8k
DoUtv6ByMp/wazAlo/VT8D6LoKaDQ2eXdr9+3hfLcD21xAJ16Oe/FeLqQIuuQ6VYs78CUTM607rD
L8LsySSi56cuygM7cd4nXut39PHmiXGPkMSSZsJdzjnA7RBDLlSIaunyxqG+sC+MJxMYs2A6EpuH
FEg7GsgdK8mD6nKpIA6/Km6iKfpa4cHUbhYUAMkCDv5KVmTMermfLvzI06adoYIpglq8woKD4NY2
ccN13plWp4Hm8F010uTIgMRXJbPZ2LkuqkGiKfQpZ6riZgEM4/9dzw1ZsNDnwR6dCPQ/FYmnut6w
SfJaofz/x30wYLwYDjMd75sRVGwh/p+bYCsMSRe7oXLVOix89IuxKICw8oIbhOdjZUuT3xqeZRFU
/K3n0vCMeUTL3gNHxxDgHucX6CYI5RB18Df5xUlirLdek62P0VK2AX2bffrx6vfPY79aIqUWntq2
HSdRP99nM71JYVPkdRhWXn2M1zjQdwTRAlYQti/iXXX4iCtmL7hglLSBDf+gf2FnpLWocuYRd63p
jWbwMPbA+u0etBzBnKdV1Cq2O1KNsx0E7dQu0a/poc+LBeMkrRoh+WmLksTAtGSBh+BokGT7ahdQ
zg6efWCxRNYgZWQOdxie8fBZjKTaHn7L99zaIS2Hw8clPlMAblSilO0ee8Dsp7sOoivBThWJ1gkR
UgaPfcaeoS343O6bZ+dm8RmQHY1BY99VzLL+ufEhFFZ6mrxdJ8NLLrrRqeAJbaSAIKiMSwHJ+uoa
5LhSUAg8AOIWZh5zvBXBIVwy/nlSPEr4QCK9PNxHcP54nTw10M9zgWqpcZD1ZXTNsx6l83Vl/LVN
JhLBTb3AS0s8wLxpoh3gsL1ya7nAOZZqwqYM+JBcUz5El8OpVLbcT0fTvl4ODqO9SqvZqmVM4Kc9
OY1UW17SxfiuapzILeYXOKbESyd76EVK1hRXeNFjogrrlAABtyTpL/r4zPC6/m44ufyDXhRg1lzP
Mwp+VS02d/RSPbpY18UPS1A6qxLhiWb5v1mqGPIED2XDGLxDqwvx4ct5cTO1Cz+uBlffo3n9s200
opNxIk5Kg8PJHIt2x8wV+weaP067lmxUe32XO1fsKh/7C1UblJHLqdSR8/MbaPMqYu80UYGb6zl/
GfxUqgn6ppdxodai/rnbhK6tZcNMNHk5MITqc9jvFQBdHdYs4tsZJs0SeeS4GFE9uJA2ur428pDn
2h8DVjPhjkWhpH0aKHjwtTiZ0PqBWmfODsuE76ezrDc+3DCkdVitVNWwmm4An8NNZXLWbevvySx9
MLsAMKNPolTBZITP67/24MN5Liwx3MppGsh2kfD/8oF73nF7uLvxkwa0kmE3sU3o9YGSA6CYc7te
DiPxVjoodVm2+hIgchil/c5gNE++hfjJ0LE/SIKA1ZGPHOI8hKdDrtrAg1mF2Nkbbf7CddT5E4YZ
2DLj62atkKzaETd+3RntKV9ZHUspzCZ9BzhkhG3nG6RJXvnRnXmvVSI/Oq8Ae+2g+fIK1HJcp8+T
OtSc+GL9hJD5EmIhOrvSPK4i+fn051yQFENkK2h+wjLdfNVCnVfgTAjdhnM6T5E5dfu109X523xm
tiU49YIO6gv8Jq6VppSiyFWe8j6ES1mIZt1oKQww0duY48umrFmtzMJJfOVL7HgLQIN8P4MjEPlX
Zy8AUG5QVMUQMAaZVyEJnTb6LKPS8CVR5K9knJ5mPJpHSvo2+urqqD4xrBQJPSn5MM7D7wLUm15x
Ma9WxNTsknopO8yg3xXd2qWMjpOVlC6THj9+Z54NR11LNij+EvIAs3RaV+0EEpRp0ILTV5NTG80s
rNYB8q5+/omQHQcJtkJMiOU60x9x+0JleME/7W5Qz8yBuq3syqBQffrNJjx+ffNWxqW0Xp8SBeLO
oUOpxXvNY11nDHYrXGlaORxNCjYVqSr2iOVI5ZfCzv6HISRSyvDoGYDSgV3oaQW3NixHnmzqwkVe
oTwi/JVqjrxaYqYE/HC1/RXCRBJiRqOOAoQE4Mn1xi2QomU4qLN+mJK6Sn/6PrS8tL2+5nBbOiOA
+IV9FA8Xiq8iABgPhYe7CV7f2TE+C1ad8ip7E9tL6J+KxGr1I+0fnHzKmpgs9azNS0+V2Q4aNjus
nX9RfCUr870SHebaa2DE4fBr5BF1vRvy/SiGQjXAUeWxoxVVH8xHx2/I8VKkhu9JPkwO0+Wv4QV0
wqOg+im7ZZCpsC4S09d+a5/iUhgCoLa8ydCYciz9pOBTFZxi+S/HVzJ7cQh3ZqjnSgnFRyDu1KNp
f24cqX8ZrA4/vFUqOHIUljsOWmZoRNpoGkSlO5KQvQezeC8jOLAvgiaUzv0z4jZwrX+IR/mZgss/
oKog7S8bkQFJwEZ8gruDrwMbI7iqSl9BCuB0EnxnpgixuqdP9f9thP9Ly3ztBcrp56r+ad+5AwQ5
fwVm3KXjpzltZHklQ8J6Qqqoq4HBhMEIEeiUrjZ7CpbCs3L4pInlNnocVZtwz9J9OQlOTd14Kwol
YbMR297BniMiZQUccIwd0a8CXAt+HNt5hl0/3idG8ma+xfO4xrHbc90rnVb5YI92VDEMow2VeHjJ
TMKZngaQNXRCHECveP4A2r7e/VPPpNtieOINW3pQXpwFH3VJJnimJtlUewaSx57s0gHrfPoz4ZaM
eK0mKA8IyahA+xvTcBqMigLpXQ688okCyqdIwhXwHFHtnQrJeNJ70+d4hbgM+aLuvAJM2AY5jb9Y
K0UhRDg050r6e3E+bjgxC9elbXh7Kt4YZFFVTX2zUe2HiH/5Di/k8QCdnMCaGGbfJXEyzyDiGkQq
lSzYczegvufukVrYFd+AnArtXupxYOGIZz8hGGm2ExcrEfxdrKiQCjRX3mLRD8DUEsNoMzQ4oFLY
o5+U4vOIwVFQ0um1xSD1C7LwqD8aReLYFgpYEc0EQIWShwn0XI0vYjwvrgRbBOO9Zmmym99j14Ue
Zoq6nA5fCX44CnTutixENNeZBKJyW9mpk1BRM2Lsgc8gaMrEht0jp2j3I3cvr4BIxen3PLQKUZKr
MFrI913iwajYpavEgcdcqHyKLYmRriD2eZkxVGK651SFDS9vBkdTr4QeJJ/+3Jd2ObanChec4sA+
UW67gkGK6hvSg2n0kFQR5rShz94w+8VFUCOvDxWI6CTUkGF0mgR5bX03AlAcfreq941yr/TN0r7b
S7pX0WFNw+4bmitqQKitnzLuSpeH1kJkc15hZLn4e6+oL3zGXS/G4eRA7h05efkcpc2t6MgOYAKI
/Kj8lU1WqWy1n2+WpVdDIsKGViqVde7jBlnKIZBlZtlzsFSTXkb8Xqdh21XzwKtjLvRmp8NB4v28
PcZVnYWIGAinnh5thWh7ddCXP6ZMVmouPAzTCJQ+GUdOTM/YKzztw8ZUNZZu1ZBjhAjKwyxtd7Hm
hLRxR8CqKtP+tmWDc5jQ2uUpw8kcU9vNv1I6M60SSq/I6tmBi6JuG4yucx1AHV1dJ40QaywCVCKg
ZnWlSFpNKG5nmNXG43N2rOgbcqYzf+8QXToUCfiXG+kRJE2ebL9PctPY4LCi/BjLdcw/4zD/IZLh
lQeXDwflm1sIWldF/3q1F0P8P8q8lyNOycvGFko6mt629xY3Y3KYeXYpfd8PWRggnUZadPGbItXt
hiYGyfCQ7QrxI/i1RJch95JaYhIkBbTOgc3HSr7mMv6yt3UdZn1UnXNIQVrcJs2Bt40uAdOvPIZ5
yvl0PdCSrZzU8Dqt3YGLUl2bCMy3KcBXVHMpiLWAtJJeGDP3k49djAhAHCQ9wLHqkpTC6BRVIZuG
8/svib7NqPhRIs2E+5VhIk2mfJupS1OA+xMSTbXR/y2rnqlZYxuzEdoRSzMM2wn6VH/A7x7Vu6oc
+IWj9laHt9z/uQPP0QmZSy10wdR371MVhlQTSsNwknAUxArnJEHNw06+46Dg/zvsVBkmNd879PBS
cXJkI3eBvhXDTNEGNp/vUEiIUPVFJrBSF8aAMTYs2aXHJfJIQgjhH8lqo7vuPUL6tjNWcBARSlZR
3gN/pV2iYMJnxsx0ZJayi+OqDnCj8C5BuCvtD+YPAWuqlOqlGToJd0Y4Y96jLYoRmuslzuQU9qwD
bNN6xltUhklhLUjEDwEE7NEP6mcDftGYJbs3BxjJvc/M+qM8xhtyezomQqr4yAKaXAjHvoiS8tfz
sLIh8E9IEZsr6kR8qf1dDLJ+exEhIZ/YLvfcuYXeNjQq2DgHs5Jos7puUv/UaHYDyIODOKKemVEe
SEd701uJtoxUbFfOhzsQQx5oOxllZKO3KBU+RxxRIoyr/RVoR2A26kSVlrDlxlxnS032lQh5eMxa
+YeqmGW+onoplwtKyVGJJIK0SelzZTboYxBVvK5Y4bjwvXa9p09kNdtM7eLADAvcWHqnBI7Kpb9g
lmEMSOyJ8flmkjorPWo2+B+T1MBJ2sWJInZUBGNlNzaF1MXTDSjpUMRE3CsgW0kr0l0shQqCrEv9
RvRlZgzTgAZ60TPo9b4WAjQNyaDJn5Q+ddxHltwo8EndeSh9Uzc4oPswCx3hFqrhm1Kz1XaILpjh
af1TXGqrT7Vstd0nKJ/ncyNzQUqfA5p60iI10yL3UasNVIiN+saIU9eKPigN45kODqzCaFSjtpTi
YrhQEZWL071C9hOSvKRxLRLHwj/uIPMeqfjAqG8SsLZzAs3Hkt3W/TQut6ktSX/t+kNPyjtbfZUs
TBeKdvrWfBBaDKDHHP3xalawTd7YahkMlwI9s8BZx2N3LA21hoO8xUxN0RbUUx/eCRCRjQCAvXtd
ww3+AMiupWjysuTjGC8TVeSDS+KYEXG1PDE0N7/VmUKGOQC6WmH6fHItlUqZaWWvHQtK5RJ4+p+5
5kVRrRSVjAb0ETeMnBoCpU2tZzRQixbUT9jV2Re9POf7r7Xh4/UgKQaOJqT+H0dUkhOS5nh7DmpR
A2tK61UCWKoLsCqM2Nl1O6/owrQrVRXuJ6XkDVLVhTTUYg+y7eFqdDdLq9tNgO6soXnAj0Uc1R/n
8o4s9J0vXNLVJSkKrV8C00CsJQ/0ivai/fj6EJcZ+3WGMJNjUiKJgYRcNNtfW7BhE1v8sIPMU1nc
zK4e06uOchHhWien0AUf4kyrE8fNJbJjf0auUnePGXkG+kFrk9GqQ19fvcXkfMOo3NTi1Ala/+mM
Uiuf6FjEONjTiD2HhU1Tu7/Allxkwu3+aorCzeZYWYz7roMMnhkuY1QorqSYxFIC5TdQtA4+hpMN
UeSOOYVo86VGOM+tpTxDsI1eN9O13mhPmu6lLdBrQnCHYDxcg6/66V8fpV1FEvzRRrgPs80SyB3K
vbtoQjm1SGDdsa7Sp0WcldSybBsHuANmICT5uSEyTmYK7glTZmoMaYfbBYAXiwty3jcJ88/aHwg2
flP6y46opqpkz3FpmHJvD4eJ+1KrWgycgTbbHZPf/bl0ZdKDMp4uaEYiH5R+Pr7CTs84qEic4y52
KpF+Jp2yNf5y8O9ak9uN/r/SNc6+djdlUt7hRFbKV77e5cWkjas5VmM5JDxSlOMQbFoSpDGVY5cC
9xg9DnbUhBSwbgEdBCO99pbNJUHl6b3Q1eVi5HTpSBx1oQksCbe5rsZpITHWojISstEtcx4to+c5
fitBmJt8mUooIrFUg+056bl4hG9uVVifvGQ9hYOj1C8A1CDrvsIpxBnfakHonHcAD8/2+g2UGvyq
D/AGcl/xa0YIRULC3UH0LO2uuELkkt4JdD6AcDaCMSO7UvN4Qrg6r0JzbJAafosYCqAN2c4IXk+x
thC5RagRHjv3Wv849rNzx9+8TGidjQNbJsavmTJ0V4FwzBJnblwvBOrABDkFbWCJpcIiAnE2tmo5
VzEonpfAF3QA3ek+H4b6BuYDCqdfDgxm9eruPo7H4UM+P9OQ0kvVCRZuVUPUoFuKnf7PaF32mLFD
Qlfi9TmLGZMfnHhyjw35fMJuPYNlNNnL0WIwFBpCxzde4r1SpcYSHM83hSkxVyHIpgbjjB9We16r
HbzE5WZusfuBOia0A7Qexpe4vD6+XXItpJy/BtWz/Kmf84IN94Z8MFt09JTnaY6TNgzVvIPjLYiR
A2sZVX7N4Bquv3qZZlYWIBK6ese4/4+c+cCkgBgQyj4zj+2/hVVOO8f+ETNEgZ02Oa6sIPpgoQ6u
TtSpnDzUXVfjAQYoq+U+GtNtIEUJnsIHxXkxqrhCCoYuZm6BFeur27hIXod7RQXRE3PJG2bIUhdz
g9veAp7x12IOp1eZ9zoDclpW1lHc4lKaXTHNBXgivCfJ7rerClq+lhteBE6ERDT9sczeiksVhvG1
yqEwU4F93umqHyKq/jrIv2mSDldlcv+Lo/zbNNHcwwE0iS1qT+xJZv5+H6QYg2fEo/cvWCPavls9
7bj0UacrAD+RbuZw7ulXSL+MqZaMjmDccW/ynhNP16gkJSyCAcIuGL1hCx73SDHYGuZLCZv13LLH
e41aKxJgrcwZi9ulZX94dW1RLdGSFJJrMj9Q8FN7vCsCfrreqVuFw9Yz9m4sF9h1grhfG3GG9fQ4
Eq+xwTJhYdJ6FznRvxzX2WoehXzG4roubtFSJLt67wnoT1bQ2Qd0nl8CqfHvwTPmETA/rJ7+XpWJ
r/2NCpBuCl8jJmXN2F6/vcaJQ50UNr2c9LOW9r5pK1/WxbIebfwU5NsKk1KQrrZvEmrXF/srdfG3
M5+EZUBA5CShEHFPhe4d4F97nX+xo3ISqqK8LfEOjjsIddLfXJYToj1yDL3cfHRl3LeS3KaEekca
pcgMh54iF5Ln5lnc0PxDO+sxlvU12u0gl4t0NE2wL5SIFB6+IPKSKV8yOwRmMguCyMU9cXWGcWkT
bGuA/XlOZ5KWZTVsbf+zM0DMPNtl5tuIbVsxSu+YzdoVDWLsf+unvYBpY7dRvG0tlh+sc4ug+vBS
QuPdxdgIHoTnEEK84qeugpuQqNm592tjwR0MFDxuld52fZSFvnDi2HbMmC44t1oU2W4YfOUC8KUJ
bMr8GRxgD3UE7gytKnUNFIT17GInjoOMBTb/Hjlb+IWHVCDGlGKH6Au0iQnO55wBdIW3BHy9tgJv
BR+jYp6MhLp5wqm1oJi7+IiAYtVaHP9RV68AQxKS07Iua0E/419wgcQ+lw6hfA78ybeOQEnZhnAt
CXXY9tNTaAkpn2je/mGQVFYvScrUazsb87F6fmwConnJoy/RCGX8BZe9EFGMr0qseGuwtyROobu1
zN4mKhefn6qxmTA00DaIrABsyTxwS3JKQzJJA5XxbPkMKDRIEABatuy53c0bs9s1GSa/B9XM1fKv
8NBGBXNCSRpfFqxiPBsyixif8CyiIWMw9ahatO3mAjOF2H52whELPJQ5cGEepYDssvV2wZRAOmDD
1kw5KRHM46UFh6XRpUASYNX/CajxVMLfa3PhPahxuBHs4iflgWlKvOFDCgi0SWzqp3F8RmW7oC6W
1EabnEZazJ0+KScC6KWFlDDLjZsuILAZBB5V55Hzcs0F0HVLEHEqnsMyRSqABmsWQWpgbNWIxO2n
8TiO3FUS2hRPvmua51/HfsMGNmolD1UtOiF7xmlJ1FvTZsx/PMF/3q+72X7yeVgbl5B6fBNMFR0z
CaFfh4xthDZ42Z0jm8I5oMaoTDjWRHj1mkfkVaWSSyHQ3U9iQ//sVjNRZxNkbucYbzcOMrIeqkEN
8UR/RFVMULbFOs38cl6NTm4BSYjZe8aKvVPxWOoLTLcR+hfe+x7puIT35shgA+2/yJAwvxDwxbun
qXu3GjtxXHnBCqp8XUQ3GntaqKMjv8Eii56CiNnGa13hrprAlO1nwUWx47DtoE9UQIEpDSX/peV/
FtOIyq7dngJSQwI7GsUj2+aBjpwWIse2NupkYwdddMuYMhWghUzJ1CVWP3z0U1QkhurAII+sdTof
xzm5TFxwSQ3PO6s77jq7QZOeiYB0cR2Yp5xsNRHA6wTS8d0crlMToA+gRCHadU4rcTG4lqOxYwsc
mXtmu9wypXezEvHGSHHLizw3UFJCfEvtVU7jXl8iBR1+CdE02WERPBqQRWL7twpce/dMIRlCwauA
D1HLrfHhKTMTLVk1Ls40v9hCHJi556jRLX484in+hvl9zm8ksv0cSfBStcNf2JeCyIpWaPMVOV+T
gIaEJUisvd21iOXn3a8MyYAJg5CfMn6gcEc+OzmYauacvjJgFvnYPHcQ6tscrdGn3eOzB1wI3CGP
PD4M2pLBS2JzzyBJrXlRG+jNBuk+xoFooMp8BfMHjsP3QbwvmW8vCPpwuj3GHO6FzUzfBtv2gbj3
+xLsWKcHA8NtKh7201iN1U7BNW+w9me3YwzkRpOvRpqz4OtZbPSeh3ieRUAu0/poyxyfg3J1k4h9
fo9qGi1djzVn4o+ytpGgYTe0Vgo9vBRntPBdXPsc0vgGc+CAJXvvxwgVuGOynKASdwJdsCtGKY/4
24NTk3hJzNn5zzW6ZlJPgxHhamdimjo1gToJufaAgCLMwQaDxUd2ye5UKCQBswfMGy593yen9QfZ
fNvuUlH2IUaqurFKEQZyftGb21lIgkNWgza4pn5l3ioK8wWYzJWPod245iCZC5fqineLIcBZR796
9JAL3hGXKeBVm9ZlLmZX/TQ3r1QHvxeM3jwcLj5s2RN3nApv9xgH5YThiq8dsWlFbyEX9HH1PbmA
j4jK3JNSucLUQ6mPnrJ5SJw8/mXVvsS9XKi3Ns8BesdZKqP3+axRhXjBMSIo5EnVna4WZAY9GM8u
kLIyGPyeb71ahveN4DuUtZhAZahDq7PTsP+0DqKtYeNJ0jAnEm89bUjFToicxLJ4zrhWtSUON+b0
zFLeMLg6WsdYtm0c6mN3JW1+wEPi376LACZm1+TkAM29iKKnMh+fFszy+z516QlvXkT9u6JajP4G
tPFhXa8QlzoLVsITRN98tLQmpwkUkYH9Tpnayg7ohRJsjb1a/yNQTHqeE8himmpSVU1zc6jLi8Rl
J+JxSa+AbHnCQ3MihmlmAdW2ob9zsqmDlseh1R/esaHhiBNHEm400KKGxvzak7VrhC0Zc6tMjkRc
2o/7TQhDyq/Tn6iF9xZaqDyL3y26AWCRQJG2+jy2j+lJdxsbczZ4GqqxQoBKFlfuSuj1g9RGPBjT
OkGza7mtVzSysKsB8aIjPfxjkDpFEBmcbHUsTplwliKdUvtJ8BSQnQLVjagcy6fs32wOrncir/nm
7fbvD3znC0eI8rhlH3oTpbo3ZM3rBMiETZcNZvTJa/EgmK4mhRAAOTcu4PUg+LFfjQgxCEHyEn8c
0h4f+Ntb//ppaFBqfL3AscI+yGvc0ntFikZokTD2BgSGhDs5ID5N50+eLLg10/K380kzugkLlqlV
mDllXFsjLlP0jNGvV0Ou42ki/Tf1UoxLINco0IA1n1Je6IqAlECDCrkIgexNXRNuXAOmhd3PYrpz
e5uTRSJ2GnOkIhArQhpB8cc6pscdEJm2L3RFbF+/NBGtIZqSNcXqKYZCQFaZOUbSTpXB0BzJcs7x
zvYOF/V36LWzeqkUOJ0rfwStUqeIDT9No8jRS27BgvzSJpvK1NqyOGNoTykNIlCPLHLA67h+4njI
KF1h3ZEflI04+4DWQqgNxzUzWKHTTYBkv0PJkokOHrAd+uRdTIqcRs7PbQKYVDq7vUsEf9NLf7+/
Q13A7i78u+XZQy2mOrVKImUNLPvHRfb+cnvODXJ/9VHJ/cvkRnym8B+nBY3XGcYJPvq0ZzUCAn9c
KcSAE4ajrikg7bJcnV29xf9tTGZQ0aS2cnlc+kEoq0G2brSWSWxxwPlqHaSXTH10Q7I+XONjH1UZ
KG1Iwej6hK/CQJNfZeqFT5D8das+UgUJ7l/Dn2OhPg2ZfUzEE7OQBf1Z2pzB43EG3ELzbNmf/3uF
I6B4xWrGOmhBqBnubPc3HFbPsIe6m8cwN4g6pV6s3zVNwD8teCBNe0pAXjrneq50wKPlzS4EBMz2
BsOrzMlCPBuf8CytCDrd4LCCLETG5itKVizRKACmR/vkFc9c0YtgWpQQJXvOJ4NBNwGu02i3EZXt
hJixyECDi023UPaalw4W2BgAmpuR2f8RMSNyuj7wdXpI3yhcoLcFFgr1rHZeebVVVMWChHCV2qii
BrnmbrXNRURAExB4ByqnBqbxCrHgCGlu4QGV24B7rnK2yWNUd4KlaOtBbe6loM3TJf0ChiOptLS4
qY/5MzJOs/pvDR6rFDi4bIJrgTxiIBrvJcKut7tMmcpQ46l8fgfJi8GWIlXBIvij5cQHXjCIIA8e
q8JYWM0k1AHkxoPCp/Lqs40R4iMt8ZIAlBZhLC1RGCCWLTlgVCw9XTgzrTD/EYpLfGYS7VFEk22m
AyvTC4tZcRy4uCfEyplxgQ6GCCaEYIeDfVJxMfoLzrSPD9DG3eJvxWeOF4+ExgVcsU7ipC8GvCa4
Ujw4DYUrg33xTkbsjE7GsZwUMYYen2kyCKHHUMnIbMSIihaG0WLTZLRXOdf8UKVumwhv0eWwMcbR
j3lBYh81KoN2RJQLxOVSQX+rSXB2ary86gTzvzV2RInnHRbKmR/XxiRz8NKt9zGviHVuPACzwR32
x61Yjhv0+bPBzQdYsEzMb/MrG3K+lhbOW73mmL2ItjrTGjTahBC9gE0G64DuEY8O97FnmsVbEIH9
DDZ0r18hwIukcaF91BWrmtHcR1p9jFxOZ1TLXk0lQIUulNBqfYfteg9wQraLVvpPz8fXXuJTOXX6
zQYQnwYXfsjIpQFNNQyYXcwH8f+K3Q9BdzQS9HHpDKnm6qRCa4/ODPFNjhKZL4LuO88Jm8TcQw9C
z6Z2CVyiW+tjOdGZwOQ3XqAGbq9cym8ipo6+rTbT0Ule3XnDVwIVt/uCyrdj5FNQwzhNaXBgJwjh
qaGzfAvFTmy1aRLQyc+ZYOpf9zEjulh6T/868dgvJicLGE8qiq8433ZwmfiwgVMW2DnOXqdlIrpU
zrd58d+5vbdK+DiHnMUxIeWQrYwm9ptnos7aloA7DX87vgPYJs+Kz1jcZRQhinmusz6z8hW5MB/I
w0wNbQpHSNIVEUzOHHHqkTfcHp1RBBFW6+1c8L3YrZqOM4pwQZIc9VzJ7gX90B8cRl7w8pH0TQFX
CeLpmdiEY2/+kSOXpL9/outvPM5NOB7YG+Bf1CZaAep8R49+hRRAyTDtkb2d3m9dvGX+XfQkVuF9
cE6T8ra5Mx3TKkX3eGXwUbv12SmpAGM6JazWY/Y3FjfjQHwA9SlMMbCW/jrnDzDAgzGG130W9bll
5/CZA98V6pElex22pAtHKHJPgS5GXlXuAAEZLpYmePln+Hi4059at7akgAMQXRe5/lj+0YtzyGoO
sr48sTFxizhkzm5HMxkyRVztIXZzxQAkqVb44FyBdwpQxXONLJ4veuOnZVAd4PscdnJ2vvowg1pO
kT9D7a7bSk+Bk+tlE5EW7jFHABwbs8tzrBe9jp9VTRdQCvUu1JNaHx+smTQ/edCjMRUmGvTp6prL
jMjIp/fmievMrj73626mQqOG3fvmGc8EWd5ym7BXeplM4jRhGaEd36DqwxBRMYPTrHwy03R5A1Cd
LrgvY/Wka5S8aOBVzayhjahMEWkzo+9iJG+ARTYdhrvkJV4foefBjt7+scoC3bACXHZhHx5BMrAN
ic9SsnBhd2DsVSarvMTE8CfyGLy0PAVN6BVec9j0Gu9aHZjWgHWgYb1q6WaNaBD8gJz2YaOQkDHc
5IbWNt4dWqyzEEYMd3y0RaJbqkrSaUN3PPyPH6nxY8ucr1taICoEbCRS9cSrPJlO1O9VQa4MDTCi
jYMT5KRoTTK5UN2Q7kYz/RvvKcZHvXsuItmBBfIRMx1pcEz0vwKhaIi8e3MbH9EYljsuwTdChlO6
kGQ+5StqDl7EEpYSpjrHZ7CsLnARl9FRysb8GF3R/siXTnhvU15WuIp1Jsr4Bw15kMgZm91Jpxy8
w2ejwCNjsYkhvHzwRfe8cle6JkSSwdNhVdWdRkBe6JzIlrezzQdWqyktN5FuCUMZ7iKMyRZomFbp
t0+QwQ/B+TA/xHgvXWh4LdDwGctmMsfXm9yItUqx8JGpeoMOlbnXvAWC1F5mLqXdnDNeHliE590s
19ds/HDji3J60TGhnzQ4gZkxxiElemXa1Tymn0+KG3XPPJ+9N0+6yIsJR7zb+DS7o6E0vSIhus9/
LYZl2OkMuVieKayIMWtGKBRj1nQOpHt7Xc5ziE1ukhD22MI742XNyqIGDngIVp6aMdqsevYrgitQ
Gk2XPjYHUmujUKOgsw8dwxmpVFYJYF0TkIRt5Eyn3q0dfi1VeI/AG28MyqmeYg3MDR0wCTPLqpmp
vCwiaoL6kMSWUCfEGKdwSDa8jP2kVYD6PW155g9+5Z3Ykk0LGbgwh3aXAVaxJvo2GxRvDX7r3cx9
Idx2LFz0GkBJrQ6QoNSp24geuM60z67sB37ocwntAkXFpwnvqRIPYj0K7mtjTxMGU0yNYOHG7mvP
OZdJmJ0Epa4poHDwkjKc2DB4GYg4Y6JzAmlfyCwnVTRanCcnvRdMQZV3mPaCumvsdGA82tlaaQEF
dZ7XKwUfwoprGX+62v/z+s5zp1N3hbmUl3H2LEXrf5kBK8Fkemx0fV493EnPMZE5S6fFjq48UDUS
G1sf0Nx9CSrVosJMnMVL4Na4zLQuwv559pasTZ9tbt6cbC9AjK8rFZABKZxTP+cSfMh93nBIGS17
OIK/2PNzMPaSKNmk6W3p6zRFiZ3HhUsaUiTMXBE7lcm5RKKSw9CW9e+7UfXFW3o14oRlKTK9mDnJ
LkXd7JKttGB5iBG3SU8PMy0cI7BygkeAlNvymapjErHWouYVp3rmpERoaQHHYnDvzl/LpBBiBWz4
rzVRAPskhcvWoiZgSkFaMMzjRIUOKJFVgkeB5Jy2y2UqmRqIojsH+1MEtUOVIFhaqMDm/JYRJGdG
tjd6XEcINHGc/1jHsKVsWAdcTJpNk5QV52iZl58Ah2sQJx1c8BN+AdDye7fodJzp3XtiekTROC38
36l9NUana/jeRJqE+hY1vdKoLefOeX53Lg1YQOXJPzO2CR7r2aPLcB+j5n/i+yePvc4jUTR0jCpD
4tDFc4W2O/hGUv290iZKzvzk8xR85oi1lbm2sqzHITw80jyqxggoghL76XNZPa0U0mnFzEFvUI9V
w1HPwu9U7xDNbOHGa526THcwHqcEJaSwg8n13pcNK77Ob5x7qt0i/FKkVGBYE9dzxagomXPRx1t9
iw7L55sa4DEuqaR2837jAaxEsxh3R40IwuheZV0LfU26Hw5bxxE/DTkrD1Hg89wrkGZRKf5r/e2Q
zh/Wu9rt8eLIaA70YYGZqEhZkC9VXEaop57NIpzwoWvZk7FLYJ5L+CztXaLAJD4ZQjOLV/PC/fjl
ZP1vxQkMNiy6Gw737D4pfiVx4CNtGd5e6gRphP2gXZSB8bCY+CL4uuzh+xHEpkQNkRIKxibSbBMR
xhaef/lB6Um9H0INFxl6BShG46hNgY+nyS0DSiOjR8keOk7Z3nEB+rFPJVYmwEEFV85o17c7DBGw
brlv6NDBfQC8KLsEuXDWob540AilNpNdHd+eeBcaL/r7s6WwnRmLSNWkrJNhgdoA/VzzCimTLhiR
p7jtG0WZzEW+IrPUnGOb0u0IUNFICAcuO2Nj1R2lKSUbomoNjGPojFjCEQJdEzAVbI9NmnvxN85b
uVtqXHyln5ttaWabTLRpR1BrmvhAQ8Qv+jF9Mb5qOf3Mcow9r7OYRkU0xNYKMofBZybfSYx08BGy
4trXakHp6EPVrPKe5X/67VkKqTOFvwrtCZqeFodhcw8sA7xVgwiDn2vtEpID3LyY94xyHiXg/iKZ
yUF/YTgI+fNrKnrif95u13uadIK0YQDJp95mIqLB2QGBQSB3c5SLz2sHk1+HisfkYPL7wW6q/+CG
3VLvZfwhbIeY7DaOy+ZeDjeLu24oDiko8jN+rgiiuwap52BZi0L2QnFdz/qjnf4MiJqTqDhqYiBn
S/HR9A4g/FaHovDdRTnLQdbhR3ls96vzHcZvDlfxOsTbP1p7d1cF8oTnzmRT/0NWYka1zVokUDYM
MyFh04lwcGYTug4xKaKPVmYSkaApktYwxeeE6p7HL2jhqPLWi1+qYQ7RSdO7kYl2fqTzD1DByE3U
KSPLfq87qMEnL7vr9kOzq89xWWsaST05CA13vQ8yZL4mhpOZ32zJmo7+ImgOAi6PNbTK4bRXT9Qp
LHaVGbn8bDcS//FG029XH8xSG6fXTB+z1LBMGyO5yStl2Nv1XKo0EJ8VKgATHSoz77vI8ViC5MEn
2phpQIarhDofUvpi8yQo5Ttgq/4ohgXplXmLuzQaF05q5gu5DT1nvXt+TtNFfA1WC/T0I1Esg9nt
r5erbT9YDbc1Y1RO4ihT1sjWUH8GDtjRkTgTPAIpVtvWIQYRTRsAgQf4ZrWBmAySIJa4eHXMyZPl
Q/Xtvi5NvgN/9fiyCi8GQ3zclZt384xJytc5xbBomUCW6j+dP7m9BW0quRtn2xAY7j16KndN8ujP
n+S4efLg5dohtnK4kxvvuYPrpf6wBGHMoAsuFz0ZIIh/oWtXVy0qYqvJGNCDv+pS4CXsUScV793w
k+A9+hFI332NCH6eCM4YuZ1tJkbZyRj+gekjkIPD7YCccEQAdEj1gEJvml29Nnpws9mhKEk60e6J
Z4Jfu+rYgHMOy7ChMlarreUssXhkTKb9AWeMlz7TCIlzeW4clgBRkh9dId/m4sm5iWV27KdfJM8X
YbZfWJVFc/s9LcBoKQeidNP4fQpa9ejqhMFHSdEtIF0Do2c4pQLH7P6Yof53w/p8xL5HIK4nRbY/
TdwsJBp2Fr2ZogeVaE+EfkHNm+QSD6WsoFTsmSWXJ5qUkNwanySy4n8ScppNP6UMUieMRuQ4Qdb6
C80+OuvIAwvwHFv/DeZRJUv++8YcdNUGtP5w2VH6J9T4jf+KWeNCfwXp9qkZlH4aHLhvOqzY6KYe
if7WRd+mMOzDpdvdgVi8br2264jrpwNUnqg9miueMLiMMDf/w1sS4hmDIBRg0GywBn+CeqR5ZKSG
h2yFm9fBCOpZ0ScziIT4W82l3wVUn8u7vjNF75SmRmay0sXINH+6ZXuVPAv0YqGqgiAhBlZCi+a5
FBwPcm8zABh0aP8eBg4juT8v1RuwPqQX0hqfx34PDKJQXMWMbC1xGOSIXh0tjWb+YFAnEmuTeizA
cqe7lFtxPSwbmvVtpPZDkBmcwFFiyue+ObbfR+F2qmIealh09QDutpav3KOXpDZN01kJ3hjI5RM5
xKdiVdvPBpnERQaUm3UeALJ62rJjMYC5NukgypX1E3mH2wNz1Lpy4PVgM2QCoJJIpZb1Dag6i4YA
SAg5q5hxPkQ8/OKk/AUw68EUtYB6XK+0fBHY1a1XsU28hMQQ5nQQo5Og+mA3+9pgJRRxOmlGxyvf
Cn633dlOTPQJC9waiIRRR++gxpseqOxw+GXiETTyDl3T9G1wsmN92c/US3McO3v4yo1Lvk5pCoaA
I/5HvmwdoDEpbRdMeCY3hi3Wqpx/Pj0V+qpldPRcGyz+iMf2MOxwS1D5266O+bfOYf9IlzxZANgF
K//IynGEqeQB0qMKLrHtyTiSyQhe3NrBsvy3g7u3Qet451tC45kf6nnGdYfje9sff/Ls3kJXu1CM
1aWq7qtoZZI7xE6nY8sa3sFitmwnE34e8XRA5Y74WGIwPjvcVuc8RSN4HHaoirYkl+qwEjqFKbdS
9Rz0sMUiK74x7FjaxKsaA266FUitwK4apyizsuLuPhx0jkPu166t+hbt31BAxX5Z51o3m/Yaspze
eAsn8cB4F5JesQ0INEA2H21Ypa4OXYPxJLbX8iPkDBL1z0JqQAe81KgLJQJTiHjUs/o7LMOajGwD
ffsIo73xHXWtWOyjSxo40vmgNrDAc5K7JiK+j68/vEMBNFA997wh2l/Fuud90A0eVBHMrM6hRsB4
eFxaw7uQX0ckbzjbN/eSqkXCtE6eBKxt4edxafJMe9Fww82o83qbT1z/CTXD/KnBI7TPEDNNJSCH
mvUfA3v6zzwpv9yJlyHyUxhaZMjTj/xWJvV6xCkeC+VqUBv8Gfmo4EL4VK5ZsDHjZN0B7FL3W7Fv
zW4r7LHFY4tLOg4raApEJlfS8EIEQbPrBzZkCWgNJ0CmsilekSf9uwidI94Ya4Wj+jmQ1H3ULL3z
ymW01HpPAynM5ThJuyMlj6tTEXTm5A3ZYzH/EiqhC6pmp6y76vUMjLo0tkhXzS9xZHUfv74/pLTj
xH0BD+piffByjOjKo4TFIr6pbByhsTHXfuWtWZXwfm3sFluivZtCjws6JClYbyxvlGGj/E2AEk0q
GAgUlageROwi+dW16RsbzDrQvndiQOPUF1iUSy2BF2W++riKH2O427T1rNzavgEND6Y8/YbOvRdC
N2O22+NpxGFBnf/ld/sYslnn8TwclV7CtWyCFhfiQWID67kEgjGVuTBQhqzt00lkGf4XYz3KSbvC
3Ek/O+EEEmUWJa4CYQNUzuDZbf0/6bg2sOxhRf1UDqmfXOXJD+Jkt0jgsWcd623vvTRzdF/azcIH
N7MuELqiSQdtOIogGf5ce5LDVNoB5Y/zdHa5C4mEczJNCiTlxHEx2bFBh9Ddpd59zfnV5iiDruIQ
lJ+o4yyXw2R2bnZuviOenIiCuxmVipkBDIH7cCa5fZRGNSEDWU48oEIN/FZ4zt4yx85sDr8h9b/L
yc+rYFYpzjS7xJCo+chM0bcSh/5xNUiqQwHDblbXNS9144nePmmXgCMIk/mngV7hF9EOZtLFa4GR
owbo413hwX/KuVIj9B6JrBIfKARRFHXSRggRFCEvAy0cM4D81XesFLzmZAeaDUkUEgBfieJpQG1k
7JZMbnnw5g6NhXeLK/RfP3p43o5uJjb0qZFI/3IBpmHevMRd34j/KXTzXRqeZZM5mmdQ8mBg8TAG
9Qqij1vtsBXU+dS9alvC2mFA/wyxmnuCIxz+e7UEm8DDg7R0CfSlK7qHZGArNmmPbi+4BJcPENce
AQg4k04D2mZlg5L/WfL6aFoX3bnGaXS3je/hsmneIe8IzF7AX4bpEWEJlBBDfKEeXqDJLEQkAJav
djiW8ZzHZ34C7lxgZvfryJ4ZhZfGVvbAZees3rxKkdjc6EnG27DgYX5lFl8vfPesog9FutepvpoO
xunN3v4ZLF/jExpMJHpXSSnoVJhGbIeoAaQTq9nmuqKA4Ev56hwES5Ye1LIr52eW4eInrHv0UzYq
hbU62Ea64Y1r7laG4xgfJ81cQH4ui+JdmqiyWt+0PrMhQfEdWVc8f3XyW4UKy2LROYc9I1xag7Jt
F2L2vmyWRVs5QM5dTIze/3+5QyE29SVoEsDAxLpZZbp6SyDJlRFUeD0RuAcKo5uQbx5BWLjrGZKo
HlTYPEQ/tBC/JvsIhsoqNy10Nj2TIhH3b4RA0PaqBwhXEsWAiLXXfoSacAujtLeiwUzBaQKL6mHk
lNhp0tcbbnaOvIzB80NGRMQxlW1BbLasOa1z+O503lk6i8NLMouXoDWXGhJ9s1TCbEVLUKVZdEei
HfeyvD06fv3SI/d4uaodWvxW2vOGZmC/y0AF4SNw5LRbxoIl+51Wa7zhQkW548cNDpCOUYRCd9jf
9KIqL9jaSMyKFIuK/lRtT1LPRArtPdbdCG2RxfeEjxLECjxrnvzwAdWP6xqiJGKNhszTuivKyh3Y
Lhvto5OhDTT0js7dlBL7CBW603fayvVoZXamPdBk5Jkg6k5ruQpcg0nLyo3lFdzcSTz7CyLVJIL8
L9PyGjV9IGzxk/STjbYrR5J+39XW3JdSBmenON4rWB9Jv+6Mzt3axoXq8KfdG5I2eD4iX2FbL6FD
SaHcIAlOVLQhIixoVfbJ/Bf//fgWGcQAGdsvZDP3nyiSMiZMiBUm4LQDGgBRtLhc5l8pNgKbxiES
ryeyjIhnlFPAjRcECGLqG5xM6fjb8CGtn4ihOro+0wT5BSFL7oKnKd+KsP+0zMDjgfleZTVmOiwG
hzJf/QbEgtkZshjVm3dBhfv30hfS3WrRFyO4KT4Jv8k4MthRtJw5fLDZ7lRU9VgNeBoZjGtglYKh
EiGCV3f66xb03nvGBbE+XiG7MHzSzIBpjHXEPhsHzZ4ixR3qrLqg7uhvJeO9q3Rd2tDd1VqyYn8W
/aGGOND8lr1xjEXdVJo1Qla75vJe9TnfqNKEHf6xmbumrtYvllMINPKVGpIqMI8iqUFuFf6qMSFy
PkIKNPAyFsP16p5LU9vPZyAbGroTo5Vh6lF9eqtxqdrFtGXKsUBxDQledEhcY2QPFt8G/gsgNdoc
rHf219+0G6Z1kUdEpUxRrimeA/ryrcAVjN/1JLReMH614huB3l9TwLCTeLtIrewsvk19lIOyWbFE
Cd9Mf/MV+kcWvzMcUa+NjD9CWa8dtQms5R0ZIFZe8jKpuj9Dlix6v2L8pg0uCWo6/v2cAcgelVr8
j2nJaAJoIbtspyOTXo5h8bUG8P1eGuq9vVbaE/ikdXv7WOg5RwEe+SOdWef7dn0wlesHTxZgqwWl
0LD4pZt6ZePuoyslTYVIjvIuMUC/4XsxvrbcjZiojdCc/Rf8GvTHch6Wkxwa16HP1fL/gCb9GIXS
isFcJDT+dtekfBNKPXJRXkOBmkwcB9ncBWVids6RljyAFx/lzEwhTAWxkz0wb4/2FF8eAh8j+8H2
PH4Ezl4Uca2omdgrjT8CjXfb7KlIcjTq/rwgCirgiQwY4uuHcjDbPUT/FFt8UnH8tNU7hFQKM2P5
s/xufqLV4YeQvmpQhX4sdPyhL9pA0Lj9v+EAKpny6rVKWJR6WjtOOjhV1367JxW+lF3Gk9fL+Liy
7fKxka/uhjuIbPd3syOkoSF+GTZQo6V7bCr4J3h2yZ3JllMMn4wtNG+Z7rX+pUXmWwNeal3VTDm9
ImNqeWJaCcSckLeL22L02eBnWea2hZU2LhDhfLzBHXqEQX5rP/g36J91L0/iR5k2UsI+LGh+FMz7
5Vey+kqqGpPiEB905D6qtr3I1hDYCcWQP4ssI4No+pkAM8j6YQgjxuOsPTah7rI7GDrHlikdcADV
D3MPb75qeLjl247bSFtyrdwFlMQ0SCifnDw4xRspYwWuBHYj2asfetcnwTHBxAHa9JfaXMAxPPz5
lkyUz+W8IH++YzhdqQj+8e95RDFZYb7+4f6fGP6Cztc7NbVrQtlEn6TSxFEQIW6G/Sb0Dh+nF9QI
eeUl8fmD9HHuDjjx0w+/0ojPajydqSBWOu9RankYV3UAcj8IZkxD11tJk8U6sacGQx/Q1tkHjuRG
RFmEiUJsRitglC9Oo53xnXmHWC1ZbKX+9tRO9C2E4jR+Wwd9bPqLleZWWL8wiFKjTPpGV3SEBtxz
asAE1KZAcbRqhtiT/edRFbxycgBmCkKGyPCvbK4nv+DRaza25unXaUg8JFqK3qGhmLwbYAo8Rf9K
ntF6nb2Jtn0hmL5Irn7e98y0cE7OPJXtHgGei4I+T1VIuPttG74OB70jEv1KvCUYzJAPCGmvptAL
JB6BD5KqBL8nsKTfRkzo0Ve2X8WyMgL0PnT9dpVHfLgcRcmhOsFece5qgLV9R8Ah50B2Swr3WgYP
FoTBgXrqFBPGLjJ+DJFMT7HqQ+5r6OsYeujAmIKwm/utJ/lkEReN7KJp6Hf7wJux7b+2GnqIQsTr
9ez/wHrUM4G0t7SfBhixgPbnvVlzoVr5OuLC5NHQzG+vKfoKvyaUMPIZAIUpi7LLassxqv4PbrkG
fmhS3hIsPMuR1IrICbP2RidEmST+jprJh2U6rcgOBN6d4X8juMtsmkNa8VQlebltaYgw4Nj0f5+u
H2RUlQmSBsFrFR1QmvXczq5lDZVF1Ws4eDE4Zrdd2rGUacpyUsjAOtZsy8N/YsKmHNGuq2jxaLVm
omJW81MbVxxtgq00YKxIFwctOETekEo51auz8lYTSivOmWkSAiIGEmJp9s/Nv43obZ67+1z8lFII
z3sXXB7V5uLJcm+FRmFYaZwyPMW+imRBByAUNwlVcVqaBILQ7tREZNTymyy4g0qD5QtCNUJFYsJj
tIobzFo74r3iOZYiuAUZdpkHlIzit2l2ylKXamlXzpJ30ufXdRxGbFM75Q/YzQ6aFAdQSU2/RcJ/
VdyS+M17JDBnVcM3wYM1fBxc1fLsdg91GoG1syFKsy83YXy9cHG/Tyf7TNTQaszkABCN3eKAl3mM
Va2V8rAk6QnDBYRxNrJoBcrkTtI/tuGrPJTkNtJZPPfoSlb7YvNhpmZLJWES/YwfW3ofX8lnWiON
tSQ5QEdEAhfPOiFP156/CsjSyNO3+SvU6x4IwyIG1drFJ/vDiO8Pr7sCaGXgcVPvCjYmP/ID5Mg8
qxrkSmY062kPTeOhphaeS6Asx298TfK6uTux43bgpScD9NJBKBbVFEGzymPC/CHcbEQgt40yFVAo
6DjSKpYsUBDUBazTwaz3boBTgu7Beb9Bsr1POqWetMk3lvFb0XtvxsyyRvhw5m1D1hPI5hRaCjVQ
SV97Bz+hN8XA8erZYDegSmIR4o6CnjwAMFNOSsNd9qdch8rxg/pOTZ9LrRQneiZbyBTBl6ooOvun
HuHfsZ1E3R1Smu/tGRxuqIzBez/4GwREiRkahlbdVc3aLIe0vU+l87SJExo6mhIjr5ZcTUBg24uZ
2xYUNU1exBxeubEK6XGZcJv36IWroPpMHqtoljs3qilhHWu7QwTAt10yf6gJ3AAkE5bnrOSjHd5a
6gYxu4iEzMRmFvStowph4VDrPyrcPMrwgwiA7QtpFtsfQrtVuSKdvzNmIFoA56P/KqnKGTE1pzpA
6aOmtLX20BCIcR+oLfQ4LY5kJZBOZCh5IpH9aVGKDoodmHxCECl/jLy9EELuZTbSF8CLwbROOjr/
orIeqGcDt6TZnZ0Q17Q8Z0vR3BbZq48qkDrygQQNJMSKVFOMhENIgfh845FSLcUJwbIwMG0vBN2s
iez2Cen15uHZuB0Lv77c7jGxPylgGM+tLd0XQhxoM0L1ZASllJhJeHFOFF5s0oaJftJzionns3mI
uVn9naP+77ffugV+NZGTv+J/vvWfoHrtEx7rUHyaSGeOfSlPO6xuXdnII1gJdUqI0vpLztjKJbtI
aSNsTsAwel5srVT2gWhJTEtxuOFFyqhiN1YOIm0AtK7Ie18yPMkcvDOXFxjDn2C4cVZQ/dby6/n5
zWWAMoTLdsnmf6MynCvfdt4A9IXMWPYmG1j3WTGejIu8DNIiAp465fJ60V56wpgOBLuj9uvZpg/o
ecP33o4wquoEKRehgD8h90tTNCt+1aIi8aiz19Mr19pEZ0ibcjluXfoURGXjDvHmPPHRe7Rq1Vp7
b+GWnkZMS6DDV9B2/f69ydSt4saHLMhYajTeMxhagBR7hB4897Eg6ZX7QpRgwkrFiUAqrdeE04m2
KvDHMKPel3231Ce07Bu8yDnzQ1yl01kpT+sqKo9ZpwliI2I6wAGxVFVih2tQEMKVclce/t3av/ba
u/XCCdklZxlv7T17pCHFjo7oE1n9PN8JxCytwofEaNf0KYRvuzR/kTYi0vcscih7LVH/EEM6TJFp
Uk5jewYK9C6beNUmGal9TkOQhLin3wVFXijmAtil9D9l8WKqjyjgjsuGHlV2G/jq/mvaawc12Nf0
iJ6eQ+QYl05qO5vO+GNngjr2VSS24vfZPaUhUE2VsNDVB/AXvzQ4bWl3WcfH8JvQ6aBctRv2dDWc
ER9ChscTIX3BciYr6+koSVCZNL/u4JYsy/Z7sw7cm/uWMCBMsUUNpumg/MR6TJGhfN81Cr/KIOC6
S3zPzeCqSQd2GAO2JLzl8wPdKueQBvkzvSvUeSSbe6/0fHi25aN916m0WLMOGd0NvvUghGXbn1Jx
KcS2jTfIDaYVByye4kLJ3wFy/PjGr53UYQ90fqa35TCVuIRrzOn1F0uLKTHpvDHSVUxDG91QEWdO
pZV4GmSjNpVN9y3IkHLwp4a9OwewuXWTpoJRZ3a6RCTgchwO9D5c+Xix8FmhEm6DPB0gkFNdCwcy
A7l8IO+SliRujCY1msVlsYxArHg7g3PgpYWxg1eF1wfwe5i6pwWzTFMM6WQoRfYGeGIzLw3yue3T
V53qZ4kgpDbmEEhy13WDap+TKc1d1HffqsAytJLs5arirTDwEjWTw8PV1KoN6WbbxWa+oAJN8+on
euiHJ5A6Rg231XFkX4BiEP5VAoS6Mv0duR9o6x793pV0cfrSG32CBtyN6+/XBWorqBsnoBdQFBxT
VcA+FV5Wwl7ZJOG+C3e99Cvm1vc6Gih7yV6F20XqznsEVDpITFcDVPslPwh3Fpd5G7eJ6LHtNg9Y
wkIi1apTniPVQpDHJiMKvZZV8P3k5gcMbGveXD/lBs6E3nWvL5gbXfR/R6cuktyzgxAPpKiplDdE
A6QSNWVV5bbWW2O3oi9Prwb/SkKxyiqdirMTUNfHWc9MG4HycKVZhGieYVaLfWZX3MzssAk207k8
haj+cVDXBzyEVn8Ou57DkZm2ljQtcJU8VkYjGrURkcqMh+bpy4VM32SZ4whzaDUax1qLvIMsZJ0J
yhMav9bxl0wWxo+D+o2G5qZVHJViMKhljWDo+pVzsMw8q4P53OtreeLoAnxvIDklQzU+yM/PEThU
1dhqUYNnhReoLx2nAvWoGH9LJgBn5D+rxqyVqkJphSN4YU3vDZLFf8aC1bAzTZWWFjXKn9UH+ZAe
gu2coUz87fg+ukW7T+scZpVs4kGc72c8hSVxvVB1lIoQg/QcxHPn1Aue5lYGe5bwMHtEMGx77BWN
Vu50AAOvdJXQxv0cGX/iU1XIpHaD9tsUGDjpjXBdw+fXOCYfbr5iuQVk5/jSP8GTfK9CcKm+wO0R
8glTmrIhcTcUkk+peofbONO8/8Z4GXDZAJo8geAxk1k/ESvn+CcirfVu6lKgZQvkzomlhTR/p/fI
Krd0/bDluM6fpCoKDWHKf38mgsnNXvkspUiyXlDrBLVvPqjlN7X0kkaPQzjJn5MjavznFOdmsM8H
VN9nKYu8cTFNX3cDIsodB8NmLKcSKSME+tJAoM9G5+nkkf+aRcvyP7C0jZLRpUnhYLersO8Fotjx
bDlhTBjmQJkKpmbyggM6zbP6urQ2nlywqpd2MA0KKLrcrKXLVh6VeCT10PUF7kGmkw9j3tXQVqiL
035+If4s3TT2tzYpeaBzIx2km6oZfkYTaD5CZUWalwgxaQnmFU374K88DkHJPmlAPOlEeUnIqrOv
VSdO/I8Cx0wBnsgrA9xpF18EDJU8IwLMVEacHRdBQ3YJVrCCiKWE+NN7lqpAese/5nVh2QM3HxA5
gBLIbEdgvHqJKM9fbuGoSsMXVljPJranOf7VyYJObuwDNzakBg7t9bCUxgQQUfBfVF2vTUotm0uJ
TkbxONgl4bkOJMwZ/mqdDe3RhwCy8EsmW4Aqk+D/WBVRn0NakN9uBNA4Z/bks2JthzB1IWm4qHhi
AyQzWNMeNNYmnqPWC2PbYD4vhoAw70RZWV7JtmWAFGe0nOvshiMmxZMlT8jz1u7DKOcvvA2/pVjP
/TWztaJy2W7iSrW8wt9sc+CFGg0aU8+9tG2UvfLY8tfqCjkUU64EjaS0piZTXQ451mOXedSIgkcw
NuLPeoFnRV8LKXQaEumPvWObaTiYUk6+hd/0rd5EIn72F0aln+l6S9ZrYTkrdfJLEJtQajn/s8uf
xlTvFkM9cS7idp5FI0uTT6a51ntBJkE6IsniGRy/9UMtobkqtBSXINcNSR2sml4jtXV8FGelbE6E
rsw4Ch/VS/iTsOJ/QcZxzXiMpsklrMChqBVjCbRT8JmZ54afscAb9a6TiAR/JU0v1ZCcotVVtN1z
Zq2rb6Fk0kXfProONCWPvJHT3OGFxejqt/ZYAfKyvEq+xI9vGeM0+tImy1YRXe/Ky6peXL84a77B
jM9qb3U4TWqyHUxGZHUzz2hihLsFWI/i0kxcnQPJvZKOif7PWpj86F9wnZ3RwjUX+ZD6Yg01AleZ
yolI9Ie1qtoIv+YPVeVfalzbozL7iYKAYh7yDhTyXYrAqLE4kFBxjE2S/1n+GQ7B/0WfKL6uXYYy
hTiWYPwdloP5GHUV3qOrC+0GzAiwchuQVVmtPyaxcmnQnmcEcl++y1+3T3RY9SsezjGhqFoV1RCs
dl33jl0pWSGCAirNTu1RB9w/TcUHv4Y2IAoZE5nA+Rr4CpvW4A2lmUxbG2+2XAsbNoVWdGTYZXDi
dUWmOfjCk+JHkuIjnL1tbhbnKYyaomYxKNx6tvALMSvxzYepBaVKLi7aARZxk7ASpn89UUKNh2qS
rxEiIY/avS5u/zW3yQfA0aKA4hzjpO75YzXJqjwaHFk5kwO/h6oEpFAbocrJibcVBat+YfrWPNs8
A6kSuypDpiowUHUATQZN1Gy0tm7TSFyM2NtDqAX5UOsfVEIiPohF9rGnZYeJctG2Ab/olXM/M4qA
/LyqLy6CL5Vtu+4BSiyeneIJc1jX9EFZoVydXFoVO/lUVk29nTVvROJCEANR1AEToc62rPuOt7ml
8lt+HfEJyAvvDrmjB/bVdzOAt6Ge/KQVLdf2TKGczlub7gLyv2AM3cpC9AewBDnp8cbKJqCJGriR
lXoRHZ3tzYdJpGCoDTLvGCfVvJzQE95iq2M9eElZf7thmLlb0WHH2CkcID2xe+zEvXFldJhv1EgY
VG5+7dT+uyQZy8qiOU+yu4F9xsUcTqcgayMK+doS7uGp3gupBYqitG/RnuydykhwfqpyziuGal9k
S0OJ2rTY8BFri9PFSDoSOv7cg76h3mgWid54tf6rQjLtt+RqtRvkDmsFUOC+ziG11Rr7GGUwLND3
yhAsdiqGtLo5y7Vq6idj80lZi/NhKAE/qr3WAMp9RiAvD8eyTAPaQqwmgofvWs8WAk/J1pPVIPal
D13Icg29Hfdp1BKc+tvytq4v7oSKOzzdfvd9/SrNpT+O/kbR5m1HLW+Uz2A3EyDwSWq5i/SQClvV
C7WImj+nRyKAYnsjrQrA4eexmLYZit1ESabHcl7Luq0iuqC7hMfm4zoi19rwym3iSoyfUp91bCiO
9K4n+li/Uuv8S1CDInf5bqfBkLWgTsdqGLMSUiAqwKJqhzbvxHj9GUeaDdTYWi7r0tuCJYXei/1b
fCEN40oS5wRsr8iglUn+klRcoy2q2P0l3XPXcv+G4nByumyAEY1zUUIktsniqK79TGj2qZsy+Pnc
w+Y8yhkUcB2V63dz/paiZAqo3o+jE7uRxCAUql41RNZoVJzF0/XO1TfHSSjjcvAj8DSy22TIi2PU
CJaRdnZm9pkLobUxo1qZx5wZS0k4CojsdXosp9vXkQbBjwq/kXbPTC+HFeYfPjYRbKfbcDNL56d1
8+NnDDlZv42+bavKGNYSDh+uY4jnHem33Q+t4Nm4RrBX8dYIBfFDBrku+kBQm3j5xQDomrjtiBdg
16v5uwKqax1fj8AMO5AjtB5pjlaUInObdLmbgcXl2lmIe49PlyP0HxhrldlSVSSCucILbbJO87yR
wNVWDaxy/9VmMcjs0e3SEXZc5lVomczhMC3cN6D88vcmJiVy39gLEGHzgoDUC/kW0Htadzggbs5T
ll+5Mu89CGt4zOUEk0CBICyQfjy3t1ys02NGj2wQeTRK5RGOm4aHORST9YONUJ2T4SiEFMUSWaHe
ZoZehRITnQLubC6u3zQwTmeS3XQo6HraRyCFFFeKF7gn6LdWOJpHvFZAoeca3E79tUGSwJS/xrQG
LsZz7VCJ2r8DDRYJkR2g2II40FmniIigTR3yoRwh6qSZ8Oe2K+0CBzQboCcT1OIxQfGdbZzdv23N
Riac2LEuhSyNQiDGm+dpVV5H6JPa8CglSIm/SL7fR83emmnamLkrxMNHUCipzR4BA9dvNnzascX5
xemCwxY5NZVYm2lCnARNZjrelHJjQXvfDpGjtXhTrrRQ7Icl+v39PV5gHF8Gin3T9wJ3NmZEIHu4
ImHpuCEfnNCTTSATN816ucBmq3hluQp3oUOUpkqtGneNOlPcjyVgTErCTiL/stwNk8trpBg1qaWa
gsHZtbYO+QKJFlbJA0S6LPolYr9iuqrLs8FFcGM86oo1gQuGitoClQHuOcM/vzFS7/sYWoumWDXo
wBqkIP+ADl+lQXUxIkfBiDP5jtDO9Risw8mtrpyjWRUJQiOLVbSprFkkm7GckMGr2+08ugWCdmFq
izeaU4Jtc5AY499E5PREeCiGLAQgW/c9F22Yw92crn4GgfN88E1MA3DietnT07GgRc+6QQyDXhFd
23U5h+JJnxOZpgP+ldW3tHL1zdFsXf2GgEXyG2mJIl0gBtu93oFLiszq/D7h0YHlJHuMZlkcFJVP
8cW2Nai4Qk+rnc39w8GzTcw6lUO2AltrN6XLtN1zFXlQgjBr6ShrRQMBThzMmR0DSyi5ENz1XczX
ss/icqJyZuAn8J96b6QIk+QB30Ofnc5+1MtpEBFA+Xtko93CW8hUp8atEiYE8iC3fCJrExgKDVrK
8moP6IpIeYlFIIE6fVfbLRKr7xK4wqOvjCySF9gigKJR5volCYBWMN4KABevNpd1pOqQ8LhG+1Jj
I0PNz1yYJScRIRzQpFPGwGDvj0p49wH/1+vnyzKHnjgY4n1T/+azdpcqc7Xu3S5cY+eXm+3GxcvD
JyrGQfYEdGpRM7EgEp6bhYXOPYvePzAZRCvZ8L/D8uc9xRpERskU/PTaPmvLglSoqAwtfWFJq3wp
YOgdJgkcn2s6JGu3v8Xr9hIxIE+ClSsUv34QTVboePGi0dvpFrJy7U3SoCZe4qe63TfPBuoH0h+6
1YeYA4pPDDAkVOi67W4T+Ty/I9Wd+xgDnPY9uhZjwk6a/XJVu+RVxZhraAa32BPdqOrWOp0UQfy9
extB22HRPFCKY/mF7wYMKVcR/cncUmiN5WVDssP73BzkfsSD8vUMKre0wX5bUYkr9OCs9GmcSLnD
u493c/lcBjYeud9aiSA3ScI86fAvigTTlnfdiPUGg26nMlz0FScR86Yk37c4GGENk1gxFJl0sTPm
+brFmhQnATA1XjrPHLFwnz0V45UQt/WaGZFOxVFUfvc9+BMnLzve5BtHC30OYPXYb17w+6PIc29G
ArSQApJ7HIhk2D2xOIwKUjDwIxVTr+Ne1CZdaL2Nv2ODwC3eNZccBPDFjNZfN3HB/0ZjyKDqCtqS
oJn4GimuKZHBBfgOpEGzkS4aywzjrZXbzbr4rWiW1FiFsU6i98P6mrdVJ3zcBiEUn5xyNVdOivo0
ut8igeTsLuTeQ/RE8W6uYaVWJ5EP2pKivgN72b3QQJr7y4r7z5QqtTYVSx33cwSWIxRC02RVGN8M
gyYLlVvQxUp/HRifADkX12iuYYUIjvf7wbnGmY4QgP8+2R01wjcSea8hKcg9X2jpYVCFt1DKu8qB
beHO4OQQXDbew3NnfSLNMqVUdjXcmy1a484i6+TLgcfiMpIn2SaRqEtXCKd+u9x0uFR4m+ql4eqQ
QbuHwaPPI0v9Cn3iKR28bsQklbAoTIODCRFVkSvPDI4kQEUtR3FQwL7F5MRYlJMDUIASldXTilPu
SiIZPXoyLqBxRBJtH1qJoif2C7jvaWN6uYNbqSF0XgK66Irw4vkXu129JIsq2KQlWf21PHJky03z
/6u8A6gjbr9g3yovvzWdTRqvnaYBK0Jwi5Vpnffh8zGzlxu4Wi3JdsN+v0gUa+rEG/yx0weFdKQD
desrRXujv/hWrksfmHFUgEGisO9T4SpcObunhcwoKqh1t46ssOj0ZESpa9BlaXZLlaIxMsebyDRC
HkWfa1zrRxZ+q68J0oL5LMlocOyrQieNIfHMo8WiNj54i421w0zxo+kjIvyymI2mHdXntOHSQRmM
SSE1HZggw/ACDLRQY7rMXBjFzfcEqdlQb6vQ8mAI2OOhq0QDoextZVegoBYqRaF+KAql7K/lCT4o
APqgx3KlySvvztl33x4Cj7qZb3wql6way5v8GBjGfHz89szUYLLJwcMkZiHlveYLXY5qicQe2w5P
NW2o/j+hv+NEXwPY4nbVNiJqdsOgPzeZgVaYgx9Z8wITAX29Woe/RFT/44zxN5IVmj8mdyxi2pkp
DrrPD73PymTu54jTnncBko9ZNF2lvLlUDxo0cbbfioYFAvHgQ7nwbUHwXJIv85vJBfSBEBoiUf2t
EqY16x4g8aaj3Kvd0yHu9cJZ16ezlGZRQmwoQYXkPqX+gKUGLNg/V8ZifLU0CYrg5D7irV52X2lv
i02pf+v6keCLBtt0ZyYA11OTe4W4pIA8/serUnnY4ZjR5HgKaLkByAPIrLHZ5XNflK4Ap+knmq26
obopClLpRyPUewVqXjr9KYIIS0GpDcO/weOe0C+SmQS5KM9xvBbEdiJQO1KdgXjsf9InM3RL6ah4
JFNLJFn2C97V25663pUiHUmeSdFEy1Pf+KXIX7E/jY7EdH+Q7lT4HJw1RofYKa/mf8PpMy7cHQfq
qOhvRu+ARDCiCHMQ+olUUGvV3o91yHBUrV7Xaz1c2pJ+gxa05eEtNI0TP/huwJnCgxaMotMg1sKb
4We1sI524EouPgKDXYQg4IKVNW6HGJPRKxm1NKUsyg0bu8K2TRir0LD0eDcDSC4TyUP/qlC0mueP
dXpFdTmF2mPE7G5fBxSVUVNGkjKQOTFwli+4244PUEAmIuLl24FhI6beqVFSaSAuIoTpJnMstZsU
jLBh7qh8a4gd/jQiE0mhobuM0W8VJ4glAyT8iaVdIRbJeplRw90TNI3z4XVh5eshAWNumK7caCNI
buX2Uv/d+paZzJB1WC0RVN97A+/QDz+YHU6FjipkEoWuAkuYLDXjFgG/c9ppfv5Jfh9H7d8ntlRU
m5VkRuHT0PrAR8VwjrB8sooW3MotmMQYX7N9njjsscfPjEEXSQOLO77PaOAm3dxE2S56kx6zf4gr
ZkKva2UCmMsThHultGaLA8m+G/JSFsQMD03pCXMSLUIpeGDIKw3OFQtk7OvdpPAxj/s/vye9vuHh
Uc1ZCdbJPHrVoVx2YPR84H+sefM2U3xfp1FB4JJ2kyG2dQxpc/sWenVL7z9wtcgoFxdfqXJz39KY
YsmcbQ96orQdfgmiSw2Fkc0Qtb8Nn9NcAA4/Y5owzag6/59vrX+mDu662vQ9h5/o+3DRPEcqzKxK
xRtJ00ZFgI7b/BM2fNsAF4cC6CHAUyuWHSii9arP2TTKDygey4rh3fXVkYWpvNGhn5YE1ofmqTKA
uaM18QP92EuhqtjQ/Eur6TbnmNYkJxI/J3VNArByvMaeHiU4HPBdSoIdAyg/6IUvL2cRFeUfHW6o
uFpOPRI/sYDrwJJ8JdJisj5XncuYhhLS4IzEf9SCRhjT0OGN94GgRuDZ9vn9fvKsbsS/JnqUsgwR
CcsyQ4o58eQnORztc6ZWLUOWTkJqFtZemugA9VmD2zcIM2QVpYHeoLWdyvF/7cmoY+LSpK9UvYHs
vL4wSiHfyWpGkk9sbDV435S3p7RwNb1xWfOmyv6DX2Uvcb4D5mjv9/mlpMtTdEn27dyEh7iYPg91
LPxihbKAsRvI4010rnqQtnTt7hsF8mjddgfB4HfzPvtAhj078H4dkQ2oAODfpu2RW3OjM0pM41Su
ajSZr1mZA0WdZSGbnhwDDuUnMueiyk5KCVi5WYjVVfb+g4JOgXXNzFAZ4/6jkvNqagWFglP6xGTX
ocVMzx6+E7WPSKCUuP1xnUydIXV4/i44QaGn9ekaW+MAL++FdO3ahfA6+stDxsG1usdo/QcbN9Zk
cIM3gF8o3UMonSP6C9jNLVkl1qQKDobwk9fARl1F/QWJJJZh3IPC/aKjof5V1DgmLIQKJRTbrIKY
W1WD4vZ2X4t0SYrselTZx953ROfc/hqqXshBvVcGn4H49wyYOwJbBCQxyULgSuUP65Gwdk/nFdO6
Gt1I6k7sbTDE4RGCCYi9n4wxiUUYhTKezFg9EVWCnZ0KMEfEeoHkQDKYrxBThx+PcTUd0xxPXZd5
Vvl6e5PfcwyICcnCqeUQgJRwTgLOFugsG4IHt7xTDX58HgA6UiQDBU7VwL1hgJdp5GQJKvUuJdcS
rKLVJYnaoeqcN41ygh3Wyj89k1TDooeh4fkZJ/XconnxjUZ/7hbBaPU2F0dEI4r53szCYGNWI/Ua
N1EicDM8h9jVK1ZYrVgh/9l5SobjRs6QG0j66MiqMTVppPahqApN1P7LznuUAYKZgBP5pH9Gc+Dv
mfkxUj1oOzGmsholivAQRrOdX9TdWjtI4oc8GUaN6bImrLDMz1QkWKoe2EP6GbDFyE0ORmLLRtEm
5Wq+oRY6Vy7zY3Q0uBkS2iYhz7XTtSsF07WR/gjXpmUMw24ok5Wlfn4Q7PFqEjtxkb5Mw8LmuPVf
ecCnncAAAsljEWOC/sRIYtiV+9+wnqIt3cjeqUDX4FIsQG8vj2HTnC54sB/bL90vX+WqrEAeOtYw
EYThcbvb0SCFuWl5eaTqbfGPafc6xX6qvgQLDUl7A8ty10ONZzLgtZ4zgVX37PqxmcuCJNKPu+ML
VUt0k8PUY0lPMF1ApShgocfNT9WLsCIbFaM2StzvVRO86I00jv9XPT/pvdOuUhDysSbfaE2bRJzN
Sx0yXuDq+nVWM7zCRLRIiC7/tpsKNy+c+FPer0ErSNvonnsWDzrPzRfe73zcVfGpSajub3sW0U5B
idqlFJtqwDdaNG1GCuLp+bohTAxfAmzJwG/6ypOGZtWroFQlItY+ptXsQ/yJHQAAJrmsEA90wRtO
/9iG5hlVZaG0tujqbaaRuG2HMMdOsbj+UMb5Tb4XJS53V6DZN7B3hOG8yTg/qWT2XhE6XhcKp7VJ
R0GtQBSbWtsrc+/4bfy62Ks7IrlaLLL+GgSTH9691QZxC7mGQD2l46HONdWP7pqCy9LBqRJESYId
NqyDLgk/x5H8ZQGtwfiRzWE+ZvRzOyCt/ddDQ7m4W1vmNy7Zu/qJqfxn+X72tnplkPIzhvcJbJdN
prkEF8S3e+r4VGWfBqeK8FwgJa2Dx58Pi86JH7bmbSvwi+j+jK0J+5euSUCEfO71du/RehndxM5N
pea4xTwt1HcCyPpXtuHniiYqZHFhIufeYuqacRwAHt/scDphMeSe0Qvfa9fXFfgg4pZEKLC4oAHp
yXw3nd/17HNKsnzFjpKBZ4koQ+hQIQmW+50IxFZRVfZjKmdOGzDlOnANA9MulW2d/ZKZij/UIIf1
nb8A+8gkf60XDQt4OJQnmN2hTK0mfTWNaDJpJ7BGZ9BZqkN2+l6q0YR5J/lltrmIpdn0cpDWBwNX
DoMg7lg215gXPAC47Tlo4KRGgZskryZ2Btkc9oibRotLAID36CCrW1W8k5sYvlEdIDgv5vXQNjK4
UvyXowYgNKDUZsDaP+7s/207/TxFV2ijTltjxrZcm8SYWLdqXdNO2ubTDmB9obi+j4ehinLUM7yZ
prVeGUzfMme3uR/9vS1VJItPhyKFx9MExzyoOjStKmTsUq5jWAbDWKNUT/FKfCJqdAGNsQblFktv
vTVExzeu9c5SXVp1dekdoI0H+DxjFp+AyiHct4jnPrgZLKK4aFRHg1dofZ8Aww+CXIrMU8zXGODZ
1+SALbuKDjOHk1wUwZUFkLX5sZUkbG8SmH4ks117wbu3IFTCyaIdFDEAx0GNnSVFgMq3Gh+6RavO
G7w576nz041rv4p/iPKudvW0l2f43yj4+6BV8vC7R1CSmR3DkrP3jN8i9WluA4zpgieoNAoafCIa
JZ/3cl0xri5UGzfAHQczcYiGes0S5aBmUQjAaBpil7/IgOPpURL9xU8SyKSrVUZQKTg3g8oLV8HF
OyVMcndP1LmwiaPGTQVkeBh83L9FRUU0yz0YgyrBaQSN+gDgiQGjlahcedPFWwavPvm4H1Z9Niyk
Vxdufejq+B5SxcgtpbPlj/oX2Gjc7wZk3qbuEkyT0C+ZWO8YlSoqF/UE5O7xGfmTXKXpD+mlxm01
7SfTpMDsUJAtmQrRhrqZtkn7BoIAnNm2nVqK3WH6WDau5/kfw8rs/+7+LJKkhTVw2r9YtzipPbwM
cBS+BwfG4o7ZyH7QDslClCTvcGWNzsdxKCYKHoy/sOnoTc+qz/s51hijZTwi+Fch6RGEYpJm0y2g
w0Xl6u+8LSofmx10abM9MVkFCT9uWhZZkShn9ng2NEp6l4KxGZci4m0Zq6qQEUP02VXD2tSdAmov
86k1mDDkaLBtQFjKw7eH6Nl6ZYt/WdCHIkfo4rSNsF8hsxwlGJHxFXVBAI8VXvrc0hvl561HLYZ6
jjY/z4cTt9eoif1Lgfb+d/K58rGO4/PQz1peYrTSWIAIQXFhXW1KvFNhx/Da4NWa2UMePbl8Wqmc
F6bojFQnkd/ER/wDHUklg0F4ekoELU/ZlmtfbmgTC7Tb3eX5ucnZxMqP8ebNhgrdZpsdJOJDL9RA
kPUU4JAqO683shhq4qWWY0E2lPpiVnjsz7inQLla6yJoVVPwrpF624Aqh5VPTZCJHreTy1De/6XR
doXLlXtGC+k0GPLbjo/ufFPoJxGA6+VbvcQofV0Y89CxOJ86Fv2ykBU4TiLd1hpPp6vbMEV2k9Rd
AIWazZPPQo2pmNFTiejG0pUS5L1EZ5qALlAqtcvAygdZxZeOsHt6eq91GgWOXVUYz9pYo6OGN2GW
0+8pIQxNQaWbFWhDciiCyuqqlSruBvdzj11Nu3O4hv+MuO+x90HcUCkM6QzcYYSw60hy7UZ1x+QC
gYdr9bOZxHOltjxOL6YyvRDGLzQax/2JDqLNXwmZvFx9n2W/DfKzprELhLwJKByWPS4Eip5F8+jJ
UB5CjIN2eLO+FXHrsrAjgM0uMVlnyNnYuNBbm0QBd6na83PXIeK1kQ0IPcMKzRb1apB5pmzlFBRu
lf6bVH0vJhN3l0cJtnUZoa+icnNHOkCrPRCBk/ou0oAI8LDiRVoccZ1hqqnz8EBATBDaMuH3XdR/
8gX4g9yq3jzz42vTLAd3flIcHDsYUnb9GqNXRBi3wvQOAmb14SugqJp2W96yT7hxsOy87yWNvdJr
PWXduxP/+4QG1LrY6VQS+PpAuXhIzunPd2fdNgB2ai+B9D68HfHBSD6sf3WmlEeEI4WQFNw7QuqI
f05yro0cZVDRibebbPa4dh34G26eqd4YUHiDUWqCCirfkK7rZDixrKxCHT3clW2JrIiFc+r+wPnJ
7KzGdhJaXEJPr0Pu/m/3YXWSqJ+ffE7HennEVPEa9pczHdYfjFcAGo2BIcVIE2cWRRoGPwpxfvNt
4KeDepcgvTHz1gTEKN5csp7zfnvXimLrbty3AIVi14saZpU/41m3gmFvXSspFJkBqShlynV7CIWa
fzwVkY8ILEzTo10R/K2qrZNpiubiUI3mndY3ekv1w9qf38nDz76u3Yc7ClDZqPcJrIqFs6sntcM0
anCfJL37n5MHTUzT01BjIEfADk1eIoucfsMqCCOCBzCVXnQpVfKOvECiX2hKdkZHH5QFTzVtWT1j
5gYzfbJZoZrxqGuxrdfvOpUqGk6o4cDYWaL7jaVubie4poTpvhaQFL8zfaRqYXvNb89meyN3Vxh3
UOlhsDeNjflGdaF8pU7zxE5xxOrwmbEo9Ech8bymnavJrnm35834ohAFXDLTJEU010QFLVt3JGsH
seZV0jCjH9lFmjbMuItxsfHtpXws3W27JzHZpwVzBSIkag7xnTeP0xvQSzW+vEAeg/5KKwgpy99n
oDW8zkY9Z7vjcnMhmr0n8RVo33c5V8XUFobK4BWx2YJROVja14AbGw546kG2dJZJfTtAp//MYzXe
iKWDydiC6BgQfwnA7bzWIqzRYX5qUlich8MSLw7XH7p5EHNkbAobjzeBOZVgnQfTZRfSil2boeYj
fojTDfJKc+BzERgWuILWSXAR3waI4eA2lvKz05oJNbk57Os55bywbNRycxC9D92qQ0LM/I5oX+eY
ShWseWD/x0+8Jp46agpDO6nsbwue27TPnfGF5l+etKX9jJidaAHhiUhoHxvIuw88GdnP3/nfEub9
vdB6OmQHha3FBD9Ru5DSdtR5gGtqKro2bOtLDMo2Cc/wxbIJTIjqy8wu6L/uHKIYQYo7n5FLKWnf
mfmmdgpAM72RPI7oObt9rm1+4qdebqd5zUsF7hod4bcc4ZKbzhvY4momwV4kEAVsb+/I469hFUNI
NdtqeHtoDyuurAXMlj/ENsoCJYbda6BZQSWcCUc17XIq7GMmlWxRCrm0jAIO+Fc/Q+b5edUa/mYk
Ln6C5/uHpm4zxQIlvgL6aEB39Ah33ZgjBsI9hDXc9P4tGzY96NQqK6qpL/QIUow7JDpscvFcnDPP
tkPMSn50Z9xK+D5s7Uw3a2QOFrGMPIqHarSXaUQ9x8qJeRGYRNQ6aFAqXjN5OEWlvDSseNEEYEVs
yFr/e+sFVYS1u/gL29J5eBAif/drUwse3NnPIL7nWgWUh8rLuiMW+UkKhX2LRCYY+3XPwxY8E8Rv
1IOhOl/UiuYMFVe51Zey8beNuipv4jb+FteAF2oxR7ScMsEmK8YxeW8wmmB+UGOzfKYZp8Bkmnzl
BGTmtEXmbj2CMu50mTFjDwmN1Vtk69Yfr0kodeEll6RWZ/24zu7cQogS2Y9pnz9A3XoGm67s4tmh
4mdorPvHLJcT3GnAi7f4F050j7dFmrSelvomntPf8T/V7m5MZOGQ8BzIWUWEXx53kj83f5fhrdde
amXJlLnyGfg73+PopCWUdrgD+HbZ6U2SUsiALDL1hdlDDMEgjvbN9sVDTkMgk8EuaEabvcOE28N9
ZmCGhdEB2mMs6cytfMAKwSgeIydNni/Br32JfOBGo9su+b305bh3D4xKCyDmephszPZM417uy+Ns
g1qAOgYF/zP0uDEJ31gv6rkgFHDGD9ekJGPV1OVQNc1yiUlrpqBr7ZpH/gwHY8YKpuctVGqQ58CN
4KlMEjik0BUkQ6Yeigzdc2strg0T7yJ4y7JFwkX0Wg8Ccv//ao/pAN2NM9ivY5KpQuZGU8RPzt/u
UP5AcB1aFDY8xExp8KtmHZKk86ciIJWd654sx54EGNdKVZmmnYT2qZoLb8TU50FtaZaIUhH7pWwv
+OFi17NYaq2i5xkpKR/N8AnwIzKpWQt3VobRxm0PKhpz6g9zElzgOJCTbpa+X41u0KVRtlHnAYqI
TiFnZnlrjMkqWHzI0EWiFVqx3rH4ErlAXA9t+SwVCvynm+F5FptVgsI6xuejuELHma6MdDTFgVLK
KBQYkus9Y1fj21q+E4OaxrAoKAQuLewCVnamlZOGPNawElSAOiyt13xDKOgjhIalcJytiLd5aGSk
IDK0eySI/ZXENUpY3tggPbdumLePttcbx2yjw26ibPeMBxT8LJNhM2+0CMf8rmsiQOzUKYC9YhQp
ZRg0c/mPMTIJneOMRpSgY2CMgvr2UNHWkHYlDzeIRqiYawrnyM8l+br9zTcxPvtpKySK+0XmVtLR
oF7Ub/uCZdPeYMFnywx5py4iUrZD5Kvq5xE7UT5wJkZ9W32gvAId/Znfwi7Vptxfdz05s/X5ZWvH
GjRT7TutdZkwQzU6suqIggYNDrCrVwOm5sBmOj5UyHD2ULJ8BqajnJkaS3lh/CQ/urGU9qNXFtbI
HaBMJUupNl/kGr+rqpSgcVeXGYda1mex+C2dbHPCgrws0vWVZXskD8SfGKqiptiJceRA4f3hNWPp
jFqTdSLm5fj9HfewFO1zp1u17uvoR2Q/OOGmmwsWM+4CgJXD3hzqah/PNHCCjn/WK1nCIH8UEn6T
Am9FfoeI/ngTDgSbJxd3Ox0+1Oq5VdTQIKbNDlnRwpP2bowQ4i8bRz1VU+P0q9mWZUudvSXL3G0S
XTUG7V5NLtqg61tJ0VhhtqhwpyFssFBfqiA6aA2NQG8h41rixhXAyzEJpi2Zw73rUR8Q1HcOxSph
jQe6Vl3W1IEy0EvKZ+wSaMEPeBPaVBueaWcMx9pT/tsBWba0hAQypVnsR806eEkN9EASaBl/e51q
v6OeoqqbkDNQVg3SRwnd59jNEUDCsE5/AMaCVHbkFcyqNzU0GQJgcG7H1dc2sOxma7qgRLC4S/ye
4jA4uLOgq0+a41XFvUjnDUIntYXqlW+zR78U8bfEAXKP5IsuD7ApZss19y+7k5i02V1C4kYjr0w0
/G2SM+xJnS5XHbjWaHbLMHKqB6ZFgI7xH+GE0N8rolfQKQ5voKusXbicxLP9fGifjawIonvtvUNC
Yhl0s0nQQTawZIz/oL2Ke4fKOFy7QPeENbPtxNzYaK+OZ3wdj2pku+eJmhpf8CMZkKINClqfe5iF
4/BEp7lydyhoI6SkD+zh3M9Fgb9xH8Nt3GZIraf6Q/5CpamDWRxPlR3yrMhRHfciTN0ggmVymygU
d4xpBa9YAqXjLGEAyU3Y2yxp9I+XFigTRK2c3Fo5zlM/wCi8w7VcZCEHeihatrLGZsFwSAePCyld
SrKY1f8fQzeGsZxWQ0UoyAHwAM+A/I/E4joZCoUV9Rho1SxYq1DFnTCx4DYhKFjNXuPKzCrdk0/R
iYLHNa/PESPhG12x9TSG2kNUNEZphyZ0Vlh56lfbNh49vrsvfUidumXTemBjGoXs8AUtPc9836/9
oJWamv/mNUH7YsQqYR3qI03rdvToHlMNLZH4dxBuYOE5HjON4fCVYk4NmfDD8j11YKIm1yC2kkra
wN8FpxOWOYfzFbM6uEmTRJIbzrUlpedXY5NPxserWCYNdn0wCxAdld044aEPtm6xKEdpf/WI54nN
mxIVNkc2n7iLEk2iHeT3EWIpleXfe4YDVSBCE/nmvar0pL39K5p5nAVkBZ2GOMZcowddCv0+RV3I
GH9rvacEP2SzYPD+ewX8WwkGEZYegseEhqlp+p5W7JO4BewuihCO8Vaa1pFBgHM114iw3PPAfK8l
MibLIq12cBUiK+snRWguzzjYtKulQ+eNa76SbHMILBO2JTkisK3OWyfObf76tBqYp5wdqczN6Q35
roRK5BbmPsDGXhE/ERI4saT4x44zy6S/1o878hEG/xyjl1S92IjUjwnn/+H2mM682rbJnWPZfsdK
Tb5IHbW1l1o2aG6CMVFMB4KzCSvaOm4jPkayKU9uOx9c+fedytd/zcwqsViiX2YLBCZW7r1JSg3X
1PfykS6g0CWcSnkK4H0tE1NF0796rcLoVxAOkJq+24kimiJ2pe6Xkwro1boWXcznD+6JGSN8dWB2
FdDnO7nC4VZVHXreByoE0f/o21KNBz1C7rTA4PLAuJZI/1x8URo/GBWxvaQqRRbNs1M3dVYlAJbC
xv2yzoSGiKm/FGt8UxKGoVZgDWPcaaGNH3jexH6x2EDFePGjF4LdtUMUsJB8feALU3F6/qtkF2Xz
kfAqOaRgLweX7rW5yXceZSZA5TIAGJhIZJ5WxDnjRmObJq/oEssqeqnCt03cqNXl5aKHsOXg79RC
hP4pkhjRo2Xn1hQqOxVtGd22yETc17es7o9D0dWo0zWlWhLQrIvtLvC7aIFx6kR+gjIdcpOBrDbB
i1LSUexLhxNwyC+R3yuQexsyaLft4wsinprWTD5uyIo1+eR6QF8AcOiYt/hRwMItHF1kb3+2/46m
a9nFKRE0kZEbhDBLdi1UtSDKezyTiSh6m/7zeAsKVa2UKmMcCEdljllb7Vb+S1zh4P33yRNOpCRU
MwggUT4It198wxrxBgLe/m4hFutHDU2JdZbhCHp9uZ9s1tQTXZ80SYnGkegixv74VnuGLALSWnNt
p1I34TVjNSVniHP1KfPEEKenZ4S4lODfX1hei3+Gtv/7+jvTKHRBU/ZHeoYxazBsMgswV53lo96f
FGggJAGoDrhBZurD0VLvvv0MSAZtjaf8LtXklE5nLkpC7jdYrr8BzqSoc//pyJUqsWO0OE/qf51l
/RmprEYkx2qdsJpp6ro9vSjlrIsrVTLy4ooxORwNu9dqrmCJE54VV5vvmPK2e+4RWpeilBWUOwRX
5riXXu3F1rCap0W0HDsVmbBeIQano9sG2W7Jp/F+DZKLwlZhk4KHwGdC6K6KcgV9tQOTXfVrxO1z
PtlCEpSuIK6SPH0VKKsO7STGvDlAGD6Oe/HiYi41FQ8i+5PJ5dv8xGryupYKic4c+shNlJcMSzU0
s+OvVWnEoaJFTpFba7lVnPVyMG171ClMtAglh5eXa+S5XjE/iIzc7ZBGTPHzemZgPAMDNO7v7iAd
5qyFvJeRGjGzD4vj9s0bei7DVrYKFlLzwJFyhz1aWEtsboA4Jt+nKc37hVECqEFkwdBo+XZg+3zp
NdgpbwAB7Xu/GsyYYox9YZcdNmcwfCz1Vg8P18lEPlu23pbICgbU2dXup+6ag7FCCKkrV/e1dj1r
UkTRxcGnGvs72LGe6Ro5zZ9fxSq054xtKWLDfS/PvJMMkpDhEJF0sH1xKX1XKtCOzAfDtUxxyqG6
jkGoLl45+KJpmCWj9trFzhD0AXB/qZKjBSYgl7LsGEqt8cJY7+7RzVwc7qMPmoUvIndybxQJyJTo
PAR1GANXo2oueVIc4H5PEQdcf8sbon0THKS4zbwyXBntnClz3RGqleZJxDQLeT3Fmp5P5vdyM/WV
INvKBD0u1K3qpxXAWbZ+NNfF0tbAw1NXCq4VhrCTNy6J7AKTX0DpLUPyHIPMtH1zqT/99/ItEmRb
cD/7W6pxB/Pfql5bM1YlsnDQNfCItbovYGheZBoC67tI9vOljSA3vmRHNZg51/pbxSZfJ7pyFeJO
SPGHZmjE3kxICJwgUrK/eBgyYxnkMTDFfLcqYF+zjBSDL5Ul0N1aKgTPEYdXO4+DVq2gikYgQbkI
W1PBhrezK9irkgJFcs3ZfNJLULjGz0qvPPxroNChbGxgSO+xL+kGzXqhCIJ00EB3YaFTaS6prTqJ
9ZlgCTbVWsjS3pz7DpgHsnHeNZRnmdfNDyQX11YnltXLL+MR0NzIy0ONv4LUKRSVir5Jmzlh7/MZ
7ZAoZJzaCAcu15U22aTwjKIBYbTNYWklhshlyfyiRvyOn6T5MzHyAlMgb9cssLLQt1iWroMDB8eR
9VVMjuGLmEDNZ9EX2Q5gpDgX92EX5+RqGhMUpJB0bXWmIEfZMFOx589YsrXvgJGs0hrbZBVj4r3o
avk0lnWSd8E0hRFSNIbPjqz5bBeyioof7jpoJZ4pOS7IoIlEHuDfXMmwXYzyUvHKDRb/XB+xCdK4
OYC+wTwrWvwn04/pbd4heEbhsym2I4Q+ykSmCTku2GpvPJ/UwkFdHESWEMWx4yQprAmYxRq1Fx6V
4DhKsZuZlUs5pPedqWUbd3OIOX7thO3jkVsMrNk2SkWuU075Tcf/QsQmi3vs5u5w5F8xiyp5xa6a
G1kf49xFTbQ6hl1kc7gq5QVhuBljTBErdLnbe5ik47P9Hxg/58Ca99Igikr52hu3zYYebBMQUBch
tenvKn9yxadmDHCtWPHbmzFHNS7qUb4xJYVSfT0yNWgXcsHUPsrObg07HaafpLU9NU/SKyXG+mbM
OWAKUqJoMqrOhojv03OaJueBQ48ylXmhTCs4rwNgOky/3am5OYrmcZpJbr4b4QYwIlo1od4LypNo
bI7Bf7SCCurCmpEbpvwPy8o4Zc2RCV6laqxp4TFmI9i/a9IGhtXwtLlIGYDwzSh19nl8Cm25wAio
W0khGbLlkDWrpqujSVKuYSHi1ZgTubqF0MtJwKd9tYnSWx9dLAFpF02hzVIgAb/h3vuYL+EHvpQd
I3tOnptg+mG6rXBXz71a6W3tpHQ2iWiOwJIbCNMIXwpZbE6rC0Ro3HMXzhyuTbfroE22vdsIAR5b
6F84/8yOfftGFMafEeeomdLDmSwPA7nzGt7QxXo3msgE5o73sQpugHZiecU6L5IGDi7F96WvJHUj
sgWQVL3/Z95Z+U2AUVc9YWim1jjINqXTejPSSZayojOwBtbSHemM25bVk5+FzauHHdfDZae5BVNK
esIFSX+R6em0SdYxcWxufrGM8fkcdjixAGHsMLPezllrlOiu+6Vq3mLZwn6m4l9qKCb3thItTIGR
kaJmENP+0rxJwcgmoijeUhoZ68DfC7hpKOwr+HBk1kYupJ/75gCkkkjLUnfhCxeFT1wQL2KZreLC
fOoiZpeiQfxFReVJZHVktO3npHpWnHXr4ZTSP/gpTHMZ1FVOY2FmWzDliY0piCpLtlItu808xInb
s+ehRhoxU17awtPQi8Mj050838aZdFbjGR4K1Inp6sitCJ1g0NEwwraGeTWeSbXfLd6dTy24oYYo
0Gi5aryTJInQO6aBgASYExecrvBAHNxW8q1YLZsZSH8X85RhBtwAI/Ayfvly/G/OHeQmUMPfoz2Z
0v4TFHjzTBpspFys6C7CRF8oSswL2JZSv6WJr4idRhPOpJMvyJ8jVSH+13PxY6fTYIZToV7ItrdX
b/6jaPixusGLfyGYFGiHFWtwUQiYgXnWgTkPPnLQ97NoVuDX3/+QmUlbOk8hxnTBy7EDKpeWEnrO
1A3H79MHprngZ0LyuO/mjhcUXNjTYOwn+4dqnKDA8KNWs7ussOwAqr2BZAq1HBfsjf5tY4OY6r2j
M8RX/RV43xsNtFiJl26Q0fqQ+ai0BwsQp7drsbS14UPOelpW6sUxgf+2N0m33SyAxurhQfsSK1Nt
Qjncfrd6cPelQQI/L9fuQPOEDKY7vtjwBaHIv+hHemKQwAX034tsCIl6mP8lZVHbpUzgelC7HP26
umj04Cw2izWjmWoYi42ukWAcVCeP5wmqajrNmYYiCHx40zxFGq50849n6jNV5FYmZ4BT0VPz4Pto
WK5kDyOGuZMZcXPvI8oK3jxxwOeFZROQXVhSzN/fNrgmu3FvkJTV1iwd5NUwxE89MX2KUB8kInU/
nEg3dpeGLPpgD8pMBOkwQRJVcJ/p1maoYVN5tlRJRu2N8mGh+Fo514SYv+xkk/DtG0l3AULTpyLr
nyNABEy44gDcc4dz0Bg7L0xie6Rg1y/jXtjGLdlaQ0+Ph+pugccuvtfbuOjofFc+4CN93kJCWlBN
cAgrjS3bK2r+PNsInP/l8BIZo15VymG/csr5vkZU6Qss6e5wxOi3IBy5dbpK4EW0o5Nv5t8C1y9U
ZbFwb0GwlYdtGBG/pHvPcGOF2VvG+IeY1iDoLfmopx45uWSZNLcFBvc15VmiNMlfi3KQXz/Qib6b
P9keXpMo0gB1lcYzeRpbXVTJbMYlN0DzRuSRR2j5JqXr58m6O36qaLEnMzy/RuKabR5+scNW4yC1
xSLAFJnUmajYys+ddJ7GfgVRvL60agft5YOYw4f4zIOTSyopdVGXYi6VseKC0p+4FJ8tgfI8D8cs
tz+1NouyoVIdjk5xVhuwjs7YRAhnZ7vI2aHSiNxMFj5N4nTeEZpgNjTQgZw/D9lqX1rnfUkDl7hm
0odajQGm0VnNcduKdXbKUNpefN0dL0pYMRFfWxdHHQzsmM1OSmICLxpk9OxgNNfd2eXc29HUWPbe
TATQuz4alWaMl9JQXLrZd1eew2u7stCS+vzIxe6duqLkfp5V6pu5vmjILGujlOcAgt/AFI8nQJ29
NUMg3oGwUqwG5Wl558UG498nQqgxe4pi8nJ0NHfMDLoIF7c5QrdS6VMyMTzrpy+OhQZe4UzObrT+
QX47TAUiQxUmxPoWS4Iga+kTpS9/K5/stzMmT55adaDP5pWtaHXTUu+wzYCW7j7wuoLCfDSy7S0O
I7F4nOVwtDvGsOdDJ3GjgsjJMj/HuRigbb75BhzYQ1CKLIPDdch0kKaHR51nYvkQzJER7P2AEu3l
/8b6csGC7UjEY2wUw5DM5I6qFTPOxsEGnOFrT1e56HD38+cvreFMQ/9Zr1HCXq/PpXqnQT/fcf5I
BF0SbELBOykIv46v4k3786Q1sKerZuRdnrs2zSilzKP/vSxmDXRA65FQawhDOijyjTbSRTFeOc72
7pDfs6xHQKpJMKaWgr0jsL4oDR4gvwOIvMPmbl3p5coUv9Q56xss7yqfK7jnGIvP5azL4VhJFhhr
KXE9P28rR3Tyym2Cayp9TP3KJImJtj94RmPvkcmSWWC/ZP3495BGmxo3TUM6KCXYFnusleVLEFu5
5FKNUNdV8KMDynKN9VER4bAlIB848vs2iXZPXQiMvYDASC8/we4mkFkbRMe+tKhfxLeY4nxWcPBL
VB6Y4wiNRmd1dZendpVJ8GoFylbZDRVPAdAzFcUNJ6tQu767WsNu9+gO9O97s6bC48BbZKMVKQUv
7Ar6P5weLWY5u/RCnPZNl4fTvLvqlgqMLB/TIe7E6r+ha+ibGKWQgTGRdhAElPc5/UB5AbBUaYwX
UP3xaee5zSq/lRQkXiv/JEPopwK+X6BZ2TeDpnYBKkshi6UtfxVKhFBPNB7Eu7IqgKnwTuOqq38C
/t/FcM+cd83tAaFAPHOazMNPMYLXnvDj07hqGNbtogd5otlyYvJlq5RdAL0Qdt8qOL9Qyh7NVKDq
xxZIDIHGCUsh1bAPY6qjHKn+YeB1HXByEym+962FLtUWS6RKy0F2RKzjLZXEOTjkV0feZdrAekyL
L5WrJJULSPByFJQg+sMqHHKxr4lqVm0/bPSWgqgMwkn2OcbPco5IEFQ0FPOHX+AZ6fjjgRoOAUFu
ZK1QAAFSGwrmAWw1cpDm7WNzvxCxhk9dedV06qi7Zt4GPuc+BPhSutRtET0F8Z2MBp50pqG8+NAU
yIRT42Ny5L18jCR/RJq9xj1H9G3TeLpfFF2EekaAI3nC9YwqrXxwhFglaI9ZxJ1va+BQx02gsllg
WU3zdeSutj9vUUzRRek4cmqTZqE4/IYTJ3NGTvGYklW8O0GGl+kC5wQxcdMP1WAwdAv77WTz8hLc
ywubNQtkE8qcZsNHplelZOdS8Wlg6JPaqgYoxenzTLFGMOi3VFeB7H/IxACQ5VKRVvGz5vs7Fq2F
YmXw5BF50hLiFpBQQMAM/t4x2JW8FIKgYIRcTDfOsjiel+hdCpmpBsNezdJZ6Sk1sqp9EYh74R5O
iGiq+RT86puvBAqnkrGJhOQj+FBVmISds6cbjGkuM12Grjxsebe9/OZsKrThRuQW6YKFHqgM9tTd
vEeG23RI5PE2a1NNyFdaKMxZv8SFwNflX9uMvjTkk8yZqcoEnik8iWbBGwKLuE81ZU18sJ5VX9Gt
eodO8JMiKIgPGcfE2bT+GH25m4W11rH053d0Vum+lqNktAG3TOpBNYT7ZaxrblfX0u+u32c1gMnu
ABmaNmpv+ncSw37XZ+bTTrbMZN/wvM2W2ps3XhS9aYNGkn4eOWRY4LwWnFlyxAvhMLfgHcVtJqCl
aQKvkbC5LXTuHewkZ7pC8f0V3ltSUan4kALA3IiZ/LE1QGxU7g3rTgku73QhXooJHkjNUIyARQbC
JX+MR4deH85rOxTE4f/iu8weNLFNYpsY1sSKMyHXuOcjDT7+Hcb6fCd8PcT4yee8cYhw1ZHRHZUf
wVtcdlMpHTy8vGQV4YMniluEzPEKiCZ78GYB1nSPrES1R/Gyv50B5onEJnQyPRcwvvECk3yaxyBz
J3HjpbICQo51gDcbzorRuftkbxQcnT49mlUQKtMlkupD5yG5uYLYk4gwymihbDx/H8+zkQcAYcBe
jB+Zgna/I4rrg7RNqnh1VQDCL8EJvH8s89fHnX+d4BHSPR3U/USe9+aOZuDEAZHx+ng0/dlslxbN
Y95EBLkA4jLG0kVJ0OeGB7GPqCKMN2vEC9zDS7HDtVAt1+B5AzmPRH7hJIO/dDhi8KU00JWAfXIY
H9ahUW9bssJdoigZdrGJQzVSxzsinO1GR5WbqraYMN6jGHRFE2THPLJIyWwVoEYXuALARrGvJsOD
laUSo4IkSh1PifQAoAdK0vWCpExwFxOsBpevvOuMlbYPefKe4gyaTkk84StspxWrEJpQOpNmAOJ0
BN0DZYvNPd5gV6S1AzmC1azoctqIKWtgqBCTMMcgPXOFc3VWbYnriDiGj9VOOuQPK6RJeioUEfWV
IfIrfFPDYTUGm7AUTXpeIaMaGel6C45rFj6uFBxBXJP53SPjv6VomGHncs/1WrVncRXWoV3f2rH8
t0TDDAGDWBT6dnc8o/S+kvfnCSyMl4QpY1RaKrOs9P/Kib0hD5H43XP60xATdd/8wf0okFCEpErt
cuX+N6JVmm2Wjbqks6CdFSwkM+Fa7/T5KwOn9vBqOoOr+VDPj/s1BTx/xKcPc8UzDOhagGgEc9eQ
h2X1kPTVBIdrQ9UTa3v2QZ6wttW0m3K4ddjVeknlFVCbQjRO6OF6TcjxPDABq/tOZ/lMhtVLJAR8
4aRA559dkJTF1Vjl+gwJRPLyBsL5Ib8Iw/zlP179499HPu7u/EqyfzA441tAy9gTYXYs2rWesBO9
kY+K8qin590mKJkaVZJwHPkpM1mQ981mYkiKt2RsS5NElqf2zB7AFov4JpUAcSV0h0xd9MfyDCzU
J37xNh/N1w+3yON/CJu0rYfVH4EkKbiuFC2GgP3kQWmdJeXlVelaIlifkydr/dF7u5n8GPudyg8i
3SK3oR5dLL0qqHE8hIpQA2g+tLNOEtzuYhDH3ir4yaplOjuM+f3IIQt89iqK7KqWAM9xOMdlp4C4
naSPzs0LbclXwy0WQoMwOeiGt28+6t1wugRZk0d+Yc5rgiGlko9j9i17oW2w6RmM/qQClf/0U454
Q2iqxnwe/QtzqkSSEakQYzVDC8xDFnjv9rx7gVc++3752OLQ58NOoUS3LhYBNnZfr+tf0NER42kZ
hhOMIoV4KsTvPggTagP9pPEmHA6wqWgd5P4YPj6XLNdmQtFokSqpVd1XNAI9yf1dPVM4U8kmccur
7U+GsO1EdyiHfizaS3zz4Fysof/LLSS33nQhLNhgk13ciNdB7H3ySSMnd5xub7bvddVO87L5sS4U
gHLF9FyxqG48V99HzPnmy5ldygn/9XwsAPTzKrtx5Fik7cOPsmnTi47FzYiT+NuZ7smbkD1LXaYe
ALqrCNMG7UaVmi9x0X28dqLoIr5pOXecfY82TYuxC9Qx4jXykfnsUMb4WjNM1Gbsj1fs5eOuard9
zfDZEWb7zEwez+y8vl6kZ66kLTCEq1q/9IdbK+WsEh39bGaw/+KLoXoohftxVEBFUNeQMEW1oatO
AXK6BtcFtkdG2BHoANg685OGNt4E8andWkrWET94jrqryzHT70596rYDoEG1vKaFqKwp6uhFo3Vw
L3WRmtnHOQU0xYmm04DyYIsntTJeG+Z5N2kCJfkNXDsCR5w1NHNy1pN0Cy7pUjrOnpobZnvnk3tN
D1DvvYaYRvTTC7bYIblBDc+Qnmn0nSXJjoBSMrsAYd3ZkeEc+ozLebU6IvVPHNEn89+eBpFGOHy3
dCwJ7YNiF9+1yw79vAWJQ/Hmv6FYuiSKQeD5fN+79iQZhVf4uuBSN8CA+byfk0pMzsX0LtsPL7wv
L6CA+0KgI+YtBHJx5JxkL4MIOgjBDyPiVc7vKHqfBEKPccXgkBKStvzod/BiZPa362o4pvOXIUbS
II6mJyWooBA+4LdMNjzbi4ZGI+T2SoQYgG/lMVgntVgav8Si6XF14HzFrsGvx2QUExqL8mqS8kaC
UwYOYhWeqzdzxQhpsrlgtuGCFGQislvpbhOUijBDHfpC4HqiKWsLGlG5mUSQWPvGM4uFOpEtV1tU
LfcBuPsWvMk5ndFasVidRUZ2rIK+BD25qhOwR13z//50xJJ9Cu1+eAXSPixe+xk2RwPi6ETiGM8c
30ajY43JchIzxRgkV7hIPQr17kYV+Q8lnQf12A5m576xPVl0XhDwj/5vHQhWbxX7nklOXrR5BMF5
DKJvyMUDUwlymKJllAkK8rYVSN/xKDgZhCv6HBCCkl7pAG1wbsVFxlXix2heK5zfcZ67IbV59yul
bd3So96F6TwP6079xfMQxc5Ho26f8hMHT8c2Bm2j0lQTqrF9mcviMZlk5faYGP3NBuF/1nYZ4oef
g/XUutbnWy5KxBMjmeL07DBdrIe9iZKn9LyXVU5ojocDXZCS67086kqb0gX8LWcnElH399RLLHJD
k+nDVP5bS5lvu0hGSdx7S3JMM6Yjqhx1heim/v8hOfQ4Rya4SDJM59rzBy1eYdgxvMaU7/glzwUS
WKExMBXYYENnqZsaxLOoDNT1k0Fl50UQnaRR9JqMHIWw01CZIxY2oiBcHig3LfSq/Fkpxeh4MIww
mAxly4RXGar0wKEMrvIRK557fQuhcBQOTJDg0qTAPcRaqmUuouX9DBakSe6XxZ7ntr6WWAOb4BpK
7jE/HpxspuYii+MRXyEPWq3bwj4lDfCaKbcjMA9/b38BfGSP1+GEpwBEcyE2/r/Cc00BbbhZ8RJi
mlUhFanc0pPStYL/5m9yq2X1KyWqqHyQZWyESMAk/G5xUMQMElk7kZPgKQ0CBvs7Bq9zr2RSDvQb
HAPnoY4egpEUI0GrQwjY7jdFw9Iq8NvYgN06Vl82RZn3s1FUYe1Ndbxg7uycddRCUM/RMG8kjW7h
two3vbLuvKgD+6T2iUJbjsHjtuJV7k/qnj1k4JyV0gtdQ3mjZNAmVRlhvppmCLGP3VeJyonH5EDN
8bhVfEsJrcNDEWaWfYll4US9/jSwRtznXnHOttWoqjGju1vekCAyQoL1iNgi4Wqtvk3koi3v873r
yPRkqYZVcZQTr0R9ytvN5d6fktkHcLFoxj4tFLYl856OzAsbAhsWNLm+F2wKTXSwg0pYAZTFaOsJ
9MsGTdJbg95N7fkRQGmJfSrnQjykrb1B1ue7VYhUErqXJXADEyvmK13v+EQXvYHzF2nPWngi7Kl7
AZTIih2ec+a/09XnFmAYnIJ+YA9GgCa2eJtzqLpsi0HB1p6g7OZV2LDKvYXg4C10LI6Xnq/CgfKR
HtfMZ82c069eBCQddkEkwL9RFrfrCu5qvGwKRiE8xXW00gg5XuB1u+GogzzgN5N47jwqDZmQkAZH
lJ2G4LoyznS5WecRqUdAatPGYLtSq/luuGRw+HmUonle7syb+nfVUkh8xxYLT/KWqBzmE1NsqK7G
49A1gG2CO86EEeFAb6nogL2/BF5PHXw+uk4NAnCQK+1ks66JeNEs7bEavYYRKWFpQRFIrtcKULWU
A0s0MsmHDaeqzb4sAIUjfUIpIei7SwNjkrkWHfo4ttAQ//SU/hz2iYW08KysgyuFssDGmJGmOo0G
VEvOGXHYUuGgVhFyZadVCWL6XxRtHqmcP9Od/Z9CfmRWPPYRf3Ya/bpW+lnO/tKVr0XVv01DoGXg
lg4crlWGKNzWziU5Icts8kne6rCguyf0CcIWSk2urL2Zvv7Seoj2Ks2PJSN6771HvkXEi40OXtyl
nrPLFeAVFtf81gm677DDUs1KdJLyeAFBkycmEd67L/r5NCluJ9vmQRUbbpvDJWIdIk2VjHeHyAHI
Pe+LN5Il8tQtUmIoea91czr10zZRvOacZhhw1M1mWX9vdKjVI79scgvN+s6kYC1vIyt0Kgqo058p
ZC36qp9p+x2Vzfxi0qEddjp8bVhotDP3ctuJ8sHntp39I4CWsy+1mQXEBEYXo8Q+aZaCDlAl2E9Z
aTq7DPMV0hqHgjW6RYpwzFIn/Y4W1ZikzJjBpw+S5g/U8XFnfCkqBikz48Cr0IJOIfgenNKh8GDA
grVyu7u+OWaSJQkk+q8KLQ/3v1b+Y/+9CxFltfgP3DPC05KBj/Giyzdvm3f/Dw9gZkCz6n0p1NM8
BttT194+T/3zdcdrMs/vHS9qkQRxBgOKTFNXoKw87+gs7C73JedWeKFndUBUtYXS4tHcEiluToF3
qzOYyZC0kYYpGQxGN4jdYr9WNe0LE/DcQ7aaaDGp71njK1a3fp/ZnZTGSr2AOPXJFblgtnCYWgWj
vyQE2OTcIMlk10uXB32QC6kS5YP/kQWTf7IeY78PAg51P7/uMpebAzdQbiayuhZ6gc9elRhMSk+q
v6/2mVr//0JQ00IlnxHt8TOeTcyTYY0/7EgAQ71CxFVFBjrN1EvXBLchyFWNB8heNj6Y5YQz1nWH
xzmcE3VhASh7HqOIAOmSp7pEhcLdYKbgwrNVJTm4Lqk/juRU4fVOUN439dnT4iRRshMpWODIrtoF
dXEr4MiBlPEMHePADLOyaDhClOl1ZgOvlhv9V7E8ufQIbxwzZwn6tuUXiiVUDXAF/jVSYQ95dF5C
RQu0fgjE84bfX7ta6A6WaE2UDKEMZ6Sq7r8vLQZkKZ/mso4zfYhGsfq1oIusuQlGV5QVHJLmhTaD
qt98YYhbGXGECWS9320SKKK7x2B59QbCwi1e6xO2rg9smnT7A+GCAmac5kieaYELw2nXYB+30fau
dpCGQSJumK8CuKvHDd3lBIe95ExIJ+PtP6H2TTgv4oADpGbCrt+PMhLLMJUNbpYmG0W6dmRcyE8x
7ZxEcMuoP2olv4ckGuaUYCkDmcv8/00mGgaoPOJZb7br3EXFYMXbT4ak9rkJNV9bOd18VuEyvWgO
+c9CQPBCf7t5D8wpWq2abfK+w1T5/BoyQOcwWapUMPhynXhDpVm258+JJD3Hcs5ZVo4EzxLQru7H
VXYgdOsfGhEXxh7r2NlxWnDD4IX0KmxcOi1Dcfhr8Tq5DQFTt85KXGQQ/rI50zTnqV4/PfMayZ1h
t7kefmfTSoYqG1G0w5swQSVFKCVJ1U/QvTSX8olhgnq9G5Ua5BCzXmNJv0ukc0qE1zDEWe158TL+
cd1KdNUwWyVm3DuroLEZGtqyJXOIXvChZGxKSD7zmEDPEDfyRQo06jMbbIVjVu+cYF3C/0CiuINk
N88pKNilPBlMXFuVoB2B5CcSFPK8MrVypXGV2jY9JHSndcIISZm2AuKR0Y5RRLNhVC2U1AbBk86T
hCFPjaAGYBt+UvtptgStRbhD6or0DHkoGx3CQwvGNlUwmyenPMKoxTjDT8wvUxiEFRRjph/hKOV9
P8c/Lg8ZJtu2SJE9/5UTjvuoHFCBkuRvs09H5l5X2qDk9gomn3ByWTEYLgkkabc59CeIQXmQ4psS
6yDD+4nAp+tAu0TEm0euzqLJdroD50LaqqytLVeizVNzPJFMtEd7+kwddKUZpfEctLGSSpWa5wvl
gGgwbjM3yLU2op+noF/Lc/QCNRLzp0bBZgjI0TkfQ5YVjZN+L0ReAEh6jojLaMLo3IXtxsVHZo2M
xcTSkxyDFpY63EF84Wm/jhyTbBtxs2McLex7QeUNd9Pbmay63ZnZjP9FLyA6Vf7bw0q470hatIFn
4FpTuCVFfmAEWhEpdHtvMXUryKQRVvEVe/q/0TBSN2HSMXZ86j9SU/quzUpW4qjNopcKQxOEn1u4
oUpE1gyb/zdS9F0sRkXz7ai7lNBFBrQCCo53Y4NcXuvRNrD0+lTBvVvyDcYmP22oZFnFdIARf9or
2U2MOjJglCrj1h1BGBnHcMpgqMgAP3garUSf5q2uOTqVJT2gSS14MbZvMS4B/ALaWYhIglc5JpjI
fHibzUI76j2SjQTvqGfAzd5SSSV9G3V3Pg226ycrGkfydKaGio1NyTAulufAiehxHlyNcPl88WJx
SWoqKiHCqA3fU+zx4Y56XPPISfhQvrfp9r0rBQepgl2WXUJ3Nf3N3lF6WHBMQY8YQewHWASZeJY3
XEfCwsTzPdFCYvYwIu1kXukxyRvzNMzIigyiAPguS1JPJC+ZBloFZ4woyy3JoicLLjM6YYwrhzBq
GDaJ9f1wUg8wjURdqN2xOD+QaP+PxzHuaVyP37id0xmb05XKEx/FedXdOPc2BoUJsWnN8p2lHZKh
SnS7NFw5RJKXTJwCrwB0hUSioFUS9g6+FcrI/TZe++mtgfA1Icx07a6vXEcgcxzyx+oaN19Sydyv
d9V8u5Fpc0nnMYOaKzp27zyNUdTc9CtUZfHfoJ91v2RrXTm3mdqJVguEKnmYR/q6Po/C5hHjIFET
Wxb7KLvZfqO0K9nQnr+JcWyem/IcBvFODTnB2UEcn+ljmDcdrjkwxJ9Wb8yfIX9vTA5B4x8iQGJn
S3Ohs8txMvHn+kzLpnnJCUP6kX2fLdDovmMF+WahV+NjeLbgGA1d2GMxM+S7BkpJKaTMFu2Xbwz6
qkZd6EAUtu5v9KMblKkT28WWO478pgIhEX4a5fKL+BTLgZ+KWdr+0dlW763e+xUsKpW2yg2FiCqi
3eC6AOBkoV4x0Sp4D8p6/TkfmZ2C/7KqT+9T2Z+EY4jZPV3J+pqmWkskHc5KF/jN2KjBf9kpYqoZ
qM2Twz8yidgzzJrNOe6kb73dVmfqGgyvfKtRVoO5vLKqT5vp74gzSkVCGaNBCzUzU1VSw+cYOGxQ
rQ0A+HiL0PHCJEEA+6j2mRE2NKwzmHodP4l3BGllHnSQTqbcIkONSo3bTIgBbEFJWk9wBwZL5enO
+C8R4C8ldCqZeUHoMu4ahVUIgIR2zf+H4h+hHRovqPQ84CEA8q2DKVX+Mxt4TBikZf1LUCf/Cu+8
oHP93vIuND2ZMZF07Lbxp0qsGZ/+ga+x18xRXAMUZF3ys92iDqK2NvoT9237NT/GcUksgOBI3j+0
QAgAktqi/3coLKa14XFs247Y0z0yAFeUUOpozxdDVSxo+EnAzTrucWcEL/n3xBLM9T+qBrdbVcBp
koTGDEBghWHqAriLjRL1C78BcPiQL2zVP6YJRZ8/Q5MWpe+4DCNJAmZ0gGcDcqbBojbDSarLf7lr
xHJJMeVlACoz6qgPhYUr87nGK8PTB8eZQC0P5Ta6FQzPRB1s3UR2vBfZl3yS7RN+Nhc6dTCR/2pv
diXaIFT/iK53agQW4IeZmENvKi97bH0UfZM1TsA+K5APWk8XuGz0ce6TekKjYEoiBNBJkhsa8yrh
SAdSZ0LD0ppD4PeeYclDnd4Tz3c5aqE/Xah/c0eKhQLVJWj5Q6DUqR5qB4l8QlJXRo405kvVWZld
PiVKABC0syotL7WiswPoRHyHDM94vF3CqJ4jPILb+0wNv83cJefRRGEnbBE+WmH2AkhixP6ln62l
DDHm4ssG0YmcqbGq9EiQUebnUv5LqZdjKCNM4jjPRb7g8GzMvsAdDYOJNTqueWylV7eDfF8MSpIi
7O5AkOiKuhUxPdsJBS9iErnS5WPH4GHXt/PCNXnAQMzkSX0DO9heWdonU/svNAAPZ6gJanBqmE2R
opt3mZWbKxRkBRlkOFVkxSfDOzddwWBGEYxyIoU7mZSv0sEywrl/+z6gwYhl+cfHhFs2J4NRMrTm
GOroqc2elAzk/dxmt3HMru9ynx1tjQhe68KMln5mdnJUhVlQdqY6jotlPEQ7i46wusYKgd9wfP4c
rgI63CT6Y+FD5u8jzRqkZBBoJfO3VV+auCt+uDC9LbUfyUhO6mJC25be8Ke1KSd+0sHVxe1vXA89
xjZ0fDho3Xcfd04gjqrlLAhcev7R6UDQ1WpQXNNe20+aAwRdB8H1UuDuKc4p5Y5Wq5Ts+RLUd980
+pfSn95RTPmdxnQo5mCKoGlm76Pk9+QjkNcU/X5fSuYl8j+6/OyUdtj6H3WUyFUcecvyRMw75Ju+
V8F5/0gFg+Pg79HIIQJ0ixepEWkDu9yNeazBtcvDjqsGEjqmLJE4f/7DUSdwms1/UPJ4N6ZTp6JU
GIkXMlRvUeJyMia+2VHTF7VHZuq6PnlCo0VTiNKfgoaUOMg/vj3yoZ18F0rCochJVuqKoLqj0Sej
8jkoGD/GFWsKH/w1lEZdNa4HjIYCQItXHGN1YL805GThHois3eJgRemFk+RIMcCgvw1RDuNbBa46
NWEA4GPlIF3RijFQB5tVlAetdaAN4LmDGGNiWq8ynZLFHfqnnTnYRTyq2Az97K5fpFSC6qKtcHhp
hiyZpCo21LaIDGlvH9szBxeQeWM1XbctHrJjy3CDrGUVOYAZECsnJ+/wfo7AY2uAGz9zdOfbaIuQ
LdyWFtC6bxMQAqBI71yqyoXZHbm2ZARB6dCbKmu6JWb7gTCsp5KOdiW2AEJzyUB6Li7zNw8gx0s2
BzQHbscp0jwqjo+6TEVPf5y8kx2DIctHRl2/mDMm+AGJEyjjLW5ua315/HcZLLJOWOtrqwybTFbb
t1/XGuxXCcZjhCjQBUMzXPoHqo6EkZ0pJHi9KOu7yDbwT9SxKGGuNekAHu2wkVoHbHTIf6O3tFgE
mPxmWqtszc8WbYL52PgFQR7NGNBSHdaB6jOD5YQ/9s6VpmmYuuUY73nnRXWsA965gmS7ot4j5lxy
clA7mfRNGCk5a9mT6vS0tdWTcdavW5H7Ex6DWdx/KtNHsV5GQwGXOVm9oYXr39q109wBDm4B9UiK
7RHmwRQG3YyDVN1OwqLSZjwSSwMpibs9W6KX1W03Uf7WxsCtWmSmTh/00sq998Ee0R88I2t+xtRR
RkS//iG/10l2BtIxKmyy2G1obvNKx6nlezM3aMNndlDZzkCa/TJinkWEOQ6jTpXR7IN+Ssg0LC6X
vPSSopza/WCBQcKix0eIcmiPm+NRPaZ/AqL/k+FO/9gb2UwONqk962LBgN1ahA/Ie3pRK1oL2JII
nkJIfCy6Pfgndvff7ByvpFArVeAMs2bs2XHjWppPWk0C4eBLiE5bnbR1/Eiki2R2tA0ljm19Daag
xAYH3gH54ES1hVAVI2PPD3zbhjExQmpRvPCxC0ncmCKdFHUvgScR/4ijsloPWlsn3Bl7mLsJ14zd
hbBQHB5DtHOokC4McyK680ErfYoqm5q1hHaikNMWoY5XRM0pogFCu/59A8cyw1wwEWXBpE5yFQFq
gtmCavwEHrbQjFpgW4DsCfpDBEXlgaq7CBJLUoPKZCu0bYG9pzF+Fk+oarK3IAI1vQz0s6mYimIT
e0hxmkFpfcjaAAjJdAUYkqCR/+6KRrx85hbSL5vw96tRORtKZUdZ4tbG7XSlw92Lw1HG2EWWvSBs
cmyDVuUfP9UxUidMm2nblsup1uBjhavTaD4ct97+suzlRfJ/UQnizQQ0cTz0DxiQDrE9BVYUhtr/
3/kjSGS9pdl8gojxdBZaAKNiyAt3mzAxC6vYch19IHEpqKtMzvnc7VuGR8LxxwqHpopdgXtg8OAM
Q0NqpMhHj8iyVEJNyRHeK3l1NPILrQEzw3o6exp94GX+aZdutyYgO+3U5RHQgZYc86gYwPQa84gU
CKDQZJ+Hsh2IeqyR2L3Jyt7MOm2NmD7alnAaM7cXKyWxOuOUS5bc5hJrT5dgljHt21Pd64CBpjWQ
DOCJQ4yZ59UFQUw/INjRLztrPqCyVZfth4rHhuVUgKRwtuQooMQQZ1OOsTIJSVqOc21fTqbn4Myt
4zgEJB2sHEbuhYYeexrpoOTfzEH5HZHuTr8sn/gnFu7Uu5WlHdwCkycVaJBLaiWZSQ5uYhkc26kh
mXON9pyFO5DRIblvbUb8qEgcvYGlwCwyqwRemHs4pbePhBr4CoQtC2mZNC8VSK06Ju6zaq+Fbl8o
o2A+h+q87oQjEKU18DzjeVjgO899BR83WCYVKwe81dZVNq/KXxDYFQIQjJ1YnP4vAa4oInwMUeFd
yTTpxYnnUHqXUiAaicRDORGfUzkukZwHMf+sDmsLIsaH/SLxe9U3EC0EL1S4BcD2C7Sptd1IcYCw
0bTd5rMJUu9MxwW1VRa2jD6lnGHeaBbOdrFdh9cQxTV+QI+6DuQUzeVCYaZXIA9hTCAMgZXBx6Hh
CkkcgQ+araYqYg5ZAP+QPawC+unWpel8GF5mvv1hGUzjPM+knsLfzOPTqP4Mg9nJJJNjME8XQA/o
WKW4GNebX4AntbzKZzu3ACR40N6EMxADLuj4XPxeMMh8CSysG4zwLanSpFqiKzjw1YW1Y+GnRdWp
c1fxPa8+aBs7V598tzVQ9pjBWGrmMSYWZwBPINouPc3yuReFERCHCnmjuP+TV5xQisx8NQneYota
a511Q+h0F+HNAytAGkPJukKIhlKrVat7VPJVAiPaKTAVwwVqKdua7osLZArhuGDSW96+Ivd+/M3c
DkONsohLht1YxouLQwTlqLAbmGhhm7fAF71U0NBoqlYLPb82dNuQPqaFFdTC3CNEhUxokr59afhn
wti0CydnOoVvWeIYtTScF6RTO6Qx4cwD5ZeTnVEh+ZO3dWx+vaF61aCWOeXz7zdm+4yVVgkLu5Cu
KfPWODxE7yIRXLi4LqTLCQ6XawkLT6NBPzv91K8NVN/sZgTazgiCZYcuVenyckuLJSXwIfDe3c8W
n4z+Dr91AlH9qW7O7iR9Q2IiexpQwHnKR1GkTv598yMOPs1GuGZ+l2AwHWwU90lWC1z7M03GOyJ3
JvXRA8+lJ4aMNJtWIZ9ao3yXSF8SOkD0hHmYu2e+GLDnrbyQdjML2IQSCSKVftW0u0lram4660nA
G8yznFcKOwBQEj9lCzFr+thZWXI5Z6GWLW4SvTeyv3rqboRFfmxqfB4RwmEzIPTh3mJAqFQeGrCR
SHfRJqhRXOdQp5gbntDBNirh9iZI0/M8Aun8zNzbzFy+VovYnfTtoCtlXuTXFdfNDj6RDvWHzdLf
bZ76btdjHiCCWkZuIN8qjachc2wYl3H7aGe0I6rM3Xeyd7aot+iAL5qL4ud9f0Wusk1J6LMW8xE4
ProXB3CJoYWkcED4qmDeQ8UrYslw6UGS7NlU3svvnyP9OlPwIdMP1A5O+2gm1rZ4zly4wgH9vXyl
X9fVt8JptKrL8kf3iPD5rbfja4g1tJPm1Dt+zZ1jxdFfP1k/Ot12r0UGiUutq9kkxN+hVQiPYRjm
nloQnrOdgQxBy4vY578j8/YHM5ttDdreSWvXzbu/rsFOiVQsSGdkG+RXRfNW+oYBa4An9JGPxTrX
Q7xCs2ISGuAI1BGqDTjsoxUOINUm9+MDHk6ajUgSVtj/kUeGU0uGH9r81doZGanbwFQONBNHWj0Y
l+ZZIc32anJWVZadrGRqZF4vjYB665tFlROmho896x8LcmmKOiGrvdSpx48R3WNiCg1jI3o9XQKt
6LfzYVJKK+Ig/CjmSrNA0OLfDPko/4ZplCWQTlHzcdGBIkNPJUJFv4K+97hNFYlPsporGaUcyHi5
WJgmg5Q2GvFsXlvBDEi9D9FL7U0KwxyOUXiEWHWUvF2ga4y/c/k/NK/BKkFu+Yy7r1eZRVGekEqi
N3ECZu2FDJcqneA9l6nqETCu3YZcbaTD3DNwNPtp/OFhYOKD0Ftq1pMDFOfXMYX73bO+wd+16Gu7
ySBOr2WEFxD58UaJbi1D7coKAKfeU4i0iexV7Tk6xndipUpDzOxRT8KDVTuE9VaGtTjnbnjqyshH
S+HZUvbSWCS2cBrTZFvAqCE8nUbXH1mVelqoXYdeGhYY/EPvHy8pKJ+Ln9wgGL+PAmkQ2rdsvV5k
86ekO6VHZqV/Pzs/kesibo9VVhGsvZx550jhjgfitlyuRXSCYa44jAYj+xBmB0jLEjL8ZOv9vMvo
e9/7P6LHnDWBfhekwUVdbQ8Mtk5yvZ6bER58wFBv1YnWJWip7U26fZZMJ723ODVme0TkhN/Xkd3a
Bt9x/Gu0tpTZ9VENVbJFY74aXncErjqMlCnz2w70LLRI2g9xbhSOJsOaW6cHPuRhZXrwOS7zqrNM
wh4XvJUwZLHyFFEL2e7mQ2EkERVbMVCJhDJHaXesdzwHQE9U/Y14FNR2u6nF4O54QL36llqRRR9N
JbTG8SE1+ygKa2KAHqZZcTbmP2n0+IeMmCt2zor+tqAH0ocpsyapybRWrcrn14pK71YieK4sooji
jRhm+6HcD+G8YxcviTvgdlZdMK3N3GkP/CKxQ/5HeyR245pPnB1CTznxIclyZvjx2l/rEkZDKHwx
t4eawSnpARf6mFIT41cQqv1taXFNz8PKX4YBEFB0IGowZPBNeXt+fnKcUk3xQutL8uaGc4T2F3lu
+rlFW6krZduOSkskFVEecn2LHbJjR1aBpS2oZzLbXIVx5q6R8gPcQV9kltxtwP1m/6vclYkw4Pfw
SX/E5S2XWkZIKG+hI4w3zf80oSrAvQGjtTgzg3gFgZGUB42KCZUtV31uQmRJFcWIimNwz7nQ66v8
gYhvQHJjIkPTKsKvmKxEGL0Zy0uizmkZZR1mNh7ooLC4jA+P23DexXeFFGWqCmHm/t7qg0R5iU0L
dUsR/RTD1u04Gc6t3WJN2rpjURYiz/36c950ysJcpjjEffshsA4mqQWjOXA8Yczh+PigcHsLWtvL
kpv2SC6GwQzzpANDe13igO7y3X/UqFujru2FCXYqo8U3TZ9orT7zhpD9qE7QnCxj5X95gUwZZBAV
xHVbPKh/N2hLuAJj/iriwGhSeJtMykiTr9DHek83Iwh91DBQWwpbWVJYEIKUkk4WbDvhRMLDD/p7
UngvVga7pueyqyl04JuyCY2JMjkoJlwt+oRozwp1OqRxe7U5KzCElXQU8MdQSGNNEqu0BUsVzBq0
IyjxKqrGDVzjvgX1/0vpbm6Z1z78AK6Mx7J927OyhjHcen7AXQxI1xvmGsFTDrSxNfamPJtQe6++
3O2jCCKavGQSUSpXsnPEt3Ld6iqoVXN5TedGOfV2Aqfu+wWRJAXrBFl7Bp9cvfmhCyDZZdgaJhLe
p4de6/iC8uTUIROMzEHE/jr8riLc7cBmvkbV3qVGj7TqcTaVgS1Md954j+mBMrQhv36jo28MOTiL
TFkIGYVlRV6Bui0P4b8rBm9nx2sKB8K9t1/8MaxEi/xqdtthABwvxC6CrznXLp3EBr3bIQrNyVqI
jlRLobDY8O1zsqxRYzi5fS65DT8MVicb2pyapnxTx5Yopp9j34iLnDLt0zQl25AKD/WCwMGFSNDh
LD2JrPgUDPxkNg8qMUQE92Bp43kSTefe0GWaXadV9iJ0XrC3ZEmT9fS+ot9zGG+KDD3l+cUVrJaT
bYgZ4oEJ3XQa/v6OrYj6r4IbB3MBN4MW1Sk1qwvuPOCq6QZZACpekcc05n/Z2Sw7ZgAMW4gKyR20
4GTU4i9Bn53c+afmH49TH+fnefOCqFi99U5LHzcdNeKOMjnp3F37T7A5E1C1sJ2ypWIgW7V4+SoI
gN0h0Ct/lsjh0nZhpH6iSqXO/VG9liV9QoHAPVfLL15mllFjCU6MoiTP6XyDUmDpJS62trG1hFtt
U1jWcsVmp3zAKun1ppCj+ANjoNTb2VMHafKlr4v9twU0InzvWOYxw/Sq+o9O+exZu0fBqp7gNZoR
HsDEEUptON09nD4VxRR9e3lihj9pnMyEEhA6IEiGZBF2fhHNxU5a1vCVwEDH53hclNSdhFe+fgSI
dy50yVVhvJflIT13DiUheonaK7K+DQmGt77Cwm17srHkVot/WtkEG3KjOVHBlropeUDMx9AFLtxG
1JzXv+zAh22mYmvBw5jgVm2UdQLqeHSPAlUK5lnDi9HHS8E3qhmGTHeO6rD5qF3I6hILDWySthlK
p0iU2K5OudLUvhF4Mtc60uWZ1YPONBUO6WAhPg2p8QI7yjaI0qDOx2F/w8iLvCx822Y4aKr4QiyU
cWAjua+N8Mjr+y322OOd5cGDkQKZ+r1vRpIqjC+dcBSiQYshWJjProApkqwDpt0K0X7tK+pz5TMh
uQaK3Z/5oBUAIP6vnetw5Lku5iUulpS0i6EBYpjcOq0MTwSCml6jm3fa2Dok+Fxdwo5Kkq6phuS3
G24k3/IHrEFlXb7idfJOi1Utzm3mvKtVxJcv+uk5kOkEgI9B8EkIDruYgyPd0xbqGKIBgVLZs1F9
UGs8Xznfy9pp1fVTZDJC+pjxaBNIgPSMq3/xox8fH9t9Zmtt6Ptj1yNokhLUQILqS8RSNSLb16pb
ZPy+omgGE2V25epC6qrrsX8bKu5xxFeazWohOWMelNZXpOUa3pa30wg8Ykg9Fp88UE+trBVT0hir
74MVGa8ip2lqIMPyZVbiGrWcu5TyK1893AeqHixaBA9+XsRYnakpqyfWAio6j7t9CwyZcU/CBky/
oYa74MlLLq7o3/qMRQT0+kWkwZBfS5wCCJMtNmjp/DMkJWEI96V+veXyMkjvEgQXelTO5a2Focic
xmkUg2o3RBh7zIcAhQXjdsetY5TBAY+9K763krLGU3uxo4bpusrlccmNyO0nRx87NdUYGse2qsnL
Pi/sgPXeTLeQFdyt1331Kvjq4BozEVVEDQsC/MLddXDgTbDSSduEt+pBFajUWnpXN0OAtdEILWT7
ys3UTvHNcyMrZQ+2cwWvOw2s/xxx3C/K+iWgHHpdiYGUxBNgbGtAJug+IwGhv7OkdvoPt//XueiC
/Ed+LXKOWqtkOvW9pHzd4XZXprgmc1oo+908Pd77Q2Q0ou4FwK5jCIOkVqCXuIXedXAnW2SABUqX
AgkEw0W0SM9Rn5xaCQmM2Uh8JVLDBIFkHcaEKdHYOY207FRknwZcY1tLLTBmLTVJWNsHCRnLSlPJ
4XfD8PiYdIRXOjzTmERyqNeAXkGMTbS+/pmsup8BXMoXyiLSmTINrHlDxZM41MfVZcpIU4wMmZ3w
urhbiVa3r5w6zi5gCecwWpS+Q+OCmxjO4+8dqQNu16GeOQf7d3eViN4/PUFYNDqY5pzfT9WnVdCB
+0jV27pOuY+FGtgCHfdfoK+/8mLmB2T5UqYR72lBWmc8iUsje74TXT27jm0GRV0VDw4DHMA+8IWW
CC4wBgeYNmw5Uql8WV0NL1h2za9OHgnPrMASqq6B4Oe9MP5T8hbh4PnMMekxJCcFuLW1e3N052ZC
9Q7zkxgqdbb0sA5yNWXEprJ89kGYD4HY+U1pJPUx8gZVVMic23yelZeblqtvT5XxEvgp/F2WrZ6g
rFW+DYsm37sW5Yt0A321DZQ85Ifjg9pFFRNfXy4CRPUw2qdSgRicz7eN7t4H3frCe5GSbPHJvCdA
uqMS710Xa1iUM71XblfIKbvCSl7h7DGr2mD2AF6g2lqFnc2X/g0ELf2oDUypB5Yt3PTbsvp81E+G
0JNayzc2p8bPSJziu9udB9FEf/E1gF2jKpmFmJ2LM9EIVbxCna9YrMv1kwkAHtgKxDhEkwOGHt4R
gjKMeK2ACEgCR2DuT8Xrmitl30KIR+J+hsjCPCFgjH0xRdIxdARTa3gZ29shMK9IlAfh710ux658
ZzB9NngUl3r/EDD8mL9eobIVyu0/x5zpucuiCz49Y35s7uQZPTOnIPyaIJpyggAUlcXAus5ZWPQ3
kgrOViY9VFBTUiPB2+anPREJ13/PKcPlNGkAI67/YCB5L8JeJocxlQg5merNnud6ucJsRqMocKAa
Bzpg9yZ+yHN9hiTQs7jHvzozzYchBJ5lAYAcF+poCFxmJOUbdg9MUxBiM6SOs9OOzsnmkl/cKMPQ
QczojGgwQUjPdTpVUs0m+ftOXNZvCT172Hm1YvuCfnmfBYoj+4Godb/hlFFJxN0HrCNERnzXAoGV
wLuS5qs5A2MyjHU8NqtG8ltTqBN3fCo/FaPqlaVbTxu46Z3uqYCMiwxF0HEwqSBccvSiLa8317Ef
59/n42Ld5iJFvutcCEm/f1jh+Fh+LFZuEEnBaLEbjpN4JRKs6rzxcXTKmW4sFbin+KDzFl7KWWBy
T5uvl4nKlmVQQn64YeeZOwdsOkvy+Yf1qydqvN5IiEooYxPZO3RIw+Upy++bRg1ZzJSEnQqowYpf
6E50v+88llfX85HJsFEczt0P68Xchk3Z4XbYF6s5xjgrdSV0j8y32cKn+iNsdnPz85eyXC+Myc6p
QdKHMJusvFnfqtAHnaiwQ/XQvgVRQ3C12SiwwgKRhLfBInV6K62k2897HpPLMLHmv0Brje1XeIKe
s4gk/kvKuDRcTi49nj0jJRekhp4kJaND/nviFJk2y2sdSsolY0tPEnUmCb/mEVD8B9PcEWj9udV3
anNClxP7k3YBOim0CkzewcRU+Ctr5d0L1kx97Eyzs4FUxFlLAIXRTDqFcIKl9TWzxcMxCbjaOomK
fE3F8iEEPl4aOVIn8cAu63QOewy//Vu4vSsTd7cOV11ygn+6BTfEATgS3iSYVmifdMFdxG4M/mvo
4sDSl3OZmDscMzLJ3mKKsSuVoHsP0wThfFodnl4QZBwzZSdIUxyCYg/qQn8hcGwV6iK2CT9/vgC+
27MwLhCRyMRaxeHUwTvKfyGW/h4lQPHCjKCishd6D25R/1+ZKfSElf0oQikGsQmJXvw4SGBG6ORV
kD0X78WdjjwUL7YcN84wv3nnq1ADkPn2ZBwmxq8VC3pIXAcY5yIavjK1UjXjOlMMzokzhYw/c51P
cw9lhqS2S1i5PGGi1kJslWOBAQkakTSFEunSS0iEq6cv6VJp/nnLM0i/VBAoXIcEYAu6V+Ww4iST
zeANQfpZkaiV6d8D/Wh64bjcwrD4i4mCCdOwfWEr3AhlJvY7MIKFgC3ZZQIJ+dIzbm0g+DRlo2lv
QcpTP7fl++0OLxFTjiSNTr8ib7ScP/VG3BpPs5RZqdtR1Vd0Mcbg+CUtNSJHG0Ea3aQVpOSMA6vl
DOrK7F/y0BepPT+AZiQxgpdY1goe1PJKUFqQK+N+NWJ/s/tdMOm9Ja4RxBYgbfS+YbAJEOCHFY2p
4e9+HQ07y/4h3OxGhskECHf5Lp77CvcDQG6bEq5Dz3BTQU7lkmMh8EJsEg9UxDrMYVz+AaqunEEJ
oOczprcAFvCE4ZHveDgfz5zVWMWquKu3cnnUPrc3bRdQVj1T6UV8ZinzjsL5qjzwancWFpEzEfoi
DQI8fjwWd72R9ujtNmD6laOjrHLKK09H1r4GREknmgrkVMRymufr0Au4as9OdZ1N96ShCIOyWOrO
U5q9W10v5NpWZz4rqdK0LHqZNbeddriajacr0jzHQJ2INCQnqOjEudaROaANd4z2daouoONE4niV
oEnfRJaT7YRnaOLw5fGIUudqFfYj/uN+1Ep/KuGXgL3TtTqU0jgZjgf9wu7JI+G55N+oUgyoP4tf
BRwB3R/eGuJvtY3MtDOjcYYxacJ77nK/i+W0LJYjwPR/fRPsqix1N0X7og/biYIbDTOQE/LbIkSk
mD5eB96Y+a0O/NoyRa5j1pZf20NNTjh6FMpcbxBXJq6W6aXt3Op6RP46P3n6CJxI5clS5a7M4KYf
RkaFjWp56wLE4meYj6zi0jadoLAvQPrNH7V0SMz33qzhNz2z/tnI6hCSyg69PFHipw1zWT8HgSX9
XZb2LxgodIOEyJ7yCBFQofWfRWAmiGA4KfL4N2XIMSqxfxpgsZhfhfHYiVxk8yTuhSkYD0fFGiWL
wMPHBQBKb64ZhJtDqufhs87AMyHVMWJQIPxRowX3wPKcCFjWAiq3swpoBPVqDqrIRmnD2VIBfhLe
GFmgBrWCMUAMVIjNMrqc0HQrfvHoT149eMazV1lEI59ioVofLtykP41o8GDBtfmy5UdAKWFkNh6k
NXiJYXyPN4kejdXOiXR2abtSPiIorMEE+7bAr8h9tHxbQXYDS235SRHiDyOK8tfEsIgfhsgb8PHo
ARziy023RMlPLZzzY3EU6Ymdhc9HE/2Z9HqfoWg99OzexRzsofervE1uFILTLE45KvM8UCX7B4DZ
ZqfMxmSVQ9xVPiF3bbqRLuPecDiR40fpx5wnJF9nhAW8hs4dDGe1bmkXGfaM7PtkoZhc+7lNtwIh
VMf4S398/OD6PWj2268CO5Qz91Sk7Tvk6ww6VuOzjIY0SDnjI5qJosVJVSJjpjzZZcKm6xNwcj1u
ufhEC0HPRzcLszvk58DDIP4uo0P8yfd+PKgT3wZaFia0jrDlBfQGFV/Xft5dBX3odcit6FEbznAD
F29ibB+4fKi8LGQn0Ik1UvrBYgk892I+NBWGsLK608hvM/zlqhtvPnORxF9CGVtZtMI61NxlWzgk
osnawivmXz34Ww/kZtnUSlWNdHCgE9F0aoRKy88EX7n+hNMS0SvGYCjEjasc4PYjxyf4xDl1U15X
OwkCnHFd3sjj3EgdEeyvfVIz5cdfpAlVjHWCttG8b27cjYLFONIkUFB2D+jBpHhSOBjoXCibPb/C
snArfvw9BN3cnY7Z49GiLbQkGDQq8YQ88WHUjLOlmjCT3Q40+X5groPalzqbfK24TEpYEwvjvWH9
3xSTQvK13aXS/S+FYWQrRB4b28Sq68jy2o/7eWxRAy3jtauBxitWybEAnMdKbn8BWreo6+6jk9Y/
Ml3c6qivkZ7qmiGuWYojhzx7fky23X+hnPm/rJGcUchOn+61SzelQxNh2sga5FSYz+q3H5lHIQe/
LC1WF8gcm4Jwm+kt7fDt6BGeV5ZUCqiUBc9f8f/A/x/zs8GGYz+zIl7PH3XQc4V6ARaxQkFeoZEm
KKkxr6XBaSUAMyZGCoogeLv3CERhbSgh1LXFH/A8HJF+mKKneteEALMz32uQ4FJz6/bPNseCkiXS
w0/OHOkO5Ga1rZwG8o+16Dydyui8eM5AP0gAWFpSsTWc0uUiE9Spmkv5DQWbMQg9hTf3Pe2D6jQw
NrJqvyPbzpRWmZvByjMoH2H6QHilpkt/D2n1inLG+ANZEK79+UJyS/V115EKYWbN7H+bI9Qmudil
hCRHt7NWvf1BWI7rdlrgltyC3bRdRx6jQqd2uflA4Uk6pO6NAsSZnJSPhORNdrd9jHr/WSWBC9JS
nc7NRpIPSy2NYlJhzPJsCXDRpia4tRJx+KB5mIls9LpSZ6HXveCBjncGhu7AKR1PsUjBipazhKy/
4Bj9xL9snsa54sf+FvlnD/XUW2pYLZvcltFpLvYCMsJ0Cq/9eSRmtVjxvHSuyty2BoNOVb1GDeS2
1v8u+ybEVTMgbwMPUSFj5mBqIk33pwM10SDAd0AhHVbtJMBT3YV8pBaBebqZ8DnGeG6m8PBoV5m9
AMBX/gVtwQ5F9pe1NzA22g0ofayulWhBytVTc6SGCWM+BJMvH/TjKtCQRY2s7DVJmnZkOzsXak61
U5gMp8TO1JIny81wslu7zMjAQyrkAV4A6+6dOJWGg10wZTibwdYbcoPR3tqA5PsRfNtZjHagHHGG
/ziZs9TodJTTwFQXebvBoeELJG5ARB7sxXIhwdMOtd1CdCwg8j1yb66tvhB4SX/CNt1GJGaXGAMW
Fa/3jFMpb8fM/zmIkcHWnuJWZY57eD8bxApj+IaqZ5FYqr/AyMPZhUvMsEaL/JkjKbuoFGrUPzky
Q7S+Sf8OJ0owqVKHdZNuPC6jSGztY/BYLv/ZC7pvEtdtHc9f2OxQq8VHYvbmtwLzy8KaNXD9hP+3
cm3g1i93eCCNmMlfJ8XlfUjjYaE6RdlvmQ8/ACa64QG9aZ1LyOh18EXR36otozi/ONQBjTtRtuT0
0nXCx+DcvaQGIZF98TTohOlcpuhLxjXIIZANs/FzC3/H5STzsE3kcgskXSch5FymIrCrfiQyA4xn
sL4WIXCOKC6IfJ8QxL+cpJOczZ1K7L8bmolnJzR4RLfgbVMe0VkTPEZm3BQhZnxHdxvtrhHO0UHI
TH7XSQApc4qXQWeN9BIjMO4t2olm9VuWSu+sQ4bFhPDbUgbCJxnJYkcmJVSU9EbJyac1Bp4Qs+2P
U17EZTx/YFFW8yczlfNy+LTzb9If/rnU2jeCu09/7UYFI7r1y5RnJHHNiTpHDRRk6CUX1sKKSFKW
fXnen4fzwblRoW5n4b815CGyW99R8wwmhFtgn8EnIvIlOMRLSm9BwuCDYfY/5QLuz078lJp3O/38
x7BZLqQLcPiACzAYjsEzVv0HIwrDHG7oyDxKegs1FfY6YHIr6/zYhPw2PipBoeDkgILuzIcB5egM
2q6cDfz6kanVYStK893WlGl97wok22MtGWXG/PV5sLtWdhaiXJmFyStWjsZgTajoW9y00IRA7fZX
04N0GRA38/skElzDAcCPx/l1Qfw/JcYRTpXcLYrRTp9nWWHLBRXIfXjWJrXggii9XunwRQGtfIiZ
lIHwKkrrEgKcVWPXUVVzP2qkCStxHVTT/s52AtRI3UyExOTQBktpwyP7wvjq+78FtztEckIMgdTB
50fu5N9HHjX9o1RD8Mo9S7EG1XaVMAoaHMkhbLCIlZ1QvSRHZEunTJt70E/RR0F5us/sS01ZEYFv
9D4xe5PLLxstNoTifNSHI4WNIWMV46MRSuNn78gZK/6NI8732A+BtXpxDcAs331wBq3fm68gnlxU
FmCcUc2FPSUFU9IkjDvK+l8Vh8YPeyjacetC7CedCqlJLnniekYy2QS/90ME0fUgTwnjQ+3e/GC2
Hb3YduEDbEPthTPOtDADDmSmLUCbT4aQhBhXpfipdftSrp4nmlViu++0ifjJa9Jz8ff48R/DMYVu
3tzDCOeNtWIDFfqO1YLAMAn+QUGVJFXTA3U8pPwLv/ZuBm3YljDi2/aOAr4tEqMcEJjrRJLKvl09
gEd/dOS/sB9kgGfM3ZexUJ8cxa6I49tkvAsMTFMKNcuaOCOV1d8JNve2kgflDRp+Rh51tW8/pTtp
9pztuRxtSPo6wiYK9DjqCrweZ4LoNjCMjRvFuiaaJW/g0dzmEDGw6yxgEB2dARLlz+zt10ikRalW
YcuHml5Zrom7mjbKmI6/6Sm77615lMeEyZoNQTMdGOyj6WlsLx9w7MqXshjC88RFwPS1hswrtLrP
BJXZLx6xk3lwK9EeiOdJHatPuKo8ofa6GCv/3nuOJL2r9dgkLDXfqfkBX8akH8gTbJrb1hrfTTah
X2W9MaTt/kZRHT9LExSiUyM8Rjv8qNFYWdm7Z3t0w4eDURHfeaelSztIut/2O4SMTJ3IprW5tCFn
Gff27j1Oj0gaqlBgiSuYL2QwlV8zO5/OpQ4+NyFi9qc1m7P53oF2TEJzcaRUEaWhY4z+niWPgscF
iIW/ezD8yBIOSje/+wAchcZNMGvYdTk7tYW48vU6JgfsX4Mj9XdbYbXhXTYUxe0y3enExyS5Wo5R
WG45JPgfa3Ni8uj0J3iApAQD+XcJ4UNdGrq2Wg3MZm699zVmOchwkBsAymnXGqg+UINxA3/F0x0V
a/y29J1rIgeM+bcuOjeXEtBYCnGuyYpjNsiAzWikF3p8UbUNDgYXKKnh+/iIV78u88L25qupZfwZ
WNam8O4hHHT+c4i+OnURGrKQE/WJPUK2Edvc0NbJ+3mCr50SHwHrH9UMnWdg8nw+JWi2P1l28vX2
Ze/d5X+0AAcgfC02bYN7xrNfx35oXjTBq+0Ba/9Etfd8GaQUin+yBvGPFX/q1XChxD8Jo6dYuSMH
wfMMK4sqYXX70+5LjgXvP8yOBQxe+s/x9b1EoEc8Rj9RKA6KeW0iNy+/HTyOvd4YRSr0AMHAf1cc
5bzTxTe50UFGFN92TlWrTeWXAPItNa8RsXeMOH36ic/sH05S3SnM/yI5a3EJXbBqn+49h8JIeP66
D032Yrxg1iv+VPmKAxCvP0C7F3BCkp70Uwz0f4/LmgzBIkS0GKvNEfHXb3KcAbjzGnpf/9LuNsHv
RajP357ob7XJZoCz2OgJztjKrtzgm1g8T0pt70FVsIIs7cuTKg/IB/d6ZuGPjYeov9mffX6UCZt4
PsQi8/qqNMIOKO0tBXFd4N5SXhLSqbskFthWPzxy+4XCn0wj1DeDUe73LFQKwhrXlx2p40xVFbo+
O5AeE3EKrqEFyDFYA1tLX3kQiImeS+jG/EplOWg4NoH27xXOBYh47vKuGkeA4F3BQoWL7uSeAC80
rjJJ7NjamyxNoxcvennjGBq1yXmjfpTOkk5mIx4fP4vI9FUNhOCU8V8isPJTLzqwD1sLwb+vFMPp
6hUa2/uJmHXwPPOdbO4eTGcfFAZCQwrSXAcvihBsZGLpdQS7zF3h66ZyLLAWQ1OaMQqqb75Ua5J1
6lGpsIEbC/FnIfAN6XdiUbAL2xkO3RGBz/88tuUXcWQFcvJ4/kW0XimKb7j6SVvkF5bTZNv3QGCd
0RlZ9xGRK1lWW3cutyJwWJk+BNnLYPE5bSnLHCZegvTvhsTmLHvvhq+0D7AKPUo6M6ehYk+dpEKD
2VMlcYH1RFRGnPH+fXIIMlEvbZHyZnToS7WHeKMsuWcxpbgpjmXocekRXu3nckXd5oOQ1IL+YXa6
36YxsUspFKwVWAGJk2sOjnSx/BoTJqHOtcYvdpqZ4nhWHCgcs6z4yk2Ym8k7Dj4Awsa0ehpWUcsZ
hNGCK3aSon5jmD53kIetUn9Bt8dQRej9yKSCq/tTiEBAyekryWApCqCED/hqzA3Mdfd6NJiBMe+h
f9L5HhQ5frCHigSHIDxLNfYzgi23OAtHrC9Q1vCuXnoDOrY5k0/nMXTBwG8pKXPR+tSkyVbsoDUv
Jsj0QQ8Wu5ySkpYum22bv8pMTwCG0I/q0btOjJOHqe2hqtsJXpnoepWbqJC/q1QLiqEplBKSjeWx
vZuJ/Ky7qyybh3eHM+/74cgKmAp+QzQGq7hpy3TdgAt4ZDuvg2uvz41tsrmgis1DRuNek9iXc9NP
Md71ZRJ/KnXQ9me+Vs57vabbIfWmD1b1WWYoEqqnM0ZSp0oTzUDIuWxotWofeKDU2ogUbzx24+E1
BJdDnQU9kqbceDniTZ2JL+Rg+X/cMUSy1wAjh5X9vDfUPoIhRIBHb8tPlFjUjOBwF5UdNDNbXMXm
uAj9KDrVJQixTvrPqZ4nfPPw9OiTPTf0SwmyQs8D/iw4+qCftqM4gveTyyyxK9aMaGD6BhSXNTDm
BykZeC8EC0SInLvi84a2gVK2d1e0/3xYv7RZ/WkSDBb/laFXJY7qALQwwBHSys2FaJ4EPITpZZGK
9Odlgz1HNF/MgHGn6luE1hNShucG78DEY8ZdwEe13Y3ERRQkra0p+RNuzATItAg9vkj+k1zhnINc
Lyg7u9EoMC85K7mTKA7rUff+Ehaah1RyIfVrUNFe7Vh6fYBNdovwymywurY9IcUxeWB4HU6Ata2X
PVkYWZHX8uTT9MKJOShmkNdee6dzPPOqv4tJKSWkGetbk9bhPFTv+mDVvI4GQ6e542QbhLDYH5Ur
c8PAaRJPrRUOrvJ7sGwkWyRFFs4GrJBQH8JRZYpzziNkmNc21tthdvyZjPZ3yLzQ8a0Mkq1H5FLB
0kckQUcpT42Rup1IYRAD4f5vJ6rAddYcoi6UINB3UxIa1MvIODruYyLKu6OoggKcvcNQhyj2yU0g
PuK5QNJlf1qGZ008sSgrm+Hybs7TiOZrNLWbGuRAcMhJ5Z6K1Td/SWN5/Fr8IQIt/l7OGk9B01NL
iEhDAiiop+9siwylvhR1YZsV8p3puf/5uh0UIF5wUTaHAcFcAQ8sRhgF2zVhqaX6p0HxOcXK9HYq
R/MWMSwiTbclzwlQIJ37N1T1jET/oxp0yizu0Mk6lxT1tr6fGwd4yjbILs1TUOJVR3mYhTpGJQfa
7BX77b4QpeUimfJJkNiq2xxdVVMh9Z5uH5Wxa99dwA+HjcMwvuTq8LFrv8xtFxoKO1LeXvhNxCIF
4qYcFkxH+m4avIcP1rEVUpOOrKVRlzy/Vwvp2NvwUh1/4xR4k+3ibBVWFzdf0gtjS7WE8MoEqY+l
mpjhb1alRdT3n51kNel9S3tw28F6tV7PjJ9gPhYmoE/n9/K7unoZAu+HxARtWEbI1mtpTDPm5RFP
ilW8vFXRMEZYJJf7LOnswsX5gAf5FUeU/bPB2+puOee5f4LY7IFUffpcUWkh+qNZycdLdj6jIWbm
3FoKI5Zdj5eQMC+mLb+xSUeeh8LmrRldsa750kh0HgZGdtaVp12dUEGDg85KPUoVnnb8fJGJ5zuJ
Q8Ih+wmnJ6ykuYIiLHK3Gl0Q/ictr0qu/NwT56Ki/XuA8eS7XxVk61DmmouoKiP1hblhWJxoilhJ
j2o9HjcXb+V47cAt2D5KqEXDgpFaQ6HRomFLI90345SlhX2PSygpDk7FlOOF3QHYsKNUWZFcWOLV
0GHdi5/5WksHJjrJfBh0AvaINE7al/uYE3mYnqxfWQPRmABfJ3Q18ZG9cyi8xh2t8bKO3hMUxSqx
a6nqneh8GWUK64h9skEQhpa/TEQqJxOMylndJ9yUH2kCDXG4CDgFnEuLnNZ3y4zetD80YRACnZC9
3mKow4ehHJZ9vo5lPT/rMZc2Ng33DXVyHE0WAH4d9h99qBV6k4Y7U1wMnbYnAGmXOhEgS+B/fcay
CpIynCOvicElZeYOdkxrHYyA6iAVfi7dYP5rZviPk8ONOraLg0qhpsqMZxXc0Kh0qvbGbq9UCV1Y
Phh5hHGwSdd/nhU5yNpoZh+4OdrU8ygb6R6D/9OBddprchBkGvUVZ81KnafyHHW8JnzCISpVLyOC
l8lRUjnDA3lxYTMrbtsuImbLg1TmfY+nzzlEc+yBCOD56JYLzKBIV2zAUzcP36GZFNMhn8kL9D1P
3tgYST9bLOvr+X6TW8E+hB59k8mBOXSjmaYA3Okh790fYW1uI5cO2ySmWiafhMRJVGRrD5VHKgs/
HWVnxK1GPc2Yr+Z6IblzS8fbfhS0ZjgmKn1ySAw/MyR12Jg+OemxxbOJjgUW+S9Mz7TP39dFGrvf
IB51qvzCL9kXzrjodkOrTbRx23SxYYWyhfUklgtr+QoW8SLmcfIv5Te3hJZXfiklakD7jZSro8Zn
WI3h8SaX/AnCOah1vepMEW2cLRIq5qhvRoIiibZrp7eoLil32RSTlY3rXSAht0g1oclxhMCZGmXv
r+F2dkMmCCLwQ8CdLPhKBn1Lu5kjDDsj+zNgfN7V4HEVK/e/YU4CcFVNU1WsCgVMJbRjrz9YIksd
bXOJBdMkHuZP1e9iycPzEA93LZ7tOUAw7XakVpmxHVrm/zKHBtfYfuk70srwP8LsXWtvvdqq4n7Y
MB964/Ocpn5/7XpORLdyNC0a64h9grJdrvvbnUJ24Bh4QOSwp37XnuIIXXCRhzhDbQMmZtM0GNUn
0H4mtk85hLdTsASIpiWXeAc4zaqvgUqtGRA3wam+BQssaKBXvwtxSxtE016Ag2yLxC4X4/1Gbee5
3NQPnSovixhIRAKBEIUY206eSVzH5nas4EF8Yzw5SSC0tm7DKkeA8MTTYNuhGUeV0eDkPhlYlV9E
HzdH9EzwtGNO0LumCHnWHJQqNCdpxPN1+PD5lF3j0fhP3rMAzFiABlScLpihyHuaLujoB2TK+/Wr
QZOAynuf4K58NGgtboLkdL0FZDojBYoPJrmL1Th3niTPUbUXSFzG6VxVu5xAZ7fxH6QmUTmwF5+I
4MIyhVt4vobH/0B0NLpB3NN0rSp0m8DaxtXD6px3QPfkNDCP98OpQOO/wSit+vK50f9kvZde5wPv
CZfc3Dyy2Y+HSfjGqO3DdUElblxxOuGsn54Es0WOptwKkrHTAttUhYQKNh27pQ4etQL3dIasnRhv
534rbJTxlUBa2s7OU7gD73vFR/SNknbQts7cNPxZla+fbNmt/3KdOovMc3DqijMWcGF2r+6Bd5tt
B570oQZx6EDBrwXxldDKEt5d77UTTuVmcvFTf6LMwnrR2IKkMvDNVO5Jq1q+H6gaJBrUUvVqtx6n
isnWY5aHCES7wgHO9dwqrJaJhBf0NHFVTTtX+GkiL3xSHFOs2PkkJFNXjRA9HUeXl/GIC5S28Spj
udSmBkvndlbDYGtWXtRA+c9EbICWo6L1/XxqB77FEaAwrAWl7GEbB0b1wtUNjjJ0VSv3dfBwQRPk
oTsCSnY+cND1LYYtgq3SJzWqHc50r/g9lUCac8NGg46DnHKrakj5DRaqHpNdHDVy5vmouEs8SgHh
xcgVx8wNCORlu0orKgaef7lV/CqeX2CTQiVuwx66ElDyL7SURnxSjCXUYE57SLav1bdvK4ziTdgg
2YisuLCYa+RxxT6T2J9A907ksT8L3D3pQGTJCrO103A0bcCCd3SQcQRUGOgOwpyexyTqI2ssxyqD
LQ2kCW7rZdjZZHdYWDTCiFYc+kqDJHMv8r0jV0pbOtPzg9L1FvtILxJusSguxzq3wamXCdc+CPY7
AQ0TliOv2fDNnkcKOH/iILVIp0cRTEGe4CgW5/M0b6pYTVP0vp7Orjp4f777aM6L/D25htr6cc9F
4vhJcC9iKNnXqx3M+eIplJPjzMAFqm8mkRU3yD0jWS3zyyj6ux8x+hMnNqPWcn6Ugx43LO1OS7y4
D3TahF0BR5I93p9rNZUki+eY9ht85c5sUNiDGhwOBaQHjMKqXeSPyemWNyV25ME9HfkkN+37rljQ
t/lyNO0ZRVItmoH8eopaiNHmjK5fVtFqE+1LaPKnF3kVIVshsnSnTKrmeGErdTz4nCcL+UNA0o8J
Q8PQAQ5JRVEIuyRvF9Nv2rSsQru4Ze0fAZL7j1Yl7jlltj9vcOj0oHVGM79kVgaMxbE4qg2gTaOx
1be5RQqAkEPXawUZZ4V4qA7h0Z11iKkAgUSINiuyPF7lz1Ub4DZi0rdWVaNHs2Rovuhh/mtGUaUO
TCYmEtlrUVc/Ujuacvm5U0DytJlm00YZ+zgObFj5dpk7nRNQShEFn0ExzGk7R3gNpaTfP2GmL1gQ
vbA6Dc8YTNZKZjbqSoBMYj9vsk8+py19nEgqAoHX7TAYmU7MV0KHOCmNLKL1OLoCRYzxVZ7Dv/9a
4LnKeMUmRmaIJcxgYFmT/BA5dnRSCIBRsTi3L/NRDoFHy6h+ufZVv5XPPSHzK8XT3XAt3ecKO89Z
rOr/ixKfaMsuBDlwSVxrkgoz0RPhg0ahduVdOR8HvKGp8WXOHttp91MZikYbfrmwxCQokWS4qtXU
pj5qyjxR9zJXyMGv7RUm+kyyccmEaYvsw23vDhe1AoC3AREN4xFJnEQeLd+c77dsR0cICHNnl1lN
AGHwpzqfN/pBNvBK1lXZSf2+m9R0XIg9ImlmaxkxraREiJFaOCFAkgfSFIIlD3e9p/veTdytRy66
g/aYVWCSWqArtHSoyINy0dEJDBa+GzWqVrXOQJGJzoe+axiUXJ4SU9D9DXB737q5gXhw5kzj4Oab
IVO0WZwQkR6P5SKBtsjL1tDONl5Mt3dCWNt8LUBkJpnPTkEb5tnR8VRJq1PVRQAwMe7iVZhO/wZO
fSfL1cjKld4eRRJ4kSXuhqswyMNjrusqGWpAtoVYiNzdQ9RPIRWfkXh7jsZoN+PDqDxw7jdD37bj
qjIvcUsxue5TCF6Usn13bSrTsN7Ga+CS9bB3ltC28Ijs0s/NBbOjqTZXX1TeC2YpG7sEicgjvxbd
yRBewcC7wdLo35bE7lVexNgEPrAoV7K8MApWIsEPsjvJq5HSEuCSFWxr5x2JTYpGVHD+CJGncD1R
wWvPduWWRIMD07r93wUBR8VTcLbK/jUw6sOEMbXUtuuvtEOcB7LE2yeFZ20s/NzAOtm5rL22YZE1
3eXWGpae4aES6o9Z47HVlBzQvLYnhA2JLOTQV1kFeNsL/4zgaW/7ad95p2bksCLJoUsXHBB225iA
G8xFcBHmxvLHh5xkRbuS9uCuti5qTYSDav4jKUsWq4KlTqsyw3rX2/tZxZEz2x5ZWeDS7Ag5MIOu
gA9XTIc4picoJAZcEKX5hLQcKC9L8fNlN7NtmbKXofPMmS4pt/mDl4zhi5BxKEsLwu/xGB8qGlG2
vTXqHco/5oJj1oOhMgduCtwfsw5CvqljCTDaDVc9A9gmr0ifoQllATk8ELgaRaOQVCP3+sqR5rnL
KeW77ATHo8CoOyXIp0NWUjpRW6soonuoQ73+k0R938ywDo39HcZldySpYEhXUsMTw3xOhE/AH96q
GzwkOrGo4mNKsGlr26sGeDYMO48PaOAsdChCr3537yEoVdMSGEamoc3pTDGbelxrydCylcuydLXu
FfH12HoEAPdgX+LfW4p1mreBNfqG/UtzCQx55K8VY6Wv/zpM8mSuTrTygnhhMV5wlQ8hd0x1TIbV
YUq07hZOzh/0wI2cA5fs4TkaqisP/dfm5lcEAHNVv6HMM1uHLVgA9OUaabtwd/zEX8899D79gLtD
aVD/vD/PF3h84NoSt/ZVqDgtXdXiuSC7Ao772sCNtEt4FRWn0It5T+Hldj2QWBvRjdxn/SxCXy1V
fUZySr3xeFrD/IKbmsuvOZf3Ikv3BA0SnKe20pTVyqmW3o9zCugWtpZaFEJJUcQRW+1cRNiaP18/
0RZYWLoWDuWmH8iuSl1Sjwt0oKckzIbcz/LTHpmfXZzgabNItsSsOi1VKGczapjeqfxYLiM+OEQG
i/zCn3PwbrGxkGoOLOMUV4+o7WkTMKMDyKIKb5PPn7A7taqolmg4cGEYcd+FeKP3JT3NACEY6s6F
5GQhsLMA4pv1susW4miEI2wz4iJIHRMksDfJU/s60Waz1MdnPpEUsiqy0QhwDwlwpIRHgKRGjdxY
EKi4VBF07c0x+OQGQ6e9awhOvcz5aQIENPbDSPbiaRBJkLWOy8u8CdYhyBf4StbuIx1mW9u0Qx0J
VqXg4bA4/XoRi/Hmn7bqHD5waEDX7dYrl7KwfRLWFCNgPJyNQgKVJRyPwgwUbdN+eEnIVOY2t3BA
9PnRwHppXGlAr/EuPhIG0MYFYJ5B6Sl/l37B01IszrGPFDNqdSCDoiWULfdA7pbFEmsiFNTBrRzA
AtuIwJaRq+9zdpVByXnb0EIbKIAnJWtNOkHamcgmzjk/vXUyQuQfFfHNwdefGOAgqFTCOSMsdGIl
PztBvvnu4K0ozh+jOTj7Uly4LH5wwCHWJCM3Xw81pXVkJivVffi3kh8Pa3NXIsZ2cNBD2XaTVb0I
i7f2qvjb6TDj+YcceCi7IHNzMbEiHJtA9wzl5eIq/vH4W+0kvucz3WVwFfItwpJLJ+Vfc1w67uZD
PSUPauqYlDmN+gu2Uehkr2MaV7fAjvlGAxTKZ8BBVss0Kt9YAouzAee0Z/7KgHA7KZlVM+2jYYGe
/0X72vnWKJIoGkhlQWHBnlcPRuXOv8SptNs+tQaO0/l//3BA8BzGccksSupCO524/WqlKPtnhHjC
ZqCQYi708SIWs7D0wPyPX+E0mB9Geznr31g9bMou+XjvW5Jf3NHfPEDB1mvaIbw3+NvFTkCF2syu
wJc5+UD+Zd8cq2PP42z9TBBf3k66MV8FwaQuGD0HgfDmTLYn4+ycwHADfSslVVCMqbuh9coeZtLn
HBnQQ0lXCO7OteRIqqggG5WNmskNUlgyXfDY5uA36UHyh4MMDay+qFVVLdR/+6pyoJs85SF7YP3/
5tPfTXg+2TNeqIHHid2xlPuhQWiVwstzFSGIrH7w6OsbQatOytyRS983keFy2lgI1kZFgIFPSZNd
K4Nl1L72vl8mOKIpatS3PKT2KH+FVWpldiP0KHzoP/HY1KEhda2OEqKw3Mp7iRbJ/XRJXET/GkVN
Gdk0IIiFeC3DB1LD5wtDO0iQm1Pb7pArzIsBd1Bms4Plkndeg/1h5HANABSRHzkhSML7eIVpGLK8
7AJCBGHegTI0UMSMehfRl+RbA12jiv0gm7YBXo29j3aBFZGjk9+ttbktwjGY0FuAmy1ID4anByB8
sWAbtZkdhTtlaWge1m0AOullddlqiuQEHffKRyRh4Igrb0lmhXLNxiQ74eIAX3E3/5lSUEQpqk6F
RaRcU/lmskIwcW6VuBNWn3pdSK9bRhjJ6fGHAAD7H/Zrh4agOfQRKRoLy8TZ/7u3ng3aV0h01NRw
nI5iKyGXiLtOj9Yo8i7BQyv399eYjfx02tthj6T5Ivhfe1riDPNjnNAxrHVKT7et205woduxAjgg
xhyj27LDH75XNIStiXTCs9GRTCg3wUevwoo6KT+jQXbzcWUm6ESYOqEyhk8MihZ29kTSWtjmR6Dw
NLGOJR+G7aZCJpeMwWBJgaLpsPT9JNsnHnRa2SssSXxvCcbq7YzZgrnbFkbh0fe+o+sd/Hq1sbCR
DdJh5x4NGa7ZtM3js+lX3T3plJLBL+ttPk3CY2jIndZPyZqRoLEOKkWBXLaq7LPz3H1EroyhR3QK
3JJAJoAf9sJ/qMkWv52TkitM+JA2KfNza+80FB5/EIwY9JZeSyfDozG1nNhmiBAiyc1PHZF3qpIB
auogWuZaywm1DohYP53m5XbEqwe4FgBSx6LBGYXVclmrF9fwGQI7CBIx1Xr/ssR/FrC9KN87rnzN
jAkBGBhYZD59w7+3hF9ihew/gNB7i99TGYZouBV8qh2lh5rn/h6CW0FAn6cWRSIAwxHdivdEXVVd
1RZduRYUX1k46xOb0EeHzzZF9ArUtfgOHsEVPNeat6rOAx/QA3hWt7hcKnmMuf0zI2SABRdnQ7hC
e42uXRV6RqCbUhlqHJCGE/6D0lTz0B5Q03bAb6r/tGCxMLBRdOaE82vc7a+qLfYkonwkEbJVh+OH
r/sMwNF37VHgD8eIqHx1qQ3/ly60dA/xCmCsueW0WhiK2C4XcvCJmwmg71JDzkYiQPYwWSqztmok
H6wcGnmc1oPyVykr4uzb9QlkG3LMJSGYEyVrHrHwCRxIQFyJgqmNNFGl5Gses4iuI2ZFIZ/JYfsG
5Fgy7+cbMjd81RE4H82GKyQEIPslhl0zLPYqkaDSHSz0fM6qPcy3v7DWg/N5eXrdasm79fI6dyNB
nMjgCADb6pBXCYo6GhdssOyPUrSavOIFxVrzfaCkYQ0PS/dJrkSz8giL5Yfn/fILlPAtcO77lpZv
WbPGOtXrN5YpYef1G1X6UGiDBzOy/OuywL/vAwgTIPHWllO6LTjLwUiwT+lXcN++lsJ2+t5rZCAb
uSjaZPW2EARyinibpvilnkhaWNxfU3UpH73UWLdIW3P0Upe1JDWU1I2tWhyycrtfKgJpRkBnUOWl
qd2qcfjtbIC+Fe/N4rhnVBArj9KaUD56tfDacPheimkj/l2HAoR5ANiXemQySJd15HTjUokdLND0
bhzJ3FJM1hXHy9SH8OkbnKQ3d+DWYhQ0dFTxDmc5u+CzMkfZ4QM7q35qNXOHVgMwOEOQ4TKYbIxH
1fj8WWJD/fRUbFEsnsp4pTEBi7WKH0rJ/wVO6qSl+pdrKlv/Q5C25CzFJkE7LuSn1dSwexuWgild
9adDd7BgsqHNQnfgxvYftRzoWrjBjCzwmf8sL6CxMa7EYsUBi37cpgYW7mZlKOA+8BtLyw10DRYd
SDst+twvsI3dtoibCS3IfS23NfNDM7PIRrM8Tv5O2qbXaDU55zvYlufo30uKQ4JhQQSEGJAcZW2w
+fIspl7+hLUcdrclpGmPhA9AItf0LgoPPBh9gHBsYHdbhiar8NJZjxpwXVeVmPkIvMaky3UVq9fv
0PPaAp4ecmsAgELgBloLtcTwPbzVIHgT3Veko2WTKqsDK/OBoORQtf4CLJAeK9HLp+Mjk5SYaXjT
FBkl4hl0eCOc8Y/Zv1QmmH1mf/tajQDagY8b24VdUS1P240AUHJmRqB9ed+zTYrZr4WT8JlWS3CX
eqgRBmyavyimYwbvohGXsEu6M6LnJD04lMMusfxk+TrpKmA4REP+yshgWQWeQBsPdDBNavkGq4Dm
cC7BMa4Ldv07TiQ0CuiOzjJt7GLwVAV+W0JMPyDrnydLJoGtPZRzNqJsI81FR3iXws7Q6ACcUAjQ
F9xPUeuwkGmMmh3z7yvAukxbK93VupKoYtdBxUGXU3J0qJFiZwz/hliawsYgLP92KeCK65LD4c6t
uMDYlDKVcBB2RQMnU50oUQcZ/4wzaulA+khlA9JntYyaX8EXjJg9z6EAgHP4pG1SQmOcRDoSGQX3
738F8FQen+aj7bjq5P22fPw5Gn7HORBVko5m5hdjhjo52HdHcTyeoXUXn7O9JZtDnt61SeGlNnNQ
6qbeJKKVLrlkGEwFnu/7vk7X0pFFW3mj5obsg78oYKhnd/D3cWOpKAidX4NzSs+Z6iAYKPA5/NDX
fzbwblvNg5JjE/aefhDSWAVcU9fN4ShvqW9DO/bpvXjpci8qVVtUzXrCc8qugxatB1udNFV8fbmZ
SXywAzfW9QSa9iRfOuhzHGhJD84NvVdXag4DNun8U7xStzsmqxT34j6/O43srhqzLfwgsnmnwjOk
v3mu9q5/x6LprUhIuEev8MIZkd+lFGR2A2XBKmaInU6TapKF5LA/g6+Wf+9oZs6RM1Kjp9RqsjCp
PzoP5m7yU8Y4t3tTtvXnQEVyMMHC22BlEMsKTAl8JPjOFQ0EhZd7y1gmxN+716wOeK6Dn/n/lCCt
vo1VN6NWXuq1Ap6wdUpXZ0Jy4pgEqgkZvyP1dbntT6E3PaJ9Bzq3sgsqxKQI55yWwzvqUCR4TGz2
tQPxdtsHDRav3LP7dUSy/kjHa7aCVUhV7oZOIfLz0wGAWA2QrHo/mZNlw2qSHTRcH4f7ZJSyHUwX
6n/0eSX4/rgwKjKbQNMZmICqes2HF3kC753M9IUHX3sDlh6sUxIuJTomn4rHBcJqWNXALEIY1kXw
NBYRylq6gR9sBc0DUXdZNpZW4fZMD8rOFvesH3dUPbSFoNNS8urk3mctvYxuRsb7HQg6xQGRyaxB
R/RqC6weAUcDT4A+s+b5tCiHkj4wgvYAZfWoFEXdKAEwbmkx7pN/sNmKxJ3W4KMUmZ68SZYlXeVO
p/BszApFoM7rpb18AjxzYC7DciLsTVx2gIKcrg1MlgrnZiOQuDjGMW4iHCNqMwlrYqvqDa05SLrs
BqlO3U4yV0/ThACm0wBhl1awsL8Mt96tIi6HTolJqu+smZrpaGEKOldOUWzvn22O855FYNh3W01U
HEiFFHO2RYBBmK8D8+mWse7Qs1N+AN6bVeksiW2qb9lXDAo7z5N7HcMseDdoLKi+eOa5M0LuPW1u
ZEsH57KUCWomqMtyjd+EPuxexPleDtWEgaGkD+FeOpHYkey1g4Ev48ScNfqPDuLxZ446ag+TIF6c
D5icu4AWZ2IJQxVRvE8LcjafuNo7RBmBl6awqSCMFo0Xm8C+wrjHN5COVT1v4LJ9xFbvYmBLKwZz
HEZd7WVBA2FqaX713pPyXwLKAtIQiIHx8HBppL09iyEJQQAWgYEvlBbQXF/DHvS0wjc1CUx/U8sg
vM2PwB0toCCt8fYPScXS5Zs3ClfWdYscCW1NVGNvdFO/CrN2U3CwzJYfqbZIvIYZ33DA5m6yLPLz
lh81euGj2fntG7u8jMDtPjy3T4Bnah57TagQW362Ei4UdvCiwNwhaJBLY0sjMCJAyeVg/UpgHGtE
qXdS/n8uB0Ft19cuqTq/wYOSdlqE6/66E/Fj5JYjZfpHdaxDdi78mSbgdzATwEUNEs6/z3modv/8
fWNuuf6NCZg0bW7UgznY1TY/K9VzlrzDmNuxSxs9vKjOfnGFdOHMldzwhHtfSKl2KAnk6xzATxVF
hCrqAd7Eic0lxu66BasfBIioa/R8ZafEzlBp44RsLYpJYMol4S6OphetkKkO0qv+/e46LYozQ18r
HmsBBrvWlitWBX+XA5U+JIPfENF0+249mGhzqsOBl7DyuQ9cHEFokctM4nnELgOpLx4cEHn/cj/s
KS8evgsGenCfClsVC38dpufLg7QT1V7p10Q2zbrsRGe3S+7liAZzhRfcp//GDQFbxYCvlg77wIM5
YrfJaL416u//tkBQRPgqTgFj1zu7x8jlzGwyFvcWfKzzyVudG+Nu+QLsvvMR0RctuupmswO4R6D8
nbMSA2rtLQZlbxV17CYHf1PY/E7CRC7VmnuKWwsMekf+TGzZYq8+pNQH3sOJCvqn5dWd0hStWTBm
JyPPp4kjRP+ehcsO4+ovPvQMX9de+BexSPhqTYwxTRbYwp8+nuLejrQBw6OVz/fmF+04pgD2AMtM
qTt/YoxSwP91NC95tWbyueHGlIo7yCHkLnNcZuYpSFBMI3I09ZpQAQDjs1wZbJ9Es7OfAwJpdMZ9
iqYQtVS4B18oe9b1OM9UucGcibaPNeOmXBgQoZslt7Xsc2cZvo1OaCf9iVfU+Ktx9XBw4KcG6IlQ
MdvsIZzGoTEoHUOdYxSblzWydg35tUa6QGtLuq0KFTcwVZasMyx0Sck2qDo3Q15X3HCftXFa2von
sJqKkEqp0ElnK3LLsOnJRFlPJmqft5COb3m1O5DWieEXDqxmpVll5qjkm+oR9Hl34iRKOuDK7PhZ
agCsUZBzPN3DXOZ/RzYRSQ25DPp4qXCww8it5rVZyxQ3DTiLCZ2Cfr7QP3rDebBaWUJQ1J+47bGQ
TBRnsjfrnn1IrKMX1TPQGOp5HfeRyg2G2PaWdyga8Hnj3szxSlxGfStWmeU/Eh9gnjS6jRGZZZar
kIkfUKxv4+KPHVhwR+Ggn5tk0sTQqX9xbUvewwFpqaaWFeGEn0Plzn0JSfLAXfc9EF4np/Hw8nUj
W8Qtit2/8wrb7ICQMAi0Il/jxei7Jyow/R6dm6NFE1J9fGg0T4FxDxaY7etm7LWxK6iUq63SGnqz
41UtCd+hJE9PVUWfDC7Z9EnsOwzZVE6XRICGI5956VfpmngxA6UonyMxtSsOyyJRfubOfI/stsm2
cPFkdwPRh1X9enW9Jiyb8YZG1dGxekhDFufgLqcb/XmWSLuU38oYq/D5q9E+4prh+946+Atw5kKu
Jk8PXs/W7BQynsMMqA6gkNorexG0oYWVFXdB16bQUH0PRrteD8AOV+L6RAwM4k6yLwpfdYAEAxIz
mNMU0nGLSEa53sIoRW+cMlWMlhvlZogTPY1KucWQYzPtziyk5YDrXzkH6ET1Ja78hT1oJOUjrK/Y
2T6uKDrT3jmTwFsSupFFR97T0CAKSWfEMigFGdBn+tkeU0OVA4d/QWZ2//Io/yo/jsEwNRmy7yUl
GdxsGBD9NyXp5A1y5xOKaQikj1/J4Inm71Is74CrmCm5AAVUPy7oN1x+pk63kVpf2qmGRRFB+2G6
siu408bmzLNBnMYCpov9DtvGKhMEq2gbceaKClbT9VekhL4NDx+0bic2QV0jf/RlCZO5UqapRaA+
SJfGtIXmG8xcFV9wa0dKLWqXFbsqRXK2wZVQXkEc5tmh1j7i0E2jz15q6/Y3wOFfJpu2OIhaDo5E
b5Gi+8R3p7Sog9toTRIq/JN2F0NZUIC+46qv4HlYQi20mHx3iEJexgMNwP8YuvDxKyce2gV3eY6d
tGDrTK+uj6bt0AG3HwXPNjnxSjUze1EET246VtEmwaWN+iFv4X2nIUlwxOS3/aOp2lC3pbuTDbLA
NCftudkMSJP8lj5oz57c+PzeHwLlQnEi2NcqZL/h7KgPC9+2IsjdaLjCA/0Zz73AKWJaL4gQJUe2
nSUiSInkcpwKuoT92mXy/2E88nTFYJDE9nB6mtMYG0C5G6l8odAzfEqQ+pr77/vXwzzlkBVNNXEZ
YZKc2L63exwGU7sf6EkJQ/DWgr600ku2iLUa6YtS9gw06joysrK4Ot3+egtnvPsvh2D0Ron3DeOn
u/klYrWpyjcExxRX3wYN6zMtnW+CQ6QlxJhqhHvTJ0a3Jhg+HrzMPlkaZqPRW8BvfKuP0X/95Ftq
tz6LWY07vqf4l4mK/JYxAwn2XATlKTEgnTEpImHxUu4cuZ3evBCU62sLBVKBI72xDN5TwtxgF42s
ppbprt92rDSwWAkvyoh20WtGqdf6iTEF4sqr4Rq7XcmJWg8JuqSyxHH382qWt6WJDr2rqm1B/FKB
iq4pMSEqrNVx7q9L/mdsG0OFWhHdkYkjzFrwyvPgdYbvKWpkAbAawDzsyiBl41ZK1O34g5KEQavG
sPddc5/qDCUKT3Iy6HOZsqzfYz+Vlw+ToJMyrc+d8iXdmYij+iZmwBhkOxgWJ6S1AloJ8fpTJM4V
X32AaspqCA9d/gOFNPqYflt8L+OUWB4mttQbHXwnIl0wR2r0RaXO06bZg5N3OE/+kyMuJtcZIW6X
qkZEWSB1IrLuQOoD3C9DTOu62UHsPZDJ+FAGYVSaEwZiYVChh1dCmVk1u+m5guP2WNFEEwGv2Htz
sr09NCTUrVmVJPkHCGNJFVc/6+ubMfl6SDwxYCwnrReRpTF2q6AUp0N7O3nDgkHVmoZvnEPB4mEi
2ENWELr/NZblb+fmZBmQpQgUlU1U/n/P9Q4i3ZNIFQKW4Y68VW0cZrwLO1TAVhLotNfq6iLLGMjn
rvRpJOlRmtv95mBXwZZd7OA5ib7wN6r5nTB0qicANEifBXSZjpvDxoz9Fnf/TwYGuA4YaBnbYm5A
4x3psYL33vsOcBnWNKtIGWTNiJQZW5Q57FrGSFFL2OMrN5hSSf14fXBLX0H6Is73bpt7lNz62kpn
3ILz1+tMcokwXyFD9uYT8qWExnUHTRK0gwb8bsl9cDGDrieHrBD6+oqneWFuqKIbn534dAtsDRx3
lJ1oGazXTRZ5WifPrS619qRcQjnkQHFwjYingmntdS95wdSmP8UZeCea/Wrs/MgZG5hSn2ACLkXk
a/SyWMfwhogoUUSuuoHTgdIPZtJqcfN5rHiD5uhMGiWg0gnJtXo8/ZBpn6rpae7fMwnFhm6nMqz+
gX3s3gwZ1TeXqdYqzzFSiTjn12Utf+nseAwP2cRvjhk5c/0qkXLLaOnWtYEozueykbgLoV8B6o8u
oahEXk7AyPkCChntxjJoSpV1H4M3gtyxQRk4g/aZ4JriQGVBmbUIBpVI32glgH+jxUOUJK/scWdw
Z3OF129rG2xDRdL0UXzsulrQatqqj10kCTSzXv5h78cxsX1ftk6LZm3m/MOaaCxOLNga3MbMJssi
59eO6y19qJuGrJjDTxllTo7OTcwVMRa0ft1GweZ6xg195zwn2IGUmb3XOGSHrtCxzndZY47mgBJV
TbDDe/q2CEmC70yeBTTLg1kyil2509w5/vs7sefZCr8BsRzRhXhPpbG6BUbUP7V49HW+s5tZaUwY
WHrJ2TLOphuFTZXKuiSHwpzGvMO6/Kp2ZTYF/VgRuBgiWilTYBuyg+tPsgQD+BOLAjpKe+niNGV5
ZIYdFJc3uIPF/0zq8z5wxrWWPspFsTha/axk6spyxq0teUmjkNQPnmPvpkwkJi2dc/+z6BhLlwW1
Y2vWMaCY48lrTazHW/v1Yr+ihfzV4ZjXkksjadjLwizIEp0q08y0IgZQNdEopp9N0va8zzWxcfYL
ql1Um9u4Dx9h2iVyzGfmTxgRPCU1We0H6YT0pGqVZdyFCpHxed3qQ7PppOvdzmcZ9HNtlBJOMcY5
1O5nlJAvPdNF8Er/JHE1iQSb6zHs1nab1zRXAKIEAS6h3VKrD9E6XautjcwP9aDKq5rH9kj3CX4v
6qH6XuJeWBA25kAIVa2fudc3kA2Zf+CMMlfLD1e6uSayDhvMt2iHaKX+SESaxADGiZtytrUTUj1R
F8eWr/EuSkUZSOZDnH6baZPfLuWvwxOGroNek4SZPI6BeoIPpQunhN8XUeu7EecKrX8ldO8Enum6
ZM6xuQ4Hmgd8DaZ+vVyuLuqC1qle9GZ/S5wv2MUT2/jka4X24bJ8lg6Jt4O1CDGcUg3bp/RXh9MZ
HulzycIYidw5275yFT9WGarZbEcI56gEHuxS1P8rOHzj0OIjZMduj4ENB+EBa5SWSgphgcCBjm+l
NfWpyR1eNfGGnU9NK/Ll/QqpNdds9Bq0rNuSgqRDsw3udbTA7lbNPBXwiRP7Mk+OySxNf5FENDXI
h8FGHJaG9viAYJOrJdtrnaBatqtFpmpgGEOLzIu0fuBNSS3/4+nWqX14MvI9bp2OmK9nhlxfIppP
4VxhAqbsv4Gjl16Dl1x41sOV2HsxJptAizZU4r1e4jOZr2MS+WuarHoieqOgCx270M3jlxqfgjCE
moTc9WZRWEgfpCSzZVJDnVLCcnvP8uRE94oZPJEFSK2mzxbKuhk/zfaDKMYR+1Id2H8OXiC7uhNY
i9ujNTlgnMLSiqh89U0UkI4iJY3HdMMMeDECjSXv/4B95eCUDzi/IrqAGT/l20NjCblINJRSYRMC
pTtRl4VX96Nd91uVCedlYPtLkc9P388qp5lHEsoHiC9yPDYMZ9h2c2B51cScAD8X9pZKsf2a13mf
nIvyxNz/Ijbhjl2RsdpF0ExleU3ho/vqGHlnpAX26Ida8Ph2RXukA1EfAEYQ1+q6ggeVjzAOUgvN
erVgrBz0JA20v5BbfhYAZLYN7y3JkIDDSjwcWQfuQu2++OZQaKan8+kqKDEgwVBmcwbqq3DghpNa
pFQGbN5YMeqzntcHw0SbIdFvnumX3Psm8Fz32Cei7zmHks1jp1bxeKH3x3/Kd0lCJmfelS8rstif
WOMGn1tBBhCi6s8zCJ3ykmweAUIq3ByJ9tMaecedQRAF/9WyhdCmUHiSEA7fhCb/mxmZZSISr0jG
khFAM2An+P94G3DWfw+RnAJs5BLs+vdJnylSgpKv1D/ES/vqV0qgqFRqqYLAZiBtZq4sFaAWM6Lx
aL8KQ8wdpA9ejChs3y5TaxvMV0tow5BK/VrMXi++WnkTbpjxufM66lHcNNQbTCt6j2ezEmRz4YvN
AHQY4piFOJfADwPfVEd5OsqsO+h1IGWwMS7OmUDLvKKzmVu5tdgHcqGPYrxMN5ht3Lpnqz7QAH1g
taaRrcB1qurWae7YR1+bCJuvKXQvrlQ8GLwLrhtuKiy34tajHm9ws2Qmm9FUZ08N1XfqTmHCmAec
WZdwSU8ouU7FJyrQN7F+28mQpmFkqnI358cK1tqhUR10M+MxOt6rgo5iHSilhIvu/PiL2wOQmYFI
XJJyOWkapIJNUtHe/GJzH98s5no/W5Of8HJQBpP7F5BR6kE73xS864P+xFO4AH/8zNlJQ1hNlyKZ
jvsJ2zRCWnLZU9XTJ1EYQuhir8CvRGZtLkNnBrWMluLsEBF+UqNxDaizLLbOij3KqUxz0iFqbfLG
ev/B1x1RQbb83dC2QXT9pbb+WuM5nVcCPobmYQU3/BP3NQHTxWyODiFMirkg7WImal5bdcRNPv14
bBKPXlwXSqNLbmuWDT0XcEj/ASMFFnyRd3xOdTMFBhLNg9RtuYVYx9RDg/GyJBBKt0MQypKvsRbp
ErXYWou9Y0DOwd/sdFR+lWoJi/sGkeQYHXePxkT9IMkSn8V60JCpZcCZfXGVN/TkvHP1aOaJ8zBb
sbFGlTyYrAsJBxqaFPgu/Mz9excxNvL90h+9CemzdJnqIcIpT+977bN6S7FklRUEFnOsdVmJ3bLe
iG1qNhzDIjKHTfS1FEo/DDBGHrCoLCMcMJwNcUQFCM7aE31Bbpmf2T2b5+0CFR5WnzDuYLhA3eDt
H9Qb64T1k2aD4bzwoK43mOH8tKWwndXOkak3T8MLkL9S+sjQpFbtceKUN6ycBWe7X9thUZ129O1D
N8ciPhMcpQLdX1JhNUbmLgx57bVtg63J+rH7Gd7bO7aSnHrwAU4/kAi6K4brNlkaD7zHrlU1dpu8
oICjMj/WSLZJDTpZIQFc/CIbg9QftAo4zS0q/5nXXasUsGQ65d2AUqUk9oSruEFuHywtrylAcYx2
7Owbi7Bht+zPQUZlffCvOZz/ocp2ORdPeCRIry07Ro3RoKkOBGrFcf8/sUb84913S5TondZ00DHK
ZcyMfOHHVUJNKzVxr4h1h3rWtupB0ovgumnv/aOqMsQYyvdthtIgGsp3aoq8+z3ZVHsTRPnFTrWv
CLbeqeqL6tHVbgCNEpIMTnTRTJ2J9dGQFXCJHyJ4yQKf07lub6hftdl8Vhu4YKc/J4y4xUqv3Elf
gN729QturDdYfu0WVBkpk+C71Nf0mg3OPRy7MGlp19mrtkzz1zouuVOqfIc/ctwLsfzMnylyxeJQ
vY5PDv2gW50w0dTpdJ5OKh+RzaV0cv0QIgQh/vtLjyViCZrmvZuIg2qQPBE9k9BW0AXDTEcz3Slc
inwBAtWUA3o9TDp7Zxd/dDEbb75nnepZPvB0y8jL0oQ2ka6HC3xoUT1OvcFx0olRyjzAGc9y9wgF
EL0gnMevz6Ud3CkNGURgwNt4Mmh/UsVbHWX76G4yxD3bvPtMIaw6ZbjIDgDbG67H4HEE8qNXkAMC
0IeOREPNEJsQCp/vTAZjCp7SEq4K1O7VhTBX5K3lGGdRm4rDZ87ySjZn+SISDF/80OCh6OapeCnh
LMfTda8WnRmY+jggWUZpPpwsclIjVl05Ed78Ug99MO+c6e+flOu8gnEYf+HJV1jBmK7WUBelvsR3
2wP2o5lPN3ux9DZgXjIBLFRXhnsDpgQAabgvjwM60jdK7bgtrBovvtuRP3eAMjhOfEmbF+SdtGr5
miIBGWUbq9SOsQo+bTKppESb3X73ROYoXbTOYuzHK0uKTrcPG584LtCVfNlKrAhGbbYk8Gkb13pS
whxkFWpb4Z0kINgHCcUc3yK5DcIudkIM072BVFtzSbt1QXpCjIgkSmY94PODqbMwSaIhmM6j4+nW
yKCwWsR8KMw47XOg++c+tkjB38UlP5NkGdJXOp3QG64xbkdsJyALBjHeqlPwElvIVPxlbXa0yObO
5EVPPH26cPCv3UOEwsav8HhwJknW5TK+KNHOpOVf5JLRiwSvXDe/8RWoWfXYPRE0Z3M4FyNIXmTS
ejh+s5gO41f/Iv4uO8nAKW1bGRXLAuIFcLHmZDbcfhZWMZHLryWpTfwwagUeO0sVzOHPeYOlZZAZ
XAPZ9rCM8L6u21MkXeew7ZYr4ImzFxmap81JlC0Dq4adHb6bY2ol6qSCThUW1hMd5o6xjP4ZmDA2
iSItUj49oYSQirqbtdtVd+SvooUTHBcL8JtuK32xYz9VKS4lRikB9/elX6vJGLpF1IhtugWES7Tc
+l8thXggadzI7O1nBpyZZ6MebiKbP0tfqmisd/dJF7Vj4myHooR6GGxBPJnl95XWWMl9Mwo54XO+
kP3kbzRwNKBOiytHN3vJ+7GnzCtBb/QeY/TNZB0YJXp7D3frqK55vc5BWg6JZ67uBOAvF3+5tfsy
/L1M3yUTVRaRUmIArFiMeqbmbt1c2HRO1DpKZY/D7vuskzhFEkLa7awpqvLaaNOzyiCY2Koq0IMW
wiw2tcDE/OOS9da6oJV+ylYrtXeYpH1Ol7nZs3zoeHExALDfzxmZ6A42vjaMHpYRojXkwTwutVzI
cO1MqLhiuQTFiMbGW/1w7rjSNGpo3j5x7T5kbBLcJII2oLpogc9qht6mXn895qKnqcDOK5aFh3YJ
BpgaSUfDpAZL4OKvkEUP9ns4bImUtHX0+pGMw7INk+tLgxok8PzLbHmUUcF6OGV5jWmxXUqc7MG0
KPq09bdF0tseL6oYISdBHP8QJCh8gf7LpCQ/UHhxT0vZ5XlKPxbHUDuSNohLRKbUaYiaewgFE8Qn
ooNQaRICL/OKsGL8ZedgLhClKu/k7ddsdmV8O2qOrsyRx36tZPXI7YDobK1OtzqjIbEeuHy825ho
xyW/q3gUePYeAcpFSEBmeiIe+O1IqLUOy6j9tOl0hno8Zi99qk8oF0YOsUkzu4BxkIKoOa5nu+VB
JdsF5XvIScJBn3nrEhHZL3eVVfcX/5yz6+jjRuLaQl+9jjxnevL+BiHGBMjKjbgXgQDeGKzEuM9o
8Z9wjDZ5FVU9IGSh5VATDUcC7U5MmU3D2EsF+Dw19yfXwqHYNrM010UcyAuYoNpmPElT+HHVN5oy
beNtjSgEvhkaQQ2Mu2THaoog25C7HzjFm78uQHkAM+foq+gcIXbqaQd409Up8HzJstNAjHH6G9RW
tnjYTn5yCS37XlHN72CnJCQhjvBrKUrAKpmbu3BI11aF16Qw1sNVUwbAul/vCZZYr6LVk/uL5BU9
Mc110s7KMhDTSZdMLYhmE46aR9ghzbUMEaZHqXes7IkK1Ag26Wn2nJ2hOHJ2PCbNFEoBYlixzC7Q
yZCuzjkTYTSte1ZRZPhXYf6EIB8kZpFaIEenvZeEr9/L1Kku4GI+CrJuqRHIUHHc980V+vkSmSqY
VZbjYtRwwmwSqM/bXGgI5iXraj5Pw+7j38ztI8EZw4xUgJhKzW8BVK7vMud3Rs+fR8FpxoSRACHG
UyFm6en691zMhJqgQH3Xst+TsPeu/ej3rOFXDSInbO0il2e5ZhXWseWEsvJgscCRt0DBv502rk06
+1ymkNuRMVo140eBYiN2T9gFJxyzQxNkGOmNxJpl6FSXr8fJz79UFUgnRQu13H6W1C/bBBapfSbR
wK08/ZXtEnYLaeIXqDrLEEQ3j0NsPrP5gSaV/qiyMeAVkd2WhGcFGdwEF+DIUeG9pHWLPJdzqtc0
9mZNPyZnSx0C8fMjGXgj3AAXU3E8dOfLFavtgr+194MQuC/ZZ0VnZmZa58mi+7qHDuA/1YPEZ+QW
AdtytCfw4N+/WVgeq8dG0jAmSLQ9zHssTC2Br5tkOk0zjKCp/VXh52fTuPzeKScqk4NEuUZI/j6x
h3ieWjnMSQwQyqpaYOduQ1+8s0ufpVezx7PTx5+qsCReXfQPvIELBNO+q7s3N00l1l2fxDAQ3kFx
r14rkxqF2EAV3g0LUMXI8+395oV53IOTOtH2r7uXaD43mjG681k8gjZbkVO3E/ORoOx4mY9RLKkE
irUP36HuciYL8bh7uN6LX1VZBwEHloxmVPe6+bfusN38xe13fscK3h8e7SE19+3+KL3Q4iY2ObsF
AtjgzOd1ToMjOCXgMphcz+PTnmWsY48j3XVT4Z+8OW2ekeT1z4epxt9km70+witGPUeYsx53w57e
i30rFEfzN1+Y7U50V9h4Oedeoyg4ZgCQQkjByFLF4JTVmQRik3VRmklkX9NYWXLmxTsKm63Un3e2
+e4dMZWGfsiumX/NhkSa9n6os9O9Sr5Ft+n8+zj9qFThPsYTNTeUsnfFahX95Gacghja8of7dbnq
zXRrKE91gZfoWVaDZb8hai7wVlIODzw4qy0+7/2N1w0t57wDtUENQM2VdGItV90A356maOx3D39D
ZeLdNsGAk4JA8MMAQ9tTkYZ9lfohX/UHSYAayDcfQxt1RDvX+ErI4AWCu01fnv9qs21ANtX7edIK
sHB2zBDUOGqK2WoMK4pTMil+RPRmaizlUAo4ajeQ0x/TMf+O04Mb9MARibcpPowXKiWAaG3qQKbK
9RJzHgMKxsKTcWHPXVtOW2ULnLRLLi+QgIAlVS7g/NVHmyBPlVoT8JphptgmUm5oBBHlGbDY1CcF
JgrrFtNsxb6I3BevrVyH8axEZMTJAh2iXYwbhC6I1wTKA/YOZzSMfQqlHUGxEIu5nEOW1AtREaHh
yXWHjVdt/kUl1AvMW0/paxAimrkZSAeFJF+m+WG3KNhwxjCpkGsGKNdQy1VDtqplcGYKF8MAycHn
yz/6AufgoQ3LyIWH63fwVA3A24Ls1Hw0rfdVOy2DulczJ41QHny0vG2xEhEQKpu1xRk07uIpfkc6
7Jn15SYloVfP82o9K6woEjO+kqouFkymFdLbx6fEvvdp/yzL/hOUOezU4jS1bv8LCTM/S2feOsVb
BjHMYNYTVlB/y12MgIMCkZbYw8Dfg0KFQ6eo7KhrvDesm8U7l72BmU0y503iZg7N8uy5nI45Qp4K
RTrk8gNTjnGv+oYrIc/QcQLyhWlfatZ761i14Ka7k6BEaKS3xhRDXT+NqoASS5JS1xrTzG7XtlPQ
X5pvSTREQn72HsjIJhDc0cCwrXQoArxNzGxBAkXBTraBYK3ZGd5eujgJ5ocznnMyUD+Q3j6uq6nd
eoc4ysRr6roFCz+SucLSIQl5v+p0TK0biAbXHE2atcShJRh2HLFgmq1sSczAf9hkBLAjhysjxzch
BIXA+cu0TyUBB0vZHP5P4k5yO7ejO8ymQHaCRkv2TKGJ8k81epyyfENuHTBeG4B878HmVQYUkg12
oLq0hP6Ju3nyHg7RQvVDrEz04Avyqmk2hB+684jAMwAX+zdl0XUjmD09+tFCgoA26bAa9Z27/naj
9eGvqGgfqRuYpxQd/JUlORHP70WVqkCDjmSeUezoQiPvhJW6x8+uTZ5KrcDGIFzm70nmLp/GgRSu
tmrYUSJ+D2BxjIFlBGyRgIk/2ShuQhPNa4QLJXeV48mfWS8wqviNxGLhl76B92DL9ZrpXvEWYG5d
u5kdtshOxvSatrU7UXeDfxVbXSdGmTepubRA2sgi423R/enGdm4bz+wOwhGvbzzEz82TEdfktGK9
NXRdPwKWsOlyXgm9Qzm05fsCzZEVQvkCYVr0tO2dVYBqmCJv/kgaqS4KqQLACxLTJPk7carhU7W/
bivA6S1CJ/IVEjrD/hcXw7CwfP1LeUozFGKvoKvDc96BhJ6vPiTtOvmCvR2Z7AKSSNxQ9KVfJmvF
2Mw6g1OIZa72rM3fV4uxf6n+AJEMGU5InaEmJsDbchnjQQKMdu3hv4OPPXZZLGnQQrzPo/QNZZ/T
DNxJT6MYsISPZNt1KAeZUQmESUKSeQHeha+6YlIjL2/yhQq2eIHKM/UfrSGTsBejunRGExuv+ZSk
1mv88ezfPTiVafbPf4PIbGM9enbQzGGkXA1xcsHbAUiM4xkj02LxoX41bHgXZoNBfMvVQroMfuU7
tE22YKuFkEtxyGBbHlvAPsu0MrscSoojw8r+hhGtrph00hxAFVpdiWU/vZ1/vPJt5YntjnZY3/43
8EvAWWAMSZkIppohuEsVllWCrkCDaJM1ie0+SiAxYDwE81VZzoM4v4OaPhPAdR32Szw2HRkBwWeC
xl4tsXndjiO8iSUAWFg4ZbPNASvZBm+uts8yBrfloMjFeQvAW078mMwi0Mh73MwVwXph8gD8YiIi
6pdhEzCVAcDlk4Locio3JbKbNGy0Eo9ThT90yi5H+ZzW81k4CXmg3SqAGdUAHd1TstKUgzrDjJBm
IcuEuxKFKozmZb80Z6gpQAiWeU3MaWeXVYRYO/6yJLityFSIGOA4FZVbpPe2FBLJ5vmlCyFjxwEY
Llu4VlPqcCzSt4u6mSNULh8gi25HXmkXI7RaqcY/XkF/IKlYWhNgpTGVk0z4EKGV+ZEIdtUUfIl+
rsr06U1QoGRYzCJUYp5Kv0dpK9B/Gf0Mb0G9+aADlPsLf8hzeIBI6eZRi276ySHeMyAwNgBGIzUR
SfsXcBGLrOl4NlW7EnkdQXvzqqCPkIE9bCqlsMe23cazecIFlZCjWhYLyz79yE+pGYDesfH1899n
lbO9VfpGoCU4Z8fxWwrpKNlKA26pf7zdVWskyCR1osFVoSZk5PvTh0QHq/HtwCCe1HUYSwM6R9GW
D/zvi03lqAbXQBxNo2d8tgiqHWzPs1qDow+se8aN+nrvZHkexaIWmpFNjEyzc0AL8QlC6O13TmNN
cOlku8iSiFXR2a9zeTR5SK3cXxHTo8XdcR/u3yYcoRtro9r6APvA2NVFp+moHssugMQsfvbCNrYI
BSBCzWnD5w0KZwZkt9zl5gH4UB+MuANz73i6GAtnidKfwrvEbMfyuIeQrfUPIQ/OW3stgSSRRZnW
ivWY1sCtC4HIpQvI3qPwfJXuRMK8mG/o+Cc8RIGyF3rn2TCMcn8Rgj41xULc7OHnxjolq7EILRWk
Rv6a+Qz12/HmzWsphiiyho0a0xwbyx8finJAdSGAod6HZZELlDCqvwhwiVNA7dOqmzPsVWE/b0/8
pmyQUxmlW9p1txiIA/mmBnDAlocwqQliGNmUPOOkYjA5UwczWjnlQQ4HRgPg+nCOJU7NX+B8uIqD
XPS6r6iiJUwhVpihqPK1v5WdDcuXo1zWTtI40gSBu3XfRZINpTs1a//kH0NKlC3Csu4KQb7rSmwf
oevjySA7Gy1jQXSVTuCSzkTrQSLfYnwRebuvddwhoNDM5lewFkJtO6fHkuqO6IZxvpMHnpsjDaOm
0iTkgReBoA9yMlzB11E9UsPzPkqLU38tNYmX57a5R1/1h2dbFoRgZsBRi53SPSewEc/NnXK8mz/F
9cp9d5qPx87XJgsKPuNOvUvaMQIiShYJE4yI6TPoaLeyrLkOgVLQ2YA6ze5cnqYrrDQ9+x8Jxrv3
Q5a4kfnjC3Y177Cmw8LqWMDo4lCQfW2phFq1mXg491EGNS6vkVGCLbcRIWuQL9qoDOTHUMyhK6nC
cQP8mVvB7bJYsGTuBIGELpsQroe5yQ7McolM4uF/jyY80YjbN9CARXcwlu+luCQbWRiMArMUMOI+
RuTxqiD/qH8FF73KsH0DoviUj/fynXC8yNKqMFyM+OMhvlg0LRo50RTXXFonmgMkIdBCUIkC2cVc
DyPx40xQw9QHS2Qs9JJa+BKzmOfucV343MoBLdgUCaVHvMk1KDPlhQLXWdVDcSdlPq91b99g3dZz
39W31RAGOuOHgSglqopw7uTK+4lEAOEidhIcfa+Wfs6L8LlCVKkFn4BnDXHtWhDX6VTe+MkGWlMr
sqfjkua2Mnc6qHQEDa7V3Pvyi08jCzKquVj0hHhsMVtp83YTIZAr0+aU8KLjHs/9S/mXrwlNJiqY
66wURfrjVfnHWPZSknX/EmIP7UCNA2+27rivvvoo6Tjds7/uFnjR4jLiX4RG9dSlxc0zFIDUUPFS
dlcbRI8ckqS7zgA56gHpTSjg5gzk5bCm/g6VwPAX8eBjFSpTA0IfPA0BEGhqWE+naXyZ3OnIA4IR
rnmNQ8rOi+OUjAdPrebOBJlv3+hhYF5EqjJ34BHNl42yfY5+Nt9sE/qlLMS2aCcEQNWHRZYYOHAA
FGCMHYKEM2R0Bsyu7cP5kZvXknI5ti4ALUCKN9GopZ86H7ddrDlvE0ODAdp8smzqb02mDFFsx2uS
bIsKn0wiNtljn+atXLmUCg417bpljawGbYBj1O5kpTMcogAPzlBegoPDSeJU5KER7yiRCGCuT66L
0V2G51YDit5MZ0WxCnHP1LwMwgVU8cW5o2ckgPyBDzhtzuGARgX0d1BRubfoUvp3PjbWY2qZAqDp
LkP32hOxeWwZz+FhMpl3KwDH8P61fxfVpbuH0azAd1Lam3532Cu0nIksFYbvkS0sE1f2k39GyB3M
ZXyWwmXRUxRQWsfxLBlbyo4DZLk2cO+dQoTlh5HdnvKpOlWCpMejigCAnz1+lVAkqTGAqzTpO+1V
8awZF8r+XPGHMcYz/icnmnX4hlOW4TPJwuKZaiKjawYPPW/IpqVxc/xUQb3u3znYHRlNPMwthA1e
WpWbxDVx9CSQndv5zl8gMEHhika2PeaEouvNlgXAmzl/w3hk4+CfCAAy+JdUfrxhBaLPm1bX203F
hMNOtf1rpHBq/iMjV2RpKF7cGHi6tpOrfUdORjPZ6ezkiHQX2Rc+0VGFWE+A9CKVesI2ik33r7Sk
az0kiIDSw8ioyj8sOlgnMQRj82PicH1yDjjIcjmcolqK2xwgAUQ90bPjOkd+B1AWM32nRSE+1grT
9jbOKHYbEyD3dOwvVtOhvzchU3AoRamd/2n8qXHrk/IUg/kxzmFMWmaEYhNYOkX6TBiBAOyk6Izl
c4IeqChlaGLofewmY2j6NziOwmh4qk9EtuxFnsyP6vnBWMaO987sB1C0mBzinNpB4AoSFrZUvZdn
Y7mzoOpoz54vmuPebyb8RD+Z30uy1HGZ4yfiJoFYOAHFCD/BhmK8b144xeAezz6V9mC/ApKTVw1O
pVsEAapUYnBrXDAWt50E+Rd9Y6wPFnx/vP7HDa8cKWVrNYPuysN/7xyq1GhBUxZZeysHxHHVyI6i
EY1ci0+c1y6IPSI7aPSotuE1tlaAXXvO8DKxf02ebrT80Y525+Ca+DBaoiJWg/b7i4HRKyzm8Wx0
7DeCjlzUfyWYalEPWO9KvNQfFnU9EH44V105Y+Vogm9jn6RSSy/oG77OQfOUhoqxgYn1PkimoNSG
DMGftNvwlOfBWeB8jkM/Jidb0pUf+jP8MDprlnx0rs6+BSyGxH+H0teEAzP1snJqyHZvEVqVx98J
O7BrTaRPV/AUryT9elKh9z/GR1DV9eGoo0J80xun508Yz1ekdGAHJY0Fnherl1a1WXmJNhCkl3bH
GWbIuWu7jk+Q62rRJ/s1h/1EWW7Q6gRckEo/k5o3dgC8v6oojgqsR0eS/FrsgOnQZ0fejnmO6KLf
RdUtFeZNuxFlD8hLddyS7nMw5p7Pk2289o9C8S4y9K9A2KqdG7BRhs6eivvUkpIe8t+wdpaeKy/U
rkCRGXrct33/15mGiwDuZRRIrM3/uvcP3PsdVtvQ2jKBw5TaRdlAEG18mCdshlLOAXtLG427tsEa
KmFsyazViGmBz8gZ2xxYofUJKD5uh/S3AR4cOEDH96/ye152u65GnmsQ5NPxx6S3TnnPNjdWbQb8
qzjRx14jlbQQrYgJPXIVISCvuVC50A+x2GwKKMJpoGrv4DTfi45vOVlHDt73KXIriESmSrIVxwf2
G56VYPamazm6rNIY2wUvCAs+IimPbRFJdwqgjs65boz9KrpbAjhV6Y3xc6y9vS1QOkFvDKYWKAi6
ZsqdocAGqCGxQFYBTzE92TWg0JaVwuwPjIlRy85UFRzKxD4oHSxE2HV1zbQab1U1PFMWyhfTt/Y0
iR9jfJHDMjFVWhX4I0eTqK9imGUXn9Q6oBc4oQv57Rsz+AgL/326e6tZLb0/a2FCM55S7yA+RvSl
AoYQiSAnJAC5s4bvOT/iCoeS0EylHRfeWBnvy77/hOZptdyUMe8d24tTlvIo2LFizAkWa6vcpsA4
H5CPkF+hqJF7vdblCC+NT8qD1ez1BXbBsC6NMBVAGttqPQnk8RjlnmK9Z0vj0DFcXgui6M6kXa2n
dKcmpvMC7o8NfImW/0nnr6p8tInTvW76lODquq56+x0ZPVdoCWhj/nQdQf0hx+3OHLz+UwNXPR7S
6Mi5e3e6ZQ7FBokpXpqCOVCyK/46HxPSRWENtkCocSM43+ptHCbaiHoWm+01ZIdwzTzBceeI+51U
KHdueGqWNEuYZzs5mNlnivzI7EZKer7WJOlUftbPEw24FzR0Lb+3nhnrdNY+9ya4pw42qa+WA1xe
TPCy1APJyBAkwyvuPRvp+aOzR9Xwk0OuQMx8TjsgFyDk2J/6hXMnakEAu4xOzMJrVoinWaS+6Qzc
/bjGz0YNIpNQJL29ReIQR5sq+VlPN/Fz+NqSqlf5JJVUDTut4qPlTLWpkCxvExgD38rKQZDstNWZ
7P100fBg/sOtrWcfT766u3l6YUMxA50TGLAFquWw+vB9KxeLDInsy/7o3zsw3v1zbcqoMorQG0Em
rYVnjpNNi330PNRiyamK3537/eu7WCEDwxAaSDFdMRo6HUBt2+BKnauGvwxl0/NUCuKaIv/QOvie
6qQX7VY22rvtBlQ9L6wdPWYIuLRfmxhHv23J6F+1soqfIZEuW/7NHMYjOqzLxkV9Txlas+0Kdwea
RQKYAftPouQ/jEgMQJvvUaSh4zYfDXrfbLs8bSD0QaZLDZi7xfwDlKXr8u2KcI1hp83kzolXbg7r
yar96DHR1nDdg4ZV8FjYAW0MZn8ps/yLR8CPuuhbcWwF+xKYwZUX06jfPSAnQVLkkjXUHERPDeeU
l6gnvgSwgcTFhPnCVm1/E9xNJoOEZB186J6Sc0K9r55aO9uDkXiH8jCaJ4d5q41SviMmftjrlds+
Sapn7uqbpG2QdLEN7tqXCRRBv5ZOkr0Zvj4hDFpOgdP+M0nKcWJBBjUJ3QwUobevmZLaX929cqSO
x/gPadxmONtL8C3B3XirvX6ubCclx2Vu1su8lMAjh1YkUYPok3LIZlg7lx5ZnclU9R5gCIN5a0WN
jA7ACThAJ0UYO/ytRt8Ikq+rDLG1gbyYQHcUemvoDEK48EYHVjzpCIpQ9NOV+8MO+1vvh0+pU1fd
3Ldy0eYvT9OqN24iptNhvCi8uTub7Gk2ZrMG7hqWF/uwGjM2BC6sIz/ae84KQb6QvStCI8ECPrhf
i7oIbI7eyUOn1j3QVmq7vBHnqJ4JulIaAdibdGAMRoAy8xCqw73cnazH3G/MFfzzvKMBTdVpFMNw
R/9XZ4C1pdQMW3vV+bjak8Rdyh9dv4xwJjqBcKfvZw1Of+xbhnqP9aNbZfuoT5Kr/jfHxaGBvdQ8
B+V7Zgex8Gc/Q998fpH39rMcEZeIDRJ2egQ4dv+lXJtsxUA2kR+bz81c1UUfT67CB/k6DtW34/eM
XHiX+C1zsnZk/NVPMvdwb2rdQmChZQOIU2fmOnsnJ1bWAxzQ452XGfx2O4lvqVbxEuDpujJ4RKKT
drmYJDLE64d05fXsLaALLKmQtxmrM6xN88ZcWvTyPhjA2B3xVIdoXQpU+XXWKAUJMd+T0JRtXIPR
ZCWDGH/AVR6vVxTkHs5uF+10UdKD4LN6Z1gdSGZ8bgJhtnuxHS0vDHlAkuy+H8H5wquM+oX4cYpg
OmigkZxGRIPdXcNuMbP9/QHK/vaogNu2aI7o0BQOKrKOGVB9dxv54hDY0FHUcSh+Uip6dDxv3wVi
XG0zTGGMNAqYU/fj9J/+d8z3ancIUM8EzDGzlZAdgcjTgOgHNQi77MvCYxzemWJoM74kL30WvRFF
NeUoaBIuxpWMEij0JSTqRKjHcTtPM8YbGrhwm2mEHlHZC9tdEfoZakr9ecZA/SJMTbXF50gWQVTS
k7CR4tt9tpOEH8VK1ILbQQKpwq0Q2Gn4CNvCH1EqKDHTkmp4sQLt9vrf/ygHuiR/327NnbsR7//T
JTCC3Vq48YmGIxxUh8pUJXOW21aFsd+G22S1Rm3PTWAosEx4F1wao86ZkNxoMmfQQw8fl3ttGVOY
6qkTvYDjYv1vR3GrwG3FVJIEZkFaMOlTwZ/uDUnR3JSFycpCxThdnk+XnqXxOpL+Egxo/lhWwEko
a/9lgXEwuerdlZK1H95/TH81KCm5T1lzFkj1G0V0FpMq/+g8vO+kUamUObzIWUdEp3YcIQ3FMEBg
BnpyuD+2w1sdDrwZz0F00Pxw1uUx88USp5Pn4X6K61uDgKxhX3SAf++da9kKq9LacpzCf5Ff//4n
Y+uA9VyHXDM1MlapO7ja0NvL7trgQTtoaeMTbxc93TefcAUv+WxzAoDzXIGxriITqAckeUvux0vk
vRhXLaPrwfXXnZHNp+la5woJzQspPDCL2pN0Z1mPlgaXrU6O7Aweyy96Wm49LEoTgxwyaT2Zr3gn
ORKYYnvsWk70a7q0ZVNfOqWBMANEFMrNkvXS13SfndjwQ8Bb0q5GmtqsesZhv9de6cVWtIQH8lNo
fT5jAFIKniZvk6K+hQiHplNzSBcmhVPfDU3VC/LNZXziNsHbSHWInQq0dYXzIImHZMvsLaTeE3BF
2ovhVXJlkI6HeaUKZ+XvO68MDk6JFXzE3K/NsHUVbFxbMmagTj1ZQOlVLKtcjuKdXfApSLpTCJ7A
9KuPjdD8VNCdliZy6LswMDwi/pMZnMUQdJPwkhfYmH1nWDQPe1cGagjDsbdjp7Iva4y0rqQ1+mBY
zbllkV2hSJ2SVJ0ZQAaI8KGR3s7FPBph08D1pkAVuzMCteqvUfR66ZqzyeNe6E2IRGOeUqWr4CbY
K7YdWvyRmpyQVlxHf7U+Bh01FpXNa8jdJgEd/6bwdK8YjskX41cz5vfma/VAaPf6zQOa9a7VOiPN
zBSVhNRE+/JWkb8P5f/JP8HIXjoa/5e1M+5JZoACrcFz9xBLJ5w+MFcZd50twLFYplTRZRtd0Lba
NRxJ0Xve+Dky6mnMcZADO+3m6xI23qe0d/P/ARVUhoagXn58KbXsJIqg9PbsFxN/ts0e1kr0ofOt
IfyIFOrufFG6Qx0yUDKQCM5cv7qiQnvviP4m58b0NTP2IOvU+qJKG2S3CzIZec0p8MmfAJXnVqAV
5cdGn1QWp8O9PAWw3Gl5qbEkz5tssPxorR0jI1C7MYGBx6JB2jQn58UZOKlznewnqP4ZWXdZT6QT
ILUN/CFsGvfsFFwQ9WT63PMgQfvyDOUWeJwA8CH/mY7JsfpYahQl6uZgeVTeKHHiyLu4wjY6ap6B
YUsl933YFHh1Lq9+zj0QY8F9K6jEezmAGHT6q8CYFtIKiWrHT6VUOh381iTQVtfGPFmGbZWN1tNH
I/n0EvpUqTUQpxa8b/aoWotFyWb1uiZ1x0B2bmXspt//FR+YN1cFqbCRL7HYR91BNGYgji8qDjbz
d1UdGe9IEW3ntZl1CPu9udM5bCvuqk4UlvLHMhmmcXDbCYJKwrTpMy5/3t9mlGK9f9AbsUhvBuQZ
72Ai/vODz2E2Nw90QoyF3RJn4JLsv93G/NWzC+Rh79Ru4dO/ejD/TNYjjVtVBs8mr5Pfl2mAZEx8
odmLSGe/p7B4gekxDCy1QzczQigV/DwPVMHpSWhJXRIIA7yVXzFxL2NQE7QIKePW1Jm6VEaUOzit
CmE0aOMWWuUh0iH7JpdOUfW4fn2xecKbXEkjP2MCb/Hwh0lGlgxr0X0da5m7jDHx+EFQb+B4XziA
3Y/FFFLO0v3iTKDW9fTJcDqoERSoJUkDF9bq8W9CCB//nPAj0ZDaEn8S8h4P0ihPOwUCyNX75F3c
vrg0sdSuM+JltQixbyrmePviqh/60x5NHMVclIzaGmiOlgu3k6o6XRwxutTIxQPOkE0QcvJS+YV0
KvW5hnCO8Kv2zXdS/NWIUmIuAd70avHR6M8tM87JHg8UalOXq2rBJegPuDC0vUgqwzzicHIen6AL
ysXA4uZMXgAmH/ihLt4QydF7M+EHin/7GNb4kCqCCJqhm2+JzsHpKTmTck75YRVu1VV9TWSquZyK
cfCeM5u3+gqbE8E6zlyHRYBq3YM578CuFKv+kGsTr6nh/atcbUd+iK7GlbyrJrti5USef+vu4bzx
UhVK9tOvbZ0uoXneGKPqHHy2ddEa5YXNrasDRIPNTlYj2/Ab9o/P/w2doTQi0+nNq52/VRdeZDGo
ym7C915dKrsUiaPpbk7VlC7nWVYvM895NNwgdtN/9nAXMy4MrV9OlnhQZISRw0szIYiUH3wYGAPV
2mxyvgsGgmUz2YvbsgS/xaahqLTcy6KgwfYUEMoUm1wcbhD016L12mCujVnw8yO5/SSGDdgofPgT
VdB/51RAaB7iWWk9ulnAx4vpaq5orpLiujkrsLpoFYfe/6GPHCPBtrdHqFeIZEwUB152kQUQbNc9
Op1OsgpSPQljXJW1XwESun4mf+N5of+uU0N4Xepumxini0OKSxpgsWKp7gNH1uTlGvihDIhw7yLh
5tH/2CG0jghVYmUlGC+9hHc2+NqFifLS+Dz/XEN7e481arbKEmCIZnzYrarNVF/Nxn4neSFlrj7f
72keRLsn8g1lMShWfg/SEFvd8d2z9mxbRV+SwMP9C2XrrrhmrfVKnv5EqtwK4j3ZK0NN7McLjVDw
Hi0EvhHkLnL5pgfmy7WWWjgqa8HPiSKSE5EZVNdeleiZDEOWEiiaRmPeLKgMy/tLjCgptWxduBL1
O+D3B/HI1MSAHK/8j8EME0GSNfKWB2LHV3ePVz+xGJxoe9V0SvNQStzMZBR1vK0tEtAlddfaYNnK
6GHyE3jJpT43fUGn76a4rmIjmI7JqvHTh4Ezaf6H3vuwfS4DLy3vVrTx8nxIzrTLXPbge3HNBhct
OjyzqR5FBoKMia0bg+roJFy2PI2YLdf2d+JpkeQexBlA9dGcP4VDXCXtgxNWwTbQAPzdUIxxTklR
xstAT1EVeNKAffPmEHsw3tA3FWLXYewDQrrVBeJ9dZi+4lBQ/R8sYZw0czGat9X4DWIo3lHhO3u1
wuId5UMvPO+cGSwvcPajAgAZx+/1nWXgzxjPPMjm6hW4y0jAqIlnJNd+A4kCyi7sOU18+5f4z5Bu
JV3nfSL/kKkmfwcfqu/SjEhnJJAKh08ntbX6abFEAN+ASQfm8f+kfGyBJCzNyVSQgSC25VmmFz4i
D0jKBjynP4NRAcPf6Uudh0ym9dwrIYAjXktCiUHhwjxDwnKgEenyayJY7sdaKFnNtn+s4LWBlAAE
2nYJXG9PoMM4n1rX+3tvFnCj+BMaxiZEPHfxh6Bu76VAMnZbe1GjXFpeyC35BhJc3p9iSbv2dvUf
QuiBczrweKiFZjYJTaC004Teij2td4wGhABVlVqjgCCjg+CEB74OMqw0+rg+cuTWmywLcenYsMkd
GWaFiBXOh7/MBh9LiuvQOCovHu5mx6QE1kfhgiFQgDc6M++AhUZ/7A/qzXCdrUE/V/kCSCSOtzuH
f3kJk270fMCSld0jbBQfUQBhA36LifygHj7OO/A4OJA0GdLUI6EhDmdX56I8sq8dossa1exfxZCD
ykgDqvl26/nkCcQqhhNthmvy/dh+Ih/vumVp1vfWfyooUs/dj+9c+yeK62ocuO+cEhF1zl+dQSxB
Qi3Ce7nj+XP7ZhSMAZi74ekxjzw+yl5hHbUmwwglYSSAZOszCB9tQUlcAWp5bDJSZlGjBvTwiwN8
RMw+B/Lpluzh5CBJTdzlRmA9sW+I9x2q8RKqx1RSKA4cGCTtKkyPsjcfyt9cvSnPC8ye2m21rQeZ
bA7hdjYXcNf51PDg9+UQ+YznskeBhGq7AEzR09bbmolyOtTzqF8ZTiMfLmEp5/LcmHyaZpJIMH/M
JZelNtoSW1v85ym/gczGOfMhONfZyKhyjhOR/eBLizgVxqzUBySF1aSrwart9F4QOw4ZBF79DnHx
HyjTw1ZW1Rl/rwDFDuPuxi74tw+FjJLfxre1Ia85xmjejHwXY3sPGsGjwJrom3DUL5qO2MB0Jxgg
IzAE08S9YVgbYC+LkXMO3ocUWEFKpqEkyIGjVnBAIWBt6MAmcpQ9YRqDz2aTqkE8olHhe3LlBvxK
cNw5Vo1F+KxGujDiQ5PZs4zOPPaqApQlHtHiA8dp/3NQGWo2G+kGfOupaw/T/SMXRnJTPyRolcBA
Q/n8oZeoQ9+8yPLJ5XBhAZw/0It5O3I+rb8te8qYRwZyV6N0jARQ6iooC3V3ZK1GMKkhA6Uxw4V5
+KA9K0b8xmbzPTiJlJnmUO55I+OFOPmG+IJrocgBWf8m0ip6dUNM5UxUJUr/x34GtDzjRxiqnvRl
U6+E1pqDdGW4yYafddYAoIhmkJCqeoqP5+YIxvoXXZtjqo9vr4I9vkxj+sfYs/x25Z5QzwwpLAsh
fC8CjRS/6/XvEY7kqhw3RysvfKqB9uCPNogZiwYpovjq2MKgGVbJN2SkgLFNXaN0nuNGiuKI0+qK
Cnf3RISHkFQL31DLFzszBgZ6dMJnm14AHV553vz7Yf9sRsYHkS+pYbxkJ6HStbTtjgy/enab2fW2
2Zag/YWZWH1XZJnTjTC/8e6BFA4SaT2HHhPrAQAA0ZWIvbC0zHLDd+KUO95VDDt2TvHZMoirFh9V
YGptzUCbDKVFqHrxWx0GNwa/HAlp5VIr2RwlDNRQvthtLzlAZUphbcJLVePtnuz2qvoqdGbB7v3A
ihkvT+CDR28pz7mMrPH21zm0bW/xUVOTvd0HBiHeMYQzIu5ho55erZG9GdeYoUdc62bBcPyIh6Zw
8CJQhG4e/1RQbEsU8GcSFZ4HJ0V2UDTlr0quaHg4M3OGmUENYoXXi9KuTtW1jaLE0YpEcJ5JDEjW
4alDSvgPV4D8h50PRD9zjZeYhDFWKZ8wDXPOGPSVdvp1MOr1CRK9gn+kZ/8ubeWcGH/picXCktTu
RAGpKUUvB8jFD4fukElWB4yuQ4MkfY2YQHW4pTvyNaWkyqsIi/jkkeFJl60TS/OsSXSg096BXNzC
rZBkIHClby1CFvufw76XsOCP2i6fcQJXu9m56WKREuHUvI7f6Q7Il4RuaQ5wW93EsZwB2ss9mr/K
dzOYbWO96QxTa7aXaklgZ9TIVIzuSgBNNxBHJfIAPxIhVv3bsJEn+M2aDWlV/gFSzKP2fzits3J4
/fA93ZG+Y5VAwfrGZwLsRz/1xDtbErBAVLOxdeLGEn0o0hxrL6pnJ9Q6zcqkQG3O8WHcjLuv+n3N
3KGmNAayKEvJUyMYI81wUIS4TPqSN8VwexeiuTSveX9SEXgNgK9yR8CgWBKl3T1OMz80KPzcTlU4
0CjfcyS+UmUah5sUGMeyOVhOKwu8CJXQdTnJ2D9LHFB4DFt+zyc5xBd32LRWiqTlLakArB3WcdJZ
F7plqq9wpQ+Bt1GRjjxAcyysLCM/CBrPu6D2bEdyRtwxt0dJ/Gq4rvPgI43tkJ9MD9dLih+TKLd9
iIgtausKy+S2BYIBFdqaKh/YiWy/kOeXZMOM1k+JYE2XCxQSlAgpx4zFTY+65vXRUtdrc3bAd21T
28Ol3SRlPy5kxtf+RUNbNYM2OujnFRNm0bAVrqnrtHZLCKJTuUUf7jm5qAylTUytRrP+IrTFvwD4
YZ4YcyrehvdKKxefA8pTkXLgdllaBUbRE3VGv5zSGlbPUpSzN5n1yxLG28WHsx+T04vJim8jlelW
vauxbz1jAJI4LRpbi/AaVECfFtejkm7KJHHT4QWwsbIwSAuXJ+6jpTuZ0dgfZ/PGGo+U5bJJ8Oll
lMDfUzngRlv74Vdi5QaE8jJ/ww8a8rkvua4Au2aX+SlCVYo6YY02rTJiVAtlQzzxvXvs6r46OXZ+
jpczqEFynd1avYJvdtsn+eYjSwfZ2NWG4HVujihWc/DBdeOyUN4eqGrAW5KVvczQSPJ7sppx7OD1
GP1Q1HE7mECGENbwy/u+8x+EhpwE56n7fzNX2ENCaxvzsQX89UenPOtwq7i4TGiRTIYEUICvV+1c
TewStVt7aehI4HJN2SNI7PMl0K13q/4tOMaa6toTgDQbf/nVDmLVSbMPkcKCGLaTw/p6YjjDfQ0l
33lSGEnCbDZ580EO3iTzKGnsiKN+tTuRnr0795SucWH9x/dpuZQpa0e6UBfBRpk1v7d0lVdatdI7
U4AG32dDwSDVazY3pjvWGHRg3BD6ypmKFRq0WRdB6Vg1WH4Eqd2yybwOLgg0v2zvgMewJuwh+X4+
RjT9tqFLK9v1k/L9Mci+PfF4pXGdiu7iL2vcjVO6Srv8/tH0Q9V9FAE0fQWVXWK63NhLMUZZnR4D
PVQiEfQzzoIsasMbxtQVeNfVXFvyR6mPkypxTnldX9BoYTEVu79qdnJ/Zw7h33Z7zftjWJun/F8K
VpllM1dQDPJU78gPLoEjKJL/nJnducoL6G0C+E8INFwb3HlReAbDzZP0mjvSrJ+smZuwoZVAYWof
3dIEAu0aajeieJGrcPQxGafo0OCI34Aa4fA15vyMJe5uCLSPxqmic8pef46RFgar41lK4FEsJa8H
ai1lBj8yG2HBfh5yT7ZIRKeXRoKigP/Urr4MCZxkbsXcLafhtP7OCZWgDCOZSlo/szLdbrX3zJcB
VGbI+sBe7wcV//5sBV1uwYaSxltohrTyuuvDtHkRjyNJFuNuJZLboGA071n+H54Mr/gpLNPC7tVg
SANl4X6BsdTnojb/qJF++z4On9aHWz2rMHGwD5qKZ9XD+VteAaP0XmWPnAroOw7yrc7zlbjhTpXT
b3RMUu2agY/Q5kmmE3K7O5AWbdDP1orqPdYcS69JCrt5xhj3/CvkdfgVqgegcRvrcWjl2SGVPC4+
wxx2uLPJGgehuqYZdeLIyDgkuOFv+pH/HnpUmCQ90p+RwFBQM+KJm4nw+ILdnY6zXONQS++JH7nX
ih+eE757bqRmqQztB43Gg88/P5EfEwiJ6q9PiogxgTzFYLNWt//DZrqSxGNPXXZtuJXEZpn7JyMg
nzDixPpT1txRtnFqMx8LGUkZbh2l91jmA4/DQ4pQ2gMIHFWdEeTbHl9GLNGwjljOU9OoHXfhZv9B
t9ChIZdovsUeU4MLCYX9vx05zHyfZWGs1l1mrYfWbkVZ1V7Xn3Nn83GgCpDSEoiZ4Pg2TGkNqfI+
NqJAWXK1MzA8GQ1SNW8U86oegBKn2GmF7Q9YwdbwjHyQ5z/d5MJhtbzFU46Vmh5pbZ6Ilw5eT2fk
x+8hqFtSB6gN3lSl3Bvii7firUPjL/aV8eq7mYosgmXmxa5N+om7u9w0+VrajxrYxhfllS9QZjLS
iy3s1WIMRENrhQzMOufutr35wKPqdFEaYI91Bo3tcGP+zsXE3P85mwSmrDm8PldFlxg99ivWQLWT
9qqu1Ghjyvyd1kfV44dsOAUara306kVHuxrmmXqEjxfDa9diN9ujLpqxMPCxYhNw2JnJsoCigIVI
2ad4NW0XbfBRcKu1VGpMqPXVMl4ihIYX+9MHlfD9/vwOYIMpg0rqRRbmOjsPNCy4wud7QpIkBOU5
Qw94LH7paERDTk+qcLYD4uQrdyKnHFehOA7zZffmkI/qxMMLlHy6joqu2w6ZkOoMJJ6X1rPLT9fO
SCkB/SZpH+15AG259PldkHr+ESa8qozEQRZhQSyMARxZkQ6TpvRps4KhuaXJqAS7tD4eBQmhnI2l
eytsgbZZeBekhimvDFAyMNxBbcStfCZNVRwNrJmAAQOtZwEHqYwh4WcFBvcndEkCuoEMlPHG1UvK
3hwe1xrEzaIzXBr2sjozHLgIc+473ucNWc5/bztyEGOxb7jDH0009fgkXfPn7uwCAARiEUhKKgz4
cDi9UzkhsVU/zmBxL02ysWfqV8BSGronxWlyLNIrlPTS7VtlDZ4nTqgvnng29XCQ2MrjAxC+suLJ
tt9AcJGmkL5TDt8LZrGbA2OdQFCd/miLj/sQEhKt2H56PxR8gtWou1KItlwFjTKZD2doV1tng4BV
xcrBDaJndKFntOnjcJnBMLa5rYDHT0uhBWiczSEEn3fTHTJBaW8OiLc2368u5/+8/jF5Ib0VO8op
24IoFPVuOai4A97wT7fipprpBEKW7+JBgyKwSZ+rFxlg/l1rxGUAGvQko6SNMMQsSELMaSawBG3f
K8CYgKO5llYKFH/FryZGoZbQkyhb2Dd7LZQxo+Q8X+K+Yv2YIjvbMzNGC+IXkQSCLD/BXlZFvmPd
5D5NAiRbeIw5+mqQ222aZ695/t3BW1RRUn7wj2g7pA+3+lWPNOhxB4RVO/XFQgW8x3WAu+1XU5lZ
7qnhdeLX3ahZ+Zc22ZMdEOp4EUjI2bAK7yV1DDzuMtqeAY95SvZVYftypZRSUsx66v81W9aw8mXj
+l7/WMgEWsPdqbuqXKq0DsbiOr7RugqFLg//sLILQSZRBawNW3Ydm0lsXvOAY+yYjerR9+pl6QwS
OIjLDXGlg0JXvKthFnu3VHHK+mtpIhWGgO+AsUpjRkDTWizLyGRKe/1PxZU+vCJFL1A7dAKmryGb
Z6jFgN/S8haGOqHkZ0z/rvtxE/iW17b1eaBnU7cK2G34V3SqYXl2gCNO2P0+WUCmR7Da5TIBmJOh
2IY3kNHIcH2ZIbcgU4tFIqK/KJ5Ju3YtewewKzbkeds6cUJLA3gQeggF4R1xbPIE+KAzVgLWABEp
iqaupEfNkBqMSUidx7Sh5WDzU6HS7c9cDr6n+6RACZZbiMOSGpCftsRaPuB9TvTYeMJB1GptERmZ
g7l8P1J3i19M3vvZrHZZKWGYEPbh4CtoVx21CbXmvSNONOBqfrMmkTQt1iW6REHmXpNgGd0JVdGD
Vf6LwqdjmTuXuIDIBw2C/EuBjoqQQ3vIhjGnSUTmHSAh2UGb219HnbnbGpV5Bs+k/YsAe95m7bXx
tPouVCLhlIsrEvR9N4aPNL8VrFe2c/P6H3WM0OEKnX9KC7+XASR9i0IJNeTSAu8lu6CTC5Dcw9qp
oV0H9xiJehH9F3rr6o5pTS9VY48cVN8EJrM6UtMs0MXlXhjeXXP0LT/ysE4zm7AIW5ayq1PPsYwL
ddDtZDK2Xrwy1CUeIfW9Yl9Hg1fA1e/DPTUtFiaG446jmauTHsU5yyJ0yJBpmUWKW4wicfN36fx5
XwxgZ02s4hhYHBOgUsdQ6m+Ji+zU0pbqG2izK44BA6a1zFpmQcZgNCvcYdkvPwMllAiRdZrG+Rdl
5QPr+zUxwQgzW85sp0yAdnV3WmpLJKyB56D4TCJ4+c2awlHq5EiRRVQ4lhwGfVtsgwsFPfhLC/6N
kKjKv3+V6ZG5Q9FDarQD7i15qlWDhj+j39nTG2GAj+AdeuXEU30f/mWVoNi0UX9jFCCd993Fhp+b
RyY3Pf+Y3DGLPD8h3ZZj8xjTkrMvJRIdQ0il+SoFhkFJkAL2rGoARU5RyY4DPmFvZUz5C2y5KM/P
03b/MuqG5PO8d9GMc4e2dCw2Ga/rAII5UKiLYEEEp4PRE4NZfsIRH4s6jH7VyFxDHSEJgpE43TQA
b/Io3R/R/3CrR5duwnN44ngSUKRw0HSyQTeO3inV+F+kkCAsy7df6TGuQrvFF/C2ANBBMpsPvM8f
l1lGe2QCWIgrAYhHYpzVZAKYBvJ59wozVNyWG7U7Kr7QeoAgYJIqvueogy16TP229Kregm46afLY
uTtRBMbuilw3ijgp2iYsFzhIXnm6GpbJNZhC/ZR6f+cZI5BVSspLkPOTHHUigbctajuoEyZNq3FV
CXsAT3U7dneU2D22oWvBe6HewBxxfIMpD9NglTPdZqDJMa/xMEnLQWM9h2LphB4txISQKACqCAtC
tMEGo2lh9AaxA5akZDtAgimDL1iD1Rytb+0dm6C0gY1vaqnZxbgYx6/IoJrdN7nYCtvk/IKWLj1T
ZDGcXgaOCxjTOjPoJPx7q0WRV/vrNCTB/CmiTHqTe+PE3QaIDjl6Qq8Cke8io22kFz9OACSvEruS
jOVt8CQuSxafw8stkfifIC43ZKeWchV5MyGPEH/tjTwE/W0wd5YwkcB20RlhcCdM7Bx+xZlip//A
/keOktEGwpKoA72dr4PTYTp0AbFNUhOw82iYsaSN7YM5WYAIkFqWYTZ4u+VQZJ5CkFgK2nJ8irh4
ijqTPnHwM2IJwn5gpEc8ILkfQ7MrIJGcmj95W20KQYqlJuvIKjupUlgRTGAb8vdxm39jc4zFf6tQ
vTeysv23G04m/QxyoXcxBpHFDEhD0CzHgyQ+1jy0Rc2xaIUd8rWT8cpCH1AR2GJp6KBppnp42UA0
8Yui5AJrSayYA22e2DuGJRcvfZdBEE36r3G3lKTZBzg6aL+u7Qw4Hr2biHyoX/RZn7IRPTXFcrKq
mYwPBUmp/l6m6usro6HB2XauWMnWWjoQabBFA3Nx1Q6uKXkANtbwNS9kswHPUzsyCv615PzoG1zp
tZcQzQkkIyXo5ex4+/14R6VXgzbuUTi3vA8OWnVExRF5N63fE2ynM22Ny1cCgAMAhvk0irqnQS4l
tp1+FDtAWXXzYBZO3zrg2Id7CgIfXgNJZJ6/gZ5zwrrOLC3WxEqT1B7jXBTEivGikrmql7Ewu7+o
D02/2v3yR+sKb3MvY0q8sS9K8JmTJtJb4Hd/wnjtWSIN0ps4q+2eEh4g+htmBV7DNCDrPmv78CE/
JtHc/dPIWvRlT3/hz9EjDt/0MlZaaUgqp2nhVabgJEhSuKVYLu+6iDkbXENNQD2ECukCRvEHRUEh
d8Ickh7gyVKF5PAVAgSb+0z24CWMKJ/oRFM1wt7EsPCnwteZ3/6aNr/sdDjr5LHKg/lQKqWb1lX3
zJ0gAmC2q0eoKufN0f7TChLkQtBqk2wJroZUBzqwzbzF/Y8qruR2+2PTcIeehFbZ3T5xUHaALXbA
t6pNkhmHyssDlh4zFjH78Hcx9Zm+vxs9hL+cXT3zZqSXxlWLljOyRe0XgXRhfUjYcStLzZOo5RB+
MULZlS/EFkiIppRp2N5txOLSpFQ0eXEk/GVIYV2j2MTaZNhh3TfyJA7VCHbKR7fd839KlCnEu2GC
l5Rztk3r9hG+42Jarb41XajoG1ONIuOKuf5jNHABvamKJwOU951EUH0+XkJX/+RRaQbej573DCOs
cJCEA57QgcMjEGmCRooR+GUc9MASvH6n8LjNF+4l3XU8UNfX0HK4Y8W2sDjDuAG8oUs4/seTl7ab
7YTpxWiKku4PyXtG2hTYdRsabCj9sctk2dCdN/XEj621Lkh4USdx+zBXSKqv4CRDHu+0sUnl7AYW
8C1jQtfzhNR9deGKQvK3A6vENRhftzVQ5OzstFqG/q89xKQ2at/ZVAfzY8ZDZsTpUdMHVyNl0nrr
YWi5DMp0/ZwtGkMsyALpFD8irpd8xWGJFl0W9jotrX1zB1jZx+4y1srw+PsQCt8BdzS2JLiLVGo4
o20OQ4DCLPgnWX5wYtg+bfBrZstkppZNJRvSpO4XaphYmggQPe/fe+JfR8Jp4GwOOmfYbMe7jC+U
L4f3PlBqVDDoq0lKnaeap6so+GQ8wQ8gjpo57gA1+patH0kyPqjuTVBPmvw8kSUOZWxH5WjSY/Oy
9+sRmTOycCIadlwh3x5gzvWLSi49J39r/svTG0f61hEbswL+JlQxv5/YNvjryRBKgNYcugcw61za
q+pm55xi37PQ9SxZsfsGR968tke7miHWVtc/JLG3DAjWlivxGrNprLt5q6PEPUO3kAjQn+tFL2Wf
HnQYYLLuUo+dX6dLZi3QC+FSDUQiSGOBjX1u77d290A6BXPpWtwBlPph7VkpB+nKsKHVIhsVyAZu
xtFWExHLWiXjutVOcGAQdKoWE0CEcOHKxy551+c2ixE90O4lg1uM+f9oAS20rergqmpzXUyx6a/j
ntir5ysarZ/U1wnM5hOWza+2+yUEGsSJFupDlue9j1XSb0BuCQv3klJia895gTfPfYp6a3B1uzM0
/ujjWzAawp52dKxkhpXbFwAv/eCTecq2ztlVUfD3bUqYSyDpmg7HduLsyd82H0v5RxxkVQxCAw6R
Z20iNpHUkRLVAfXY2Z8Z3/rcw9vaB6AQ93Ka6EZr9yknOqworEx7qgb5UH6A5mvXe79ix7AcpgH6
S29eplXXEFISYKSrXoFG3ny5egz4BdlRMrCdNGIXOLVs2gAHppNZnf48DuPYLq04cfG9QwBTc7Kw
YCohWa+tdUVwEYflgdvk3nRR6lSaB9MNBYIKbtmx8WOCkozkJkDtkXKg+yN9kBzf5S5bAKbBieAZ
4gE92B1mauDvl1qqnRZBnf2y6gNnFihw/Yz6MNiLF3+uJ4G/DwluGIKw7Z5D627QsVrmwLQUKPzn
BZF7e/pB6eagnZCG6ksyGQawiYhjSNYGsbQnmCmY3TvZRbxGVXC3/bJ01d8ujeVw6Bhy4Nz/5eRs
poNbM0W4TAk1MTJJn/gwZG+FKdcvKlgohEaPwGc1SmTVmc25gHY9kDnXfAmebZJ+R68EbvS7jir3
ukt6/jq+PXwts3JLjvaC9yxUhw4kwdyP+Z0X9/VZYs+7AIrMsWLR7qpdRiMsCRkvvdT24GsNlrPW
1X6uXbz/JkcTyicB6fRZKyJcs+3Azbzg7ox1dosM2juOH1lQueCNerZU0dLfdNvOQK1gzG4SX2k9
d8zmIcLlgfnMGVfFwK975b5MI5jG+8toOQh6DgtQnrAs5UBHLeQUGFc1rugz6+DOkKGuPrUYW0AH
n22RtwTBGZrDQZlDx5j7M26k/izu8iRXohec7FYaCVzoagWEQgV1hxEoIUEDkHly3xp/1fuylzbc
za4VhVfUISEuE8pnqyzaf0NZsedoHUr9kz5slOckgyKVz4gzGuy1yxGoC1KkvE+KY1sKh2bhj3K7
yaOSlVhzCNSDZ9AeTDarWUM+cib6KCwBAP8oIBbig0AN9gVPufRkQ4H+qyahnzqx1WUQhuwwovE+
ngg0HFIQCscdPNEtc/+DXFoUJAhcHDDXUbsV6oRmw7dFYtDSOqA0eGP9JaPkT01joxM81Sxf7bBA
ZH+TqmJhpKvIqjONvJo4/Sn8oM0kaCVMZlZBDjwaBdHzswxheGVe0gHz8gwIrqESHHKVMm32tWk1
B+198QORsQtuRQBnlUM36m/YUaK5wphBDRau6ctvgZEiQNLFPvx2R9bImNIF4SDGnL071Yc/O5Se
g4re03GamegOPuQjUxdgZnYR3GIM9yOlESeHoiTffm6iOhBNiKvg7eEO4BcRy4O+k1ZLU5MAQKDN
VAfGQhSXo1eUiLuj9OOxf+a+672CkgeffNBc+v/VB2PjvmiqxRfx+rgJitp6PTpKK+KpXCV986Kw
0MsIAqflrC8fIcYbkysReEtrJISzK5tLAVV3rhdGf7IX5Z6hSSEs1ysmNeuSnKOVITsVcFVTsD0t
cDC0XNCKWRecOjL6l78oF9OrTNeRzY31id7fVee9DmCyaAXufa5VKEk8G2UDgq3MM1fTOewMBYte
S7UbFLOLTJ928n9SfQO3ONjjh0eTtQmO5EZ1EVUwFX2iZbhmcsqnjYkPYaD/5i6VYv9Q/2OGji0k
r1Q9JCQA+PCXCLOPZc1qTzAuU62SRhyPOUPiqwVQ3vaDntE0ehB6vR3vc6wKahdcLv/zwE5qtnDR
L2z0auavox95HONJjpiTmoI/96PtXckVQwRHMziWgkHiEsMcJxQigLZRFGH9Hl6EHBHCwBUpQabl
0e0e3Ayp1Jhe3B8jYcF9A/vsKPgI/aQP4cnuBR9z9GdTmNn4Cuoe5SNKdIp7o2WELcFM7Xqw9K82
gT17fhFIt4yM/dY4ZTp52x/AjkhJFbPjbbtX+yXgM37GryB/p856PDw9qwfG+NyuNncwOFZmmkQ2
LBCWuGAL6PPG1s7gqyPNK5+PpluTjph1kda3oJzEEulu5opUq1cBo9O/9INcC4RlSv7Zaz+DJYo/
bJds8C+x4RfW0Lx5t2iAJ6qfxVxLSBY7MbwAJQ5hDuep1TzaQXhc3VYiveHOUlmw34lul6Fy/Al1
0+kf78an08P9e4KM7BK4RavEgri3axdBILCqn+RLFtHjH/xsUppFo7nt7mZhwRv5E2pdvT5JXoiC
hDcV4XChf0Y1yQZAVqu5+GSAqKirG4tLf6ZHEbBRupozcMlNAuCmwlPGRzmiA4HFKHCC3ml/fMQP
FuPudbKyXt7saTuRMEharekbQTYn8Pbf8cKS4RvzD/UEWyC+ragzeIqj5YxXBT5aAYWMHXWASGwB
IU0QwZlvmjZ6QqBVso5FQA1ADWyUaJzX7cMysckmvT/drgOKC2jfAgp7GfEvAzNQVy8GIq4vuiiA
LMC8S86na46qK2DhsJlIxF1aOsrlNZvSCGzyvPw9KKbPm0YoeV7CiBcEdMRBOg2pudtpKwU6cb/s
J9AabBEEWQ4pz6m69rnugovyo3QnKHN5C5lW+flzT8kvAQKQVDJ7qyEm9kH1Ua5jKv9DevlfVrm6
KfXumlsCLNgCSpJOlmJpbjof7wauIbeTGxA5soNYMKBxuSPT0ATi2Qk8ZZd2MO3/0KnNTZwfbchw
xavEwtgSzgcZCrHisPQLmLI1ZqFsc2RM8c5eSMiRO4pjs2DYcmafshynvnlfX0cLctGOKmoLTeeK
GUok+g2s/fwfESSYtONCMlRTOWNgJ1aRf5+ETMwcC109qrjFSY3nednPn4mqALUTUU6ngfhjv0Yi
MRQNFZXzHHJiychqyfx4QW45jiBmMFSHZTBrK9bKS8IqNz2ha2Dk9vh56zNqnUI49clyPphuEMxS
VFePxruaQ8JWxwpLBRRAdhJmoZia8ZEHb0rS++xfsJ/rS+KTdzWzOixC8RDF735Kd9VJx61N3oRv
WUwWnr5bV67ERqcFyRcbNx8YSm86w0e9OBuFadJUV6H39McPhk0ytLaPx2SBfwGQocC1xHGC0Ce/
9AQGhYw6JTmFlF8FL412eSPrvCkkXkxhos23pSawokrSTD/RphXgGE8ldseX2DZzJMVnySGBvaJO
bPBNZjVHKrxPYezAtwI+hvAs4lUYv+TYbRIlqZkOf1cAMEXLOk68cVkbKMQRBXUkRE1ewHB5+q/4
/3HaWOhiUb0/29SIAsHYO8LE6YA5DeDDr9OWvxz2MhsZtvq3Hq1x68n4R/s/5W8qb5SqM4Yldy9E
vLAQtXvmO8XC+L5iOGLG0AUBvzarFEZdbdHqEa/hH1sB1+USZ8EoglYPMcC60lj0bCzhUrTtGLEc
95/Hm6bldWiF7jBEphIXRHi+173JvxGm9Xkf1na5bbagExF0elt/RDEsXXpvyt4tGoTEjWfPMDxU
COlhKlECgcs2hfe/z9Np+cl5AlQZLvv3i57V+8uiTYb/V7zc6Z/8kGK9QOgC/5wHUF/Nd8sbYkyj
u9+oFq/pNTmdtHbMRav3O5m2NBTpfNrdcDYT2OC1KA0ieZxQkLgcMqcuJ3L7XwmYGaUHBygKOoTP
Akitasut6FbEcb7B6LcBwTRzRIFIT+kOkRyWchYnxAchHRlDVheHfKQGqVSwfR1oAloqOz5fMr6Q
x4bkViVh5yrRNWZI3mzqTp0G0m6zzy4otZLYV56IMJgUva0giEqfTErPJdCi5FJFGauWcTqs8y7s
I1LsSTk9Bt2tXPW3LdqfRdO7qB2xR6pQG23k2IdfZZx/jjLQGYw+4w8uj9SoA3NjcUKolyGSr/dw
95xGic72Ou84eEoeJbh3eIhxb++1akWby5L0XtW/DU040WYMzy38LNAs33zF8y/AWGiA/KARz8WR
VQmtamBpm0vw9ngvkkp3FetfMtVnOXoM71ZhTbisVgbbda/eX52NzalLkvAwEMGAyEER1H/eOnO5
3U9m0CZof1y1oO0nRwu6aUAl4b+mj5JriwRC7A400rDbqAkUjGygiy2NxkUDSrUNrQGCdi2iii9j
b676v6PeQY7C622ARgKeh7I5Wu7zg4w7ciY/y3pMAbErJnuRyxX1+nWSamTLS2Ed1/OWw0rC9RUG
D0T39JhYmkmtf/EAEzOkf+UBKCr4pGU/76yl3GFBiJX3Kw8YhJAX6UBHXNW8q9jhzaKSGk0qfKmH
Bcj8hVAUnztDYwNbFUyorCYcvZhldfnmqZFa/BSrE20cT9lEbzNl931/et/JulBYAmEuLybqDOpI
And5UiPokknDMvTgU5cqtw/ecgvx/Q8fY1kVPIHQniXXkEekwzgWC8uH2NZtWxQKXWUwtrsKwHnt
DQVfUM2O9CQ1xA3LKpYzUEb96fssW/MZSCulhiBuQTLJZJJw3o8wXMLnG5daYMw4rNTY0ZWWwIp6
magooU5Net5nQQEEyXnsNrt2bth3BgfF7NYf6/H2QBrtXrpWMxYqv3RoP2S4zI+PU4YIqc8Odbk0
+PCY5yLMpv/BEGYv8P5YoNx+T19KQLJBJ3qffxnbhbKz83cKQahfXSRiTRsGhlvIDcT3uFS6ejHY
tZclVQOc08dCXcX3UUJOmvk9lm3QMzj6eK8pgOJZtAtI7zDi3OR0/AwYltGo8M8qrTPrSlP/mbmG
7+HdAwIm3SGDo7EevoQrpAPFhO1/AOobXBbzb7xklCWsI3IPGtp9FfiqzOivyorgiHOUqYNqnErF
GQxuI3cr+Pg8Y2NKrJGtVNZaGMYB0nRJqBBXJ64Fkn0YHbqVX6v9QAXnEU7/zZ6OljIv8JRYgj5d
0vBuTnPRrrdCRhgmRIlAMJ/ldw77WIWbkkcwCSr9mYwQGXftoB6bLjJS5pmFaNDByar1CWJ3DCF4
x1sCrzTkzkuDdp5HOGSy8N6qMhuD19Sil2fu/61y8DRJugKy9FINFSZuh9bSjumyTDeQFf9vQrx0
xkP9ffFWQa563wLqHa1uLzu7egySI8vpGOfJX2qqWiezpBtPiRLbTNjDtEX4Xkmx+01TcZldaWni
qjquAHEd8M7k7t3EgVZ2rXvbBi/KE8HM0e0bMJMOWA7q4vQCHQzRryjAldLAGKuR5Nhp86jP4i8Y
/60/V3zuFXjPvS9Ea0mhnsafp3P23MndSiwKj2HWIYbmnIMPlA2Yhl8m38uhUDtz/10RSdfNNKtW
QHwyjucoeg/sOzJBUFyI+biTqhpTvpzQUmDwb3nx/21sZntWM31swz0ytKSDBFEgR64RCRB5Fzo7
nPnfxDsASquzfjlt2+o5w+y4WUxQGi4JDUjGjlr41W7h0K8VusVNtMzcuU/qJ7sTb4rsNv50Pi1r
BUB1RFcuWu/S5/A7fznbYvdDQ4Z9QTHo0dJsq6xh1XIslsCzLPzXaoxYIdV7wz40wDhdP3ariiwN
tk3TSoW7TkvNiN2Boo+VlY6adyCugJVDXxbnGU3F0dqrh2bUn16EkHY5kOhmmvXhL/gXnG8HHLxj
vD+6ax0GtUikJ+wsQpnmkfFeE4zgcWgMBr0P93a5rhut8xX6YESDSZshVRkpaUOoQAlowTZqUVP5
LK6bfksX9Yk7hcbARlhHwhV8nASKbsvA/qdfDm/NU6Z2VGULG4ooNm4r1oapePLFAp4cbvHS1/O2
Q3pTIM5cZYOlFmEAMhK5bAnYEpoVk2rsJafgmH+h2mbVNZ3qgw8Fzm5/AT9gAOvcA61XPH0ZVD4G
qxJpWnTVbvvrCHznPC+2eAMQblNmIh5fnOInvjTM/Bioq/hA1Mo6/euJQMPNPlOv1OfpuTatAw4K
FS9UH5tOL5tJQbNPPt4jc+R6YFKt25hnXqRFYoDHjLyYh4pzr6M060PkbG62LEzJru5Ft7JgXi2W
yQm/SGcIBiQhCL/jqpywXN7M4O0EJP9ZmSuxvnGFM2nc8wj4vcHn5fvfSh7Ta0EjlPsj1bfiVqL8
xOE+TZJZ0HO+HyNaWb3X1lyvEUQPxwzKxXMj2PQOvJlF5Mw9zbINIzIJUjp2bQQQx8qmqrnL/hb4
UEzPtUCS1UmrzfTGKgFexwfw30+akkQuQQ3OHSDjH2Zm53HE1qhKFw3nleEkkXZqH1/Zgqfunnwx
zQo4+jze4M9IaK64DedhuOhAoyiUr0LrLV0AvEGtasErfTW4pJUO3hYkI/OXTQyuK+KHDazgn/zG
VCCWtZQTrok+/CWS4xjPXtLlG5RhWRHm6LwUDu7Kvc9WU7edDODdCw+3DaF9fIJTCWLHth3xMd3Y
Pi4z4xGBsdAXSIQlIu7R84hlwQO5osIn30G7sV0tcFdrBJgEHIgITlqIFZuCSmsya3ZsRNRk0CVw
5KEX2L4eH95LK5W7RxqE6h6GcIgZku8bPqOfJ+Howck4tuy0YKzAIsK3kEwOnQWbphRe98EpiF+N
5IrYJBKW7+YDjqP3DBbgCT0PwcCfQ7CNKenmMD4BzRiylBqqK4c5iT/P1jlB4QSTU5XnRnzdeLd9
btXyCFr9pnFy0AqxOmGXfYnu/gME6SezDV023UwMT6Yh/Vz821lfum0ETq3+aBN6h4FPB9cfH03C
8HhFSz8BuGCCEKZsCr+wfS4PGJ1zQZ8rwJWZCRn3y9ZW9EevAyzMhmln+REFRzYWZOJgnXfduRVz
e7zY2EqiAAtb9Z9U3ObxhbDXrFioFd0AaJoUMQr8AkDyN5O/twE4HsUYFL5bDKU+O4Xa2psnEIiT
LWQ4KBed06qUH/hM+MPy5GUXRIn1jY2osFHMuczNE72a8yr3mQcMwdkRPQ2ONsILj7ZySBziSpHv
fKeObRcaoV7L63MX/c+tZE8aB3uZTl6ZWZoAeU1iMSLsVxlV2ZmY5yrOPfn7JU2T62bG6rrs02Ie
9kz5OSglaG9SFLuF4Q1hLVx5lU/VTjNtw4+ibH+mFDeQ9XQg4E/QCzGzj73AvjGNFsWVP1pNwCDM
pKACTIHinmpyf64w3eTv1A75lV4bxdAhkfKc1A1n29Tt7ZAk3/J0mUGoIq7yaliWtfzIJnVRw+wr
t9fNXFPpfiaf2dttOH9YNHfKFEHfSJQJI+dUfofZEkKvJ3Qfz7EU5ewVOeVqXpQSSU8KYPz/tLpp
W8hyfN7zZ4JowGIv9FLB96dSVADL5NiKVm2lv3LJWddGYjVc+bONPy+fGRrwXCIjLZv54B0vlRI6
OKmIOjD/c9wXuQXGe0LNzywUh4NYrKT6VEjYbQpCnZ2KPyQ8ISwO/1+Ict9nPtOD5ImX//PB8hfH
PW8Lg/o3B+CscuL+OsVpgpnUzZ0df7+HiVb5V37V1ndPeYKq6zILQC3k/a1QTmS/fIn9GbsQMV0n
0H5dzVnJYfDcXALf4eSseWJt6qBIlCGcuDo+dn1Vrag0UqlA33y28wbXasEm0Rr4HnJJOaZQI77D
LxkAxJUvpqd7bKF39tPU2oQc45joSk0FQhzOZlks61Qd7j9Ac2512XaHhUdDkLGl3s+WYfcdK2NC
gnDYoprIFgeX79xooonGh5IJ0WjdD59bNFPOWf7/AQXe7zAnzEPkFh9rnTIExiQzyQ38ggIbKiE2
/GNm6INLOHfRfNSznO2bjd3HuDRZXJX9n3JQjcJUZAaiaKxG7tMQKxtvTolhTwecLdTrInuZPJvV
Wvob3ZgjKTNDuwlavNowDALF8TGSH3lFT4cSVollzFq2m5DzuuJNG+7flp2GxYW0Z6afAt+YMiXx
uMI9SWBKfrC3L6lwsbxhUWc62dgpivdCULMr33PHfLQW1i7O93mWe8N5M1MAg4RLSGKCCWMc64ml
ymgRUCAlLlBgeoFb9jwhbJZLzezaos3tiazZaQtSZcvjSej4jrDOhx/cSBahYHmOyDFkHVdmBc4z
MLI/ihV1vPZVEAR3pNj4q9F3MgLNwM2tkN0j1G05s4S1GZNp5+MpPHkaCSEO0OEIWXj+hF+3DeYR
lIU6jKVT6HSl9JObSF2/SXbstNCqqDTX7zDdIn55OswJu+KDt4lCZYkltdfoyU6AjXpLQsyCk8wp
1qvdRjhw2q+691YC12+ERdFsBHYUOKJHYrkWMLoo/FXKm7VdZD/gFx07HYrcTFkWS9+fwvNv7LUx
MDdpNYG6beTjEeOjlOoNxszad6fd6e0RnfFvM5JM+hWMguRMnMO+aI510lqM+0OFsBSeYaC7S4se
/RPR+LZCGkcEG1P8OOtuTKCPL2HVFujpw1eAGd4yKo+9esjPxRMwztU+jhvSJL1hYJxD8Y3p203A
Bc1oJsqKxuCSzzqBJINQBnlmPM3m0hNfZ2hlAnov5nQlb2//W2KRV3izX/Q6gPWxR++FFMsTCf/k
V5iKIPNfEg+glt8MCXh1OA+3NralwoEtA3GuQOfvdcyxp9dEPCG+HhzGhbDbDs2jD18zBrnkLslY
tX5wQWmj9tEWhbjdvbLS8lYgwl3U7t8vvdCOV0SjvB7TrV3qnH2N4ypgH7D6NBp1VIez7FXYcxpA
H5vws1gwy2CnyKezYFJCXKbmSi7iqN9jEm6PBg1HaKGOpe3RYPd7iAhQNmUKTlY1Ljn/HxNMUTbn
o/F2w8aw2/+cL8OnQSk00gUs/S49vwvjXKIlj2Q6UK5mEyi6cA/lJMsrEDr8QUyw0ASBsIlve6l2
TTZjZRvm/H6eQ9mGxVa70AjVXmY5BUWyHQ57FTo9GVUja3tptmWZe4UUpXA00UWnGmzC0SEIOy7c
GNUXYyctLycSv4rpaXy2SHu5gWZ0NqRd5RfxsOYFlD/OxJxGE2lUYuBTowQN/FdhfIYFLh5WIdO+
HamOXfzf+JwMU5xPwGyqOnq0QLY+ImdYNDDkvBTfs4vIVbnaON912wtg5OZqa7+ADDLJ1d5rE5ZC
5GfzfGNBLbkC/0eRkhHi3j/NZzZs5770xqyNLovxqdPAlSEV0wLc73Sd0+cmw3qzlz2Lqub0zXF2
GHlgou/czo3yOXHMfQcpDnlCBc3D3ULRuux6ED0R5SZywmcvfkdUTE0VAxvqDY/UI9Uheaq/EW2M
df1aQEFTaAkiTYv2sOcWkmzENz/MukHXuICNdJ8DRoKQtkieosiMc/QMq2IaApK5xci/pqB+PQRQ
QCuh2fSgsSrV/AADtG6/ZZq5L70ScWXTpKqfiGL3yBYS5SKtmLC/WtBFExW7ClKHc75SIHRXre8U
KZvEy9gse1uPTt6UgV0f+D1HewHVZ7liundicSY9EnhZF2r/G4K8ZpqmXtsZ5wHQM0gGwPPaU0Gv
IGR91UaFsY72WcHBJhd5b8CMH6Flxo9khwHIqq/Hfq+1wGF5k3zJqTy66AAsGm+OqjKMcLlwYDp0
d0clHpwangU53oWCTrW9gWBGYpYYVhN3uFFRBWhj8zxPV/FESf/PMEGujoZI0M5Mi5UznKFkvOq6
Pphfmd7k5y6bB7U0aIszUCSRqvGGyVwPefPu157pOwQbx7zbfdQRXu9Zlmrkd1xz+EcrMwnYLCSk
IsTrV1HEwYRA+KFgC0WvAIWviR29qvd1b8g3sQs9NNlINdm4JKPphPrgbvw5aDZTA8rLsMBj45dD
jDZczgow9OaTv0KjA1DLKmUIfUaO/oj3ZfMMeGP6ozW5Z+GPF3Ust/hosvALieiMeTBM5PFwdath
o21SPOkKvt/+8bYE8GsxyvhbQ5iZ5H5VI+OPVsMlTMk3DKsLEs/0/CvDyOub54kJRMflrMACGB5C
gxFOGtMXLOvfe2jT/VWuffnY25hitDd/b3aXyuPC7GvhUcdA+l4ZkK33fG9J33jcFDVFRhRfF3xW
QAZ1yCdxX8HcTUbb3d+5/eCynu5m3uoiimhzWcnLokFx+02G/FgYyHReTo2ffD+GVi9g6+xGio1L
NDCIiYPLwJ5WJqz3b87XhGFiiH+d1G9qk800W6ueRHPQIpT6gYK5WBsEIY3RQLMuNtUsIVLMKQiK
vUrrYOvbidhBqCJadby0tV4ITcQs14f0UUiBhN+fBjpaQiRIZ7qkSrvxUEhmnJQvC9NHYjf3Rmjw
HJzdIj2L6yuI/mLOV0UHJOHx+fHVNM5Ujio4jRZC28M1RBjQheC68uSlL34TXuXzp7q9WJs+/2SS
CP2ekG/uXIayYYKEpfjeTg98eSfPH12QinBE+AiAdsbtuz1C0Z/lAFhW6y2aVUuXUQcRHoHhjtHo
CdF9wf/V+mco2F5OV0tYqoF4AAnC72z3bTFoAyESr/GTCoADbsk24eSUxS/C4yc5Y0+10ahkpT03
RFUlA05GRw84iiF3elbwCpNwl5zDDN1VczR2NvJM8lPO+IGzqsbGa+fpcvgTSNl6FroTy3ZYb0/Z
FNTql8aGQkeDeJChfwi09c4sD1SL8Si2fhgSpSoe5PK3p4Ft0s0Nh/r3xBSPWuGnoH/rVGGQIkD/
r5tkEElJYQmyHH9NuelbDaxX18NA4FMbzZyM03o1MP08RH3rjk5XFvOVnYfqcmNMatfY+NrjSkex
kBZs/GyYcsld2odWmQ9hrN2jND4DyL+WXrGf46u9207tyEPRk9zZPeVUPEiLlPDctI84mgES6ksL
OFQAz/zbAEAHTCPVUghW8CQOtBcBLMXCEkmbrxfHFrUqog19R7UiXoSNW5UK7Vo7NMrvgawqULDZ
EX6HMFYtuj3a8yOGLRT/Du4UbY7qikX7WOI4SX8zuBO+7zBLtQ8Kla9WZ1iwoqs+UVhI2uKd66yZ
Y9FBvzugZ3i5Hrv3i0YacTTdmd4L2s3JWq8ui5WXR2Xg+OiUptoX+eSwplJXGlRw2WAbnnOepVzK
aaiYqNQH/fVyYO5M63BDbIUm/MW35SjhnbSf0CYVgIQpgPWH7aHDR4SbQaig4AwxQnxv9SN2+Jpv
SJ4jVNY33NawVQLB0LHJnhoGmdyEXYhjY2OeIKyeiYA6BEWqvzME0mr7YDavBfSvZbeNYsTVchAO
NHTDM794va6vqsp54M306yekP5LR0l+AOHEoOVxHER4yyS2kOrSbj9UIenKQBg/5OSCzopNJoEz1
xtTsiyrKdTYYlsfsVBYjUxX2i2WqzpBRSVxlsnVGlMQWTCUhIeI5uEIJmUE1AI1mzavtc1iUKCED
2ELiiYWI823EThyNSZHy1UD9/TSSPhOabhYUDpNJnX1PX3vRsfGoIobn/Mxsis5KjxEKjoJ9UIoW
vCkgW+hnAwEuTWfgq4LWajAK0gdmKd6k9LGil96k0n0CahIp7VBy9FgN0XYZwI00+rProlO9R60J
MBeXAL0mcof8OlXNG0jwDi83EocD/i6pAB1Qm8BId9PgK5KJ/VBVgyy1QyIFICWSy3wX+fJH5V+h
C7fFHDu71zdo+skaNX6d01kYfFpzf9Z9YV/MEVlkBg75xfjvLRUMQQaL7jXCd7jqxSLGnrDwS5ad
bH0xnVkkate4qFZ5SEOyb/Sw9XS7yKIxqj0k3pc6VLnTSezyz57R01S+lEDMP1+A5qKPHJ1K2eId
2fL9UJAbMA/8Xfq6wqTUsTBxCsqxT0toEYEmyOdlDA+ZsgVd4Q3jJMKtuaMr9uu3U/TGXtExvNPD
sOZh7h8LzDtH2a4WTx2iDZ7znW9ori3+ymgCs3OMGqTZXuPxGAEASDd/ty3Zr9DvN+l/un3NHKgQ
nKA6hjOtEa4ynUtd6qTzeA45Yjf97YkniY9Bcozhhbmr8gBudFy/PZMmei02+cVX3LyPZ22pOKFX
ZyNP4FdI3pQfEzo1fBUzynXkmpayj+fXMpFcDY9gQaHQIUlzZT4nbdDqlflqvooSeGbJq7K7WdVL
xT97bcFeok7h09hzkCIfBdY2d/ad1rkcGMrJXEWOrMWhFktRaJqJdrrni8ozi4CqEln10MsXbV76
zvaWGWim4MUVuWltczAAAKPLJYw4H5KPXntCHdczHCnJpu/pG9ZKx+zcPyTi0wgK8tpX6+AYk7Em
sB6/M5kTj/ZX6SGGrEjCHGtA6fP8jJdb2fAWP/OSaoMJFyly4reONyCpgvC26atsVsiEPLQaUPsw
kg5Q8LpcxN1P0Znb2pO9f/ewZEX6YlC98yXWNAt0GcpKhAnF/RDZFJkWCUPEBtsxi0roATxWkge4
8TmQscXw6DSWiiZ/G4Zl2XKA6utF5jvGmfO4nEllRlEmFUbTSbSM1PdUSRKKxVBv755qQaSmAnwb
4v2+JGU4rNvZ1kZuh3WozOL+w+j7YZ/89H6v/ez8QoUHkMJKOCb3tZSiizupvqHE6oegJxlkAjJT
+QXvEGGXtHPZHLsKNMo4GaiDtem0aJ9ELeLe+H2eES0zOCpOjSXnnS6SVXMX+LdAgG9+4dzDA40n
J03gbcX5FNHexvBKscyL2ssU8Dn4sZuOAm+ftAOpjdbYRVaVOVz+4HHyR5t4zdzE8Ul1lUpPH2IZ
f5Szr0rIB6bRPZDB4YV//u6eDeM1oIf7sKiXDLAL5LiEopX4lry6Mn2uKHNM3cVR4yLePRH+qdWa
T+ST57VO9tlHI0TGWLdHP7I97lFCIGYduLr3Fhsyg/0j94NKnUPpEjnlwCKkI944HpmgwMR10eG6
qSqa3huEOu3fHrgGhstkP1jjPbxHLfUvWM/ona3c2yxPohGRljihDiWVD36sLqojnJNpAKe4bTtF
xXSU8IsNW5hRvAaVsEp0WbvexmhRI8AQZFeJLUxxiNv6nPj8PhNEgejpwiLvH3i4wbDQwL9vg5Ku
VPUpEs1cQK1p3czuD63SmD9RaS86ZRQhwqQZq04XTS/Drpo7v3Gpsu5T/+x+ZeiPCEYMbt4n3daT
MG3ihQUMMO5Oi9jvF1lajtylyHliS0d61EOAfnn09mVFdXyMHiqxWndkAB5GB1iEpznpkvE2Rwxx
M6pva3DKD16UgZsTEOsb00b+N5kT88d7r04QGXLR4V359W5Ik8n9kxnhNa9m3huotAfLXg1EFuk8
UCgekjZUsNSAzWKCpkXkgzH7m+akorPzGW72tRUNu5vH9OCllxd6uCgV+ebnp9xW0gs6X9eTIE0c
W8RDrKtx4fgR0bvmYIhaMvxzskGQcuhVdd0yO9GT4DQ0ZZovnXNvUuYmnZWUjd9TOgsC7HKj1SNO
4FbPOQWIt9WyXcApV368C+93eKZGplEKz2bRhmYmjT32X58f+XVZZypNKJB7Rl1olyZ3EZG9VV0r
k6R1Gg07S469EyU2SucRSsVHMNDLDXqYAwspbHJL7i1nafjOCn32Nomke6YPdTYvI1uFmzRNh6bn
NPqpeE5p7tzPuWwKkEvxrS8gQUXczUylgbtiFnKBkCuQZKOa8WQCjak+omCPsstl+Jg7SCI3eOMo
J1qBA1r02j9iGllJRdPu5QJuC4xn2+B7WXF8hqRbC3rpfiAyYKP+Ty17r1zEfQlK/Ra3EMpy4IXZ
i90s2Zr6RGWER393QD+w7kCgckChXDEPvc41zckUc2QHz+H+UO0IkIypfcL/ih/mgmHwZo00SSrI
lvOjw1o5AUBZtP8fLZrvyjunGyv6st3gZUBPixgy7H8rQTgigD7Spt7hKTJe4fU2lWc00SCr3ZFJ
60gZjHofnAr6FJ+B35vxsOqZyEniFT6ielsQpYSdSVVLIlO+kT+Qhs3INyRQpxvxTX8TOy+Fpc3Z
KrfLaNEQIaLIhWaOOdzksUwLtCxA33Urmmtbm4AanGvE6jpY3XB0QzfnxY0s5uM7799HA30p1Hks
4AWWrtGYS6utuzQLnZ6RCAUyfE1dp8ZJ59Pa6VXS9KiqBNK2v1m2dR+YPczVTTUbgHY8xud3bpjP
QdLw4PB8Z6XCuNJfMcx8V0JbFe7tuC+yjk4rnPiptRy8LNsHQQhrdUojg3WSuiTtEmE+pjkIcipe
d1XJUqUPXEvlxXZtBQPhsy7/AlYQQzSSc7Co/om2mRObibLB10Z5RAmWoA1QY3tMJ5wtAbA3zm5a
cePv7Is7dEH2UiVsid/4xzDhDd9fwBfWRa9ERuPm8KucbA2qCoQ+t6z/icDLZItlQ8ZF9Sea7u2s
MGUA2v6ENkd1Klcv1ww0c4YO/7OmWRivs6rDerqmRPVViiRVNXrZr4YDKCPvIhJ1vhstPYC/meKO
RTDlaXTuTItjJqMWJ1jWU4UObGsE46rFQ9CISAdLHrHDSUq/fvG9MryXFQzKV4aS8/IDZgnmEZoZ
j6zvO/hc68eOfv/f8YJACFES0L8d90YmgVrZKOiluQz0Gm2FxuTfpp+dlH+ha+mLAFixsOOMR1YT
zn9wQRAmOLcTypVLs/UpR9g74XIHj/hNAm8URYyXLY9lBWtv1iTiQjB3aaHNTnP+nJPGiYE2FsoT
7KbbF+MCy81SglwK1NTyp1SCkVwLXHtmtTx1OnJZp8VlfLFCwWGMLs1AMriQxsjCF6OOg1V7tizl
F6m0utFeDHcfToy+EOispGFw8wp6iF7xn62pQdT6aRZGmkQibab+hlBB3XDpHKiZ/YhWyYRKgKhe
elFOk1DMdGfncZx9gRANxVZWOZL+Sp7I1GEBBZNnd8ACLGNGb2+ziEMZ0yH3dHVfj/7xkvaZa7P3
zRPwkmFvQO5GyD1XysQk1KSMfaxQqCeiJAquLRKcRHSqmL5HHRFDM2DwzOOJM7flEE1xhZ5AAsPh
ldDvYhQhbtvxdRcgtkCoB+laNQ7g+hS3TWUlbs01KLtRBxS641c6258uCtw3XGubraGbV312XSO5
IHG+MeJmJIPWrJaxROgyJkfVSCwq5WG3sBU4a/BShAqpn+O72y88o+1KPH6Ipb/O1bdNTz7outKZ
3PtuIPTegJVkaByoGf1X3pe9OcaaNcAuoSCWHyAWuSm/pu5uX+kTyiA0PuZYohZqN47inbdB1g8I
AdniF/KDeMQD0mtv/lZmFf/EVQL11nOHLJmCdi5UyUI1eYUfVaux0Q3Jmluy69H4uDNv6JG0/wdG
Jm5/+fdqCszQuUhTqi03Ngot0vGN8x90/WSZe/8NRQ6flYzWwLTiZa8O3PsUQ0XDEde+jMFhS2o2
OrQhJOwFr8cmbS1ID5CXzvWulLGOGkTA1t1hE2hl/GGgrTY2F/+Su8Ro2uWgaRZfYU50yXcTaa42
PU4BoE9A9bWz3MYLpsqXeyMqZp+0BrfFHFw3Vi81P3W/4QhNev2k8w6zk3Axw4J8Ihrdyw5nKERq
3VXkNhZ3RigVf5l9vV/nUjMiaJ6hwPQyU/io/cENs01koWKZVwYaYvo6Evu2kF6VrfuGpG9BBVBh
Z1x7G/Lj33Aa2JGBwKCxko12Cv521KDBzDiDIWm0mO062eKsFATRUcV34Qi/zL+pfXOYVxKpA2f5
AX+Ssq11ujW0DW//EyWRNWaFphItkFOwv9ZQd681+ZyOH3q8krOxVtvgaacaXUzJ47H3YuOzuF3h
7jB36eKZOW6oHMesXQYB/CD/ZZKBeR2Mn8j7m3CLn59X1ik9gKqlMtMZNH6rc9UlVfstaUFPqdtB
y2VARO1V6zWrlvud8K9vjqPIjRkYloLjtrp90T9bHMG2Lxa96Wg8yQ44/lQszAvtayqtEAuxk8Y+
LYjr+2InHkjOP7PiRwCd/7dpyHmp1hqeLL3BRf2p3V4PKmof/Lx8sOPrSahEhBB8rQ/6lOWMeTAy
4W2Ydn896Vb2Yd2/58UuQ4OH6gK29AeB/kZViFvwOiHnfGhBFd6VY1RSw9ZYZLZsYu1V4OLDYozN
S6drgfdkf94CRV8i9rJh6jSK8zSBGgnQWZ7Opxo37L4A5Ue1mTfwXsV0OKUftm1wGBty+Mza3I1p
BNHRtJX0imh+T/XGtm1rq70BzzHAcgHfOXp86Ko1HkI4PZlKU0CiYd6OlI+ziDrlei8XAVpvkhEq
DzHxtAXV3OzCs6cRr24tiIWgdA7L0B5xO+ZwjPACKg+TGT5QBYGFgVVy/se2yljCWrr8R131ff5r
6VrGgxY6LXQV7V0zM87rN/SEPJ+mhJUhVs++VzwwVhHIyx2L8UbuWoO6LlziaaEqCm7UTmUELGCY
2UFo7UvCFTCfL6istLQr0jQ036HGd5jzheZmTy4UMOGT2spOZUug0mQ53Zw3hJCZ84xgS7ij3IbQ
UZOYRk4MWmE/3JBn4QovBFOaD6YF++cCGskTUO2JcuEhcKfEVwU6Me69vWl/fvkv4ubljD4SI+Cv
3Wsob3kpZq23b+lMz3I1/ilBVUDxIhOA2m7g7IEVbOva7WAmiFz2z30RX6SZMKJLSeNpAyAqMtC8
yVCb1How62x4xKtj50tdizsscSnSXZnVis4/6y9G1qCR0sbgcYt0p9rxWNM0GLS+PqT9Fq6ENFd2
mjAbi+BLVqGqQst5O3rDX+OxzFvyX5R0MKPIl+vujucPU0R5UocsHEuvEtHLLXPTrK4QyDPgSX0F
GdoXECQVr/roLPNQ9Uzb3lsGtw2syPWlpwQLrq/YtaMbcNtPM/QfzSvT1uTHt+bj6k3vCOH67sPu
wqfSPJTYFQACi8zMLeel49Jd/EuawzLZphRce4k5JUTV1VM14iGIFgQi1knNo2yDrQ+ysUA0y9GH
oClRdspA55d5BOAqNDeHtxw1p+ZOQgNa9D3jsTIxLM4U4eEbbyvDxVmCCKCAbpuvB1at2aEFItJF
Wv6njIN8KEDqGrD1sGgPWw5s08RwrfY+z1cpyjSTjMQlwKlDG9EekvcJuaMYckWy8ZgWBbTnsAdL
bQ0ZwiN/a1v9NaM+O/eCz3GaDPk5aa7JDRVBK8jf4U79MaqPdmyyFKlIGT2wMbzEp0/edCXj2GMZ
q3Qthcnh+dCsRv7ao8iMmP7f5aHmWX85eq67R6dHlRWroHXTLFFhGMnRpNJoufcWTH6wjpgFWzRT
zXJARHoZ5CO4JW+vh1FAYeYdmpxLTMYRq8QEA6bU/svGn7Gp5LxBpPm/pF9ErjzsJfV2auga5uof
swC9UYtrXTl63x64PLVhvG4gaTLBQAWj2RuSpGc1NzoRpVFl7aV6RpP3Loyz3bg3+3/gtCrwdWNw
i2VhcVSlRiItqZYhXSmd/+Sj7dAWkGV+jWphKw9piO6y4+B8xY9Oft5FHg6WZeboMpffaXWE261o
MelAupoHFiFc7etujZgdVbgAZsHltcAD9Oc19VBWNFE09Q5UBAOhtJ1/V4Xv65V7oREkq887VAgY
NqJTKu6TCZzXoWZXC/9Pe76CZlEA2Np2MUp9WPGMpT+grdSYVzw1UI0vxE6krft7LjFxPQBx73fR
Bo7nkLUHswn88X/y5p88dgU84s/subr7Oh3F8/fgMeWU1YW+y9nQ9dUeRYDpSr3vv/6wXBjFJxzh
f83f/x44AO8B421ljvPUi5zYLkUsXU4+oAIBG0zaluU9fLnQZBqDfo4ozDY+SWuON1zxzNExcYrv
mB91vAb6WNqgDHZ79t5C+Utc+Fa1otd6l8Egz1Rz8jBPrLuPo7xs9ct/RyDQskyPOLJObkK7TXqW
zCGWn76yoV6P+mY570ekTmeWlNnUQyW2Y7Xub70DqrWfe1Gbq4x+pFQ85Vxxy3japk0YELmfLL1w
9fxPUOiOcLmkBOz3MPoVtAbSNUsSvWH/3kKGcTK6B5UBo3kn5eIyR6szdCZy+51TID1Wgd42bLDg
ydCSuuvYmzmH65soQkGBmLpcQd+LPopv2cMuBsn498AQUXViG9rrTJWctioDoEGTE+nAtbvi+GVe
xewHIIIeluj0oKv0MuPuQ+gR9mAcW6rHayqdUyyKI3fncWzpbz+G6FeKXMDBkHptYxzYyxajzKA+
G3WEI9NTK9l4qI6TJJw8ES3cWAI3JICxmQ6o1ogukVcFhRX7Ilzxvqp5Xb41PNV8QmVa45+tV5ue
VREF9AybF8yY7FzYJfwBj3aJJWgmuyUlJBI18mRz0IPgCDKb90VnjeN9YSxA6yuenACtcrKafjBc
pXwHsGIcONnmgcsmbV+YZIQELGc853RNx8jakTugKhihek5Jl1GmzVDlQbp39XmYKHHKi57VgbP7
bRTzQIbNgNbVK5bhRbDGtUPC02FVptV+IXRQH9jSOyX3XObMlO2Lvj29j4wbkFaOUaDXzH26orfQ
V1lCnY1rGgkqxJ+zZ8gTpQSVoxYDEK0jQg0b+RDwJjeOF957wdIzivA9vQY6ZPSaHz+qq28pNTkD
xIg+/sFipa8j5wfcSpbBkJfMhLonvcLGJe+/AmlaNx52sNGfU9EM60w/15R5yN3ZuUWXYPrd4ROA
E3JByPYVWxFK7iDauDhWwAGezY7DHx5qjmtvNT19KRu/q67pUgmBWlXN3MMnQDmu93fWclEh+z5C
joWe+xau4eT1Po1v9xPB0WqGv0kDUnHiZ8/05nyAezX44E+HzutXJPppoPJhNw7dlyHjFJxhSvwM
KkAxtMF8dPydgAPJxeqCUmLVkN7sirsa/NXCpevNEf5iBIHFX9evmHrZ1uR4zePPOcX/ibY4gnps
Sd76uaUa0cfSl8oHnAFj79O5g4SpoQeHiIxMnFs3M6riLUoA8z5wRGuCuH/37YCvFc+CCmFMEY7a
iVBf3/8YzHkRHAbHuswCog+sAKNbl2uZURp80AHOMFZB2NnLF57KV6OsSfOSIdPV7YEhoZFBt2gv
NtiWJFzHT804Chgf+4FZEIUL3bRuJPvoHFAWHz1ot7ONPqJwlOdpjrKlblgQk2r9mUTE5Qfp4C8N
ssEwkDjIAY6SM3DRo3nv9z0zzZL050rgwXWYECwJrpuYHqfo9+F0ILZHKlFSN7mR4h66ZaAswVuX
aaIwIOvtdD20XE2slfBoX4+TnW0hg0w3mwx1ofJViKk/M2Ds2uuacxPQQcB5v56YBsFRJYny9f+D
svKh/eCntcaLniJLgpwZ1oxNzVxwLy/NSygK3IONaSW+k6ieStun8txWROJW4lC2fSdv07Ickula
wSkSuf1LDAc2hKwEcU4s3yJ3JDRsxFf8S5rgTRBnMKx6ZJn2DBxDVlrUqyukJwhb0tV0yq90QxhC
F0a4Mew76sZ9fv+aBYCtRTXy6JNr2K/1q4sgc0Ouer7kz1SWbcv8WrKBDmo1ZXnwWQ+ferJaJl8V
HsteTPZmyeMrKMYiZCi8KMzPiPj9eWED1mVg1FhpJDRxqX3/gqgs88YMVexcpGkFq/N7O8LCba5U
POpExqkuajjmJuYT2rEGqb1QFhN/xZClmNIvq5VAdaSDuma7jrGb9HGSeE+a1t0CIra9kJrZgJI1
9rO0meKGxkfpPySraUkfpd2mF1IE2KOBOTHij8wxz4Ddk0pRXyetd4OJkneyAahtdMORbKWNNnlz
meG4HCsctkvP4aUcTrJqYSaTm6iCuGJdJMVdrBvUxWW5A0ACbG88aP8gbabX8WGzwLubrJuTlUbW
4iJcJc/PcEuieRINwFcVEIxdAUXj0E7TeW0XDprYfCv2FBI9b42E+9CdrVb/1MF8gWMMeHzUrnIq
27mSL17Fv8TlpKptHP1rZdcb3mG3Zmdc/DRYpySpFFKteSYeGcctSUsgpFdPtDsItZKXiGEo7aHU
gPTeFfojwTNEsp8J6xUVrkFWZEzJ+APS57JNdSzWXsYEooiin3UV9+SqEqLrANsH6vb8wmcNrJwD
1Sn/LAJ90ot+NpZxp1cfUEJr/VoAlF2ZayH2EvHff8bHlCptvDn4E7nD2cllrjmPP7YWmJtFfPsO
CCQcHcMODovHunQXNI0JmuJvRGfSdz38bFUcY8MmLvxkYkjINmtFvs7mNmhwmNgB61WVbmLN0o2V
1sghbdLNgSFTCXoNX1mTHzrLqS14EdRelQdQFvmuj9p9oCQd4uqk9DHaY0/YGCn9P8rSpgM9HOEW
5B8MM558Er5j/3LrJ0SgNLgTQw79M39hY4vEe6V2ramnRnMrMrXxIcrBF+R5Pls91eEIlBIdUtnt
6znK9z3Qv6Ujg71GiTL93eZY9/9ZLnHF0VE8LI+Zfn/2nHeXqTL8N3VdFmvF6ZhL2XE65x8KS4Om
BIz5deUhqe02Ypfvd5Rug0512dsj9aXTCfB7nyYqb2b6LMoT04f7crx9FJVVh3gp1trm/dixh091
dwQaaRmDNITM0Enap3f8rYQ+fFlTrQzlrnXz6NIbtm4m8C60XFxuwKW1hzc5Pn7Sg1tv0qc5V6r5
TESsGx8L5zZWpHSi2KghLcwWJI8QvMmSAxs3I3cohnh7ovVOpVCcVdYe6LMRKbvaLWjNbsdvbHyO
kbF90seOhvhDgdK9hgIBiDWhS7WEwTlus3v1oezWyp0mP87xD/b3h+iVcjoGO0tutFdp5nmIp5LK
IMzw9mQGexEIaGn6sxtaD5d7VE7vUgF1HCKli0/GCFLKhuRTDmswGcjj+CEXq0EZfb/Yflh5tkA0
r0+4zELnrLx3PPLjPEqHbkCZb21U++7Hhnx181HMgmB/VyD0Bd2/0GCYCQzk0YAZdwVSb2CKYaM6
SQTTN/QJ1tnV546sPZ7sshbmDghukGa77w1tFRfZ7LU8f4n0qxXQlv3C8BJALrkw69v60WSoeA7Z
7weSFIGUbHi+c/fEg8COXP59p6LtrGrbHhKdmxfwdodkEchhzdD25TxqJY2KEf8DhtavHlnZocXN
IpU4zv7Gh+TAcNF2Ori33mQwr8eNvQH/1z3DwhBqzJKUxma0Hdv6maQvD8W2bejOifKQ6zGo5OVt
sHjZdhXm8FOS5vm41laTNIkAbROxOoOQh2LRXjNrOB45Op6jd4vif2fWkV+7ge0xrHyMTKHr0kjN
dzU2ck6RcIjqkzfjgMMVD/DMpp+oDrpJqKHwDX34/qQc+cQxJZiXMecyQmFqTIfOea5508n/l9yv
uyUDX0BkDufIpJRWmG51IE08cdhk/ydhrn/yqYGLXeaPnrYNzkeMulA3HvtcgAes/eXXRxMo6bdl
W9OG/rus1qwLU8cdVezm0fetVXl1AB7dVej9f+65vjkEh3wowddwvvwYsmch21wuk4/8X/kVgzjA
fbb4rSHteTxrGc3GqbUejs9NZU64Ck1MfQT81lwxv0t2NhP68d8m+U3o6yBUpWv/b+IryuJJltJj
Y18rm96QbP092DYC/nRVUI6Xyy/nI1qm8qs4NbcAH1sLnlK9AwG/Da1oLWdN4TVw7RSvBwwGtbcm
7paC01+dOcuPX20IFq+6H4FGqlsLNXH0WO9PX2XaPItPP1pWmy063W1GJZWIDz2iwXVUC8jaKP70
+sY5xg/nK+fLjMARo1w2656DYKy69+GSTv1UZq55c76nxf0b8nh7kksrTwa2BfxLFqKxnAG/9i8i
VS1wTcWLAm/atYuufTJu8kC+FeLxllK420SH9P80kCULk4oQaEXVw1MEOCe90jSsiK3el2eCP7wf
JuSD/seQbsSehIzrnRfVuQz52fghWDW61k0hbkJfY2pH3ows6L85BfIfOARUqSNim/gqf+UeDYII
TclQnnF4GcQYSc3k153uEHi/iVWS1UMW2bJIs9fB0wGX8hEnVntgSzVoCC0FXw8Wws6QjaHfUt7f
qxzMa0K82/NVR2Qd6gx0cvMZgjYnwN5kRs9RwuPfgNq7rQTHdEJtNp4QqbplSfz7F6jFTzySMQ6n
CWEdnKXDKJJfHxmyMm/eKCZHPrLO2mGmoj55v37ZLaeg+YZHldlVz1dPTvYhAt/4q5/QoRM8pd57
FjELN1Pd8tSITktVyklQRr6AuztZHJ8OHAOwslw3h2gkV7uytqdPwX0qClYU4+U1ZDjYGTkMV4z2
7Hmu6m+KukrC4Cr8BsqtF553hygLISVHzUwoiftFQ4PPZuEilMD7KFrSNVEHCyrBNwiIC8XqF6fD
XBIYkq5jappanurF85lBebpQj/fLuv2EonEnpezcjcdxhUw3VN1ImX+IRvYQ3en32mhMWk6i8Fyl
0sgnwJglQaM11S98ZnvmTB3wTpbWODLJ3CzUEro2ZH7agJamfE27a7CsMAeTSCasBJEDVzXkavNy
u7QCQaEO6GTnvOyCe17OvZK8l87P08KojaYdKOzMYs8k0Iatitd/PkCEkkgqAYGZKMTIkYoMFoZ0
ecCMuGv//rjLP5C/IgK+86smIqLlm/WmuNPBQMtV2V42xpIdPGhmfxKd0HqcOz17ejhgZZSBIhRH
F33Qa9xthmOBrbxLtgx+wmtBffP8SneJar7oSOe2HKT0X7I5B1nbhgAXeU0XUxml5Wari5qxnX4M
VsOw0rphVq2p9YXzMJ5gdrEoqzbTsHKgIbmwHXWqnmVNVTCGtPUx63FMHcMpBeNop5IrGuvZpOyP
x51wUQcMNITTo6EqjGnwVHpdAKR4DHzMs0spIUqYCLF0ai8LkKcnqmBWeUzD0yqXNyTYmGK5v9+y
RGKosqdHTx3DS2p6oU3iNAGt7MkUBn0j0FxDRJoNaZS/pgFZySvZjIQe50QBa1JruZGh4W5kM0CJ
jenox2SwEX+JCbW5gPupYFaOVOkDW+HZS1J+UYc8jdGbiIc14lqmXSJkabyJwy8Yq+c8Waj6B6dY
PE3iaYE+ewG4BiRw3XXoJ31n46d2aATE+YKwOkC5TtPgCGMx02rFjn0byCyrtQ74gn2dxqSXx8h7
bK4TKvGLszF/Z+H7tAro8VdtGUd2mvDpg2lGUDi9G1MNRkJVhmZn0Pb4uGYn7sT/PqtlsB3FYJff
RRPE1Iywr0RVlIUAYR9Xljw1b7a84PZ/y3v4WU6xTuDXjYShzVl+VPLJBTjP65A8GwQsUIf3ptke
f+bCEeYhmRPj1XZkY0kITlApC6yQHOhC8IA5yVcnVg1N3L7jlucumxR4Tpc4Qj9EZqPG8vs0MO35
sHkGtiH7SyKbhDoFPrb1wtZQidtJjvkkVWVMechtwlnGgzddGo4Nv51GmA5kHvnOpDtF+2Xa3KEr
2kdRy/UwEQyrNGDRsHRb904qDDEOQ9G7Xq4G+a7WcrVE+e8DCzS3/ZD7AitunM/Uiywc1VS4CelZ
lZ1huDjLJFDJrxZahmCq/5aM7LgSBhEQ9vV3Uue/e5JpBdv4hmHA9se/rAJW5qZ1qu5eEn3aAfob
J0pORR52eX/oSS5pDa/K1n5Q0t1QVa/PQplOKeKQHD4aE/RaK4E/zdpR9Hd/vqXJFSRjEnd1QDVk
UTIt4lv4utlhpMiu9dZSxI5EnXcwTstubxwmSs1flOpUGj5RGGixS2yyQQGBGnAZx67ccLGDs/Uu
fK3Vy4VWTQ5A1jD1KGTbBNh5fBjlIUHoTHdozAHb5Og1pUiWsP1FXhySveMz3K1R5XWn1Vtfoesa
GNDCBh1lbwwbfSQ1AhUzZ63hGwDoTh89buPNQWsMNySotirNML+XQwnM6/3CPFagWLZZy8jGbCFc
XtqDixohyyK4DarmLFupW7C49QhECdtHvint9PkdCN449C+8tkRM+9jnDri8UIyXyxjtB+A1vJ6+
kCCR9JXxKg1H0lzZrKssMUoEVcLUSixXLgzLNMPP0O8T5hHGx8s48AtNGS+idVy47EsyQYW2XjyD
HUBUNDwgsZkPgOvcekGJQC3/RaAtphXbVzZ9+ulCIH/ch7yaxcYMaY4fuDaj6/eL+dMVQPxO+mrv
KY1XD2zNT1j+Hul3gkpMH29AOH6X0qdqnfZXtNlpZPPHB9GpkvCc5e0xHQtKHXCWavnYNvHuFx6l
D/abCeKRm2/r+yGmomCyj29taf/TtENT0ShLMOzbge0yM/VTN0/QRHdjlYKowW4ELjel1oVVufwF
nKHvOLIYelosFsGF+Hiaci8fak6Hukdjs1cMntNMCbT/pu3r3wIo5h8gjMQoAPskeMHGTEgx1gnM
7bWK4JlrU9K9ok5V63i3EtqtvSrT19xNoWjHBRq3t310L+1k4ZBM3yFLMpTMyCtMouZuPJ+DrtgV
zQyDKJvnsHC1SXFQViFeoFNSFiZNZz7Qytd9YwyWUP+yjh++gUqKY5V2nFEpfDb5xUdUzGDpCVOJ
1ixcKKbqkNzIqtVeamA0fcOlxj80WqIKz6LYL6ld/ddStcr0LDEWefJ0OL6TcFAqeLZQMFwkTJC4
3A5Pxkr9Frsdsa84XGcHcXOtmeKIq1QsJFbXioEDS/zHjzFtTJebtn/OgTchgjMVcIglq/DhLvX3
LKuf3a6AefOK9FqfmQBIAov/cHtQbnK3YBCura34le1PJSVVTk6P7u042wQlHx8LqIyionPhB1K3
EUPCZV+MoaBsDdPQqY4ZfnJwh6m/xC8u8jQI7IkDWUhUiGUCmVVcILWYwgodumI1eoNMBP9Lu6Vs
UbvIsTahHK+Pgl+evrwCOzgnc5LHoF/Fq4Hm0V1tvuVUSAktwOVqpNwI3ySxmHm0WsVn2RUS6jMx
FzdHhCRVhsASZsE/tOg9rjInvnmikwtl0MjmI6A6TuxNwH91qyJCWxbZNDILdSt6ectWO3SUHGzM
PdC0obiMG9Hf0BT8U4HJ7JzDMcUqjfj6VS0n/oX/6kgkV86VcYUHQDpFWJCaQuz5+wmQzkygESVl
BfvCA3FWhHQ1DIGNm1Th9o1bbOGgrmHz5cgUNwxKuJX+0ARcJEXemh2qLrRT83OzzFZGZoG36CUj
t9WZIDTFbhiX1rvand2d+piNCdzsRUsHyo4nLxumGTdD/vJcJylqMiInng5jmuJLzWDkWpAt1/yk
1Hbxh1NuAykP2MAj6d1RtPDW5lkczesqfNteHL4MTB9+O5MeRfemh8oRzXk+YKvhDvwzNrmmOh8C
7qrTGHVMAnaVSYChs9LG+x3ZRI49bAJum+xAJCrxgWRr8+bf+pBVrZbLGPWoP/JrPbmzNYZqM8kh
aBoMrWtMIqoWdo9L9PUr5oA3dvcpqUNQXc1YvprJ/qXIZOGUkcqmkOCl2nxmPZRN0IA8QSmJz2uP
ySCQ/aXfbGAvU2h+VGq2eoIeulMhOrjZpQcllR3x1HLGqH6M8wypJWTrLCu5aFPHpxbF2CtI6pmo
qJK99DGJe6XMP9y+HWqBkAkqyf2lm2cBc34YWgsKS5yGgbKp6NcVFBAJA7wiPiTo79gKFnD8s9Xx
iPNo+6LqbfiDov/PRP9BO1AVI5faBud7+313CMzaHk43GrxpYcVq5A2y+YoQLlr44aTQBPpFriQo
wVwzXG8CHYeYo7OeMgZz8JzyWDtg5MBCz5ReVQ60IzVZzt0NEr4/1keHa5QkqDeMus41UVyYj02B
FrTcBkOeZr0SzRroOB+2Wxt8U9r+0wcXt/VQA3KleyAWQQu3tkxcqKhBk6W7WodT8tPSBTnYNkW0
qy8/lefh74txMDUPcWzCx6bXNw9hjGdwqKa4jndjGcmCT62yqv2PVe1dgQJx19RfxLSc+eB+kOWW
Qy7d9yGiLIE+p0HH+iXxmzsutA7Prc323DbDmIUor4EWC5rH/bsjWDeiYOxbe80OwXzG6a+YsdP5
5taVqfUtYScOkD3enHWoH+bZrfaq0IK0Uh88J1YWb2tJVpmf56pwE6XB8a4gUR4zlFrKUEpNHP31
JKxFBmr8y+GWre1d4dZ2aJpjYPPiKNMbt22gA1RJmaIINTJrKusu7t0UXOYATBwtwxkuYl0dgO9K
4LCuwt4St50PYKSfIjfIUTr3Bi6FpHtmzPl7RwkAL3YS91MkluxDfuqJ1VQiuJ+eXUV8bxDDR0JQ
MvKpjcS+xCg7MrRrOCzEHTNjxPmV3RjuwnkoueN7+T/YR0kLSWwHdr50u/EvuK6hY8AD7+22OtfJ
4J6g+mKfpRObW7iSC+39IkDU9CFcjjBCNXllx6HAiK5VMqh8IP+EvEV+HRpVquZNvX6R1JHz8wmY
kUns4mUDvBkvTnTLh+3oayDmnr8YyE+BCE4hkNirSX3v48bMRsiHK0+Kc/NTPd7BBY6dE5uuP6cY
vUHSCOUvBEuwanoZ4G/rDR+6NsszCbj7m3zItQMKp5yF89stM2rTEbyaXwFaTK0A5bfYHJhARZWS
qsRd3UTqdbVzmswLQWD/QIGsJdnbaBZp24zTQOEa69JrXcAi0JsqT/eFAVI4UUZOI/PH5AfCt7ZF
St7dbk5jZUaQXlsui2NCk0960OqGZkWT7jcywtIvOaguxin11LV0OxMH/JbbyZBfh1hWStgLIkSt
bwtyRfXjefI85lawViQCrcKydwABo1IyRXRYsYqNa8w2Tui3qjXS/vNxeMbX/f8Qbz8OpFrvuLUJ
3Es1X4aGC0bljr+E6VGdWJ59AfeJyejhDdfaT5wdr+x41i/mlJ8/kBZqUCxW38qAceo7P9Hi41Wx
4TGFYZfevh43BvUG0XXnQm4OzMU5wUpBkXqEiLXIThpG5fFVh9/aiYoPVgA+rSdzc+oZaoQR07Pe
AG5Y19BkiQaxPHLvmyhYQVOlbIDN5ugrjxrz1nRDb6ZvJTSDEhHIRTcTkDfOJkUxMevY44wq6T0L
QyTFkMjgmKMfU3DdsC3bO0VkXhBGTb1wiB7A2S7gJB9VbJcT2yFktNiz6grLQCT/KKbglYrdfpqv
astnbaHrsj8I2RuD5ueZNLut+pVBvW5r8z35zy/3Z6sg38lYup8oGOoZ7InFBNWE55x+YzbeOZl6
cbsrY9DmtlpiLtQHsuLZpVg+cYKr9/L2Ml1tQ5WsjdotIYU6qLftXv3sMj6VvQl6Lm4vwKXc19DN
I/PK+CHkABR2AXYjDK6vIIb6j8tOp4SU9ZmgKhWhSSM/YSWDxas7dAD9UWn94oNF9vwagjGaK/HQ
0Casz4+czhggH8QaNpsNDCQWMhikt4rK52QKhhaDxUAr7r2LpVo228idB7DFnsydNnXcd9VZeYKY
pg9bvybYp9yIbK42mmvrIxOOKGI6YCBcjOYDQIY7KH7zStdDz+j13ujPdBrJr+nS7HT39B0T0C5m
GshxCUQ644C/wcPgg8Mfx5KvnG/sp0D5dONHyOOcsXNxj8grM9DPHumjlNAw1kxFt5oMz0B4LgVi
q8VQOJIyIkqjlJ3py54+BgIHTFrXdfz9d3cmHk1fwnoFQ5U3lptURKHGStUhW+H9kCg04z5GYtSk
+b2W4oRKnLCJ5eM02Fp+CmcgfPmcvU5FKVz7S7TtuFBSNmcRtpfztrTRzKEC1vRrt6E2j2QTQyAf
IO08/jWE+Ls3FNsP5mScnc0beq5A3lDoWylrasGR7yxuNnu4UCXxE2v5bhP5pfb75HeYgtDQYEQF
cT4/AlNrdA1jMl77w2p+8wGvLL2sWBW/qLahsBHAn+JZHzoxk09i+gRdBf0NASRl0yZ12KBQWiii
EIwU90t2DPo4pHT3EE3ewgNmEsrnes9rPAwCnTzmqxJau7kumEcJtfJ4H5N0PdsKeAGSuf7gJ+YZ
w0WnOLIHUJEONhM7DefqnbycONKlO51J8MhTuZHx1kHfs0/FOS4sUAR/6yfraZl0XVJdlH5k64mK
xEfFlq8Fx13TgxpNT1KeqyllQXklr99wPlE2NEmKZA+ixW/LAVqcjoXQEqCaAgJUEmap3E79e3tm
ijG2fkVGWps+bAZaJ8oAdpQlEFjWNrhWJPzYfA5LpPgUw/u3q7UJEvYl6DncD8EPMnzZwj30rlcP
mB84+/S/0XertBXU0A0HhTJky0Lm03ueP1idPLENZ5baCHZ2ypFYhrNJnEUFbjnN8xf+4km+y40O
lr1sO33sDmJneDqrygB63583eNDvOg3B3fv2Hw9uVwJkoiVon2g0DR4+fx1tDdtrhzunmMupIOSB
e3kQC6qDx2ovZJPNQrkNYA7rRtj75Q//oHTd184CkBeFu8UgkXxGwc7UC2Us8V+NE/PclMIMdDmX
VodavTvP/PX2mNZaKZxc5eOMxdLv8XFYI1kM0cJ+5A/KEXstL770pZsCl+oLP39+bI+JB+lRhW9u
mprQJZgLDDiO6jfOXjtLuJCGZPs1zkW631y9QXbH8iTP/CDBsmpE4NOTURc4oLNwnCV/hjuA9TnI
fkz2VoeFvTUyciJNDME2ANYt4U3t6vHXlV5Ot6UQ22Eb234ZABHIEHrfI1eIKZpR3EZYJndP6ESD
St6P5SQcqrxgN4zxOJ+zk7UIvlclVeg568pG0ivR/4MfKcjITOPQ0UjeHPxnaiOEA+VYnGWHSHay
CqSHoLd5xiN7GEk1uuDHuSSweYvuiRnv/6iLv8yHyu80fHrvFORJXPbxSajm5O0kaDnHq/RZumwV
bgzwKTgUuCFcjdqkvoMJUw/eI3NNNxFTnOLfALj+Drmo968dGjJ8rMwViH2cna9/Hhi1YnX2Wreq
IAEUn3Yy8ohklZobL1bziRznM8lpzLxk/TBCGBsPcGJK9rYj/MmewWTZY5NyIXuDeovjXvwf/bTH
kJLCrjT4Vx1Zrl/qFNPi1Cbjiuw1Q7NKSWxasIB3J42NDpICWy/uYLQgoxRWUsvZwcFsbR56cUeX
E//e1qClDMkG5n0gT7j79HwdIDheVJ+R3/8PfnMA+5uJeqJtWAa7wZ27jWYsvmGa/EPR7exHlQev
FwR+lk0UKv4Kxorw9D7paSKCcPb/wp7ki90EfcLRh7d+id4zRiCPANfpAaT2Hslotl+mZj558ptx
zsPyc8o5HRkAeH8+2I7J1FwTnj+G2/D11O5OUc92/2aVwCQAlQlE4ENEynIYNWBINjQ4BOWu7EhZ
S06MAVDMlR+sa1YUFt3wVljP5aPK6wimMznHRlA+4da0i9Z0Oz0fzFkuDpOFHpsN85B26LseegLu
13alYVW7GpXdXuxmpbCA/8ohB1gniLy/OTczPTOgB/UJviw3Z8sUJYLXPKn+5BXpkzq6NqNpNYyO
EFudMU8CSn3LPjTv0qfhmgVljRpenMT/jg6f/SlStcdjANCUkFYemPvWcUQ0ZQr3VHH4pl04H1Yx
H5ZDoFH8ZJtMwv1beJU3AxVbAcaFYaoH7I7yUEzgPUUfIU3YIKf9Bo3K9EAhuzGK0sgg5r/OxiZU
2/mWEpSdXIi6C/zDRI1cCwET41ZDU4seF5v15JkKb/cbtH3YUL+cgxc//qKRp+posezuBdhiUQki
fWeb304DvIIRwmNay0K2Uk+Lr9+DcCHFBEr55PGE19trKPoagICQhmTrFxvicF+fiC9FdU8YJ33M
DFhzHwKL2HimU63BjJbXRveplItNB/5LYl4vkZobAXJa6t6RWUyyjARya+95Rtgc+/xlrjtdemIe
4FPdyoyvpTCFX5GUaxWtcB9Z3796VZzmoMakP1sO8sSCIG8oWgGac1D8pv4WKP6wWvr4/7N8VGYf
sipEqOLplTBvwLl1TXpPjITFHc/ZTgQ/P4Pp+9LZsBtLC00fWL2TsKTRJKV/6ejpBWUV/w48ivFr
PmpIiDeKxoTSFbxBvVivV7TStIFXuTIxzt4OFh7MmdQyAX7TdOh7QFJXY8CkD00gHqUw/lwzZ7lT
f3OmqPOaqnPMcyAqUCvIrsvHpjUdS+ws5TVOL97Q6Kay/QSIaLYRVrtKtIr7U5Pswgd+zUlkofyv
OvSdfJGRsYoBuYe6yQ2Cm8cHCut6CnzhfpRQTSFcGufbbzIsCFs6nydmH5qfB5N2117wsiIkpmjz
nT8YjafkmfW9v3/qeEy4Yl1b1M+jnedb9rSbrIKE1XcL8k5CcGYcPsw7MCXn3Hpk3Mn02dqUlngk
TCbgQcqddVtBqN+aCY4Nbb0VytlguS2M3V9AXPmzJLFqLlawR+comEJ1Obkid7ku+8fXn8cANf9l
iWNv2ABZYZQ8H45tlqJ73JUfNMP0p5EYdT8zJ7Id94Y3i2/0nWxvv1ERwFEUS5UdJG28RDPSwLTg
+fes/LoQegbzzDMWQ1DrJDYV7eYE8m73tIf4FdqzAM+7ggqP+ej6gwRMdFoLCPRaaaqSoLm/WKJ3
7sX3aIYn8FRg284nazLcV5TJ6tb9LBXVwhINYLxCpjum9QkOyS5Zc4cPP6DJzuBnPjBX5pSxqA8i
NtmTKS8Oz5vSy7V908xPjKgR1aYbu9QtG7AYz/H0uN6rBJBPjl/1Kx93ITsK2Ig7j4IFgDndAUv9
n0podbpzfNdqdvF+ZkOkcIkQ+vI1L54dlYEgQ9g3Bg3jx15/0B5SFsEkM3WcFJN45rGxp0o8vt5b
uGHxvVyaPhaBVKJ5O1ZH7z0ZLAIQLXe+JN694L2NEvSnq8KSIUNaB0aZtUdygP6IdZNMZEJreBC9
VyGiAkN2IlAavHAMcafvKIkqF/VmRpo8jnwEKEfdSr2IiICiP34NBLbVRDHDSq9PINP5aTxXqoU1
UPIHgr02cVvrkginq3s34mF15tSFrk6/9qb6H7RnLEiA3D4OmDtjPXmdqkvnh8sD7OdRmtSnQBa0
LHsjDSmcdnpItrDHQFbm6A6D8EFjkpvFL0Ebl3caIaQTVVAb3u+Os705A/T59O7HUb2wPdkxZXIh
aaCKtyPaRWSgzUUSxLiHcvHdzQ79CGCE+hbe8TgEmQAqmYcKOFnWLzmQE40osVRzL7hkKtaCpU0b
vSWlGL0jF3zueRqNQSdt3pwLJ/VZLQpXIgYrkRxJ3uOLpqFLeEeVEnjOxA8oK8qyIWAmKAhAcbg+
MKKU67yyAJSG6rNz7ftjwsQlF3MUJyxSd9ttSjvJKfFPMLRoKqnnkTXwdU1w75/mlOjXokoqgEK9
8LqlV4d7VlMDFvkpsiRIAJaCz8PLm1AzMvTaN+myhOhY6mabwzcaTEEHm2VSWSShMkpNfKoylk/N
TarTYdFwoIhviLk0FsBt99eQ9D0yUzYdaWcmT/0EYH+8AfjajrveaWNDqza8UgmorWfWoj66HKQH
mq26eYLfwiKgtVj/EN4wBvIJDXvkAKck/Idr0Jo39rhfzTrpA36cqNRChnfNVnBh2hNVqVp4NiBv
w8PZRx6Ol1mRoSldlY5FYcuuWdU1zLxIj8iOnDvZuVISLmyn9DOEJp8CzekwNLlaSf+MsZlvub8X
y4ZWuI5XalmqAlqhWuFp2moRuliMJmn0RI4cLZSM66Ii5Yvcqw70YVL0VMZmJ+kC6vRNwqbhVmqI
VoeQaWql1YJKUF8DPieBVj9oqDbPybZUQjVEY3rJya4XqsmKh1wq58met28N/gzLp24xzT6PKsxv
n962ABptdeHyReN/QFAQp9e5r6iJ3kq0JB6cwos0/6yyRGCn1cBZqAW6kDdLpyjWD1o6XliPf1VM
OFkRwYDvcSBFPMSFTRwiMH3CZVJqgHEhm6vVbqT0xQl6tUcvqymjF9W+MxZmzBo7Bk1VRfRN6YEx
VAq8cHltesHDrILhATmN2/Y7GfRHFr29HDTS/CYR9IpjkV4hVDpfsnyituBknAf9vOi9nd2E3GnA
9mMilg3W5nERv+q7Y/fZbYvQSSpqkMOix68lba34LUTBQESnOfN76pUG/Yn9vB8jTt0Y0JJRu1BU
Uhgair4z8vBUiRLZWb0EqxNhQcD8+3P+ltnpCzmCxOyyToxucS8nJr1kDtLp10HSIUBgydCbDFSs
gzWjTSCcq6cj6vnu7uhK+HGNJ23t/l/L7nEnlDDNQ34TBth0Z63bNzKug3LUJ9mDrPsGFSIrpHeF
cCaXjChSsFFtRBVRzdmSIAM494mW7a2JWo58SWyjAPVdP7EDU0ZIjyu7tqQD/Cn11aB/dDaPtQ1A
NY5z6j0aJ0LmNQaHZjpvS/Lj0tl+XT+XFOn5zsCDEmJ/W1SY4DIuLEk427rZIpzxxUXPyETHFNws
cpDKUd8jXCC79/xrRKUiLHsQpvouVOduvpSZF2TFNH/q1EVeAarRl0hVvWTY/jKYTqB72ZwcNoEj
tkeYKqjdKflsNh9kRks30K/so4ifuj/2R7YQ/Nl2EFRjpjD8DhykJ+Q29ZTcVsr/aItnnLpYZ8iQ
sHLStQfGpTGwLD1Ow/uUj/ZjcR1OezviVWhWacFVom8vfoICvtcuBWdkDUrn1iHcR3volKtzb9V/
/t+56gX+Nky2Vif6IjjpdJKHrC00dmfR319tipTdsGv0aliyvXRxJIMwIiK7M2mdKQ+OhSQlVsXQ
1pK3OqfVNDOC+xvc7jnDDVwwPpiXYo9HiX0OMkozAAIpQmx2LRHKnrXffrlWswZDS+xRigaPBAql
uWkHPl+m7JosJ9cOSEFdTzAhX7AWVTzAY4qKDUFZdpLswsRiH/C23/6/cmbFfSCLbI8k+5m1bUDf
NjV817xNMloB4GQxC28XjgOarzL3FcJN0k9VlNNPDFM+iZXfbZL6jxLrUqHrj2D4gHIDh5Xlt1qh
/8yWoscdOpI3Pbm3AlN/huHTqmIPjawWsNA44ClZokjY9HKuQ/tLk79Eziq3RbaDIKVOOvcCXqhV
JzJpKrF8WxiAPPA3U5JraiBvW81TslXEwjOZa5KOLzuQSfWGvfiwyeSwDK2EfB71oOtxa/+IrRhB
Ul262t38ZFF8WwhTUyUlIHgs/JhGYWba8NxFEhoJ0nAUDexF6revSkdtyclJJX0HIlfd4V9Dy8VE
/w5KDhg4ADvKKpg2+5B79hcgl6qLOI8ZMspCVC3isrbAJ8UTbuV423OUg0Y3qgdV6OxryeQQNE9X
f75ph9U/KLiuimDDRJca0dLFrv2pxr0tat0mqhtdCfF44UyOfH9sLBofsyal/37KEiHBtuEFKQKt
Gt5VL7pSw+uWWOrYwIwI3usMcRN9XMZlaN8jYbFVlxkQ+xDyZ5uqiADE7WRRFvF2l7mO6K9NHU6k
uoQVx00A9pvtwMv/NraTOzjMxqeVVBBKTzNrL7pOUl2qp/6a37ffSbhXN6KGmilrQfC5DNRi3m22
dJPwnUktMjX5dg8AeOrqXB8xx+Un/29ORVXkMzUZ/p0RYhfmy+9AtqqLEg4jG2zNGOMyxEZ/CGVB
U1SZfPKEmHilqHd8ikZ2I+ASMrYcIYFMYM/fjWFtA0GUW+7TQUhpzqIPylrE+h5tQG6h09u87NVg
nd3SJcs04ihVMyz5Lc5G8lsgW2YgUbW0LJoOXJXZZ0j8kj0NbitOdKG1iQGLdAsRWmalEJkso7lI
nXoSFK+/5UTJvdYAbF3JUe+Af527pbCsXvQOflLJo3s9I2CL1+yraQgHgAHPT68GVpE0gI8ntU4Q
tWavQJv11x8pJ+bDrLwTPsgAc2b2KyribvG0cSOWme9D8Tkst4By6ex9F7KX1f92v1cejM0rw5/+
OCcN6uSQML7dHGLS9jvGHObTUtg4UObhtNf65kcGzcbaIi8Pl/NzV4hXN0lVzEZahWzTj54zUHpC
dtidvgMFRxElhBrl2QMb5ojTFt5F1wxsTegVnfPdn7szuR4SzY2LI8gYko/+wqsR7Nu540ww3LIk
psT94VHWsibTnkhtVmPaOPmb/C++wC9qCqkoZLomxPdkJmsqh2NE48wb3I+hQ+/jMgmc7BhLgYDS
9YkXPcoBjy0adAie1/ipHD/Atib2PbaQj3mCJqrcJFaAqUiyhClHSXn1VKLjYISL9j3n2NgSUjAC
vlq1288OyiA3kLcsJ/ZH1pRS3Mbt7wp4FmGqOedKteW17qI0Mu9xQ9RfuiDyPa0XaddURH2n1muA
rlT0VO7/0/DzlVaMr7mZZgIiIFU8Garg53Jp3RIvY2rXM1DpzOKgGmmOKy4iUkI+uu1Kio7DimMz
MPbSWeWfdt5DKIggCH9sGYE/omUsSd1ViQmUHBGTaWsz3TG5FQBYC/zO3TtSiKxeIBLHV+1V8dRI
kmHGWf8kaF5krw8l+VV7QshFp5iWnNJ+YOFJwSTIkLKrfuEHM3rJIAqPLqkucFpaE62th822Cjjd
KH1fI/CHlFamt7u9h1t/zqRATSDGffnvmUKp99Dd2AkXHJprLJFecEZwOy4i2f2jqDFDvGVsnV3J
UXPzuJTVn2ZrJUPGFVZrIJF0tKdzq5fJRX1M4770DX1gTNiP0hq2ZVp0gB3Ssbrw9bjoVi4xZBbQ
x4QtNRNmyyKHcQN/ySXRmQapj4nQnSPhKbZD5d9P8N7faOHsT6JAYCPIpkE9/zxPDqunytpk1IkB
Wn90Q0jw8OMVNTjPPnSsssuhaLgUIHmpvov5zb3biJQRcXPAgD6STJTRRD6Ew9dtyBn2PUb8eqtf
OdU9Sz42BotVC9C18ojvkFtFtukNZTlypaVk7pX4Q/QY51tyiN5Zqa21ChhUQFn2HRl83G3ermwZ
oQimpcFI3fzMHYMp8DKpcUWC/EYFDSnRD2+lQkbSIK7/kMwFDOrBUonOyU5jgTJg8w7gPfK8lpd7
drAtcSCwSE0ge722FXs9H8zAanEJ7skXVK0FCQLTaaMBvw/wCmLLb2y1cummw3vBPuXy0qP75lVL
+Z4QGoDqMA/PhrretN0YxDMUWDGGx214z+82HlUffFkiJNAUgdAkr5VIw/TqsLZlQ5kgKz5khlKm
txG/LzCjOoczDq3d35VVqqrF7TFz3o6815CPZ7H32s5BZVfI20CClmedPUsMpTzIsHmdgYJMacWO
bUNHCUUDp+7d3vxHQrSjHllBLmZIg1bQGCQTZlVeaTCmKhZ5kNM7vBlwotSUcRuHSALn4LblQVr1
xeRBI7AHlDfCzW07V1Y5oF2WJUI0xHqOyV24DeeL9w17eWecbhWzsEjG20sXbU99GeEiCKS3kf1P
016V3WiHLMfMLwy+V9mzjLf6K6vcZ3gEAq13VcWS5nXk1n3yAg7VhvgSjfz+eVqGA+Uykp3x5piD
h8jY7QwEMvqtN4PXmHNFsP+86k31s2lGTgz33PYDRPK2dqdzEpK9qJKBiXtYClntg+5UODV9YHlM
JBI7T7m+dtIpAc5TyVIWb14QycMD7MBQTQqxp8azedI2xpiao/QjI5vuTiegQ0AQZ4Fp4DAr7o7I
L0CrJDhtedVZUDO+JDD/msLeZfsCGeMmYW9qcBP3abrSEKSTVfUF5tycIEf+rfs3DN8IA9+tgn4G
auRxJ0hVpM+gqlq3vDil+u8NMHCVWWI1Yw32/2SGdiQefQhix1P6SFie/u4gMwIrwb2xPTO167wq
9h9f8ahLnZhd7WdvSaN979G6wQsHuhmwZ6/jW5iaRWeA3jUWV7fvgPVrUNjaigHN2eePVCqBjBdY
BNSU95ygmrQfx35UK9cWHG1DQmYMDt48y0n3vJgAgGp9Xg2gUp/DVGszPy74rOxuxAIeGNNXHOij
4Juar60fM0Glkp6AL1a+EJeCVCzYTZbV/INViMfvcuRM3JGmyY9PkV7QJt3qO5jPzNeLYSDJJmGd
tpOWNIp+v/ptLP7LXtam0sAF6laHXbbP+rMMcC8iNFMY4aJqax4Mm0xttfaKVJMKLeuP+/9VHGlR
TKyNfp9ojWrdAcvmGgFAfaHLOsxI2b+Al4PmI1N8Jrl2oQJzQS/bnExgUFh3guN2r4WsEKage19W
YfsWw6tjxh9norxB2oQJL69SNsl4T1+52bZib4944aIOVgPAwGuedJBf27+mXpE+2Z2OUdrbbWdp
ntvM72iLKuf7/ISq8io4dscTrkoHllYm341hVyDey1/wjR7lpUb8iitypUpTISg4s799OyxprS11
fd1dD5qBEeC/wN2tDLz4v0ZSjc+2aEzwuOlDaZXKPvxG3rEN4616EctIc4GPGvXihsTB1Mba4mFA
6/W4XdsQF2HFoVOAurkMVN9ihkPYe0z0WaYVHRSIRr10VgMY03+rgzZHuf9sSACltqShJtSUmg19
L3urrrcyCPwnEq1a8ujaknWiBosja8OEpEsCpN2GjIcA1Ayb/PuIGQBretMLWESxUrBuOLFrKKwx
RSUBe4fnRRjbdJDGfkUD1WPwKz/NjNBfx3ZqGvgwmY6y5GUb00j7ASFRo8lPVGG6iJkFqsTdAPfg
W4C9nJJ91R1stmdgL+4LD9KeUG4DreDddSagTuiQ6xcBiHB2N+md0U+rx0brPhkVC4nHMiVwfgve
F7eXFbZP5HFQGajeFtoHAJ9s8ZZLGy8Me3lwoHY+D2WUTOU3SMIFE0uw6COKVR4pabVSiMLVuL2S
gj4e0H73/r+4MBF5yjbo7NcTzaPY8dkeoPu78upICnme17h4BYlig8HeScynqTgs+8MImWbshXNh
HqRaAwJ0uVE6GT+iL4eDK/DSOuW2Y9GN+WUEhyWjycX/cQwDmGHBABYoEzMhzuY6SUBXvO5VFprJ
rXkDbbgZrpEstuFZWty+2LUiqdzfLI2Y5suZpsvm3j6P6cD4nQ8ZB8Isy4mp9elEHD/wv5U2f4+0
HUa1FP1cktCkFoF1A9gKh6rSMjqymjznICOsoLFEyaEgZaMWcohvcU5xvRDZpPTTA87GEUsMQJ3T
h9V76WMIZIMn0gWQ7ScGxnJk3+Eqt2X7zKJOWLR8OMsbH3YAj1lxGKRqKXCeriejh4IHyC7k/F+f
mT4wcVJyYa2kW2ztSQCBECCtABqbWTTYsnpQXcVX3cYtkf33igKsvortz9ydAXm2FzIPcjX8C/gS
BSY3WJlRVUl7aq0gl8rfHG2llVJMEMQEexyBnN/fuRetAe7MLMcb7v91rxcBMqks/CoFAQJVw51m
Gcsg3qx0R+YUf9Nar6enoHY/HV65qip3tewAS5Xz0zDxOcjnU5oJiwmDu466Q3Xk2W29XTyy2tNz
maaNZd7lW8DCzId7ewaJBpoxEHKLjotH577vL0FkIdfMb8SdoaG5al312En1hzEnKLDIOf4t2sml
KicMHTIlRftZZUmZg5LZ7yHyPNQA686ys9MvOVg61ExoVUZkOOOTs5R39sYdNlmqSsqs/4j4D/pq
nUz8E0luYXkzQAzWLdtersaNEJOQzxe8TTcuVegTUqzQhilcF4zLwXPe2dalzUG4QxRTHQ2WB7M3
yOgHN+yOHVElDAymmBGS2OdOzBJ8OD4Y6WKjt7eYna/qiZujuy31iXnX5V2m3otHAwr20Eub4T5B
0yTNGPrp4hhGzBV4HlfVNSPiIyH6O7qzJL99F2BqVpvLPm0krMXr8TGfLrQpELouE9KLnfCG6fjj
nuwvOVu8GW8BsXvVkuIxuypPIcllOYhHtc9gBjX5XOR0hBlGIW7WUof8G80AJQVBFi1NJPjwz+VP
lHJMiH7+iaauE1m1h83YnGlApescr0nR0Y8chOWEUs9aR9dld3/w9ktHZ14Q4F2audb3mtklHOSN
Acjy41ph2edW95m4xyf1DQi8eosmyJfUnBxH1Lb6k3ItRxUVH7tCP7Tx64vcWEQvs5ox0li2RJzw
wCkDaibZ7Fs30X9HmgaetC2IHzmlHVoHf5YtDtbWSsrkZ+98OfSheZKP8J9YTo8zZ5r/YOpRuEyx
Uui1mYha45ZHuI0XXqOReOlT0CMPa3ytgIyCFlBBJsYeToh5z0fESBH0XfUrFfBrfc0eV4LK2RIH
FBi3cvacLtTLqM/HK9LwXPrEK43xyoXcx8c5s6qB2Rh3LAoPj+C9R4vdyTwzcgkyaNgZ57CWxe15
OfLmX5CHJfwNkmZjBMu0mQ0FoM6p4paX1/AmPJjue3TVsw40i8gerQgBxLgksjRhGmZ/cx/eOH0k
ovkie4Oo3AoKMtC9arEGQOL8+Q62MmpIm0ObVecaacyx9v7GKq97mOkkK6MK4WsjU72yUJYhWvc2
hvln6Vpp0P6zBc0csN+2BINW5HwSMNPmt9Rpa4N5FOIGtheQ71JeICFVyRSLzQpruEfToC20oH+n
cjt9i6OgNK1t0CxMKZZqWrV6puEasNYFnplIigrRJX5+To1h/GjzDQX1X9/O6H4x7fFF1lrpDzIz
g5Xpvu+M7EcnstWavHB4+ZqLpKFIvPm/xUCstsL1P3b8clImDsgrRy1apSpaNc1zizMzOviscWQa
4WF2SmI6ZyaDlVjM4ViD8SVrqqr0cVZQUWM5miBZv9qMlZHyI3uhHhKIbF4+W3qzmwPySrNzGiOF
lxSPRTG2vh8/ZtOEbFrFDqU+OL95uAdDLDu6BNy9Z6bNwTdygZPhcFnywBS/1x8QiTTLo6UB+d9X
qfeGNoSoGaNnrsgdlpjNEIe5kEyIDZT5Krqb0Y48Y/ajuWr9ZlAmBFBWMYZelIumauy4RuMbF6/W
ofSrOlAy2AHEZzq2AP/0a3dfGNGaXnoJVA1icxYu6LQvlrzq+8a6Q/0QdPFNlXI7bH6GDxq5PRda
9pqqR30xdEA+EjkmwEibFZHXsotYiuaT/+hQiw3X+7nYXOClS0j3DeFM82IhFQRFuVpCzdnUmd4f
rQrslxuLqh8fw5VSW6bhWtkg+RPYO3uTNiSlgn1+8pwDB+Dksz3to7/4jSeRhBLQE9b1x/wv14tB
2W9kH6q9ACCQFzHz4eYrGuvwbXHkiHuhjE4OJpNm0dEmmMvkhL6SBgCbtuBgyu4Fu+RKjjqxImg6
FNb20pQbHag8IUI8FgY5+C0FMjbODzZq9XKg44y7Hf48dO5Jh1gW9onu6lV3yXSdrggZutyYmphE
+UTLOj5RDt5fWtJIM/7JbT6RrK07LSdQLCStVLF7oGkNcXJeUcorlCzkIleiyNe7z7vRHgAzuCKw
Tv1AdxhZ0ZURxyThA7+cr5PC1M05+8sqiGQ+ywoQgQaO7Oy4mFvJPnLUdGvy/HZ2RHC4TEvBBoqT
QOyQujGaB1iUIGYBYN3mjrlN1S1tlmyQN2sG6A03heLY42kyZ6VuRyQ1FTQfg2emGvtPUsg7upki
yCxfqR09mG+xqtK98cUf2F8nBlUWptnoAA1cHtnHsenjCP8W+EnHCFd8WxxJbbQ/WTsxAQDPpvFF
yNV4zZEwFPWlOxGHxoHTn6S3wrykMYMGgOSyJfJ0U9jlt4va/pCzvrKous5SlngHxeEm7bu5BEtX
NLr5UvpgkudvvWL5x/D5DZZEgUfmrNuKOoXRklIhZ+lqWbzJo6TM41CyLJNSC0P5C8cs85MKCCfN
ZdwxNH6x4Qb4ROE+N6BJgkeoZv5Hk7aQuSTzzaw+1sT6sFzY0tXQvteg/Ea7ureuFO0OouUn1PIC
XVS3X1LdiFq+4GVhrgj8+0LtUP9stMQAY8tfM02J2YOnS28EnR6HrtXvLYiFBZoGoOAPH9NFLoAd
vk1KNmz1iliHpn1ZhoX2Dar2KpizsH/ZtJ4gHSXsTD9s9HfY3AlRNFJNmhDA9onxXdiGWSQCB849
MMd2qgvbdDY1DdBRz2xllUh+MipvTE3YgTGeUm2HHuUUsyjsVHhY1qHw0wMC9Pf/Dor9A9KnBdef
V8YGGC+lZ8ItHLymQxYCjtzaN5CtgZUBcnlZsnTMteSp9pyW7/InR7t3btnXVN7CVlZuqh8ZsFCs
ecAzs8hY00L24GXHq6VxjY4Jvv4vkaEdD44bKPPENr0mtvJ64SqesXEC65NnA58debDFFnCjvfEk
96UUNdmVCCi8b9SfMRjx4q0IO5FumID/IKXvAAgzLaIXSLEN0w2GHbWKCZjWLxg43XWmywSH0aPF
7/pFJ9RTdCVkSiHRCMPs0Sp7C1pjYFWAPwi7eOYEik4wJZIJ0jEq/WuAnb6Xh5uGacVyBHQ2dV2a
5iXZEZHE15RVJIncoETm59krFBSUFDL2JazLyZ/BvvVHja/WrzfSkm60o4WAqrZGtBpNqXV8o0H9
y57JD4Fr+I8Y44qHNebN14bdnsGK2ukKOD61h9cISejyORketgNS6SOBETYU7IiVzFrb46ukgHHD
Ly2zHbIMbJi3lqjycz5L85QMpunQd1MJGVLDHRDTPPvEWwlk6PA0lYDZ/97HKxU1XVHR8uyEl5PK
ecfK37iHUrQzX6m0L4EpO4O0WE2ObYQOo5zSQcDVLsFdOtBi6XfYpztV27Tze/R3Cj3kC5K3PeIL
k/Wb7Sd6n66dOfc3v2gyMdtsViQDJz2WGpj6PRvMvkmngTfsPVWXj86BiYR2t1jtI00wxdVikHdP
VYm1uTSXfv5IdlQu64uxwmLMjuUrN3af+9AghGcehoVTjQp4pLaazrhBDoXPo77dNYAE1qLaIDTS
8IZngPClrJ2PJ7aLahx3wkNqjf1PmnUY5xOuL0056T5bk4+DWi46KD1e+b0NmXI//OgdWEjmNFwV
Utlh4K9cEEisJiEA66jPAIuXI0vIQsWdyzXyveZ0knwGrGuzH93XIQ7WtLIP6SClkWcepaXoCLoY
ULJetS53vSAg2B8mQ4WWZggKfEceXi5qRqqyvuhNiy2q+bBiPAYmgK1v3vmTnuzlkZKUuK3Dw1y7
ZVVgoa/mVKzB5y1xxs+zLEGr/paxHGid31ukGEtVoEsyUxOLdfVxOYtv6aBpJ2SppxYHYD0oCHTk
3R2+rZugwtum5BmCYITnvPHxBmvY9AoZR9oiDltrMnsQHtAjnSmhwmwwwsC5DIHhxryB7xWynjtS
Mbi81Wsf8fWyz/0K3dTChhyOLrbQ5lPULJAA/f0LXfE4OWYB9E0N842oyGBon2oTjD0Cx6kg5AuN
R/EHpsi0X8Rzb/Flthcz73IIwFWOrc4dU+ztNYeBiUd6xKWmKMuQP+xsJV1BJ6F7k3Dz8HV6k6jw
H0/mYgoT86QFPyteE8ulThgBr6vMOw41zPE2OfBqIAiyg8HkAqzrRhWqcBIaJVWiwToC8kFJlnFg
WtiYfZNMT6PMvtoqhBrthgj1eJuDyR7vh/LjEtKB+rxsrZAhAAKC2ISMq+acP4U5zHAoojbIyFvS
PKqM4ykNrK5Vu15L3cPjxynjXQ62e0NbsbPo3zmKEKnhHB7mWkGwOMNhtFhfuF8R6zm0FLyDix4y
6hLjL7diKH0x6/t2ow8abkJtqLcTJ95hTEsRyezO7H4M6YT3ECGNDnbV1OBGwgVb68Ncyl9M3wZN
FIgcnseyJ+wP71Kw9rQfjlI1mO3XBlwriBANSvoCdBGCmg5djdfhBMdcKZR6Xhp9Axm5yap7kp82
vWX01pgPfAvyGccleV8yMKcnkSMvpB3EmvZlKqQk83zmQhenfuRjz2ma2bxKvpyU/j5DDEUwI3rV
cYgH/Y8Ul+EtWLeS64ofJuXVUp6AYFgXmUp22rKG5rm0Ju4JmjwzvFzyzmfXXV2j3JsujCq5/Tah
U3nzk+pmY7BxBOj/QbbNdwFnjusWjg1eZXu8VR4SUoysChZNxQYn23wSofg4OgqAwASHf8ckexLo
mBnCsdOXyHsU+ohuaKifWe0T3AEO7MVp4YNHWAViH2bIlIghXOxhrPRnz0xiEVEGUF5Nn2MPlavK
xwWo1gSm3zsVL1a/6opvfM7akxaeZ6p1nGKzqheQE4239HqyqXTRbe1Uhjv1dcjtbIAawNjlhbIP
U2HOaea9chz/JmhOaztaoLO00YaU7howDjcXkiZc+DYZ9MPGm32GjwmHbRED1SlCE88DGcRhad1q
eH+RkoBFoyS3fuNjomRyorlON0a4Fk2y9tsahU6OBB26tcLQPLtj9UtqnG55If1NbkoMycFFtscP
Hg1kee3aNo1hNEVhM6iaj0AVqeWw4ILO3f8mm70oxUxrlqcgjGj9t41tJdyScoa8XwFHnei2PGaA
4V710QFqrOIhmOMHikb0FxbFwMdZmX7tzx5IEvj6W8ncuBeAjAkLqf4iwFepvZgJb2xzOs2aN/l6
vj7JsZE/PSD/x6vaAw1XoSNWNvsNOlba5yxWuKqoOTzCJps8z56IACEkQlVHA/zkDlJ5PwmMykH/
uLX4AsfQ7wqnnRjg3gD/aD3VDU3oX2pFGseZ0OvrkyV4a8rLYNlrXgyMgf2/VPZCw5knyJKHbVcp
u4jMrlXbyPzQw6UTgagUBwdmMyI0JXRhAZGR6H1Xdm2M0+EX8vGk/n6nxGkfmME7fLu8P/6ZjNKS
QONbo0mAmTA0RpFFHEc0aUVblkpQEchsZdor8BLdYe7AezxeZN+HES8qX4WaW/SjZtSdpFS882Ip
sGNsWmTW8peanzj9vPgsMtWt9f9IzDSxGPDemzsCpMva5bTNbhVVw6/C7kd8SMMlT6ZTZ0movfox
ch2sNqW/ZMWMFyL8nxvB30MIB0DEctrMKK35Uz7fJOCvEo+QL+qC56ukpg5k5kuj/jgczl5qFUkM
gqmqNb8Nfs6xTKokKTgiYcVdaogS7rTXsYdydWuqA6Q1Pl6CUZ4QJun7GQoV+MAeo+egb2kwhsMy
zmkm4Fp2xmbyPHYyGPwauQAmgsmnTTCnfqTRX6nwuX/6ARrkqqWENdVdgWYaSO2C2BPuNHNRupCk
rkAufV+WP80oaQTBuYRa0AyKoowA6CYPHcVIegonyVHNY7Mj4FFfuYeii0hnthK6H5V2rQYX6NnE
1nhjSwzXLUPe028HiqNROK7mLJQZXW1RciK0BSPlrs69e39TdTfsEfRjwW+zHJey4cSQkj1W0rMy
j0LjSl+ylUyL/HyD+JfbLs1xzKTxkJ/mS3bk4TNqO7OYgFrNO7ZBfHIpctHHYNurDh3kJKdgNWQc
3tOIj4Fq+Ejm7gy4j6fuwfGaMMT9BgUbj2OBeMLFIqhfJ5RmaotLJgVPRJ3b6QKiGyhlgyh9y0zX
5GTfjLieJmuJGve1738YNFdnKubSoU4N5lW/2VwB7vlkW0uDPb9ZpFKDbq/5qM5RJp05iIf30+1d
kmSFyPE48BbrcWEHYXOe2W0kNd1JttJ3o7fQXzQWh5K4mauIXPoy9kKkyyS9j+0CIIHXWZtVYYRK
sSThfzhINoK5z0odrzpnLI2HobSF8RIS1r8Ccy9tNTtk6VEFcMlPVbSDdRiExFdErBboCpub8jJr
BCXu/6ezEw3PHmKWJ7EpsrcDXlvPlFZwNgmMcEg31ssUoXWV+/RiMSk/Ptox0+jkA/A0VVc+bpJi
Qut90K2NgbYt6qBKpsl4rP7g6maCL6wUQlqyZXQO8k/YgF8oTL/EOfdR+5aqmRAwJJArLNFdVy8y
rTMPUBVYHKvvqCo0A9izD0RCEjL8OUeDtWzxRb8TpW8t+bauXf7RUGR1p0d3G56iMTl2mw3VQ6/i
4T4cW/Kp3XeYw7vFNlDdElTN/mdmdPD0u+uw7Uetb10Fr33GzXE/hJys6IEhBm0LKxURv1TtU27Z
4Yl6tvuVjBAliajjgPJy8Vw/bipJ0xsHpWieBvGjp/lq2Ky8BaIbGi78afhroeYzLg8No3r0V3DO
5wPkfYG18g3Rbu3CvUyZVMZm8Tr27VSSeBlphEL1+Ym35fOxlWP1nQ1dDO9TRrNdBKtYhkzxc0we
nx5xotSZHo+6wt1jjrNQbF1jRgQ6wdR/0AfP45oW8h+Ih/SBLisouAAAcKHY1EIyL9YoopVVDuU3
eQAtsmK/AEI24V8wbARbhFdgfNIcHG8e6SG1rEb6Kwqwj2u7YJ4xyatgkf8HoSWsGiOUjNZNYCwG
e8wLVxNKOrq6BPMBX97MnUvrnxx+FzCe0X5OGpi3SVhgr+lQuc19L7BCHIC29+/pk2qexhsrKm2S
XL9mwzOcUIa77bR32qN4bkYezNlksTOqcZ3FNIJdrcia/T9SnvvyaO8r/f8RrtxPm9wnph3YPAF8
Cgj1YAL0vYeXGwffZQx2iNdhBMcpYQ93BmWovIA8W2IgpNAGgUnfLTQWcktD6fOLwaKUSt7xPua0
ZgKzCZZr3xvuk9pa8UA9eXgVxExTosrRcVU68ubufg0EBZGxpTRO//HSNlAzLjN7eaQmNzKwdH/x
9o2rIM03oiuELhe5/qBTuoWK+zlGR7E246pXAuh+7DJ5XWeeNPdOg4zL8/AEtS+vOwuus7PEQWOp
2gm/987IEI+hgooX4Ei3BVDv29pXDTGuZ/1t3vvucLbqxuuaZs2lAjI5jOe2WcojG5vkIT78SDZQ
BG2fvcJWrCHOsFBqgfbfSiFiWa2B7A1y4i6xClj05sZDtTQl/5Cuw6MqztmaYS+v2GxU+1d4FRST
8UeQR1Bc2A5N37VaTiHwBFQwVNgXveuTZHPo6l+YpXinSuTVhi+fgABeDF+um12+0dZbp55m+40Y
YYXW+rJwUpA5uQSYbuZRRKchM9Jlesy43IQQqsRNsMLKdD832ub1CCUJOYwlYqcZYSWMO/BYgBAP
Chfp0rlvREAlrl7byzMKOqfhtaq3hIM1hmVaJskGTTqxPZ+63hK40yHFEfcWGNTtix8p6fhPfKCq
NaF7qtvBtlB/DJR/BvWVQSPaV+81N3g93rrb96xsM52mbUTFAPU4SSRRkVIPnqRi/91i1gb6XmdN
gWCnEKQHglnt595RCgXPdrveii8ufVKSRPZ36VsfR0569PAwvCYhyy14f6bG3zpRyKfaARafwGH5
1FvPMBHh8Xjua4fZNw5jfZTax0B8tliSBRXizgbc5rfWdKN7owYhs2VDyWnx3NFWIJrXYDc1ZxgY
1dxMfmuBwj0fRYArQdjLocglvVIpDp3I0Rbi0nXFgibMQTcsI+0yrvXQ+MshR7FIziqkC7oKbo6g
Qkf39RfzNdcvNA4mXCoEXRd2sM/bRXPCJ1QiN1v5VGxJWqrGL3UtbVAXk/PBGtlhnpzDW+R7q3Bd
48JtJY2CAdsgIchTlCZOTBfYJc1n1xqfNzwP51KG8le5SR6sApkeA29aUcQccD3Bg/1sLuY6k4tk
gevJvEbWOtt+tkDxgR6NvkKwYxxz4o47yZMU3+p4KaJrhDpFKDfZqUdts67oAp08YLui/Hwuqa8d
EhD4dbyzn0iYXFodsimDcd0Ueofnb0ElAySch25qesrGcaEoGGPzn6+NV1FRoOv0xNov89rCNXp1
eVbQRRzHzttD/FDqhgjSUxITw1B1LwvMwOjoKV2TutaqSdMxCSZswUZufdxjd/v3w8v17blllPcY
k9wJDm96RgGf5/kfSNkW8moumsOEFdIkWC4tEbeqVPsfHI4aiTjpGLojtFAqMDwpcVqCi8LhVVTt
Qulw+bvLTudO/3Rw7M5Kg4q8ipTB+d1rvvAwmHBYnGoWiViZFOf9FCwwCw7rHzIea7YaXz3i6xJL
QFrEZUJzuu4JSne24yO7K0h5L3faAFvZY9/ji7Al7evBtpdvel6ci3TSR4gToHasZXfhQRHCd6Mc
xtQWiFAUct0VIkEfIyl+LrwRfd47A1gVREty5M8xa/BH6HRUzbawy7ghUYZ5DnGJKN/6vL1tINS5
vVBC1y1c06tvVWR53E670axb0IggzCCYDsaSbqfL6R44Pdnf4J7wnObH2nZioMz5fflqnaVrsFte
uqJ3yxCkvqKSd9we4eIm/PG8TMLTmhNXR/YSgIo4CsTnmFBjuDeDBSN6tCidoblLUTPPtnHhSGBL
1AeY88PVXpIvx3upoPFN9DHDf4WVadsjrbWfKnQFHmHzswQCLi7pxoIqhEzc/8d2lHX5Q5xQ77+N
ASIpHDZwWN7jmjQUleKijoybReHi7Wp6Czr4hyW1T1AyyT2O6kXYhHBFew8fDS8/JbxH7g7oLJvQ
6FHSsA+CVHtpp6sDKyv54aoc7bcRhmDigHN6t7s3yX0P+fJa4vFf6hJHR0uF25e+30+YOEFq26Dp
A9OUck57tqtrs8pdPr1pUfVY6YZW0QHA8MwtYMragSQs7zUmw3sStGlkMrxODZvK+srJ5FFfw+MU
jnJrEFEWl3wzFm65eFRjv+KK1IzB2BISt7WCJZ6MjHtazTbQJ2VDz5YanBqtSPEhRvM3QGFrIg0q
fA851F+fivQ4bWKh254neSy9javgsOYUzBrCazQBFdkteT6s8Gmq+P945r/HvQhz8A26VHrFGbzu
4ZOtDA2ESb462wpF9cVL1cKQuJpNSt99H+OUfEWciRpmZ1dV1oOMsgqN+lfdjcjn76AIngWoehrE
Q7fjsRnbU9jTyvE2/Q0obCUS9nbeJ09UKBQuOTCeF6/EPG8dq7RrPA53lQUD7979lduruTIYE7Dd
MMMfNjSM/j8xyO9zu+fVF1dtA3aSikqbrAXWszPaZb3TrW+m9Pvd3NL/GhNshlPJNmz13CxKZCsh
Ep1rwrMg6qaMyL8HeBh11/jUTRNgHfifDUGZiYBeOqsyKAWghYek45I4Pj4RgYvk4uEH/uKOwgAc
hgTq7m0HjOh6HsXTR6NyMyLBClFBPXmGiDzqqAqBn+XCUbbYIP/3oDCJ9OLCkKWtYI5rsLmIAviz
9oSi0nLP7S6fEZScmfliYJc1H977NSC6ZILFri1n8Nvx9eEGfUv8Yo5Nu7Ve10Y4HMkC9/nl336M
MyUr2pEs4ls32+PfoTZbibxryMmUi+adzxLcucTp/JO8mBypLR3FdVyoKYOyIZK1qEuVNT3jYCZb
b/2ElCuN4zhW0QGZ7V1hJX0Cn9RSJ+T4b1CM1CoPbM+SjGBNp1Q17QfeKJpOjR8t1quB/4K2IuMR
kWODW6w0aKZiyP2Cqn0qM4YmFvlhcjogyDzUjn/N91AqmLtFhU6DgdG7dO5j/FrVxu2UIdE42Lkc
LO1heDQtMY30M3/7vSQw19AS/0d7UPmbg7oXseaWN7Qr+49+40HJn2jZAI5sQXpBqYHq94RKQgtA
kKltf46d4keKKSqXhCAGdaEg1jf4i9++9BNW0M7+ZjUZ+N35Y3JdF1lyrtL+aRExG00SAOBqlP8k
g+xl/yyVhSsHG+VtqBafneTY8TBXy1pMB5WYOzRbMo3kW/h8Rd1nEr78/CHJD1BTpn6ZGNM+TVL4
QeuTo6ZtfElbEGLNH9pI03jgD6zJ0dWynN0avCa7EtCh6Gg93npH1uMDVTk2C9H0kU1MvmWj+oZB
CqXg0Ro/lw8YMHhPyIRz3QW9qtVpIp88RTNW9YBvE/HwbIdtWa5rNlXfHu7jg104TL+su90xJ/ux
IV85OjPlOVdhBuf+DxPA/El+coBZPqvgSRrcKlz+f5NnIlkkkHle2B0v8xIQpd5UGiyI1+dafXNh
H3Sa1mg3Xw3dN/ung3SoBoYdmlbNrFZ3yct505NfMtGyYXMCFScuALZQ8hkxCV72fMxz7d9k5vMT
wG1Kh5xuPnsh5yq8TQ+KYS8tE77XT5l5S3wA1lGQ7wPV2Zc2Omip3hEGNmabco1jQK8UqK1d1qXL
uReWr/NSbD+1ldJSkpUXC7J+79VfdwQTKL9/7Q7XO4jN75MWWYCoP0v2c2oxRRRbtVPO4cfyxh84
GoOeiXKKdgQNjYfASaFn8CoHxyXnqfi4Yimj4Mu5TJ/XHcJR9pCcXAouMPi5IxAwqsvWU5iBs0Eq
vyaRxqHQHzJ+gdjJkdC+ivnP+1V/GOcuA4nA2clEq5W1zaONINgeAiR4pnNY0t7RD9rQMHGQgWTR
2lNZar4nw0g5TQLqoYthvSOCAlWadZ6igTfEZX8F+IpzGkC591TaGJRfox0F514+4gIjhnC/IUZD
3QRttkbDzRgt+lonH+S97Wi6zZp+Jxi2P5zzcfA9lNPOFovZMeXekHfLMPda7OBN687IA+nVNNCq
b3sQcjyVr+/L9NcNMQT6GAmXt800n6KIHKBV7yNhLDdBWlCa3WAE7tgc6Swnc2NceECuPGbqAbGT
a4hAaPuS/ORalaSW6rOGTD74d+lRvJVE/eItmBIFChfN3LmUKds5nOASWNDpQHMa1hmX6v1i5cEY
bWCjzlyj368EnuOvK7A8WyQJBq7m3BFDhcAvLsyVnpZYxQ1L4z7+UVmuqpRxjawcDxHT92H3H1Ye
YCRhw+2ZMJ9DdVdVqnRBjc31pagpRWmqqwGaLxc02LwyvB27E2lOqTkDpVuf/5ih4EStt5L12OIr
e04dylYbmTzPc38H3Vbw1OZHY2X8PREjbKPkw6JEp9THiHdtnz9/Uteab3U5wPF8qYvP+L6rpl8U
gX7+R3EG61zNqpV2cKVeBnVXw+fv+s3QRIQruV2GOe2GQL3ToeT34utpykkGuVUneia18HR/vl47
/zhqBegnX6jQxydrjbHCamv9ZiGurlE9QNmhcW4i1Wy9bgNZ3aLga3ATVifOFPq0+NKzu7YlMud1
a+ehqH1g9zKVhDr+rXDCKykXbxNg+2b39NrIYY5xMFImvCnWHS28JhPragSDbAU/GBnZiyIe89BH
rn1K9BXl7jUSga6cIxl/FsohCArn8/xGmHytpsJNkFSzsf8blTkxgwCWEFmXDDNQcvLCawUbfTEE
YlbSVzdgNPZENkiIoMiOAohxrJB4EJNO26BFwiXnMQNa39HXYmVPSJiP4FL7BOgE9Huf3VI7jV/6
LRZ0BVaMIBJNEl6fa7wGZ4CSaYIiJ2Wy7mduTUF7phn4DgV543d2b2WT31rJX1tV3zxHYHFkH7jn
b3f8mvS1h6WBVi4SyaAAwy4y+xvgGzbqfBJT+fLpwoRpu1LzCGlzvCVedDBoxT5QhLoDhn++Zlb/
Gz2teA5qnDaxvV/p8iZKlLAl4crpumt2ZxwJrF+LE2SW7PZsB0MjhOwrNzaJ/g9SWPmPFKfpAeAq
YjliXg47zt5jUiRawDX0JOrmbCoAiARHY6nB5U4k3vT+jrR9YLh94muOkUqyThala+LzWVyMq0jo
jpF2+rl/4w6iStrnbMrN9Ej/szjcTe6/O2EzxxhA7ozXzs2nBhI8llapSbgjv9/0ek3vfN2txaej
SpzkaECZEeVrRuakHxHb4K83f8aZtxBaPrn9PfgOEcmD2+jeg9SGz5Pnu0/E5dBZfRqPIAnhk5gG
H/q9neCKDsRzRND9hPNL+URIpDDHOAT5WruVtggNTyI0uxgpxRSEqM82cVCeKMl/HIixXTcNGy9p
WNre8gOTNXXF/d/6U+Yd6jyM9+8F0lmy2+7dbOk0j62Za8RUHCVLRRYPBUO18dXBrxVvtpAj5N3a
8C6iCLteG3KkSSBHbEQBKsTm9J/+f71PDzVxve4OoYRm+S45okgQsm/2arDdye/Yeqjr6BPSx4BL
lcR/AywTt8kfinkceFghA/dMKTkczSZVrLUgESvnyAN6FnCaLYy9mnidHwajcsJLtDqMdxa4Q1ZZ
gCBqnLiEIWhy63hKiUswwkzixz0SWFgmonqUwfoHL1Ue+zYRdY9XCwLNpKaKshWL2h/H9c+3F5y2
vafWmF6pC0qEdBYAm2hpTM9X9GLRGYQvdVi/MgAuIezptqO3W0kVddWkCwWwmi3UoipwsSXH0/9a
f1osFGQOKx9HO3ZrAmvEx3n9rML7r8j3ysx8sDLzj5rOrTWdP/ZKGDmPPFluRELM1aox3K0EJA6X
kqQ2FdMZq9JEGU9h+oLEZu4CnY/ERhcPCN7vMA2q1evdrIwtPF5VswxkKMYwhQADjEbuVMzyRaT1
d16OoTj7bLqi0F3NlERkJy/EHbg5AjPf4OelmDMM/2Mri3Kip8D93OFS2RiwBOLaWk0tTkD/j0Zb
GwXH2yuCo8+rDsTvvqj8uss0eAEIaptn85gna7cxngj2fg/xwVh8CyVwWZmtHUp2nMk9udRFjVP8
KaVhXII4hM9DSQ1I0uHk5xrnO7nzlmOlLQQUFBYdzDcGTkkFKBhJ7TBeE0x7ltVV6U9gERCgMW8k
7fb7NXE/fRloFe32BqDa//P88sFL/9WJMS/TLIuazjI05MxqO4QPh/24dQU6fveLRNATqxyH8fqq
GMRc1h9HJvhg1ZSmuikFDwd5a4IVJ+ULrDsIkYAglcyCRflyOCncB04Yr3WIbzZg3RKY/O4Y+xjU
eepD+ObtmP/QCAxPLwTkyQkIKtyQA7yDJfhPIuuUV4QVgDCacA9tocArs8YjHeeZKdquSaEPRlqN
MKyIOBz4sOVnhE/7BF81zW7ARICmfNffVX8X0k+szcCMfEZIBR0BhtJkIek0PEDOHK3t+maJC4xF
Vpb+l2q6cPS1z2YNfAIEBzxZ1rwRozm5DPR0C5jDRC/dhdFYb0uXh7l9HMMeO5SBCxdOX6jsAtoA
4OGn4YZgqdtclQ0BkWaPhMYl2/NEPF6PoGLLZR/O+VMAohg2t7qmMTE4A9UdbQH1zwjLcPHeOZKH
Z2H1FXfPH4/r129YGlTC+BJJ7hu/MeecQHBcvmGzN5y5bBQxAV6PfWcDJiyaFIlmEwc71EyoC9Eh
hHkjP6Fx6hMXIWmBPOVbU00EHrOF6/O23Y+tARNJfFiJWRjDdp/RVpdXaHwCFhZ56Pu5ZBjKEto5
KEXPav52PNr2k/YdgYjpB7WYLwZ9OgQ7Z4B5F1uUGykhz3x7g9m7EEF2szys0pCWdgoPXKeI8NfS
2I3V9sWMxKsr4eelZr1GQb246uYBKUUJGddmApOC1jcKaW9T01cMLVkxfFQM9lhai/LpeOXUiQhr
5fp+AG+yzZDaxbV3vV9zXAvG434uPMCvYt5e2E9GBrPwsM7XWJp9cVc7229BjpUlkNNhSr3Z0Kbj
KXA/9SxGYQzoyY+Dprc8JDw1GFTOgbpryeWgPoE3DWqBEeP32xWxaarBvijmG3QUsGCr5jHSfECt
LfOKaYBp9dPr0uPJR0AkT3DAHV6MMqt0qAbfTTcRf/Dlbys1HzZF2uVYma8JqjN4dsLzg+XZ1R/+
LsBa5Y2yoNKBDaI+Nnl/QaGWc5KmgSgGyDvBqSQaXIK8skWymLaVgu1NS9vJqABrnGY1xetUDFPy
dZsUQ4+Pe1vDOzmlYrBEx0Jh4kcRtxkq7odvlyb8krNP4/rN2iBTaSdomEpjx7yqiWwMMSCOXXw3
EcLHw/Lu6Qr5JRUJb52O1XUSS0i1MsqXxCh0kvtasucMnifMXGnMF2l0E61fl6SOcHkSeJczOB2v
ZGW1xCOvyPUJXtto4v/app0zAucV8zhWzRvIvKz56yptyQzUV/wXbLYQYobniE8V11KETLj0VoYv
kyn895yWDRoDdP9ORfNp1GsI/hcNdPON1VNh6COVHq3Jp/ucX2SMu1MtapgifPz4WFLszHJbnsOz
TMIGrj60Pbk0v1jplbO6OEFwlArOobW1BVXnjEczNxzUSMszrzSX4Zl+barEL1g4o90234HdmCI0
3S1D3PFLA+jm7+xXeEVGuHsmTLdxT+5sdeGGhZ2zZc+HH8VXyEm3H7vyRC/9qtMBwEhWbMQXRma1
dFiyw7WAaKxSlCV1rwVo7DJ27t/1SPn6/0i7n+EpfinkpFh1qHP+JZkwFaY8ayhTQaeiG51AxaFG
F4h6XehO8JGGne73tSNOqRO99eEuIedNLzZFmJQWhK1wnoXCEr0eFzXIOhvU22bkOphecxzj4JYE
A85MFAVsRsgncusga9nO7tEX5MbM1tSPdnqIxkq5YNH1Q7hR9uC/4Snv8wkBG5ONSbAJIgy5Jbdr
8lIF3t81uP8lt/+rlZb8cOfrksT8Oqz9FXMLKkzrdaKe6lHbuZlYQ+StWSw2itP1kCaCf7KRb+yl
lfENI4PM11rDzSkjc9pyZpMv+sU0xap3p1dD0aP0JYGICJfS7TyR7YyFXZ5kaJaZF3fPbs5yDXzu
KA8r2yLOX7KzcBSIbLPg363jkMUzcW0CI0cehRZP+F4ZzYia/KnN+5AIw86lFjFCTN5NNa50uwHp
+AK+W0DqfOqZlCpBNVTSDZsAIBS/0YtOvvkUBHZ2FcFzr8mnSG5xCS/MSonTbgfuw0jLlB532+/Z
TQBK/vc6QYCMuucH+k42EWG2k+fel50oZEuptGd7hJgG1DPkVZ2PZpFzDHSImgFcUNUCmJwqE96N
709aMPGkYKdc8GcqZfoRKeZngFiN64aD1RTWY+KD9MbejZ+zamoLBNzW5pKjo8zwb4s66X5w8oBD
0bLtxCbXd1AWlVAyFwtXlK8KPhcjWzxMPfqillkpAClawIcnnqKl4bn2KLTAPGlB8EIjy4OntDHi
sZ6wvKicUuja3tZ4DHeS0XhbesUr6UbuMjNxvezH6lymz75iAx1bTqqmEZgHUraRA0Jyo3avTTSg
bZmdzvRS+qAKgGzgbgJApmNFxlayogOgnFlsM/JYgZ7+ACP052CaYYyQby3iDl7nYVVAv+7f4xCJ
QVkXrSoQBhmHPSK6QNFuMISSkK3Zhk/COx1P/xwdIC6UOzZKNCwuli3w2mMcTWN6tO25mPcPDe/X
rzPC8hhGPglr6Y8CsuDrvHFZ75mSR5UYuQzHAA1RLC6/xYy+cRhYJv5aYbpnnfLkaCMAWkclosl+
doXnx8/V7Vtj+CRT5ND7JYNWyIpc6ZzOnZrYYpho/+xxneey4UrepftekWYOpMDvyyZ+GFgyzXYI
68ndOVa9SUFU6CtPjjSL4PkKwpV0LRehQDIbH0FM6EBaFvzojJGSrOmnUIfeHe/nkMDC/80Lw5Ar
8hqE5Gu2zysUf7HkxzCrTtebUOD4Wa6sEwKO2gIvFoykjaUlhEpm3rAf0hcucu4teX9saybtAVFf
ZMB14NRYy29b/3ZNzK8aq27JWi8hGJxUpPDB5vNYySbQmT6iz8RCLIcK8I+vWA5ECOTPuFFMUld/
U07P9gnKLm0QKcx6jUTU8sTf9Dgn1GA+n84NGTW4IK/ZIlAZawm8tfKjd75eJk8oJdF+hD0YwbOa
QihRj24kmzLrSmPfLVDMcyDliKGOBjxOlV7yfcg5DKmNoHTCqy5ziFdVihOoJis+GFoc7TNnaIG2
E86AAbcFPJVkTrqpz0AnNBt3Dp9aCp3b7Qoev5KnOSAQvLoULpTNfQAg4hN+/c6MaGP5xhS9puiD
PmO6kiCBHDZdoUbFJiNOt+r+ZrhLPnOv6hp7wCbfvI3bHl4SHlnB8w2KdxpldbS36tzK1rqDc1nQ
p6v41X8VKWKN1QbxFHi2AqUy7o0IUo33WVxi3ZHtj0l8193NobdRkoNqBkpYPG0X/Vnyntxr4jmh
Sf9Fxcr4yWmx1dvZhmT5lCZ+MkKmcjD3fFggc/1cMC7qY9tKILWTWtLCUHaPnruisuhqtzDcwkWz
/Zb1sk+fIVvSsGEjv8RJnM2NIBkYkYUOPmn/6s86T10Iunnd3m/fSWraqr2PhlCJe27fzqeh6xEG
FKO3Q1ntQ1pkhhgY+YyTyWAyx33sqG9uRMe2egxoWMvCr1FMG8CvndToaptLNzToySLA6T93V2bW
8rlZcWgswYn05rHJuotFO7xMZ4t8rXQ/Y45y9pgakGqNEQIrWys6kuxbH3zuvy5AE6xO02Aes+cZ
ef8flueFqK5Dw7EhDfK7tBGqb0ID/+lJgjthhhBRGTVfYEO3EsFQ9LiVV/fj+bCoSgTTXmKsfnFH
r8adNmE8QTBtr0bvBXlEzq1z5fGMETiPaQQ+QvdPeIYyNvIE2TApg8MeECT7iGBleQB2mhaz8GJO
MQGgIvCjRdm5E/Qhf81CLTDBA2Rs2hZVUNaoH9PYjZ2yVtR2tiJF9x6S3WUqq/H+kjTUG4iAeKlu
WgktvzkLNae9hINsG5tdupfxnqJxcE38u1QXWMtfrYf+EqvduvTmsTQOq5V76CKNYFWuRbF5Hymx
DxK09s4VibwVl3yoUr1V62gthcmVtR5XfKn3zOND8y5akNlETTc21W/W2a3/B3XKd0uP+iLXTIGk
2qVlezx7JPoasiST0vqGsHDgAWYds+X5tNraj8JFDk8OKGoNruuPmHUwLUy6UwHqCzVXbXcRqzX9
XhsUSVrhnS8ufiP+ismk/fj0o8Y0A+TfjWqRobsoHWP080RQMbtuM7N8T7fPpmy+klqr54Zeg4dD
6p0sBW7xhIuK2W/Ss8OTygx1S6ZIS2GB+VuRtd73S5MSAY14BZyQy5oYxfpyzZSPB8YpRVKWksv1
Ir7AWkxuT6H1B+zkLzBSsZbx1zbUtLRnL9G7ThYv079QgOJ+2Fo9SRUgYjvLlqMvybRBB3ObHwJZ
LdCmwkge3ylZwN6lKef79M7fVNBY6m/peSI5XuVQjy28B8YYSbgMWKksDDZz49LXMntPBqVa+aSu
eclXYh3DKfhFP02FfGThoAUPkpk97nbqVUDhKASM8V1gNb3HBMpNfjMMEbEilmgJsYwsw6d36CRX
mQ7wWJRfHA9KRaIIlrm61GUQgJTSstQUxnG6e8oKS1bTpX8rQHABCDrPN/y3qD5iIFSMnBppqhBy
IuVxoeEQ/6kUD+0q0dhWl/yZ4I4fQJlhE1OCdKyYpaPjaHHhvIXFKCdYXSydMEhIJRtls7sMw+5w
WxbJah1i4Ph5hjnuRRMia0d+ipN1xyZPDRYgxBxziiXnU9fLFmMcfLptRtzIuCjFeEjtOwIHnFb/
UbtiYJAs25CMqM13GJgsl/ZvP1mDtSTyvBbADqG4Wpnr8qdpbwvDardOOlJfK5tustXz7lW6GE4h
/s1BLgr8ATxGJGMroUgM+BO5EcMCQPMTJ1iG9JgfAT4UhAM/KjDk3JKj7wCQ24jBj4u/uyFG8Lcx
YcXnRoUZ0QErOy3Uli8zonYOU0vcjVdmszWOpWY3fbdiVMAcskIqPVXVungm4FnFTX6VxhFnn0QL
9oV6uG2g2neVwJwwxMlZ/dz3utbwCZ+Eabk+dwNe79idAOjPIvizlHtYDjlm00bBxUgoMZFT1m4y
U+0ltnwiwdx+s5/kEDNxmuemoCnmnRNRlZYy09zWoickZSQsl2VHzxxR8E7qHpvoLSOqewry/S3+
xQwUABIqjDKz2Ies81lPZwDnMmM2sgDdw3EVka9ef6r8BriHBEfzm88taQ2lbNrhRQaKMFmy4Zza
EQ7VNUPAMdFQC9YrOffHVnoRxyFiRcrDFZtjp+elNeniSlekQAm6U6lTD9ctxHb3q9NS8U57Sj1T
vtBZ+f/ShjxRSrYQY+6N6BunJJSltvIeXlKTV8ndFe7gynOYy5CyfTvJq60qS7d5Fua8h4AUOo69
9iC1rMtZwQ4dyqO7xKNBBstFM27ByMRpYLdjAHvHGygCR5PH+19mDNsH6Lbh+HD8RBul1mqc9Yuk
2LD8PW8EjrU7zKl5eoZ38CVRWt34VpAiiDwIi0TTTyLGjceWpgSSgMlWZDhoLM4beBf40HBWDLjf
iIMBKHtauuXci+YfFFnMJUEb80SEUd41pUrwwfIH71dgAueOZVKbpPwsE2HJe1lBDZjE7CkGqo1N
WiKK1mn5620GWLDFg0s2UpBHFYewM/s/nRAw2mE0yHfWLimfgqPZVQwqac2cxb3RGZms6VX+6qLS
1IxoCWK6UcU6JA80ZlHeagpQGqJ7LLpQyoySu+6e9iyIMFukVVJv/iXs6hZFQy43YPOvz3acFdLp
8z4dOP5sRe15Lui7JvfOu/Unkf/5+cb6akvJGxDR4VhdkGrdwMgIVscbSEaHT+CTenKEhs7PSBup
dctmEet1G2SvJ2OuiHjBkKYvb/uT7EhWlT1BF2GyfzWQ4SVBlpWbQmiVT+PcHkGnLwEdFca1c7us
/g4FP29QUqEghSFKUm2qiNb7cg3DM6dk46SXN8NF3XRiVPuQtGpO5KDLwfaHkVgUf4zuO2mwRrcb
u70RLWwB7zIHhtrXJ6JBos5yDAiU+av4LLO1rypmBQMwklGFR+RIf80Orn9/XOsqDid10nV7eBBg
yLxypZcFC6i90vRnR1p2wlnAT2yTOpLRqEnoSRuvFRmjFfcr9gVBG+IcPVnr0FXErzFMzF/61xgE
Eajk8UEEQu7xxbIPPBmkRVZmCGtYmneOyO/xyjcjB0UvRUaHxX9tfzxJ7mBb48wi/2UzBFovBGdO
B7HMRvyoitLjuEXJI23YpcwapiPBrI+jIJOyCMApfmT3KtepClAEW4GNg7ClSEinyQA13TfL+1Vi
N3OCBfkGfYRjy8XYuWSwcEsWvGFArDLNkfE4SIGqZ6JDcIEsx1xwp9pTjPLWFKdRXXd1FM49MVUM
179Im1qQHo0hOn90POMFgTbrlT0E7yHj+CIos3OFX72b+pMLOPiLU3ZQajIUVfEdBQWDy5T6jRqM
yCXf0yEMUthxNVQaMkY2LOcfujB/tO+nsAmPGUvMmydQAxUGYv5pm8k8wtojw4xV2Wju8TiTI/e2
vphhvyYWFC2YiCKf5zPVbNHmSZMLsVN3OBmYEUNNpLV6XTWuwxgp3FA9MpD18mjdqMNiXLgmJcIj
2h/RLOaa6ICMIUFYGHJCZ9XNK534jsbsrkvP1uVJo4hsAQXbHj5O+OdlADhhUElD1plIfWDG2Nmf
ztsv2iZod37NZAJeIoJiC4RdNCL5kPcgS9vhA/UJm7L+muFT7jsY2LNqSbCgU82p2LOfK7eHN87+
vq8JTmdObo9LMeIjwM1hs3rNSKZi7fs7BnZ8G5Xqkq5zee/n2jtAZiDR0XTNhVjce8xhCwS+weJv
oK8XynS+dfd/Rz9NM3GpJZN9H3NfArIjmr/DsNz25u3uFFpCqXiL6EvZNHEE9mAmvwhkszBhqne1
hb3xteK+sLoLkR9gwcC73dW5urm5JElVyc2a3pBzcm0kzPnpfKso5nqgs4z4b+Juct4S0Orubzg3
jZMrv7B4/WlzxhvMIvI0XXgZKC8lDi8w/xO0LNiVAsRdW/CubyGZIfigjUvKEhk5MvR9zk7hJElS
8kD4vrW5qDAW3nq1zn3ba8Q85HgkZuFLfqorbWUo7lhKBNGNY2rf+9al9XvcqIUI549E4rkQ5TzH
EcqxaVL82IuuE/0/mlAeOcYFpApszQNf76vKn+f+ZBwVe1c5VSScROTcaExWMPdnkgff32OZ/Pl5
8lDEVzOVOE5DG8Zgz+p0HvCSwsBHribEXf51m9l4FROaSBAcVKGvOL3jL74udJ9mlnIrFlpu/kzR
HLMCvJUdhYObxJFN5Uk/WhcAHQa8PCR2Il330Htz7m1Cz0ncQlQZlXUO1mxeSuyJbiLCPvOCKchA
tyJghV77xIfYNc/zZPQt+zvzW/geNCQIp03dhmA5q8uhxxU/kqb/h4BCp9hNnqp1quEa7bgBiFyI
M6dYHczkSrhZq1LZq8lWSASwq6EdT88Oab3mxrKx+ma53mlHFGz4ZPhYzqzh7qOFLR60IP9gEM6W
CeNvu5iiiUfnMX2Tr6ZlV+A8AzqJe64kGQBj34xmEsprVlUQ7W71VAbz0rFcc1Vt2batmhBxIL/T
0+w/jqktOfBBC2251bTyK7aiMQU4qXrB7IRv0slS3/NjOem0B7N1qZ310+XNf6hvMN1Rm5Ujrw3/
gTmobsjmTS6mtx4800XhnbJ6MLYg5Ac4ZiChNpOvZjxSFCfVwTZkUzrVElpX0dh6BDA2EPCMbwn2
pd60gByvP3LJRWUzL2B2FZ8vB2YpEguoeKjUzwQgJuKKzeH+haTDecSaLUsiIx7cUaiKvBzCp9zW
urxcJ4cA4hH119oExhY4wh1zlEnhOPRI2QSXDHriuN4ABOCc8AsIjP540n4DcaRuhV/UHTSAKl/f
49wMN6Ohlz7IMdyct1bNmh1z7n3rietFxFKvgFetZCwgdA3E6H8WrF1MemFb4ReY3ty/lFqR7xe0
yJGdO8ilHJIOgzPQ1gZZ1gXPL9jIS9rffE3ig1ULpKdV8b1aWkDTQ0aeye/LkFXUWokt1+K/BD7L
N5arsGNjGCv9o/rvqE3eHPtlGwQCRqEDnpYrRpOidni01N+QX/C8uAVpHxiRN358WYOf3t5AWl62
ax68ndgPjAVUgI+0DJjb58KZHPdYhClGZR8c3Qwsf1hf6fBrFq926vPyzjISuxw9QZOw/xNPeB70
uMcab5f5V/RxrKHqiTR7EjLyWdLPPksn+nbcWW4RIgxc0OgVZy6MlmjU8NqO2yXuwCl5CAtEgBGM
raYiHpqrISfLfEgnB3kOTsWlEZXLegiNqKk5r3u2V65WZi+3d9nmHIfHE8F0/oJzAq+TDe7zg9NI
hqf0u3u3Mj3GpFqNf5PmhXGaJi8xsWOxr8Rd2OMRn1I13dKkWtq9gcXuM2DJtUKLWleDdc7QQjLd
sR9Rr7XzrDAmwmoSiyc/Kw/TKvcU+rYz7CmfVzrjxVp4JPKtBXi2iX8NQQUhJIgOKAKjyRB31SCk
i+tXrPPU7vbgmh/jGfb2+A6DJwv5tJhjF0O/LIJJ0dJJ7+uhbqxNhTslP2gMEru3l8weQzQblXij
exz7KhU0F4CvHxWv+QZ+273d48YxKqyWRPjL1SHhIa8Ezz0kM6lDY6JxDglLK0sp/tDKOpeHxDiG
ZNVGWrdKwqrYvIIc2BiNRbPPVf/68ry6qHhOE6XZv4/GhG4yw/6GSahmj11GzDiiorsiYGr0lcwg
ZRtNQ5NdQfZa1A2O2lvdnwbuyz74hChLvt3MtZZZf+eT5kXzGFsucBIVonKoEA0EDe7NXTq3pF1z
KTP/p+3l0lTacWj4iXnMt8Roqhw1Dq6ysqQNCBz8Nzek3Lxsvae5aJQ3nEhKlLhHc4JY9uJtbjgP
arCcsEHfyzF6rLxOqLHQ6WYqj/9fik96yFud9M1bj7Q5ewQsa++THWLCqjzSK0Deza9d+xGaCwFg
JxglltYQP03QzqaGtlb75Zc82voj5Mt87555aCoY4WNvslaKOApQXuFoYvHksAtIOT3yfQU6FtD7
2v5rezRhsD93WAU8yqORdheCUJje8HfWPmx3qHTOdZ8eLhJrJEOxZdzOP86SsFGjsyc8SsbeMgpy
u0QSmUqiw/jh6Ut1/2KbjslI4Ssn/Cadj1VYoRJMNbfNaWRXixV0aeYo/trZjnBHP9QsdhhNVGfH
N41T2mwcYFqkmUY75eorUCDzEMZ783RSaXq83ePDBUE1EyKZml73ixImrmHMkzv72LHiAEhPzQsh
wRUWnyabOhCeIyPDJhhw7zMsmg1U1LtBFS9WWivn6jN9q1gtIzKPKvXCsIX1bcpK8Et5Pm4moklg
D+wC0pKSXCVrO2whhGxrCDZVSyu+ztaOu/VOGS5QsmFVb9lIKv3GTBcD37d7SSgljzNlInmX+qnp
iewGrNxmFotiEzmcq14OhZlwiHlmcwUB9PyiKIFk/Aj1OkgR7/rjrElD1uIHFat3d6NK/JyctZs3
5/6Fwu4ZzQSxdeHSkqkWO7Pht05HGkFBjwRK0MkXYMgiG6cntOm7n4RQ40PSsVEz8J/vOgmC3kv3
awPNeG0qqnZMj8PqRWNVlQ4hFVMJ2giGiE9fKLbk9s/FnwoDTUpXV3Rll24+MrkXuMF1Q1vOZkX1
I10CY3lSZsl/cL51/arz2tKORkM3LHFNawtbvMBNhZFJhQzXKGDQr8lokblJ7wxSUzHARw1alRf6
l99JZyvHQgr9TtJ1x2E+vpk6BVg3ka4NnFJtrPFJdP/Z6TyzqOoTRPRuvOzBGf6UKqpTqJ+OSwQq
WLItE7TUySllxWhR8mJvG3D+5R4PxBnVYr7BiAdvbY7OCbA+/jFPMX/TVTwN278satWpt2mO06xj
4NQiVin9P/Ii4SI3bZuVl0x7hc4yrfG0bG/zundp/CmfUyrL1/ld7RGJbkqjwu7mUcqtdO1f4U1X
5uSyKDl3X+cL6FVPkoI0NKO0CHprG4cPQzOk6cW4IsW+YUfpCP+DaBoR6gHS5NyS7o+M50YVlPao
31adNwg16yUX2kmJJI8gFI/Hu1ISQkWAZN0puJMOOXlxNpCHcqqqMZ2hv5GfYhb3Bv1jypKwVUVJ
ZVCi6u9XQmXM08wVPmrUYpct0O8L+Qbk0+PeDG7jh+uAxhDoWHZb8Shoi0LX5jaGsaJjzFVQ5AsU
Jy0yH1EwWDYFHpn86ZgMCLL7Og7iKO6A9hCoNqUy3yHlBkVOM+l/DGyOpxq5Qe/wagEZq+BVKnYR
/hMHVpxlUIrjTCSaDH02NHhL/IDYR0yezULY+O3ALunjpzAaOOnMw1Nb+EZR/Q11vhJKBk2XmB9g
rMQASEX2Uz6mtB3gzia/73ze20G5a8UNJsJ3MakFI+sF0Um3fIzaFo3hYfoPo6njdAaUCyGixGL4
ZsiVkmsx3OGorbEM7A/LowUqG9MhE8Fg+ZkywyWpMVt9kFieY9pcFvh3J5mvdCOjEXiHMS+JHHF3
Ko1piXldNuY4RiDsNym8G0finA4gUaBaxkrzdPVIxdjInm7L1KIQeclcJVKaLk4yniJPQSq6IJE0
Xz+T422wn8Q5qTkXYWr4AJJykCOKFUuqDvc1yPEWg9TRw3+ydMNvsRBCKsP4ruQsScQV52iSMzPy
eEvJbKb4h4791c268fQwGuvtlhRd6aPW5gx8Ay1TcLXYv0WkqpCx9pLEjsUhv/lQDSJW289QePun
LVlLHv53PBb65bL5RGHQWQw/t3gIK4DrwrUfQFNmfilOZAA6sh6k1a/VcLJEaTS1HwATu3KXyY++
SdzVulKcINXt5NjKfT8HxAaZjgow+CBBVlL8KPbInQxsiX51Nstx6ojQYQzumbCgXN8UMI4zKTzX
mWgtSVHk9u+Gg0iK6nFbjjNkUUJvDLFabWRrfAhJM8ryRv1pNZZVhm3tOJi/IFy3pvnnYMCgKgBP
sw7fFzdWk3qC+f6/rKeZKozqi2xhY/LFUneXhCgDqZHJ9ux8LgEfacGQTQd6+zhmVNAwDimCWl3k
N7j77ROixfBqCYhTjtoOQSC1Z+F+PfUgR1CY8YKOygWD+nap1hczlTLCctR0evp/LmLamQPvQqoA
AQFTgYcgnpEZku6JKHzWoQGI7nyvGn0sMAen0KAz/Ww25FR8iMNB5pNZx4S6wsjojFTm6TYyipVg
BwpLGy+Hyy59mB2U7APLu5W30QUxshmwXDOCXTgm+8uLI4EmBmtS1Or5a7PeHk30REMxQO6Dck93
mZDDZ8yWtRo1lJIOW+5jpA/dt3iqX1EI3R2jqD0qM2xWpneoHcuTQSB5b5PmBlPhzDGNSOyYx83M
lGNVRWScx2W8vSdYN9MWttjdU4/gi7WFB8rML9SD66R0Er2d93QM2AlK5ofIO+IFLg2jMHhDu8n7
U6X8BJEH3Iyv0hF9Gci5zZNNKGcRemzI5ZJphhXCf2L9QnuXYzcRpKzlbFb/OvP3C0b4f+arruXd
4Sow1YSKrjhFl5a13OV50LRUqcZKaezmTDDvZRv777E/XJ2zYl91S57cDB1nBrs848v7UIo0YExx
zTyjqqGBsiFqQW+n9j5gjPAxrXK885JsnB6GRBZFzlPX6Zk7SHnOrSIfvOYYJkvSCrUdU25NRPEx
H/WJTs6HXfclPgzWg/acFubPtANd/gNHWOr24tvoRJtP5AUFMV1JOWmLr+Z/iV8tVqIdEgb/3Yv7
ATUk4Ou8KGwWIYr5BChjPSGWfhwFs9A9o7NIHlcLvpUyK+wTSJmKRHNypqD23Nh4SQE5bqatWE95
qX/VPNeoPcaENDfKDzMmpfciMQG9IleZNsFIAYX0MCnVy60dRvAASSnror+erf/oSzz2uNOGnBqf
/hXQdiPQ2wUr9ThRU/pN7UN0dzQMdyhkkA9VipxET3Votxcq8W13jXnhSBGBDqouv/k2eNXHjKRS
cd2RwIuTCGDQoN1xVGcidZFDl1gihYUcoPjZeHvCAjF6k1matHhwaHoS3nz7dSc8Y4IgDtiCZPGT
r6YrA08UGh0v+3Hjl3SzLYbI92fEoCF0T79yavoTu2eWwZcGlfnmIYgULbzMay83rbA3GixIuCAU
/a1X3DryFEaruHpDnU1qowBhYx863LhOsdhdLh7P3XIxkBM1VuCk7KJFiHB0/G1InFFsKH2eEu4z
jDtYopFjVU9fPF0y+zemszLu4o8g0Ui9JINpZoTard3o9B/idHSHvozIIU0rxgm/HFAy+MmoF6iy
H1BT99JVU+HGYlfItNTsiURPIMqy5ABP1MFEk0P7anJRsaMs+wtfbzdcBkvUXmXbJgwI+694ddiW
wtDXZX62ZDHEkOYtl4NOYXTUCZdJ48wMTyvWKlWzyxOI2PYGC2W3mqBIk3QJNazPvh2xIcnIjgfS
5vs7hUjVLVxiXw0FedViCmilUXcplvzVoqFUuF/Eq6gT+gh6QMsBHBbhS+aOWOGqjrF67k2HNKHj
V27bBNUylIoz3mSNWGCU/GaUBugtiMf40WdHgl9/ic1yqeB13g4RZhdjktHESH7J1mekSxLiKJRW
xNYAYCe+HH183XisIGkDF03d80MGCNID/6U1TFgoqqUjWYhVSyuj9tIgS3+xKrE0JXEVtz9BWlJx
eHe0qUZf6kAfohawA+bfght+uEDAhNK1vHCceg8YNyde456HdC4H8zcuyG1ctjxLibsnA12s03Cw
MPDcMVOcYBaCowUmcLF5YJdMuvUbnz5pxcpZS2Gg3hl8mC+Xxw9RBjZXEhn90c8h44HkClwCqsWq
uPFmAjRztNMLSHh9RCO34ypWgGs1bLgQDNdT3FIwxW39kZCl/IpuL/4uM1n71j98HDeg9OVXlTQY
yC6rXKBA6oEluZwrwBPUO4Sib2gQL5jU8/bqe4tO8WlgGXuzJqU04nIAP7ksTjoJ0/Y6lgPe3vhY
cTDfF6I5T+lJCyUBQt5EhJAf43BTCAgBTlarGQfTXHBx2aYdjciHFlY5zMgzoEQKFxiS1IW9iW4n
XsBqtqJUS0mWCuypNApqoL4xiz0pgjk5fThO8xegVJ/CRiXbWI3NtCXHzY7MTYATFOZNMEj+uS11
lmoKW4GFqRKTxBXb/g8/0iRvehHktgW+17X2WIp5jVbeXYSEcgviJ/fzZPze1mvaY71NZbTge4Uo
8plYqSb61TFDhGgU24M80wz7VZ8gZLoyYXjrd0dhbLGFoqMLRdGZZIFyypDSxojm0occQfQx1hll
W5Z+ecAieb/RUITQ3hevEypwty3+x4Km63N5uOYBLuhCLe8hUeutjZpi4YpRejAgMSo1DuHrBe9N
Ds8jN/iG6Gq46JjpzybkTaoEHVcClAPleBzA+b46yHPUCKsrFXzi6JVk1o/SDXk0H/tMF01/2NYI
gWGBHuM4yny7yZV/TuBWBpl5NCnrdACpwzDfXSAGaWUCiZyGsbJYryPJ8dE5lQyTmn5PdmGZLASI
7JiM3dmao2z4eRq1apzdpnIb38j9mBEkRNhEmwl4zd+xuTLe+fRT7v30DTU0gfzmTzlulgZvTq+a
obahYfKNqnHHdUC/U7Wbk0r3NM8QE1cZ11/m7y/Gf8dLihi5lFHWsJQnFK5rVxSllrgLLnExmq5o
7GyVzlaUCaU6JyLXut3CJrcaoPEYzJo/VzHGllkv7fptCuIveKf/oScLcOHZSXAFJiQiyq3SiEPS
s+arCGuDINHD31X2x8ggwgq/sBCgfuxdexSm3LOLRnhGW2VPyvHRRvkIGmsopjU+mvYbLUjcZfZs
vG7lBVNhPWlsOfJB1AwPpONrFeumNZxzCMvKEPlZvOdxvwPPpZC/tpk0qTvv2glCeDCbARO7p6ns
WkdCJiHaL3tLwomjLw05KpiNqfHWmvrB7rr6tubRQNLd/rE/J9AIr3F8HuBjcszJAdnZKuhgZ5XZ
rZVTVsiRlpdywAQNDX7mKlqvKFrsqj2CDFeGuO2jsFREsS+DFBIrqiCOYUBh1l/I6Mj7cFWl3yIt
kgU1If6ApUmFxTkwA+hLbvdm/248Tl+OG1W/4UhZ3OTlxiKbUe/upztVPInFN02OX3DMxHP3UdPA
fNMzu7Vu4aDJYbOGQ+jBnyoJIF7nvC5k/SrWffA45i+HCXCcVKS8mJEkAq7gF1x3fRLSGA+lS3UP
Fyj3uM0WMIaIi6srjt3v3PDGLhCdzrqF6csQN8L6ckQYhVIdX/rpvbY82hiJUMDk8DhQdL7C4cwS
ZMaCx3KUeqRQdTQ9wq/pAgHr8lO3s9BRWZLyijU6cxRf/nh9doPIM+sjuECXIx0Jo7v3RocyiFNM
WxgK8f2lkdAeksqZ2b61M2WF6yNEMaagmzVG89VGrKz9dopkaEzI3MLN9mdYT2/EvuZJfF9W9Qju
pBcb2x8ax6/9FWT9h38bUzQxDdA9FM/bZ9XRMOH3qXriC34iyFZ3ritS1sVFpG8Uh/MCMV9wvN7Y
Ygm29JMfSBHsPjdjYC1Hen9YUR3/iLeVLpf7mH3+y9RIa2Fj2R4MNaGrVZCzlDoR0dyObA4cgpb9
o2AEZiiDKUIdo5vtS4TH8GSBYHwctP8lBmrkHLTPN0YJpZzPngqqzmIU9wINUXAGVqLU4b0sIfzo
pPgDfcuksd70jj6xPxOLcCv3MZ5fssNC8zrrPGLHXT52h3kSzD5JAcEq4rgHK5JG5curKRxxvwgc
Qrpda6EHj03tcVvpBxFM33tQOyDmBBgXrdwYhPwb/mEDMD4cXSb/dkvRuNs72ryGeUbMIfPALtQz
czxPd71GRobLH7bKxHPGFkNVtoRcCw1N8e5x7ITNZKGLkQF9B5AOIUCosqz9k1j3OejXre5/bgaX
FTDBRA3e82pJrjKZVV4DcMSVP7w4343RSiLIesg9075yLoMwA5ndLEYU+mejHqf7FcZPfEM5hSAV
Ve4ZOuUpwaofX/lbHwyom2fZ3CNrY9fP58VAGCAwf2AhlMPzAP7XsMZupWVQPafPyF13JAjyhokD
X1S2G6NgWuW+ZRjHRGw22IoESDLJLufekp2LdfGOsDKqkhX2sj7OS+hXsK3VEDSeu9wQGK9zxyx7
AVoM5LYZbAwCdUGta5uDjBWCDThxO5jI20Wy2iCYjM8eR5tcZbSnSu1XmzTphSId6DkgBxOjLvFz
9qnOzgOz+QuOs6ygoJt5uQD3obz4GOds/Z4SQLekdnng5Z0FusRDr2c6aGKAe5vAXZv3++I5Oacc
XSIFZ3VKKIQJwm/qOAGL1F980YhuM3d1rEUmagEOkOpBawBElmcSAdOdr2IfHIOG6itqXIhuXYcs
Wy5pavHKMIyUJYpcGGySRbZg5nAmpdr8IqwVkoTFq1vl6E9WweWKPvPskGKNrXOhimvVFpewtDQc
P5a40d3hzJu5I5KpV/m6B34347YtYnL4YPfk8uKjqqVBOq5ypWDv1pQhSmsXK/aNHeatHxjXEuWs
ZRRRs1keHrjtgelnkA8tiyZyALffcHLNo8SM1n2NgKPpdy+JWE1qUg1/u8cmD6Zj31HQdtithvf5
SFJPyrUJ9K4zonpzuhwPZVj1UUQ/62/bMvDNoqsPNloxXkxwYta+IgKOrjtUJw68c8RoqQ4kd6yO
WffjK/o1TaenN2YnN6LiH9DkV5awy7KKqrxLDdcOJWAtdyg2tHUxTc+E+1tgjG4BVJKpaX3hpvzt
K/EJ/xTAHd2k5bMq6fa1BCdvIzjxrMLi0no0+cyzs7SFjegIA1eIvSiFYQnAt97TXQbC+qWsOtkI
14XA5WC+ZY7SSrNPZ0E806mEwM9QjwPy6w2JnfXnJ/OimYhf1L5W8+w8tUvjZmRdELjpm585izib
flYK8zzjD54vzfea+H1a506qjV95C5rgC9RFCGVG6PQhYSPkBGxgpNxl1LbTo39RsAK3koKoVj9T
WUcpRzh41/uJtgtinjyeXic3jMiRcDE8M4+Vd9L3GNIVyJMTQ2/P3EAhAgGXsMZuFwWgRW//feoz
EQdW8JAHipRWvBL6sFdqOyMcEKAWf96P8bmnf9MAT2e3lKfNp0xJexrM9IaB9AJvKt088NbvHBfB
NSUZwkchGUm0pZegugVA3ESX1ieq/cG47o7bkECWhMqd2opq8Y2vRDjZJFR+oORk1xG4XzMeNnUR
ISmJmqztEtTFgcr9tMrqBHuoHihhu3EYBQAcaNXpl3G20yipaLyha3PZTxpJTMvm08f+phjqzasg
YG9waM9ZD1su0/BcbWqVcJKFBrdXZ8SXSgOqHC1LMH65Ze/Udb/xTNbLY8iXENwTlRIwQ0yxr1T1
mlGih14I9jqGSCYEWopkoyxNFwLbHYJxlQX0ePedD1J3WyyjzULBXyXB4lA9NNBl227WBGnoWaoR
hWhrMVAvkCRRKhmYbmQB2JjsYtNVtapvjmp9x/AKv8QCRYTuRzFqQv4CcOKGSfdMk94tzwOYcNMJ
RmdSSMePORop4TYCP3+HaZnSpHg/laIUnNIOvehLVnbfaVa7BYnwi6eWEb+3NndhyAzwRFTR2uB8
XmG3pPDV2rOveeyDkEwYrIfqyc4XhS+0U1XMEYllqxWLDMdywo6acSv5cHKJWlANhK/l32RmsJeS
z9N/JdFlTaJeCzO0XF2f/S+4dV/TnXORzb2eYqdVx2zFW6cDpkG6IRPWeae3Oi0S+DaYuKxapJaO
N49cbuoXxpXPVskqN22Xh3eEqGl5jNyPJXH7tCIjmAWGScW6EEvlF1fZcT+1dD+uiu70AAyc05tK
xKxg560neuGWCUsFHC4w6Qp5msYHNibLmBCCDu0ZkNi7D+g8rVB3RDfN/hdNQsohrmYzWmXwE67N
w7VcGIohGGvLQn7K5MA0rxUABwcFmSZ+cASFL2X0WLlgxig0Dyvn3dcWt883YMDVzoyEQs3UKSgF
twz5W6T2I0GooeKyWyzRMlYpMBggBeUnQZLQWGzC4py4qEyuAo2ZGAXGMuSdKaZOxNYI4fz5r1Zq
KmBYQXlWKK6KpquzVcbonmPLcxHZ6/JUQeytbjJkJScrFh25MhJ45V1xKGNd3Dqk08vJyE93gMd8
Ub1/uRgVUdZjeAIHUX9Tyj5HdO7Z2aJLkjhKg8fhk1pS9xtCmmQDXvSIqmWI21K394f3oj6ewmc9
FGFk0xMGKKWKCfNAtnBO0UZPG8WWLN7oN5YmsxIQ5CGV+HZVOV1kjPO1WM3Ls+uDZvyJUHT7+pim
bwBl1cYPpXCc2Mc66BzGcu4oMxuQIFOOTDLy77JBgzlLIE9d1nBbv+Jy7lCp+glGz0eboChvzXW9
Sj+L2z51Ldn+4XKD/0GdvnSdmJHmsD2MY6c/7iiicdf6tDxlPFc57bQKETf4GwC5TjbI9OmJ9dod
gitAVxuFuf37SDZkgHZ3mD2ar0so1glT6mELSQqwpMwKJoWpRSUs2E/ihDh6FKYORwCxXVN3qAwN
Zkv6oStupLMrWcykO5gWHIlers2LuIFivku31kOj7yuRX+IwrIGDOqvxttbLtk3wX6BiaBM5/pNH
afyhDt06c4vwDfDuiuJjY8/v4CcApSTwYjK1cGEkIRqP2s4YMMysffq2hjmzGrO97+ELEhwicUKM
CBJR1Bz+GP3SoV5phDmJTAIkzarmgYBkA6AWSdnHa9dMtNquf+g26pNSdtBl3tiax8aumd0WQ4Op
KWhqJWuaue0suw4UNmtBwHtq4DfjWrU1QJk+LcDFN/0wWoP5j/aB12xeJ37TDsdo0VwbF32gbdUR
CFhqim9U+uCAo7Ozb9WUEQdE6annkR6wpbBLNRreBi2lfywtYSa+1mHLNOF+/4mImNfzRNvNHrUH
IGOaSj2Gq+YMmGzBhWeQ648q6cPOTl0wpJ9MC2KFI//8W0f0N9eLUxLEMP1q5D+xN+6mawSbkFsM
Ct5xjCssOf/rdcyM+jL6klLkysacHQR7kG9ikwpWtlzkuhGzgG1L7RO0zGlTbOpwcALFehbIscxf
qB8fzmrHIwesay84oESb9RGMkXYjR/Ps5KfDJueln4OH/qbJmbqWXFuiJQ5u60aoTP7CUvvt5+Uc
wjO+kP+XW+BWuv+x9TA0mcFUt+o7mYUxtEKNTjzMSzqysTyAE7oaj7nI0ddSg9V+65VcPa3dWiWn
SLh/IPhOAwtPdnFibH9CbBRV4lAUIQZUd58Xd+Vw7gXSlrjC1BPzhulL28eXT5d/rZYc8lNKJg05
39srhgQX+x1wb67ZMertfdqrA1kqaWTGqwGc8nJwyS47g15RBRSXTt1FGYSFsFcRX2TZaeLl3UBI
bYREtQjqeCN0IFksXus2nAyls9kWWCYqiWimHRC2fW/V6Pdh0XOjekv5idj17mpcbhwMbA3h/NLe
NObz97MF0/nINlr7ONd3BVxZatgWi/IoJHOvsEWb4xHRTx/7X/kyd0lIeVnMhbYWoXuK4tq0tgEO
iMQJx4nAlOu/OHB4iUnF6ZqXsdmWieG42mY3MesEE35PImnrf65MSgCOJ+eTcABj1hBh0DViDh6Z
OS2dq04ljHgONh9s5gdrLBT7zmJJfosf9QhbwT+7ZUXKNATpmVGFlFLFA7TZRBayOe3cBiRnrHsK
ZPWdFCK854tjw/SgL9lAiNMK71zVVcdvGI/udXXBB1FbVVNXaumdE1kUm0p+Aob7Tbjcve9vhhJW
el+MtOyGMxiKLBKawQ+yGFFmKMaeDYH9ClehKCtHMw3ZVj/ot4mpmNOUkj3fweMYwQtB2q/i8k0M
Npm+jt4OQ2uWHUF16LCNnPr/KPFgSMX6b5CplwjnjAWE32QVN9NOOt6eQhyVwru7UAZ5XSBhEWTx
DOoO5kbiK6WlNCS2+ISulAwSoxU9xWblyZzvF0yfdcTVVVVRnDIyVqjiKVuiiYEV1HjJodQsktob
2Q5TZms4tyUoIjZ1IgLIoraIHXq05p/LVef4oryEYGvwB4kK5DUnPJuc9Rhe1HOA/SBw0LBzHYWt
R65m7023GoPRep0ae0HF2zwClY9ZrKhl7PyCwDsAujIzxRRwt5jhlmH4ioFfBeeuUhIWzE3iJSbT
ZD55q/6DAesXNyg5RBNsjBFdxYtfe6bqH9wZb5sDmxlmDFa7Fm1z8hV08+65hvuPs2Np/IIVZ7Yi
c8NPzyOPhF5P/JHhNcid4Q/1OrHE3sVFiiz4V+usODpNgFVMv8V3Z5SeMDOh9cThJryK9OQjuetb
rs1uG0w/+2ULqGmtDFzw1EON6+6mcKuCxx/vOHN+sT3kZmRjpNPiv9Eo4uWaGV7wuPw1WryUrEou
sz5ExvdUPyZ27SllN9QhNAUVYp44VfcCic4E7k6aIA/R0s3vKXQueGUzZFNtvhipyBiumUIjs5De
Bw6C9Ys8+4EEaXM0/MFMIAhs5Kk/9mnSjRMfvG1YklDsQCsR84HrCZzVOaeAANzEvjciihv2Hnrf
I4OVJb50/aKlJlW4x04pTXa6IWHJHiKPlcIZuWhtxRJADBd2JDDH03fGbA+ujtrog62k69T+m0u9
kDjpl0P3cQ1wpasR0+MW+e/a3tzyAtbnmcU/uOBk9/L+F9L6g8zrcKpC+bvf+zG4KQY+4Dd5ncKc
lX+IOlTJvNRJHMXOKWpJwz3I2SOogOHiOfRBR/LmbHwEQTt+yRuxHACav29eVYe4LXhRzkJYUPEs
PAQZGFbWb5hiV/qFPep4SoeFjO1nBNNzhRXMSMKp5jwsxUpEwu6mrTjzI7xhf4KX0BUthW5Idlqt
CGJTP2MFG6qr9+WlhZL4UHkqLGDu937cyms7xhxgKD49a0RmfvUyiP1Qz0yNo9sjKgHVJLioOUFG
euPpJYRGFyK70A0/vSGqOwx93qUIS/VpWsBcDeIgE+XO+Vxc9MRhM4kb/FEZQcn5J1J4o8/CP8r1
fjEhGxQGHtM6IiAWbw1Mw2xrC9H8JttETRiNCdenMwUIfougdYQvKF4nqEdHe90zUfR9StnRO/Xo
T9tjX+lzXchrxdi4TRWP0Za1KEJGSF4tz3+yltkatV2OJINzEdA9wHi80m2IGCQKJwPWy1gU8e9S
xoRpd6UcNiDqP+UEhMt0yTRm0t/1xbSKTdRTcgZbSvhqX/JpnE1Aepz8YBfR9DfYa2aLHXYW/3Xj
H0y06KeZsiO0TBl8TInIHupdK7qRBg3rKOg2XG8++mmy35Ks8q9fvkqysf3egyikCMd5VxTLnAtP
QJZwCqOIxB89WP/7wRBHP4myMK0hyibO+MihK2s+N/CzjLjDb6/H9wHDmg5HeoM/X+A6Iq2RoBru
pRofoc7YBRnEsVTh7/vOs8xuc/T5YtxVKHklU1pVIvXLC3GtjLFQDA6Kvre8yjFaiR0TdpiP3hCT
eXy6HC1pGTHqJrLts5nfKDYl7GINlL6KPu3SRB3PAr8n61NTKjFr7Pq9sufCA8Ugvb40TxmrsCkP
SvREiXmboNSbleisaAeGPKisoMyg/19uTDswQ/AdQ/k5fQk7gWGpVc3Be53bx8dtHd4c4YfhEzxP
pORQSW0Z4yR9e0+gxZBedWsTDhT00pSCMwRkPBkqZhRlG+WOJepYH+R70du9i4qWYvXTWQs3c177
iFJXDxwLkZpji0DSD8iK6P+1dE3++cml6hA1Ov0qhIXTK/pTFWqLI36um/o9gRILmsuNxxMI/l0c
TCbseb+4KDzE2krdxeyd2pkpS8/D1jC+O33P2a+1PucdIj1WA8q8afmobzaH6PTjFZDrnNqj10DB
ThO5G9VwK8ZSwWQgsB/OO0OqTZvb0onM2WJJAh1NV0p/klFEs02iAW0IbWXFSFuUN56CEiNNwRIQ
wEmUS99apqE2v25pwsF4gMzY+w072YaFhXeRASUzC3upGk2HlFzq1mRqHFgA9GKMEPmoa67TzFHz
DB9MaebED671XsSbMSW5gqDSsNMDhwPSjxpK2r3TlmfH9YVvPMOAKJzt3jhmleqxUutUEmb/sbGY
ecYu2snpGyCLsJEQSy4DUBubM+WrFxcYJHjBqkZQ/UqQk6GNJt6vvEeeab3bMJuf+G2+Nkx643es
2IxpePc7O/BNJzi9lZXr6qvV05UY4r2ZYJvTRhievBKBYf4oqw1xeOU80jCCEGvr2OzAVWfVrN7g
rGr3LBSgj92rpbjk6rAcch9r9b2Gwk0SoUFom8tj2JHKCKBjDrLtjNrbl7YUKRu2BqDswg18tcpa
5EVIJ9RM+4v/ZKaxDGmMUBYtbfsVO3ITmYEDKUKY1zJc65gO0ECrkW4r+1qzwPB1n2w9wtK+ifO1
SGBolmG1pK6OgVe2On9qg89xQohC21txM/Ii9MZ5ytfa5otCdRCCba/AnvDk5Ud0vQL+rGgOyHNx
q0SMNB62D66l7+dLMrrGw2uODeJGjDEEFyP6UOoRJrlMoF8fJeDHxmVWKPkFwBwTU+1qbkFn/rhY
GAdR42Niirj5CsvlceEHA9y1sM3URNaGdgJZcvth6bQHr+0X4EsOP0nsyhFCZETgvvhfCaf6jNoV
zuAaBzXWq3l4iX+kMZc+cgXMt/Bvd2/92+D7lz4tsa4eoXYmRVHEin4IvSfkmOzepHBai5UXAPYY
VehXjWImdNXkBpchQByKCyD48ijaeu1WkPmHmBDQ4QHlwE+vJezNE/yOkYSyZqbffSpv/kMZeJCN
HUxOb3ihrU4JH7jWi6fgIzy4xQKni+K+YEueEwVVDy9hOlej8mZAf1uLj9N4r/LfKueckIAacuTE
l9vkH+DG8QlI1qMpVO2G3mZgRq1KViD18/vA3f5z5CGIxfgz3w7yxu45LUnAQPlZ9xb9ASLo7Z8C
ZpNl1GnYk7DDTCtRM6mzK3Snw1OiY+vgLh85VICNsxHUPZlBKtDruq0vChCJtrwCHu20U8XiCgHv
ZwrNfNfocyGRmSk9UH5LK72T8L6JhCHEEzvHc335pVDLt0QoNFZRZSMFtX+28R3Rt4r+KysrgTG3
WOAJzz94jurbz1V+cT7SwJFPJSREB9bXjcpba0sEqCx1q+yMMXLRkJfZX4GVW0A/qdtifH5PQqDa
hmGurU5P3ddUr/M0p9uVHrTuylQ9JwhxhVj8z/MPWSuAzqvaq9PefQwsWwgmcN9udimZQ1YC/z8t
zlr6N11FNo8l1RhSj7wIT+Rfrz36mjbMRKXW4b+LPJtvrXhnrGt1DGt+/onb4IIGa/SiW3gpPkSy
9txzfdpeQAajKRl+Onw8/n2hnFxoMW6aXsO+DZ2ySa2+W1oPFPQ9q7+i6VbffU4GLxo+S+ZPTzOE
h1Y6H526wZLNBVCVqpUHScanfg0KdYQzTuL6Zn3+FCLxdx/JfGnwjhZj1uuFftbZ7GwNoHJLjFjJ
MQn1gfCccOJTLUQoYox5tgicLOmGFK2PcfgFfcePFJiVwtXK5BXEXw2x4f+bFnRWWvx2wMj9k0r+
TbLgmPalvzNyf1qIyHU6jOU7UDbL33Z+nPCln9yjWqHdXXU1GXQ9MUg3JfYvULTxn28tDJBiobqX
QArs7V7aXWNabodmUPZF9n6RjZ5kWWLWUD20gBZrh9FhhNvnf6FVJMXFeMV99ty289QdWkbiHKlf
XDTkjgeWucAdwJHHqJu3XDccEANcujeVE9U+iSFAwSIeDXloTSLg3yZ1gQcxhBOE4Xui8H2IKLDa
jOkNLgFYz4j70kyqVtyv/iEKqbsXHyJ3Lnok1ZMUzqjXrFfH9qKOAxyqEzOAc7ouS9tNn5EjQwDZ
ag7vgdrV4EiJb/hNqVmDIvwkTJFfwZ5aQdcjdMluFT05CwDmwQTSux274M3Rt5SgbwTL7ZnIAwiX
N4ZI8lHhuspbpSZQdfpSongA1jNF4NZyLr34mXfgMRaF5gv+Mb5vzGFQenT0euVfYSJbVKXjsk2t
wFIeBJBcWSCH76znfHCapIoEqMr7aL5J4SAip8pystPLYmH7xoVmdigD/NFXphoq8E0LAsNUK2MV
BkwXxu1g4hVgo6XmgGFVclAitxJVgeVm4hwD85GQMTVSUsPfouUk8oI3gbsPMkX9NXNLJbndVbnE
6N8V0tLFmD+EiickH3i0HcA2VdGXqV16Hg1PT7Rnae26cW8KWQxS+vYV281O2QLE+UCIEpQCo8xc
2dQFhyPPHkU1bXEE0UweEr1f7xRuKk3ZOjC83CBxoh6OZtDfA79UN06S+Kci21bb1OM51awtg6dH
DkEPmITbXiCNYJ8VFbJWzqmeo3sRP70VOHMJXZhEgGYx9ruPFwDgjTD9CSWUYK0MkHdryhWFFmI+
2l1N1SE6qI+M2kIUO5GXhpqgFi7Ru4+cFdb2uZsMXSsgNmLZCcN/n0XA2q+oaGbHYKFQTAdy91bR
lFgaAjTkHpv+dZP7iIeNIq/xV7pF2F2hb0YhpkhL1qoJxREXugqKROOzzFm6k6ab0rWmAi3gKpHm
wVmFb1ppjPvosHXSwwjDXubLTZWbzOdBvz6XCXLkeu/L/40WFXcPOxa8V+5vARR6izfwcpxZzY/f
50GDbJySZXFPAUKAqoKijQRaTQ1nAZJnFG9GN2l8YTDs2EssEg6Z6ti1735s4PqISQ+gB6Zkdgt0
fS+rzG8tLAV2gCpUpeg8H076rSdMWpLprqoIRATtvBHR8wvGhqJORqXDP52qb9Tes/Uwj1EYpUvx
E25pg/ycmla22VVYUX6aw3sEwt5uKDDuedyb1PwDts8iVXczuYwQgrTYvPZ77fg6dLx8yz7CpMj0
YUcQ+ZE4CxLGS29Otfqi7JRBjLtpAaiCOOZnLYZfjGqW+iFzXS5Ya3JO2c2hsL1Jefo59/YKxjzm
OwqIYIjY94GXVwiN3NCVm5GwaIwq/mVUgO40gIdQDEGXypsoZzJQzV7AWnI4oq32WgQ8Xa1DwRjM
6/MpGezIoGf5MEant95TOgQKmGH+rxoZiAudnGCQYXPyEKcghcFXDUhfsEwt2ska77IAYyja2wYx
FcpXq6DqW7YVeU6Ix9rW7VfJfiSZJzrCsolO+YwYDmQPCOosuHrQZ2uQBlRQZd98lxa4XtAXq2GC
Sw+mOX86xTBO+Yt3ZZ7/Ic+48CLhL0H6LkgU+xwL5ipjhgBbX5jr/RmPI2rulBH9vn8jqx7MEr2T
R1FLLfyqfk49s9eUCKBNOtccMwjoMqQK6kHq9dJ+hiWteQDDIxGeU6qXWdAoc4JjQxmeqiY/9DjJ
UMP6/jl0beuWQreqJyAjhio5oAJiw5SRv5BhnHr9w8adevzr/OHDJoik+ZPb5n4O1nx4w2A9z1wk
6w3QG0QO/3Wwf4EcxxM7geZ593APGmD5AQGynRzsnHx0Tdx814xAjnL3zBPre9rwz6abu8/dbAOR
2Ka/TxAaQSPWVlG9JinH8xxrZzJ6SK7drs8wa/NlrbJD/1YrmqWpjOuExpYB6R71Oh+nd13yPVEI
N/nFAqTExkU/8za9AtDQDlhmvmjThydQb9MKDuY41vyvIMoCXWjcyntcJ/oWHYTOR9GXJ01TYBkc
X3rGVZ+zqieRDug9/Mv6bRB1KKHSluc8/y3itloadGgi8GQi++aIk5DT810lEdvZoezMBgVBzlc+
bqnDNYLtPY8cmVscRmxUXdhOENiYdIBeJyjKpCfw2QDjZwArPPZ+BSFR/gVMoLaHe9WzmKrTEBYI
wlYCj661Iy/xa+UDZnbHy/kPIWDD2i0ZWpcYQdSLzc3j9IVLy/dQJdHB9PGNnUyAy7yecTasqky1
9QywSE5vemNMhcko4kp0bhh1Du4UN5iKJ6LE491USW9SpL0v5HZxJ9zz8p7e28YlKxVbycUy8Pmg
iSOtuLbgu2FN4WBWt9SpCQtth+dkvlvBO32U5KK8Hshrn3eOD02bgoHAD9YJ2hWaEbWo0g66EbIG
Gn2ckAL6DBSkUKzlX5i63yxikJ1eeJUlzDsbijzPWsKxTHysQuKWCIk1R25pKgIHi4U1sjbJPc7h
Qou3ZUGjRfL8OwMlqGXZb5myQaWF1KsQT1/yypu2jhiekwMP1YSko53KHYjqpvTOdyI4gwbiqQ2G
1+lG/CUFOy09fBWTurbMVhs2EiHIbtXb9ALP7yxh/dL6KfWAl2FZ02zZ9p3zXDqSHn/rAJDHnjSJ
XoG76AhfNe8bn/D4OX1FcR20JyzMZMFPv6rq33vzw9cUEVHS5IqD3V50TV8oJLozQRX9QMvTBUTU
HHCFo+RD+E4imASjqiTQp1sF7sK7RBa75TTr3mg+xOR56FJXjiPfefb0F+wEvwKSyCg4PMfYf1/3
cKI+9UiIE/SEajS4473dkbGZK/3OEiyOHmFuyAF6cwsqWP7xZbLLEcLus9S2Ove6lj3YZQn9HxVq
SKgDIgw30T2eN/HpmN8Z3CdSI9p89iT0FuYRGsnNjnoNKHOCD6fKuhSZciMUp74xM/n8dcV40utL
rGGD5DoJIveNZ7PzmfoAH5FHgGN1Kbw3NNORaMiOZIRLrxGsROPzrclrP3MRufP7odPQRn2oIQg8
mp40jweKRrIKSMeVHfgTceAsDYGdnvd4/StwijhhsXWW30KZtdhD6BHh165VW7WcSremn9Gidew9
0iSaFyKdYSTPFSiPvRC/kk50Bar//qYhSLa2DD+4Hb8vmxv/JqQHxiTrun3HRu6DbFC5eVl7nUXr
ilU5Ncoo9Csd7ZNC8lCUcjphasiFTpTbv+6c8RBjS1AVYpqMmryYTnMNvhx8FXovCGnzEstdWtBN
c4YCi45vIQbBZW4NREGPJU1UflmBUgcWrjeOMH5xgpzIAEa3YWzBtkdvxVZomytxL1qTBempNGlu
ElJiOKUg4gl7HbfQ4513GdgDPoqzOpC1tsWFNyI1XB1kGrfs8OvHTxrT7oqX9WvZBEwWt6K8Ndu3
tQ9M+DgAe0LoWvYbqGvdxW5ms1SJdCGVj1hoZSFglCXf0Ph97X9KDGmMOr0vmPpweW0ZW9Maebe6
0gBmAqnwdlU5EOBBZaTKlJUo9Pb32TIavUv5+oWmPPKcJ0ngS1M+Z9nFA+yK+4V2LIYfRQwV7O3W
GvSBjk/OTSOa+Cq7/hPL4/Zv8avdlBg3seg5kGTFYO0bvyPMYEfydrmJRMCk8JHHHHbTw2Km2gZa
yvI9ESke+gL4U/GmzKDjqCiaJrniyPOHeIswA02FbQSB5AKN2PvI3nLO+OzmItTkr2ZcD0hOg794
5S0sSm2iNWm7jCos78PpC58U1QWVpna9L7hpPvQ794nbnQ0L6NFK9wy4C5IOg89o6WGXH3GBBrqH
u1VLVsO+MNMsjUcpauTFQfCOIsyB4wQ4rZ9QBvHYEafiEOkJByuJdxcd6JtRoi9qG6WzJD+Rp2tl
53uQTdtsDkhCcsYgl+rGOVC6tQ/ffcFDVS8Hg4jP6RqUgyxMd1Y1HhOJMNMEKb+Fya5xNcBmbTl6
plo+Bd3ilWW97dmgNJCuOvBcsQPxBwA7kU0UBne5uGJUifrKy/zqkM4mWsRkYyMQQVelBXJt8hqb
pAPLmMpK373KnN03sSzZgIr6sNHJncg/iMyZ6o4wDSa9tjP+gzuvyxPrrZPI5j2ra5XHes80OLTh
2mjoQyvtxbK5eVi8ARPzAW9KvJ28itekD77VBVptJFOeYNXM/8fH6I/a5C6g9usgUXYL16kuxDw4
5k9mH4uMiJ2Vnnh4ePRpWXh+Gc+HQZ2v3eakKj97T3+8wGgvE+Peyu9yoZCPAg1CJPzR0cza0uG/
6Oy8bIL8JvVO6dRDOfeAEosJVyh0N1POf5DRXzGEsDcQxh527YO+2+iB021GG0dHCy2J7Lv/YI2e
v8PfD/XNsFO8nG2QRy5IksNrMpRAdkxIaxYzvjvAvebLfYfrk61qASSAe01VJx2u7cpyUZwzYeJE
ZWU3VK4bo+Fxxt4rn4fxdMXMX+U098e1kWm14IyOqZpVSD0zTDG5UTYM6fyx0xsmRVJBASq1AwNf
yxU7ZWuk1tVaL82meFxGfikVK7UOYL4/5ZA7YENFcy0WJ4hqKMoNlIjA2Ku+c2W+xtFJcLeawYqn
enEkXEcZD3VAQH8SoMcLltjBd/4nrto9hrvyvUCo5hNOOz8FW0/qSz4OHnWjuXIRr2w6Xg/jzKm9
99WXYiRNrYHUI5JHsLZv7fQFXG3BHXdFujsDrd1po2mXwE8dfFUq5aY0YVYAxQtR9CDPlDgl7gpC
SXnCUixu3IuOnAQjwWf/JOjTyRJIo+MQH52aWAqf5oEx4KHlIah4FH0zyZjGr5hZbVXETKRhbb6W
xQGh/71uxFLrcJfeXD6tDX0qHNE35NqMrG0J9edJcM1tXaKTGHhi5eyYRUzV++IePEGGz70nYsg/
YH6+sXRs4A+6BKxoPoMFKq3pIZvBavbdD10raV/ZLE9BwbDlVdOOoAHk9VhGCJtrm0ZMrj9rjE3B
esiaNwh0A2Bqmao5UmUP07k4Bws/COunca14e3lIs+JclnkYXmwlQvDCNYMkEbcu8gkTcpU+RKu5
e/7qXbjJdMZkZdUEpl6eG1vG7+msMKa0BPnLOqGIbW0gGKkIqh1Qq9hT8II7QghzxHqh+9JBYzHO
DhK8dCkBb0IavQi7xPgwSHbsGxKakvevHR0hW3e5uiwIq5OOxKL7SnuHR+NNJAmg3n/hPRmjKJPr
92wiUoao/aUgx0vq2Kx7MqedexLBl9JfzUWlXM+ipCTLHlK9T02gzxhNzw8WEXKzfJ3oS6Axrpn0
mGi60eiRvizVZQQhOijslJn0nnc6HAb+wOAbBiedcndBQcpvq57PEGj+aj8jCnUjgF2ITm/VLke5
ZfdkftXDPYl8si9q7lEh2Feqx5Exp7TnIikVR62pdMdN4HBIiJV/hdzQsDazvVmDg8wdPVHP5YTO
QiSsD50Mn8whxncjOUPNiEbuKOxoecIVU+c01uCDHtJHFkzjyE+evDnyTMKqzF+1taXClpv3a0fR
nZWdCoM299LZ5KRU1UW1rucM7QmgU0cm4Z3NzWc2aHL+MZRfvdBIlQwcwPJ8ueseoqLz+T8wk36z
2Z5QYuZR0ZF5Km1iRn2wK0zGdAhk+wI12ik/G9KFDqxt6Rtvmtma/VLuLKRV5o4rz2aY0fR1tjbu
8zCRanWb2oTWB+ed+ADxaUhmFi5/+Km96TZxQaJcLlHx5mLw13L6m1N0T9N66+kOTbkFDt+LRVE0
b+4nPb0qiYz9taxL26iVfrQYIPrc6eSz21B6stfpmxQm6FFnn10fcJEyefH0pywVlFULvVxriRar
I/MrtzX/nDnugiUQd2sbMe/RFidtZOccCPlCyd37U/kIyJcz19I9PRlZXQKatKqMvIqZ3MX12Tsa
bYpIk1nZjSjyaS3zYB9iOhzgZNKHlcr2tSeYZQmpp6Kk1m2T8cxGtbF6AYiUGy6FPPl6pn8e6OWT
ViSbdw4XLayr9JXHe8wYvtJrTKQj4Acb1SbgNNGw/sV2oFg2EAYOZ4X3BGXDBy+iWQuk8fQZ4ySe
Y3bril9TJXqbMJkagd4uYEbI4elIH5VbAai8LwH1P5BtXaYtJlAHBqeHz+oFVNeWbxayREC8dBnU
QnwAD4+Sc7vN/6pXQT7ukJIS09cAo7BfeK1yjWTsbJme8VqH6Z4IZNrSP6zrtEC7bshfE0kcIzpL
Yra+a7h46Pv2A7/vK8nI3lDssbJ+Hz98YDt4PxwzRXaDvFVMTdp0FQCBwFACaPqKZHrfVQoaVnhm
qkBGr/8BOny9qHbD05RRxEEpHtAauiXkv6sgJTmeLiep7WuA3NwXzsNSSyhaqh782EuTIvpX3Bqk
QB44pDUSvC4MA68juiccHDgPFM6xj7WG/E9tMad0KvsgA1r1QSDV+yKzgJFAjB/pJNf9rQtmY9kX
/rkSLRMb/rBL9/QaeHdW4A2HX82DjpejqnkhZcvY4N1uUkI613Dif/Epu4paXlSbq3/NYrPNC3eZ
GzyHkrogLwj0fZ0jn2Ekdp1VVAZbhT1raAIHi7Ju+E8a5hcwjdWsEjgPskJWRV4parY/HHNrnvlP
28UUR63Ul5tWuS2WJyHaUeYSahx1VS2CQ1sPHIqaIaq0/FMKWS/Wydx/RN9biOWoVKXMwB4nbPDA
UBloHvyyIRXXfI+HiIGx+meKX4giww0z3uLfP/wLIgUAeCTz7v2IncSHNTuhY23vvKTLfzIUFzp/
Co2REnRrwgMpCkG8YIbc5lXRnzhuiWisaGKjlOrwJBg+cHP8XTgauOrv2LN9dwxu648BH7EsMTnh
bXteOaBIz33Sz1XzTUNO1dx5s7Fuuh6cQLI55NYQuLm5C35YuZauNBjw+HfRdcS6Bf8q6nDIsMpf
K+eoiF6odegiDS73TfpIPBZsyRgikYcfZJaJl7zALVekj8dM0nevHasqk2eq4aaYlM13+JDtJst+
tgZWhUXLPA6w3o6kL+67B+Mu2yfsk3MZAv1rOeofTqGVwHstQvzg3EU1OeiSIiHIRKtRCLmeWKkt
LpAS2px4wt12Zk9gd6t/+KGX89OwzWc3JC3SOP6vo0HZGZKAMVTYG9s7S1j0sWVJNLvaH+YCrKfp
PALiDkPU3V1g+RWYYoTW5Ku/QL8+VTIjIAwDUN6BvOhV0RbPaYlSp3l9Hj0aVEjDysdNiKA9Zmug
zTb8rxJJYDRZcnvEsZBiV8xrYCJDloBe9Wcmp43ahiIFxb9hbUJqAyZ0RPYvQt3ozFGXsxON88sq
rz0USeevIR301swGLRqzEhWdkcGVVNOH+e6jilumt2QH2a1Vdf2JQQ+4h26bXrK/7imUby9wJYJs
EQDX8AvHedr4bnh8up7OENFpWk90WSu5t3U+1CvmtVn7ycM8Qxh8rdv+XG2PKhPF3djalNtWnVIb
g08H1fnNynAQa+rwqtIQbuCFxVyOUx0titWxLB6NN0pUhqHz9HcFN1EotdtmAA7e5HYN8jDOyRfB
1PA8KQacc1itgIyki4Q1Faqlfs+llipq4LGimaSa9tXQna9Khph+hGh+fI6NrSnS+eC4WfE7VpgN
pqZv6fPEqDm/dS4UZcS3qXZMG784uhGe18hAw6La1uBhrmRaWB004yHoZ1k+mC0dcHFTkl+rSCdK
WpEIgdvgIiYJA2HYOla85/CEBa5KdtiHTOERgD4ZJUSl1dBwLy3Ma1sXO4JNEfELJMNjjy+AnNKw
fXoJkna9gZRueJtdaEt8T8WRBvY0rnztgiVhZU6hwRNeLAsD6koRCVyjDvcHZrj4B4p9iaKMwrIH
Evf97/hoZ7rsm/ZAzZoFZuR8XGBgZH4SRGbc8LZxJy1EYRVpHcEEm7r+7hFQHFa2bh5h+fBu7VoF
ZfDMtxesnr/+kYwA9nl6FkjfB0NwzbFKKuPHBOWoNjY2ZQ2L7Qw0xpM4DHMSxkUPVB27xQNVkUR5
qHOYxmXNkDxIwnDIg0YKtbCNO5lV27B42xYBDaAaGqJZyGBc8pRKhntviv/V/i8nAGImxpX+ikzf
twa4Hzn5aTF3Dy7fGKnv91CX3RkpGNQTsXwW09owvvb74ito7fcn3efLSJ8Gc0Fb0NGD+V8N0d9m
D60h+81hPgK3LTfa/RGHd8upf8LzqMBcy+Lv1XH6On/XVQA9nLC34fRiCIw2vzCK85QxIMUTiXHE
UQqVsSWYMce2aDSeRj2G7HPevr/GRKVaPYtlt4P+emr1LNVMoOQQ1twmd2mzyWAd5+ZQCervHASb
BZS4lhmXhD/t+eYr96++9Mp2/RtgJZ87TWdyWKyZRqOWK/N3+KqbBk5DDSpuD1z7i2rAaw0UdS2M
3oAUSh/jSrwYPmUkq3FOh7RUZDaPmAPjRRvZnXBfPNVIddsULfUs4tuXpYpY434ibhxDw2D1dFSt
Lw/ylMxb+7IKJRcJRuyINj8cJ3+x6+VWDHc1lSba2ltJNmcKd6q+tF8tfQ0mJYVzsAHZO6nTHXLl
EstHWiQBSFOQouhGOTG7Evo/Be0oig8DvMpYjMMqttKqQM7gjnCaQWRa2R5UfTyLc6fDEemG4PyN
5N5QM4HIU93NbdLSTHsB7ooJc6G6pA/HxqNBWYOjlRlqKsfuzRfxQV/1BZWsu1TQ2YrbNrUMbE0s
58qXvrnvIXPC9hDo6C2s1AYIWn0+8JQCdydrPDwfz8IzT1zv6SwsECKal8demYPhTK2W3hdG1YYZ
1VdYR04r5R/IaDAvMpvgKD4Z+FdAe+z6Hp9qWIOSlbQZTJOuVgKI+VKPtT00cC6LA+4jhpt0pH50
wJ5sCsLhYMoO9p6QsDuwfyqjQqfmGFxnp0H8EhUkvz2P6fU+xgRQ3AxGCWOF6+VV2/Xs5yN2Cb1q
/mPEYwMSsHSBy0oeJnqYNoc9doomh1y7u2a69yQuTRhurtYz8N05XORvQqoQ4p0KGRGUR/q4y56T
QffrSNOeZhuAy6rpHmNjSbSXdHtCRR/XZ2ILB20cEGtQxvOdAhhkjzbRyuvhk6AVm4jWOH5vr8lD
xLQrV1s8Vm16HCaXR3bvwb/OPKMuy9WsSFmUQ8cWVgeHogkz0gD6sKU8F8o0NfI5p3PlCwyeylMA
pwpoagku7FMOgiuLR4Fp0Y/Ia8k2PSLuhnutceI6xjXZ5gaF5Jp2YcnEoG3ngG0H3TqIQtRjkDdn
RnBOiQQnlsr3HSaCVUDcBlMWiRiq1O26xCWGnIgpP7IzFvpT3n3THDbOBUrz2TpoOY/ygU7wblX3
QhM9sB3ochFBs4BgMEv5hqvLvEe+nIJ2XB74yl3C8MzaNCPiq0sDvJ2iaMw27RHRu63yKYwtYPp9
V+WTUB9hDRXH005BCOIdpFzEj7EbIgbB8lk0SilFiCGsHoC51mCK9nfLD4DvsuM/zUhT+bn81nbB
ULTXCllyd5qP1KiC6IXH0bSs+7VaP3wYsHLHBVbZALGvIzJ9OoQg1T7Z25zpT1Av3zS+jT9p5BOW
6vqPZVhCPm+USFylJ7p9lTvWFt0V0ozcfzosX6s4xvi3u0dgB9y6pGBAQWnQF+SVqPSLIGBMfFMp
Wr/oHbjLSSHr4RINqWQJdRX+4jsvzr6eSIRmY27Ee9mg3osBFO3qytl7+BBv9BVO0+lWFs4niSLc
mZKvsEYwah3EvKTKFqZhdNb2cp7l8gw9IkJUp3Ngc2hU1QRPSQocVR1DsOEKYqpKQcZINTABRLO0
oUplQt1O/fCizjnxsv7Uw0lIduxJdMxIBNORAAmbqrkVDVeXeLyz8YuA0NYFg7UsAPUVRMXoGUzH
Kq6dQket9Haq4qhZIeXru8PtD/Ecpkf61t6UE2Ljqz1/E1hT/mhdW0/1jC/XegUS749MqvlDQk5d
E5Gq+Nvvdo3gXe6QPOmlCEV7RVSwphimgzrrwj45P8Cr7RkvpGZRaeoysSBaCj+bgRMySVWa1jZv
vUeLl8XrScqjErxjBA9mvs0uDysY/Bx+VpMQsnffLJbECufR3DhW3ETLRczr+wsN1DUbYFQsauCv
WDgcXMhSPnQ5NtYyWpgVv/SQkTCcjv3M+FUkLS+6Fdo8geDZeR7i8JxvK9S+EGLEn77538mdSPTY
7ctpLyLCzC+UMK7k36NGfjJko5l23aJ5Du94Tr8jAnQ6iP/VlDAq5bkpP7f0Z1viiOvOG8PVW+2h
N6Dlq2le1rP1LEYxxbg60gKiHIHkNI3CpBrZLxhItmExDPGJsp74zADal5fhwx2crSDbONujkJlX
350tD4tmPQkNdPS0/reTritv7zm3Z3s6ENlKaNpQ64Jl5LvaRrdBLfNqwA8w7OaS6aeadp3v79S/
4Y40QINzDmrdGuFqzX6hkXEbO3dO6MyAvF5VWiFeCSH2OJxZmzVnzkM73PESPK1A6CDOm6TqN1HD
i3JzSVQyLEfeiFJqs+mjTqVyHkXim1KCr2FCc/nJ4ubGJkUv44mS07agjWlqPgnvUc2eQsbZi9Qa
uafngaLldTew0TAmMlqFjWNQtmRThglQIPcY9f4mNqtIL73SGuuKO16XlQuJDZ3uh+5mhXEBfQDm
pmLisluR8ceZyhmxB1YpJK15blCM+paDsHqeL3tLP63RnzRQw2NkHgR9y4xySeTbl6hpzTRxXISQ
nkd4K7jbSm3/Lbz/MMeTAJs3eWCvuiD9yrwWUphZtePdy+7xQC3xvtAlvwxBMCvOl/2f0R28utSY
c8Sosa8YRTE9/i+c1GxuWM0UgBC9d71ww0Aw8JL9yKnzN2v98IUe7cM1QyEF8NbPkh50ZEzF7Qth
mno2VODZpuE+TkIKKQQhIqVt+9Ifo2UkUWmcL7Ha5fNpRFb7TA2ehzRzRQw2F3Icg16e/4VWVL3Y
7fg5Cd5t5dSEejesrj41267dWcBtLuq6iaJUEhtCI7XGnhNoMw4TL/FuIOOiAYSU2eR8EFyEhIGm
GB+34VI7sb576I94yfzPQZODXfc3fJw9fHGv17ZRGDpZRgvh0VkTdzF5AE15zM9yFhpbk6xp1W03
wewbKXwU1ZiL6IAl3uCQ11JQYW6Bdm1l+5wjLGr7pUEJjxPn4uuwbHKE/R0WrvhOwbk/qy3rDqmK
+9AiVpPB4BA5Ew96diELVFmKRQ8e1ltkYccx4dpHWmcMnQ+INFGHpCMiSa2ERQCMcsQFExotwoLJ
8nxF6MBevQGBeBk79ONDinjxF2GoLtUwLqojpx3jASLHM5DAQcII39KZJ3d24u1+gvYHdbxv/IGF
Ut14CYpX1WM9fJxrhquip2jUMRUiwFJHXmKvMpmwHVONibXsQ0fOeRzupf0+nBYc9sMg2vLHxZH4
rPmczYR38M36wIRm8hP9SOAykTeij6zulmL1dWX8Nw9OlV/JX/6EM+Yhk+MC0HzbmO4tGbpibsWL
vOjfV/nvjrTUK14I00BKwjnEWgz/NJTRPf+Q0HAdQFiEKDY5fy02EZ3WGHsE5x4mAEWbQuyUA6zP
7N3fv6VCjOONvTXg8U28DOeQqdx2q8fR64czlAC4k9RmjEmwlnjUi9XiJoEzV+YXfdt/OWqFiAmb
gwQEr/+yrnh74M6QPGhgdaOJp4K/gG6Q8aAu353Uy9FCBPJ32oet2WJD+Oc/c7+C8IWc2LMZeSMV
KR78P7OPz4D8a5QXbnLnY01TXgw+PSkd2zez8/RDMlUKN95oH6u+O6ee0afgUPV12tY+BhMs4dsu
0XN5Sgwlt/6Am5hI8Utrkb70hlrOL+CnT0CBtsk6xs6mgWIzGFSVfr0XxQoRDDnn/9fuCB0GNvSA
eCkM45ulR1jHNldtQtWqpRAtNfQUskrue1yBAkAIcutnWl6Dnt5OBjVTpxR7k2n8VukU5IKmU84y
REseG5wL+jjRv/H3Dy5fbe4h5RkGNJFxXwkYMPJZ/po2/wsszmM/wYZcdZzRIM+86lDQ/9sZMhvO
jJCgQjSqQzMuK/T4NbDBtEU+PsbO9mN+Em0GEQD7fKx6l/ZvgjyyURkjuK6XnmFPwNHE4j/zhQTk
YdYZxCDOKV7fnMtUq8wg2dA5oDlTm3rEvjYjXdh7dWlSBqslC/eoZLikOaqFzfPUUxbddfZ4Jrzr
fPcxMYY2UBZUr2M2nUhkscclbfZux4KEB9++S7oOcvhGbR6AKi+q495GgrBHFm3usxNT9rETK66J
7y2eSF5TSH0u/mZLcAENiu3EXe5PWN4B2o06rnB116QbeL39uiWBSTKmZwgr9t/D9YZZdEo3Fi65
Z79xb0t7X/oZ73THRsVErTcRKzorcAaysjvsdmASQaldd7JwpuICd2HMLahTWYsQsbsNDhiGcn4n
0jcKGzl37tG0pUZ+vbRgUiSJ1yD0s4T8xz21xrhnjgZoVAY57hkqLgiblkGSu1igh8lUHObkkSkR
KlKPUkB1KiWadl0eyARxL99SDOfmtQdn3etta7DPgiPBAdXlj2KqwZvA4TfTe33eKOWBqbC64nCE
q20wlYVc7B5yWDkYkHB0BwAz/5EcmrE9RAzAZKaYh0JStq/04edL8bjBBLBiXberoFud0U6VHw92
hsh6GuJRwfUCVtc9mMO9oryewSTi/O1xEcUoa8JExgEiax5aUqL/N7VaqU8Y6sHgp4vHaDlYCBHS
lp9JgrtOPX6RGYX1cRFz44HKIGxz7Bfe/PwwBbxqN+tbxYkduZBV8mmiNy3nkFixDIC1Y+e01SEL
fkCm/TBZeshKkOdjoufLLw1yl6FRA4DjVnmASCkseHb6sNMuLVBYbSZvkiNw6/MuwFo8r/QYPFPT
iuVOy17oAzxihyl73pyrMUOlTBvM+OZwaUcqT6sD5hBckiZWsOsSO8FSafzg3i23KSEEDWfl3wRN
ap8T0VrY6QDDP0MfboWnUJ9wF+B/7deQP2gWyhH+2UPI3jOdOJHSEHVl7TdGGbVdn9Y1BsIm4Awe
aTg0hWyMn5Don77/cxUBZCHJsIcz9MGb85rMVGo9PAf+Ej1Xy+IGi3zFH+EKedwTTIC09N7eqjkk
T3jWGiI+LYAHKicbQbm0f9vQYjXgzDQV+9LIJx0TWU007mRJrIbbWiRydws7sGXwZGafvZd2bCIa
3W5Taj1yq/yjVqjI7hmav88HpwGPFUBlltykl02ZVTQBgqQKpeRpGUq4/NBzNK4c6TqOCZ5aDzo4
fUBy68QB7lnUFTu+O/Xo82F7wYfkZuspzFYoMDozS7T0I7x8ML/LSfZloLwi1ZxtSw+3YTr8c6Wm
umYFuW4vd5wWKxYjhSjthByPoByatTi52yuTs8XsRCbBng9caVMfLQFQXNPvKCkJyhax9AbzYcYj
qzzERFtFEYM+bkR4zxqhIn0yiF0i256V7xVt7yQ1a89rNVFgKEQa3HGqhaEKaFaZbe7DM2ZjU7cD
WtDH4i1G/E9kFIYzXCprvhLdHtPuEzmcCzu24ZvuUPIQbAFM3uxblOEb08FpxGVq13fHa657jKCe
BI5umiZ+l4eow2t4UsiLzDiRRfpdqFXf7eC/gUhiWaRT8QoTlYg2dGt0M8+ZZAiGNTr4wlqSvx5a
yaFxRpq+b5og0BuHsGp+sULSCUD/+41XeMJrVtXmDE1UnN5+z1y3QSj3hOVhx9ZdYPhsNF3taEhx
vbYHc2Zc3yBOUCnMpYLPnk7XV337lQJaoRnCQxiZtzUf/uphXrqSIrMwnfCtSHLPtF0ORbfe18vA
7LHcoLD2ZGIVCYiQMpJkAfrKhdDK3YcXkjFAhhO25kYcYSdcfqj4YLRgspILZzjvfwwvTrarlzCW
/hoW7+yEoupVPJNfFrvWGTCUfpnUwRUzorK8pr0eTIwJdpr2hvttf7S9EBgIcW9fxi8MgB7cFeTH
Ki36cn1PeYLP/1hd38hpIrCzdSYvfdqFF+IaZHtOFM5GCxGs8Gen+NrIIa72MiHEKgVis7aGrXGm
AiEAGCZgEsAD1JBLUcgArfDzoNsgydZMuEFr99w07Vv/P6wrHWZfUDvKISYYjnv7hSpRPUfYIi54
HRI7E19mRIZsE5hFmYZfnekTTchIoaAxTU7/SGZ03+2fXqta77fVpTysB0eDDzam/bwhOSvj69vA
D3GJlwoSCY7IvHEgp26A0cZrq2xGAtvOQT5jlH2ezLFlOfyNbN5htpXn9hwonPe96gjVI9vvr/9L
g6rC3PqCQruhnaffjenkCZJ4D1cj4Vs7BCcqrD5licS+yQVcmxSRRDy7uU6iJTCmFtU0OEDnjZf7
pRM103xMRNdMetDZ2hfL0zI+Lf7guQZIMcfYbBt0bcJmSk2YsaOGGT9UUrn1l0wo5Ftk6JlH/mv6
uC8E3L1Nz/jnn9Ru2+Cp2Eczfql7ebgTeu8QZRGRcETWqd8ODGGju0nbn89dymLRAzV4HjJWsQq5
szyY2EZKgQa3ggjNJ/8nTPPqg8nngWGwalNfS7AEX7fTC4hpffKOkU0vX3AcAqC/2pjGD6codvFE
safhIk+dnqCbF+qgaddeAhYjcrl4Q0aLPFBpWgxb8Ic1Ma1xxRCor7QbwuHhhiZUVk9s6Di4u/RJ
Tg57x10rhOtCYYuCs9KBZydrbymV1DuE0goZs8NSJcyghfVkg/TWkYlSreh4fPa/D98mpMPQzDkv
aV+bxlBI4CBcKaT2Fx71DkN2tOg67gWs3bD0OrlwdvPVYmNK30WgIsRdMyNIo0i2DARp5PM2ozSO
VM0NftKEsawclrrYcyJllHZNW8pS2RB/Rq5lx6fC/+pm7MJ5bHU2GZTa/zcGGMPXC5D/EpajdwIy
63R3z1X7R6WbaAiN+PDe+hrAOgpXl9U3HMpPqYoLoYltOpR1wFWAeziiNdt+zRmO7pAveWs1PK9k
az3qgFwR/OHzTXdeT9z8TcrJB9fWC7AtyYDcsVOPNidutBvd/eQDvewR57KLP/VNSOrGl6sfLOTm
NGWz5OtFyzyjSpnTHhCnMtSJJH9uC4YvjgdB5Lcs4tQZro+ONIQw/OW2v0wuY1xfFvIriN1bU67t
OFtaovjx9MNiVhMIa4E+e2snvJ3wrc2iclqiJ9IcOzktBL0Eep9Z4EIisubl8vmlUyBwqXyTgGnl
1KgDxjWRDPtE3u3z5c+7DJvt85idnYCrhTySL4ftZPDNnd0ak2MoF4F+3SsmDxLKR/11tc3vF+32
+9pLzeVVWT4ZfF76es9KMVkiFo+166nr4DUEI9mq9TPTAGDwSCEBwniVims2FOU91NdQg8zQl8Of
bc9sKztdsfVKuIJ1zLar94YX99FllutwTixUCr+v20iNkk78sq8ZWYbB665mMvRJE1Sl5IxB8zW3
sqakEPeliqeF4g07EsRU3Clu8KErzanwTDgy9yD+iZS+Dg2TOtZ5b3u/ZzknpXsOneyyq+rVbPWX
rSL9kp/fjVGlNMU698qkG1M2eO8mLche9oJm2O5PDJJTeNePRa8Ro9PvqsBADsUaYruBzV7qWNcS
0AmIb5L4+fm9JXxOOIsRiOv8w9HDbYz+0NdTXJa2r9G5HtIntIkiwERrnTeB6fAYUJlfcShK/UtN
ksZMjOjoZ/lbMMetfx7Cw+c4TH5hMgPqfFbyspUkSKkJAAO0XCjWVJDELCh2GT4x66nK4njIJOmg
XJdw9TgQSC5+qYloJxb1LHssCOt8eGx/muT5beHJ2bH07itxkXtTl0kicCmCjw8PB7On0gMP3j/O
Vdk+sgU4w5bu2BvyuNLIjSjcFGptcuVOqh2HB/j1dGlRslQKsz9UOjyV7j6jDp88a2RpmxCLMrxX
L9RHgBxIdbtfJ2kvqemZpUEXfjfHArorgKdc0ZklScYKEyts340dgMCCb8BhL9AcITiZ1hIDv8NC
dSYwO+TsOvEmtGeexQ+tehd7wB0e2AwePAggH3pRq3eu6WQ/1rXkw+z0xvFzOyLG2QDr0r4hIGFG
In4l6BBIoH6NYRRFsYyAbYXyp58DcG+UtAWUlgUF3ufTYgulqrBIWkH3fVRf3Ci+fBII/0w9EKp7
Nepvr59xevgMbjI2PtZbgbCNrh7Ve/D5EVOmAjkY0OOuqa/haRspNTROhS0jXwUeECrsT9iuvFt1
2UoShoBJa4h+GfwoPl41mWaIVMplsDNlweODbHEoTElYsKpQjdCO9s5Mkk225TWuGd0X03IJNyxR
bI9cct6jCMZAb8K4V0q+CBTGBXrZfIIATk2BfreC0rfymSND72q6b/tLie98Zf4dGzpLZpsNONr+
FzRPeyWTBIInwqtKn3RgygiamqxL/nzMEhR3IlQg7+gnMETPnA7qDdla5LF0qU+ByHQlOPJhmjGd
PEKZ6hAoSkRLKPGJuCOEeql/MOdjDOhK9ayVNrqIno2VTySkT7AduCNnPr8d/ROkhbRIB9h6QUBO
3HfscW2d3jcMpYskOA/l/YKrhzFV+XAH3kRmW4T+ZKSMkZDcW2lX7sInjPpDX4BghH66EHaY56uk
Z51N9p4EUwn+EB3Z6nBM4mXBRSoDtaZAUeb1N9NkNxuSQnBsy+HAF8yN+u3Gvl44pXNfewwkEMlE
qhCAj3OypkomRB8sJU/6QBuAy5QccZILvvXH4NEGj/C4wUqV1a+MCTNHNp0EOR2w1cCENsOnxjsY
Cic3J/27QyEzpNBV/tS710F6BtlFLH1KbQzB9J4FngBAlJhHOybEPY+mRgtWZyg5t7uStDupXN7C
BrUwl1Ohh27X5HonoRYB3C/vanjEh9mSY3iCr4toX4Rb5cKro3exdB5BQZgUTmxUfEGF8zNiEemy
LK+824Yg/Vpxf62mMGOJcgsNK40OVg+nNYl/isshXFaDaz5gexOmdAckHJgij8qqWO8zMtvzG+hh
gJCSfs/A1GEmgIu4KSMWuZOKIkrMswoD7KvVYhJcRWCe1mFZhikI2GpZoQkXr4QerVLGsrSlwOTk
cCNYFcUkC2PkB+M7Vk9wFq9oM1VyCKpWTKPdZcyL8Ob9fOBVe6ysr81ePmlv1y/8IeUD8qbOeT+D
TZ362x24jpK/jakWukFwzKOf6VpeM9dXL09Q4yrlnSBVm/rQ0ZYRfjYcbyDfflgD+XT+vGGq2hgA
VeV0OYR0oLHdIpA7itm0c6X/BEyu5ehyHkNIkJr6OMzdp4MZhiO1cay1wIJDQdmi1UudnTvI472n
DiRsX+qDZpd3aE/d/sFRmm5SwsYN75j23VP3emTiOWKq3optUInd5ooN6TZ2h2LarZrwxRa3GGk2
UzcvZY40PmBDMJEWVuVSJo66PWzo7DQJxukVg0wEerWO5QL2CHbqv+gTLZS6x8u7Pf4QmapRKvSr
0vLQKiQkEqKaxs0JH++ND/veHOo350ib3Kn7FQ1Dg2kCj9QD9Pr/RW3kyU2mbMu/lw+yGmc6dtXY
w3JDUTmPqeUErgIi7EyaeNxRzMTvjaJJcNnXZYTguPqHNY040+SKYMLLvza27YtBkdOMWmUvlu0l
AIDvrKLQlvwvMCU2zE+X7QKIM/m6KkKvBruj96b9sA5cdhjMVg0duxbcr8hwWIdH1nk3ak9Yuf1M
j5hoGDaZSP4Hv1djApRFa8+xyV4GEn1LIs+l9aOcQ08hhKRnowGyiqkYtTmIsmPV7tiYh9tF2jxX
TKg+colYUlfdpZGeUZBykyNZ/suKGquR5F9mweZhemEGje5iXLRAmFqm4tOmnVEJku2LLZukySVt
hezAmF7Vv83XYp0lIu5pMLeLceYhs1sTl4Lk5693lNPoaGbVmHfAOvmWwBX4U+PD/8fJOz8QEKZC
hvdOQhgQU6j9pVpvNbn8PUTsRHXDCIFuAq/G4jTqv9TAtlon4ckCCo2vxbnhiwYCdM4U49rviBxj
ijjgoaVYu+GZAbRnpc7tpacuBM7Y25uuPUEjA9fqgR/Q7cU9pVtIDNTq878ZNaZTAuT57m0Yppsm
OnNexiMMcRhtp9ctWj69Vin/qPpfLDzy3xVQGtnCSC5/2C6pNE6m7x1PZJt9dQFQj7+w+FBGJDgb
588B7LAoFuKrv4ooa2bbkK+jWfBcFlu+TK98KkHaQMqmFj4LKmN4BcigZc3uneYdnnDEoUC2s8sH
XIh/IOWSzFcFIe2ePan4RJq4urs1lFR9Jb/X0VKFDHhMlRU1txQAF4xLjlG02xPguVCbpvCTCG7n
5nYNllWf3M+Sl9sDBZ8OwvuTpwRCtvW9d14G0hJgyeTd0HgMok28/VfuenlRFe2qx5w1HG2CUeQK
dY+TwEXOimDXbRc/R6tpS3U3hEgYace8sd8Qnm49ZmL9deVKDeg5dU1fQ0ltPcQIp4VKY2s6Rfnk
coaw/XB6imO/GUC2gxvpg6Pss/2r5h7wr1sySafepbwpN09SGTT8ISPSrsWHpZihKi88P17kvxB7
jdcALZVHtD0SuJPBvHjgw2oEeezI8qSGx0lvj739uBbVzOO5Zksap0D8XW4DXoN557CBl0qpJfzD
KALUhKJX8is3634g5u4vA3S96YGqvRJqLv3Zs9/SMI+NPUbwKp6+j+DLF65teXLhSYXOkhqLuMKC
+dQJQv7vmsYdfLWdRTJSQBASFRqnQk0HPdGc3F5N44DuknaqWhTi/li2JB3U1kQfHqOCeGG7vmel
CLn2hEMsmUDa3DFmr0j4BjHZcShVKNAXRthX1Hy0idUAkaxvldKuvoivYlKL5inJ/GVYX72qt0sI
/XV3aHQfuq7OB+8IxbP+JskH6nvNfOgwQcyLp0/lmGrfRL9herZIycBKIYPW91C0xN7+dsKORiZj
XpioBgeZzjS974G+Ct6aLOYkB8ZjOgzUp5Jk96vxo7yXLh53jXhT3xTwwVsPlc8bICrNYWkFt+jb
nmokWvbey+wbKfdbJ48rRnUSA7APYSvdsysYuGyn07ehIi9uHnqRV7apEm1zJY0IJxfpr3VlV144
X4QjkfygHujfvxLtJlv0JNjFwz0oBMZSGNDoSZag1lPGzyNvTuoQojH+IMsCTqNzM5PDYRq5DcGp
Gus8ZA7iDEFi3NQVxoLTVcl+cB9hSDsYa25Yp1mKnwc1KEs7Qi2BlQyNTaGeo7zC6mUJNFW7UH7/
ftr6iCp3P+zZJMD55G5kqCVqZYTdCxgFLT7CbHuGG7EwhwmFhLBD7TkPwxvRESR4pUN0MoTqkkAR
Hre75Qm2syblUQ07OGv6JtqRz2N6g/JYp+l/ynq/syvYCEe1hrod1MMyaNRuAcnosoNjab9gP+5b
TTE8hoXacQOSqb1Bief0t6z+o9Y4g2+Zh0++9+n4bV56sYOeT3G7KH2nfUk+9AmGtSI86NMUTvxZ
9Xhre6P/kz+Zpoxvex2IFPFCXd7b8oiKl8HKEurH09YldM5Qbrlr1uUPSuf5RbKdGeLI1yRb9ppO
vo+TJY0oloWNDJ62pjIMONwhwNwIoTCd6ia95La0WY/ZhJp9dcM3SWBCLKCmNCBo488mgYUu0Cbo
msXYVtKCKUZ0kKvZe+83X0Cz4qYpkWeO8OgBRdHI+cYIC+kHtRtDWCS6AnELhqprwQbjm34tnIdM
9lfeNIvIfiiFh+TYzKSyHTkSBcL6pfPXhlSKc/YclRYJdRDLBg1fRaocFgs1EPa2QjAdo5tGkpo6
qYpLozlY7DXR0xS9+PaFXqk6r/f/lyzz5IjtvNcdwfn8PiqfmXoxrjouTjaoy61G7Dx1yWCk6cM6
lWFNigGt+iXhbDimU/t5IC/D5ZP/gSmETvAqjBmxi8eIUkV3dS8Ak4UexopgMOZXPkp5awbHqZSg
EsrSud0XKvJYJAUN2UN52vBbOSUPnhJN8vEH/uMToNLMCKuoeqE1H2H+MagvRxsXk9htLy9uCzUa
btcW1XSsQUCYz5GQT+1bgVh5Abk60ltVN4DfycN25cE641xds7LAbhClfl0kMPT4UV2BOgyuXRyt
lvJRQj2UJO3Q/YYmtZHkVWgRrG5pmMYTyFXTBOJmTkSMnpdb9+AxdA+VPeBcyuzshmXm/H8shRtG
0sAeT2OfOvsLLsoVWQ/7cu50efsYpQgsozI1SsTmQ/3WEmtCYol2Npu4ywmHXk1anNAboZ+LttdX
7gyDpl0uYN3gozwd5mZfLuhXKY8BfyDAO28NsTYHgVCkQWctuZxN/UVooalGWWIawmwn2N95NYGR
Km9IOKcr8IX7H2EAiS+YQsuFQM/tg7rYhxauamV+UEfjjWEr/b/VBIVv8sabQm6FQr0FWnmnfQj/
XrFVyVU5ROojdt0DiexBqE340PM+wT5kd1mzFYPAzc9xCcVr7DPBOxl2p7OISIpc107zWhXaDFwS
JhCgidLpOqcWSelO1BNhskIPEE1NP/eQoz5ntEJ/7f1QOyIe/nqKFD3QNsIadtwf1KI12Vk45uyy
uPwnu2qdPgKcCmux77W/JGtzBuo7kCKvoaXhfaUtHxuWLHBIWXPLxuYtPXmfH4gllEeFcmvRsAF7
d3DrGwraND5u8zKJIzTv/x6sCQIzncF9o/7FLzcfaNHldFZ9KvyI9K8V+HqtKdzi+hFSwZEqm2NP
zbg5HAHXrgzVHteeYp/+qD4mBkUQ/e6vtOkD+QAzEdEixWFuiKKH/l82JQajaAmHy5q5ZFjLzpAl
ZlqyExff91ANUoIoIF6WXXxahK1FNi7Q3thvA/Z87P4fUft9kWeiENcrgyLMKJWfH19Zxuh6MIo6
b1t7KWWhaKZZsYWYKCZWwcI4UBmndzWeN2Zzhh9qCoIYrpH87i/YmCI16Fw4ns7RVFkpDna/VyFD
mION4MicyoyL793Fr6NMb4ozx5czCSFkBjp/grZkF8llzKwXVq0/GaEyQP6UvUsIZ8Enyrnot+dj
o6REwuMV5yh+qQ9TsdmTMVc1ife9ZCX3eG1oAhECoC1RGpYKYaFsJxNjmSfVsfMhRDCRHpcR6w4N
jvE3d2xggzoYXQ5C8SbVtWA+iPNMUyBr67WOD7LS5lQHnEOuVP/Z5tOu9SPTp8T7Xkfx+UQrG8h+
hNWMahT+txxlXybliMRO3GoXB5rkS4GVk7gHhdpMzvEV/gvMuPrlRXfmapOXUG5CCi8kQ9Kc+ZiN
jaO8tQBgxcrcLQARy8YpK7hW4SjJrBX5OZjQATJnq9bjUVznWHEzeXyFPzBARliISyUXlagci22T
/gsBlDLOPANTSHbmfNZ2b7azLe18oVg4OhJuuz9NPQBJ2BqXaUt3IT6Eb3JgCaRAEAHNaHd3Hevc
eVJHIvpQxoA1aooJrg6sLnh+s0ewyy3My7x4HDGCXQuqE6jVOqXCrRTca7ZwT9hNS9XbuqYgfic9
utvFk6VfdONBdhAqFQmPrx7evrz7EdA5GYCSdkslR4Z6LQPmTaCKBl6niNGCmubA+4huR1PX3TEz
WgQUfmgd56lvHXOQhUMB5Z75a+EyEGyOADDvRbzrFhq4Bk/y8GdHBZdowgTOCy6EI1MLa/e1EEux
UT+4DM3FC3OAR30QMMSU9ZincL6EPkDVeluvG9lIuABNIOAYZBxrBimwqdcaiqv4kwbpzIZagS33
06FMyiBMRLFpHCIFt/w4bN31JNg3O63YiXSwQrNYuRLnq9WQ+pkBFnFJwltfMZ/A+NSkdVUDKvXd
8UBJEGd1iXOtx4G2IUS2cMdN5arznq94P9XEwJemWSaMe6Hh0XbWNxpgUcH7ewljFYdKts4PHsNp
ESifUfIHqwSZltIO+i49XmqLtwHQFdJzpeZfvNAzRfrKCUD4rjRH83NQnwMUWV83fZTXJc4YHhP/
r2p6GRfiebQ+PDBT2xbnxJB6DgHkFF4zGycQfzRJILC01YVqpFcnzq3Iv00DxmnIxeQNmLvnnQSo
ZzMp3Xs6YKhvzJXLMj3XexElVGFO86R0Jt9Ug6wwJglRsV2HNxnD2Y/VlkmSKbY0Go8mHHJszbyp
GZjM/5PdqSq/f4xLiFc7ory8tLDvd39aIiureBCqFVAOfgT+s0E4+Rh/TULJdMbX11v+rgmn+0Lg
E8oKw62FxSY1lrgusJAaDNKhMYFvI/E6DAjd5kLw2ZKWNzj6VKXjM+yu1SyrYWuv+2YTAA9uvQM6
0naM85bcyYzlwMpFcukVaFdS2IvwcmblXQ0zVbWboxORdo0w4S2gZFnVpDLuZtpqVLWbNUD/rlV9
Kc58a+idef9Tr0ozmp/GdMJqjSEICEebsF+IiX5MaJ3h1O5FR11x27j7M/jsznO90Pl2dCR3YKI/
8KNZZaDNcZrfqNPqi0eoXjoFYJtiilu682ihj3teSfPlexL8LwKtbopd6bbWresyu/PEstB6tll/
EpHEo0pSt7BizEvibjchHnsInw86vHL3M8jw3tHdLBAqgdvDIdkCer+czsrDy1lFtYW8FAGZPwJ1
ySIIplraSB6KZ8DBFznuGNtIsY4zvIRDp4jg8eUKT7obBHni+Uu8Zt47bUqeBGxcyb1/F/Q5yUMX
vy0CaAo3x6oQ/f85NxYX/nfMBTrRy/oX/XQxrdG8sANAYobMUwVZBtopQh1S3kaCsxp1FsuHBes1
ttFpmipdpX6bQGs773chF67suULy6M5MdNQZpIsKRhTF2GFE37EysxoZVQxRdXWNfNyx0JI2tfEz
QYzlYBCdMMhKMcQKCODqJoe8UXRd3Da58j/UD0FEQV6bramN++fz4mxAv1/MxIaGvhFsVoYJQAMM
CEOci6Wi9GelQ7VgpuZ4KyI9qnoKTpO6LbvBm9bat/9gT8cZn4kG/LE7fbRmf8WFz4RL4XSSnN0Q
yzWxgqW/hWx/M9FlqB6HGpZb1RCvwLUW4aJLXBhMepy1yhGB3MMv0p9dTL7rg/7PTI2e7ML66Mbn
Obc5OjcyesIV9N+rnlbxKU2ONGH8um78lwfux2hLBU7isG5y+znBNJ3rJC9gykzxTBAindz5JLAt
Y4JxY/5bjxnC6cNnT7Xv6q0nV9hspPxPJKNOiIhpBYOJD2nZlFmkuP+NOeSggaxa+H3FmQvLvs/+
SLrw2ZYSyMl9O+o/wRxIg7eYSQUOVkkwKGYGsNnpknQzXhURAWMosf2ra5Xmrel8WjXBr/sRtm56
NKVUH/jbip4mRDfI+08buksO+JcQaG+Hc/hzCUiaKq2cEb1mZgrTna8BvCx1pHA3uT2E2BazpCOK
lK150ybsVYuJzL4pfvb2aAVJL8/U/wCxZxdfxxxI/LIY6omSOE92HZazjqc4bq3P8/mZ0+gzhVLh
edCna2Y+YY+Md7MMd7C8Bf/xWj4xUtx0PWtOvMIYynvHYRuTQmfhEQsSmNFnYXwNYvosle1He9b4
ml3KmAjrvWwX81IMC1dKPkvGMvTAUr7UJaANvc7ayAiGzltBEfcD+Ld5Ma+Xyb4YYKy4oPG3HT4U
l2T7yfOgVgRaeTLqx2I0tBfhT/NM1HXlSS4tYebrBMgpypmGgb0GRkvvXrX5dRqLTSudpPIrii34
9WLZRsR8JlqkmGSGlSqhGBynb4xK+5OEhMniXvhOWijPB402iFns4ubrBvnzLbbIZv5otmpwnGkE
1iC1MbOFel7PXtUjUbKUr6YdvE9W6Ml26T+lOxeOCMt2tW7iKmz8ElQ7ZPoRnoEpiEJGRALmpQG5
LP+N8uyhIEeaMwJHSpfHNbbNNFGBqHo+eDt1CHRB9hi0VmSXwTnNZEZ1SNe3Ju/cPT9sFT1XHHhq
A9OLnuh0H4Z/mBeHEX+A3ZD7h4++TC97LaQJ3wxTYE8tX5Cd7bJb1h5wzO8fmucZzHarYm3VKrai
WkWHskeWxTx2y6jU4SHKxFIAe938LKMLol1QHr6YJ3XfZxSL2pbYN07UhahaFpAS4e/DpJSw8YQl
05rm2FRtne1/S0QWTBeLBMCnBO6nFaMT/hVJV7RYEUWedKM8u/Bg4rim+y3eMce245zKIFj/kmpP
fE38K2Sl4UkYA6ScnfI6o4a02Ihd3HrBGqeaw8wyPOtY7BonKhW39DGKFAowudJp6Pn+0cM2P6ye
wUWcRcGEnob2A7z8oIZuyPzuWjXlrDQY+RfnZeY+ucE9vqZjk/0gRmfRyWiJYs2HvkdBGhEdS3B+
BRgLPD0ya9XvNDigANf/NDacdlRcONDKLv95GCJOnBSmmN4EvBFGrXB6RlYB/8ucDR/6xwsZuZ4l
nlQrYd1411xkV4L3Gb6D2lQ9+goRNMZpigmw4BGcnkDXiiW0RU6hoQE3ENyt2cYLvnBp0Y4TMJiL
3VNlEpXZzh5eaB+CEQ4F1Y4aPB2FfjdRvw6bg+LcddoQVk6erMv+7kWfItA2SL587FRtN9hEJ2Cg
BUcJxOuopVBhOTMemPRBAzbxo9mhzSOQBIKMNAoSM/smqI/zxHxSy20DzQQJm7GbOPVXytn0kRV0
30oILz8NT2tPSRID0cxzhzESivixBE6MCncJKsXMjCY97iw3eXEAN7GHvfb3KxrobpxrNgZmXK7Y
n2S2/DdLvUiS0vygNqqvD8kjg38v7+oR2M8aP9AoFJHhAmmos5mg/Y4jPFoEgmSE6m9UOGcTl0PT
nlpiY8KejRXjewqDN9WpADlHsIEz73vjC5e1RW+oj3JWAAKgvAcdQym/5xsThZqFemDdn3dx31MM
HOdWJ8z2mEsbuqqw9hs7JCsKgoBgcAbGYsfJtlYm+keMtxWSPsDtwRlJ3965cLxFh9judJ7z2liX
zMMc0bx2UpsuZlgqOG5aBfCL8Y7m5umCG5ezD3udr+Om+ZEARtwEcPGy/XROrZmA+avv8MCsqlOg
/6EsEfdUoisDxVmYLrJps9lm8F6pu70D7NN3RT/aQxfJiKDbaZ/o48YaqW4NMiCvmAejZj65EWFm
AP+4OhCwmH0ybRjX2g0Sw6A/y/c9XpbqtyESQ11GqbOu/Mu+MhwixRjfy+NPnjcyXqKUlImu/9cP
omcg81HVCQuKXXQg1Segw2XDEGmM7FXosmghTfgFhJ/NbfA7iSHq6fzZz+D5UBrK1b17y0dDztj4
3nqEDnkT+PsQMKpTCvPwa9EwSWBfRHPuOIgklqhV4bhr3+OSTW/EHCvw5z8zsAdi7rT8jqHC59VY
csnTDZjigpjNbuiPwOQ6B4Ff1HE/EQj/PwJUX5aAFrQEObdTQ9XCwB/RLHcIdw82AMiYQfPT/gu0
XxPmGOX9qviU5ay3fwyxVjMQQljrJtcsyBg8+CIkiDcRYywC+FgZ6wsYMlL1izzQ0P4+DbA2iPMk
VtmN3L8j4YpSdwxme/IkIlHtXCyulQxfvzEEgRnKkLjG6pU/uyuu2TnSzh/de/G/J0kyNPLPPNe5
1OFH8yX9ZviEpg/nQ4YYZ4gPCjRlrMglQWAVS3W6IymIzg37Q98s88FAlY1fL8B+1HFvI+8UgqWC
ZDFRH31NTjNLoMtKVu8KXFjGBvoqo/WGSMSVoyueC45LA5sUbfgScMhJOIRCLu+ngL3YK7SFWJHL
iXAKxqpB1TnGpmwFd855ipv4uZ5XCT5hX+LP4M6ChdaLY/yCDk1uzji4FCIfAVvIRobZFe1ox+RK
fGGP73wnialZydYdl1G0ykJAQagiVH5NNplC+H94Msg03g1g57glJiRkF2awXkk/uac2xQ9i8YLK
IdFk6LBSpQ1ir4dA6d73d7ZP3Agktk+zyEzhF3odr4wh3c5CwyU/i8R0iOsPx2tuK+G680si/b0i
3JyKW59UuWcbVqoZrd7+M9Qlpp5gFYAEiWXniCkb+WXMkQBQr7CufMrgB75dLcRMPcORLOOgfL2E
Lv53PqrXKZAECqZaNGUflNKQsqANv20xsQ+Z+Sroejw7pq0Ba3dPxGj6mvbtRSLRrc6GG8CRp+e/
T6VgzOa8vhGCunIuyx16C/vDJzZnlN1gOvaafY26X5zY5L4gxpC+/5RgSxSkJGsyZh1Nt8EYZOrn
UWBf1AM8JY5c0ztojXo/SxazOyvSZ+wP4OZF6keWZco42lSbtgEtBvh9CDoWx0u8KE9+4iomdz9D
XLXQTP+1dmrQaF7kvguMwSC0Na4lRqoyRlviP2gTLJM10KdTerxqJf6K29+NgiSoviA9tnk2C+Tq
ajXF1yKieWki/kjjZA/V+MCV+8iDewAcpIOBF7uHadKyVGEIE6RpgrTw5uMRkGmL3PoP84Z8unXt
4Lhm/zn2rnY23HNhePoKva9oW/wGVNBdVTZC+UeVg6GejtR15MJ9hxKUTlMwnqPi6hufM99pvoxz
2G5w+hN6q909TT/NLxc+PiJAzgk3BbuzeefmEtDCrdSTR45GXOOXabkXinQChbLHNJO9TDWtj5xf
Gt80gkEClK005Irk53H40JQ9w54mGUl6iedjVOar/IGHH+qW5PdG7Vk6+sRAOswFuZnAi6RIKgVM
h0KfvpKHjR+3PeQaMG6shNdyuGmlBZIhpbski7dUHGNCP9hKoNWOwR2/y5pp6av5pVBkgsReieL/
0qqtkNkJky69jDeFJz4h9sWpQH13URRuEcAG44IHdb057frPr0ORBec5W01MkhB3e7gSwcvHuYRp
5KIPKBe9ObZqq6x+iXdF0Ftz5+M9n+w/9pzvD6rH9yAjXI+SiArpmmAlkHrwjdHxHQxz4/+Nczdn
Q6+uLTVhlxUPN0OAEx7JbPwJQJ5GJxAFilW1byd46uL3ARHafcVzv+GNaBVJmJFfPBrvJBA5cvd7
+TYiXqofpkRnE1arU4SWAT+ceP7sfyogHcqUfS+EG+e1pOQNgvoNBq6nOWk9UHzJGTdUJ0po3OH5
sNiBBnKmLeIQlYfZcsxVEtOqF5IWV+8qNTSD3UnMrnbnVLGwm9WIq2AzG411+hm1vF8H4Mpg3bCs
vYdLGGHVVjcM97mwPzydn2pIvfHsSgqsv+StHbm0VzkutzpBRfyYFSHNTQTt2YU7geI+IP5zgdbs
/qPAwKd5L3CwrZElgBT0V22JLFCIPVliBLzGr8E/KSUMtv8zHc/uTRi6tkEbDjJXHACJlSVEMqQx
FwBM6bHg+q7CWGPpYWMhkFAv/omnDL5Dl7XzSEe1YtvXQ4bumQRikU20JnQUWX+psGqLS7DisVDN
l52kyOWQrXyqIJXqe1nNPyk9AZuShlT8Z1dOY2izj4GPOvOXgmoKD1feMAI6qf7jBl9UCAxP6N+K
S7CcbvjW0cog98LHwmzuSkr5ucGMp2woGNcFH9cbpzzIEyMD2PZwnX9YzrD5Qq0vbvqD6GykAMjb
du6ynr9KEnWjw5kutKAOMKJd50/4/qHVCRx7kTBxve2VRQpSVNbloEZ01IF017ETLOeiimRg0Yl0
n+sU1ZAi7zbZlpU/qMgmgFMrRcyisTLKwFYrE98dT1aWwTwBCHWq3/3J6e4+5ra7s9ZaknuDJ2nf
ef8Pl9ZI93x7CH1jtOCm3zSl2lNH5ARaGtT/rwu722PkTqyy4fd8tVwOJFfsM8ASvB62Gp87sQhO
Cp2kZz5KnnNmtDIqR/zgylSxfBVqgNSBsHXovD3q6f26Zwr0Y+SA4etkb5Kv6yvZASmz+/cAJPix
hJpwZZQ0q8DlcnT6LekA/oydZxbjjo40IKKQMnB07fD1AF2xRZ0W3GOoND8nbyxfuCSX3PLDxW3U
upJpZVlGaf8DlmwbPMDrDCTnFx6VmbbkThS5anjEmCHxXuVGVYgUtSHXLaMwdBV8x+YpynuhxD13
+15gz+tCy0cwtdnyTSI+h1/GnAP9MapuT3MN52PQknVgcAJVHuaiA7xD6Rutno6bdtvmxFp1Iwj0
r9mXNkGH/GeRt9KG+8bLJGKqliFxjepk6j5iuThbd199rGhJEQV6/kdmXnBbREdYhgI/BVwvHSIG
WpttXlNKDpOGU7nLp3I+F4+MVHMFqiWjIGiHWrWpLlRXePZx91p1VFnYf634N6kkGe4KtaokOT1j
vtWWMeNxZ4hTA5nvNYr2fBUdjAA8atuLNSHFVT6Aoe5uE8b4ygO+GHWjJ1NnecEGvUJIYaTsLTFE
YJB2ClP00nVJFyuZRc8t0EqxWiCPjt4hGnFgL90MUZrViKyUys867fpckuWAkIxYkOhIdntLICVM
JrVjLZ4t9cmtXJP/X3GXu8sIW3//acsPFnjqj1SQ2LCZHvjGKRv7VFdzSqKILk4iTyCMMFXMEKIv
DTw83HnG23aRsfshjVBouPHh0HPOovdRKn5B0OJOsjAAZNe532BDvGQ2zYBSUgYbOHL3W6gwCg7i
PEEOqn/ArME3BtJLgZbpqJZr7j3PXXQYy3VZ7BfpGSbUuK7xWKTFJOengdgxzqDRLSj052LJz/ML
0nMZhm1nSRnZ7bW6HsrqP3xKUXGnrHpqq0Zej/5nLlvHfupRS/FVBrNgEEjbuXA2vVBym++gvhIi
uhdrdBHN2hbgDmfrvyA15lVvyAlUiRfWiW9E/jKgp7JgI0F0VWkSvW5OXfE06VKOwQHhVtF+O9e3
oSIzVJuw+biwUUzvhVw3pClum4uNOf8e1XJRP+Qd2hImAwMOCasfuVDsep2+4tJAAzp8gfnOoIfB
TN7oTlJiEmzVhgVsSRE4A6vT6zZuIT+/ESieH3ewDxNfLXaO4nSLSKyvJQXaFEIUGf8Pw/Rn+Oc5
xUdkN1mtLT2oYXeVnpuIKBmdEQpree5KTh9TCwg3nNMpc8bB7jiDGemeU0P9AfZts0QD0viIlpAs
Sz/ppVGBZcaKkOab1aGQkoKMV5Pq30dXm7/c1Ecp/tmMUQnZDkN5cl6yrr+fgtBI9izohRcCpIqI
gEu+QEuV0faCQRNtr/Zdj/F2kQnp8zjDuiuJzMsMqGpx0i+bFhUUkgbr+tlJITxvAmJ7BS4awvhK
xBVB6h12gY5SRbJn/HgWH7HKal48mNK639lRRba1TLgL0CHna6T5aoNHDAPRdYcshhg/SMRFEu3E
/VwAvL8SeoN1sI4Np6V7ka6wILk8tSDay3DCq7p1IcHKG8ILSAieqBZDNfItXfZU2npkkzYzzaaN
J3MyJTE/SoolszzSgOHdvqnu91ompeYTVU9P3B9GOk/gjrFLmRUdkYWXZyQDWtjvcuQr9bbBdIo+
FFyyLc0nbYhzfmvEZMoJicAtuavHHLDsdd2LEciL9UCKb7sEuMbJ4n8+C2gK6jFzj0+EY/ZhdOpB
BSSHHGdr9PhuuAJq6JVLZ9N0Ey4eVs5R32oQ/1Fe2jRa3EnHrXaLxQr3oMsTE6k/3s3oWuA1CGhJ
IQG6iAcax8Q9cUt/Eb2b6yqvqzXkyiBfYJ2EPN8DXtqXECuOrpxKOs/LhJ/nkdyiHshvdvXODEqQ
lZzMh1B1PjVwzhnLiQi4+aS/i9zTi0n57nm90wIYMYpUlR6yoqqR/9GJaWuHKKK5Ali3ofnJkh39
phjkmsgTt8qj0r62qNmfpEr6Cl0ZRz3nJ06iFoChiimv4cDbr6AZSJJS6fbTOGZkGVgilcheosrC
cpRe+ocbLBIrgL9/WlT+dxpJPRHQnlR/TRhg5XDlEFcIpsYXdLlVIqUMlJsda+d9lGO/UTBKymLh
1bhDKy3NUkoYQJGDUxoxBfZe/QaqQCqJ1iQh0YCpAUGr1gak1A0MQ+oK+/rMIMyttDzHKrC5wmcp
kc95fxeTVRcqOqE7/Cueu3pvAGpxZHtfqZWGBreVWB2TcpdYbpJvw8I+w2egefzV+es+kH2ZS746
8ZoryoRMghzllpY2CfrsdGmzpiYyG2IPVy7Jpd6Z6VggEdc1daBO8FUNUAAoxi2+ghuwTVTOoHtl
LvgG34g8P77E9AWL2TqH/nLMDkRbyIh1zmO4NJuf9wmLHVyLjJoSwHJAz4m3O30LrhRX3hTfv8qC
7qiMCWleUFqH3KqUF8/wHsg7nKxzC4aExxPol4OCGJMqKf7QskmPy1BrxRxzHF+ZuiZwYLu8HK4I
KL50o5Uf6F7zMxZ9ae9YPx67i+91qjCeBD1Z14ONwVwW7at1OsG8jrKWFARXNMaVcF57jEJQYq59
qQsZWJ43JWvFLqOcRSvj1wpPhWzExn4PsLcyuoEaPNxdRQM6lAn5zyQY10M6IWBQvle1LTrdSetU
w6YueTeaCavLHzPlSlorJRH6m9I5mc1eOTGj/ELkxRd0+puPvwVKbj8Wd24xv3i6Dc3n43AzqHEl
dS+c21USsgPnOS3mqG0lpHHY9lJEAypRyqi4/PFgNJeZDav6j1iKSVNzMtc+Agj/6MHhZ9+rEJ9b
yvHUhnW2U1sDrolys/0JHZPBCp5qVcj9LzfXDhUf45BBoJpXN0VDx9aqz7otVpRehlFo0GJaw53H
/8fy5gmWxRAr3Oxofl36HUKfg6CVmcF9u2GrZ//Uvo/4Z4h5Oc1YOSTjX5MVxWoQyRdiQKWHKou1
mIxbtrMY5PIO1Rmfe5Qb5/eyBXr+8H7wyLhTmMbgAyN63vTKFjF8UljA9dTaMgA0Kg9snwKoTKxD
rw1/QCqwnLJ5UbixilunQF/4QKrEi+6BXP+wL9/b8lCW+M8dEWXAXfi3AhQOlrnJdgCUqvDloaGL
E3w8gAaJ/a3wdzqRH6zT7xU9Q19RneKyoh5jEJ55rH6BQ8+8K80+dbWtivWB+Fyms/yIKDvMnbT1
vyLwlMqluFPpaCIVCBr9gObYr9EEKqS5n6o/3kOQEXYE5iZzGJU7uT4Bo/QVhJ2UM8K6aSw/wGBV
1lOBMmL4eIU1mjNyl3LAfv3WlO3yr1p3S8d5KWcF5FpsynglfunNG/psUUn+7uKbLtMPRfiFeu2e
gOrTXiIGUzhFpBetyr5gHE6ezxbl/mdLH2ZKwswrc3l6oemTg5Fw9RlKdDDbl/+nYd5wC8J/AJB/
3yva4+nYbP83K/PzV/Je/tbmPDzt3TnrAtAAILxqfxAtXLSC1rWw1whUNJaLJw8w9RQQtd6i4vW3
UJGYLrr2OfnXU/yu5FXLvaONSASHkdHnspiemKpncgFj5jAhWT/ItDUrON8LfXJGHbP1jCJIvpLA
R6+SozgNX6KiDyFdAE7oUw1juR4/7wwHsw4SecfDyToY1hOWx1ev/yBGyq1GWKjS6P5TpUE9ysy1
LWJO1VhlX8Scvpcsi93RZAO28i4Wn1D8BGqVYsQwuNZm6DhkP8RWuHMKz3GDUMvnCzuPRzoUniMw
Lb+AIQbxbCUNa7ZZ5B13PXxbhHf6MoM+QV8jj9IwMR4VgQ1oqsxiJbXkoUw6XAyvlMA2kzamjjp2
wta1Pxf2Efhh7b8EAi7W/IgtNTPDjf6e/9oAIEGlxYxMw8vMtL+DNWJuLox031CY28fvHWhmpiPj
CkgwjR3cS20PfplnjjwVGWzCErln+nUL3P5hltoAR82qRxj3y1XuqpmA3iXXAUP0T+3DQDCPJLJ3
Jl0OMMbbw7l3mwY6FhQCFwdL/b//iFh9zu/SpDwICInnztRUfAdp66ZN6VGB9AL0YmLf5tB/G0Fw
mbmvtVyUPBiS6SO9uucQ9HDyb8O2dVSFsY9rrvshrxdWZCti5bucoZgKomrIycNnbQ0VW6uxCpyU
alO1R6loU1HC+CH883xXBgNycdajTGPJ7m/bTM/stnJJ/SnzFAjedtlnlSjJ18cFj0Go9+OsE5PZ
NsSy/kW/OMVAcmblJPn1MJEbNg3P7/OuOwuGWdvCz+kMBR1uFXJ6WNgy2j9wdyo/eB/J6aoRnaBu
g1KqmZ5law1igGo5S6jEBNRDQQ43qRU+DGDCJ0+34kDzC79gROMvm8vbsVdsMr05rbLwe66Bs/SU
q2T5FhoHX3d5m1gqLpcS26xFUO3I3LN2FZ3CfGTmu/Xee7YfYmqGmp3MYEEIEHnfjEavvgBAgi/J
+OrD4esju/STYaN+90gyLhNojX6X9QhF9waKcFYC/CcUMNSEJprKt5c6LlFy0wuKBMT3il1bmFDC
eZzCi8dH/mb3q7lon8EUFkBpO9M1T0l3k4GeEWzaf7JTrCSWa+yQrwTQOczZ1UvELswmIJwQE1xA
jCB5DHJhKAHCdP7zJbEdNPZbrDCZ8CCFIY8iC/1NoWCF1/1GwyMfBKFw/k6ZUPg7VHOA4uDxZkjE
CeCfLD74pyZE8MpljuOJLRf2SpakH4yIH+2QZ0aux6Yk1FFdNcUluEU/U77qpgbXEqlhlBZXOtz7
Twqh8pU2zPnSGsbtDdsoyqEQnZupDqba8uwHg9FsmiKqR7Ad4aAlEOqwDNdMe+X3pVPBhJCPbeVK
Vu49ZW2j4+oHOeLQldlBCK3vuIteDKtFFgChPtKsTq3urjZs2SJVjhiN9DWGAj9AB6ZtA44blraW
K84os/2L3i+gYpQgnBh/6DHU4FjhG0kmjjjYaixwMO31nbfZrfR5zgxD21jP7bs6XSoakARB24ul
XDBfKuyqvcwmCjmMqj3X0zx0rAJdCk0opvlYpZc+0vlOBVF8UTiBxu1mXFdsbIS+giamBD4DL1Rz
4O8r8iNY937RZvo1NnqSyHhTbfFVhjrIT6Av7elNTuCkHMtad4/R92ICNf/ihO+e/MgGMoVg3OJi
/JF+q5hxmt1pmA3ewH542loUXCYYD/xALdEFYLn5RlTxLZtskTk19tGiTt4Ntrj+qVnch0HVa65l
8uUgdtfI1L9g7XFNtiruXuF4IAi9oZ/pbiXHKME6wwqv5+m+6cphPg4H6EnbJKnnDiVwOGDUjCWD
QmLfSp22JG97iot1ERlQkqJzzK/1qg58C7+QNoI3rQxsvSyYzS3M7vxyIPx8nPpVxChDwMKe5MAt
jeHIOwWMOTzpE6IePaDIE18kDbRWSDin9HnAzm5pWGAgxYQCfYr4s58eh4UkW0l6ELhL2ABkyTKC
LttIF/Sgygp8grkiBbTMNvpFP1jkWWgayhGBjq4cgCXnOc2BjZkFKb+1Yh6T88swwbVejRXb61G7
CPfe2phxq/DgHRFYCuD3y7yoJo9szFKaMVXle05LebFnrcxaDlfrAc0ymvegPegZLhFKF/GtWqLt
PHXui5N8skqWsu6A9JGtgcT2g84eKbtKhhKnZXwIKD7iEa/jY9vOMK59TNpXWKrEBCXQNjt1q6LK
DPeABnVFwct8bCMYEzp625jz4FwyopaYcHzIfzqms55YqpYqtBi/lUlWZjwU4hiwykn/23oT4HUq
H8X8OJqu/7/urBsgLeLqWzr44xjdSQrgtjsRf1sqc5E31bh/VY9Zm2NdqnW1VmtgGvCSLBlSVncp
FMayrPqbCTaQ9iNeIgzeQmPOm0IrLfAgl5d5QwTu0tGufODVWQNOhDCVhHYX89lmm/p3M/3WfsQA
Aa6YchTSAfjrK2qBdIDc83q/oediUJ6DSrDvkOzlMcgOWNt/DUi0KglDVpNnxJGBMuSClpxrzc8h
BY/CfKQqU0nW5zWuLFt06u07aAnJ9/FTJwYuzurgO17MLY8PJOl0dZWbSq/6tKu1dkG0fRbaUmdE
0YDTLWjOORFtZDnQe6sAavYO4nGGjrrOjH6ZkMDTTud4kpV9TwGT+lXRLskLVSGF1xsTLF1m7ZYP
JpV/wjMfS6iWW7a+uCi5aAjrSdPqi9SQK8A0Tlq9jk0wshsE9oPzWXRMWzZtD0q2FEgoFNVzjipS
kHx7lmvch/+1CaaxY1XjnBQcwDrlC6xqCKaFbo3+v7YE4MO9b7JC+gPYyl81oXwpSpK+FOPGlebB
jmUS0n8REsK7z8OrK8KwDLY6O1S4QdIg859Bg6+XnV+6MkRMUQpobnqMGGD32juihtsHO6qClxrS
iUimv2sYuCBHJTeqz/Vng0p6UYSm0FdoO19SHsdeK6jKS9bHouA91p3kGURaOdUW4epuG1FVOSnO
kSEVrSl3G3apbWKvJr+GcKV4cRdBvUjhRXnWhPcyZyz1QjgcxPXfDY9/ypxwOB+umsPkeXCW4S2C
+XKsa+zmb+3Aub+P+xCmsHskWSwf2R/58o9PjN6bmyHyex1bJ5pFidef/z1B/BpdNoa5ar+BQlZV
MsuiNzD46ucylh+1UT2wYDNNw1lNFZYSp/+hca17RwdmFOJ/ukAJwHlhzbDC6SqGeLD9AcGARFib
J6+a+AOMrMXgHcSgko6rE1ZwxxoGD7L67j0sknyduXeyd5ZoOejHDhP6US30a2ZcBvqE5wOhveA9
9GEZMXs5Dp/OZ3Ho3obV5rPeiYKoarqRtEGy6+eao00do7qjhUhO1PEZkDyF4nGxR76xjjUGkE1l
nKDNuay2nFshYx2L3Z3bAdePfM0QbGEq2xFBEZEBkujAFwWRsxTN3K3E5Jc0enK2geZf+s0gPQW8
PdFVupBkMWNExSfCChE4K1RKTRlvzuHdeBAecOZx4zMsr9eCBSC4bes2ftQartuRzkDqzuSWUpsT
MRXeUbXv+Xx6oHMytry+PTd3U8DoLnAN4HLbG32AYr7HMcneZXBPOhruWI/QsgkLiRzhEU+lGozN
rOIKZH94+dgquQ/gKzDKYY3wzHhDKnXfENkd3PG7r2p2IDq+6O6qwqzGP7Wt7HNxN+IN/RAWijFu
BE4UvwMPf9G9F24yGO1TphOxVrnvi+3CxtXuKx3evkWZUc9QdGMxqfg3R5oZLVYmYnNzc2wBiy+2
gTV40bhxjseYGtwd5tW/n2wUyJlwEXYQo1gkmsRPc/+VrlZ2WQyPa/PRu6DrHRv5US7TIYBmLALl
w6Sv6xmDj88y0yLqTFHmyuX7cZ56zkiqiMCb7V0MvkYpc2Fa/2i53Cz74Eg50WcaArsISyoZsLfl
pvhjiBHqVYQgO8r9IAV6YVVHpppB8h3xHhJCrRBf4IijUrk3nO2yBCGOnvNEAotXcc9DMZi0TFD9
zhxPni2q4QMOOu0nPd3YZlXWcGP2kBBl8f5hWtPyh//L9q48VmSsrpUbAhVj93EvWVesru7Tnelv
VvxbfrpKuaHYNqLR2mPsx2SI1O31TVulwTyCzGXU7up59HDYbbSK8506kH9oINn1i8Yyrf+fIDVt
A6UjhQDMhNXY+Kg0/owzeRxDdYuyWYPnULAVDQdiWTWoB2avmAT/xeb9uTZSoSpKzXib7MU07C5i
x2yHkHQgYCEtEETmILJrYdVnaIrGIBmm52MmSgZyAsWknAEfLGXuIU/wPJVtWMN4vIHwTngkb02V
8HpkJIXL3MCf73MDSgti3kC5p2UqqziH16ap1JQ0UIqWBFRfeNizb683i7X6ZJWvoWou25V+TmVu
1+j8Mgd+ibAvljMFgvZvzh5ypPfW6ur6+BmiwQ1ewG7/mxx4l/+rbO9XGT+nlor7+9Lg1ZSZJVB6
9Iw0dAu5T4dXmx8yUear5pVkquDqV0+4dq2oF8zvmlC48hsfzY1mxpkpYm2gspmZaE3ttMOIewjO
BMp0cBolnrKkn54EZ/aPayMaiWeHc2tQe1PCWqC/OJ+kgabDWyOl8SdMTl3pWtrxbcCYQK2E+Cwl
YWofS7tAh0goEp50wgFpK0uoHgRbohR5TuNJzXkou8BXN9lwRjDQ5uMWwofqCZqwDnOvHkMv3mFe
Nzi4lskC4Far6qaOBMd5KcL1riwNgqvsawkqRY3Vx5LS+wt1QhTmCiaOsYWnI61P32k/cXX36j2o
bxj7nAvwnaqJ2sNGQ2k6t8NA1AfEJ9WgrA0Toj5zFeFcCB6wZMRz3g73o+W/u2PhzpkxvRCE6YGl
EKDjaHIy7yMIBRUhwaq4mJDGhfWoyO6e4/qdxJhTunqqYSER/F5Um/L3x7gAJsLxcVa8NqSmlKvk
BZT9wUDVWzjNt2LgRTM+BJpvkIYbtFCrK6kXSsLf+FGJ5ey/nTAA2bsbKqKTZSPjRb9+Ja7lsYCm
Rqm1E+gmrCrwHJzzglvcyKwP/AaoKJWyNgBpGB21Fk3ThmJ6a9pXBe1BiMudcmkNUKhRKbOocg+P
5u4LDUOpxWf2+LqIyQQ9M34QVi+4KOGpA2zejVQaZyX2FjPXrGOQwIiHT7cx+C8QrUGuMHkJmW8a
N7QipscIHt4OQTdLHrOSiHyBqWLcApGcMk1IMhemWneotuD0gpNogFMTvedV2KidIFgF+yvOTgyn
4TUb6T6oELK6bECIgO/wSANcUCv/zN2H9ydII0JPkooyEj7+ZLcobxYiHQbFNiOrEjMBPvrr3sr5
7L2HCF/GPfZeBzv0/9A0OTttY2PJ3EP4d3rxslZWM3P2B6bXZX2Jz+ADcfRYQ0f1sApfFJTa+Qab
iGERpydn+GpdKPb4wB6YiMFPaIX1StaGQGMsUcRZllIQ607fTOXz1+9Tm5/t/+rYl9dvO0fjYKkj
kB5WLhDW+0LbHb7rTOEHn2TrAJHQ2tHN8RHwrI9Tnc401TlO0XuXbJHVnsq7l1GPAe93kJKJSs1m
Wj1Dv4hLimqfWJ2WqQjDQ611/yLK5k6FXYv1oH8rpxF099yVuVsgqpBtEKeO1Yf1Io6xl5HXql8g
pC4XLgE775pEJBQl8IZl+tf0RalMz4l8t1NZihDHH5LQC8f7jkhYUu+uCgPgjtB5MA6JwFFwSQnO
Qx5DAe3Spq99EPDnHjfTHe9NoFBps3C6akge7wLAmw72+TZ62rZz/xiGaXBUXWWd9qAOcNXgm0Ub
sfZfyNcq+n6Fqw+vwwROGAlSDedWh5ggUweUIC1cu9PaffL+7Db9aO9RWnrXOiOw8blFQtcHHJzV
zuBInXuZqA1Q1dN6gRUIXAfa5vzvO53Pi4xNGPjdfAUHFSlqQV46s32L3wsoQeFJ35HPCh3ksF0T
WkLAy6ZRCdvtbY0FJbiMtB7/OYxNnNm+HMRu8CP21EsfONnTDC3/spciJHTgigVRb1nvMqTxvzc5
SRzOh0IlWV/QANalfaSQGu4PJa830rBQ7VeeNMAUFY3Gznv+7LvD1zlDavl006gZZMEX5B3fASdT
3szZetR0kziai+9NVky4DEUHKBpalu3zB4M4D+joVtTaIwi98Vo9W8jRkDoX8VQGnKtB/YEGzWEM
Mg24H+6fWBTL+nR8nydacFyqb6ZHrwKO108ui6BOVBrtc/fMqJEdpghVFONFy/Os0QZWztbBgCsj
1UA60cAE7aRBXA82OqrhVn/cgkZcmydPbkJcUKZbioKZKm0qZYAuPkKsnmrz//Sck8O6QIPF0xZp
kMm17JLd2Wn8weZO5MGvtn4i9aLL24NGdJttaCeeeopbGyBnrrNZXJ20ceot7NTBy2DxwEiguC7l
5+++BoqMDxhrMuBFvHEsCHJMHoJGahnERdv5U6cJs0yMqWhPzqD7CSpFMNg5foD4zaRHxvkpJy4V
1vLEUEUeQqZEpkfeAC644uh4sN3fTbA7Q+1Zm6LNc5KsD1zLtkGrxo5ZbkkGfauKqMvoW93xMYeL
nSTQLqabCDICM2guuxVIuOOg3ZSkAIhQLztHxwwWqVlDrP0aj6UqjLRzh8JGen0J7amTwEGW2foy
44I4EQaxxrlb7FsWEH/yFsJs4EUDRVl7txjQwGxKmBH4OlL2D247HlX2KYY+RhxuKHlJQWRT4TuP
K2fn9GfF8h1mea6VtO9KVBYqX+3EdYpInxC7877/qcGTKJr4IFTn2IZr4ICqcvZfh68zqWs4o3d+
xBlzjOhx7IcULWFATpm/KsB0ledcXjpk2dl6QQt8lPnPEpi1iDltVzWOPt2TiuGrZQJaC4YoYBMs
2yDmhdZtFe+gxdJRM78U6tJQ5mU7U85RFuDuaemhuCrw0K9VXHeoQyejyc0fMfqvlfVaqJjCguIa
SCYK+crdmjypMnRhEgvQL7svBjN0L1cnAuzgF40hLhJLFu9kcBoXdhW6lPzSw5b+mUGH+Ap++wk4
7CT229/YDx7QVToGvQEl6BS9g4sDio6ngpgQ1fd+6p/kuDTByHVkrz3WCVHgW/7jd00Ur3vwt+sB
FItw89CLw3ZgB/LjLXgUY97EFMLDa2tQllEsipn3Gg1rbFkQgjAppANusA7ypj3yzrOnDPz08Rc4
SkIzNx2739ZZvScqSEsyre3LIEOPG0DWtd2O9Zawb5XQD58mc9WKQJDK6wLt5XXd3rxsf4i8lzIR
f6rmjaixhuCzkSMESyQngjPUXUaO+jNDN0SV335rOikzMpWrXylH0WYG7hD319Ws7Vj/pg+md9dL
/r5G2X5aT/DML/b4Qedz5m15TVNRzfwnle683VsBxo+VQlcMbTQc0FJNHTfxz2mPBjLgIHtIBm9D
x260F8Nv1sDuqWOx5L7coPbxXoaEfMvuFRwOM9rlrchtGoUHTeUbak4oKTIrtNNPt89WOaT6QTXq
85vhigpObj30a5fw0xtfz8kLPeQYHGsVSkKtIlcG+I62SiSE910aTyHAuwQe4WuhEDI5qBwwp8NQ
InvYdgbYmUPg7K79+/lZXX20agOcTVeHCH+mVOlzoN8ji2waLfQVud+o7M6BWyfqS9sHEOS8Hpxm
60RS7uJxf8SoM8kjOej3jW6bo/bHAN7EahD09Fwc5BjmTw5NRPR6b8CZ8J/+yZVP70wzDOHbxoQ6
ADd4CJR1TPwDtQqztrjq/t+tdDag/PcuJDbGx4AeEu1uWdGlKzP2TRzHpPZNfYpRlsM6FByUF/8s
aGtOc0x35pcNnbCIiGdoXOuJGem34/RxSd9mPKFNATUSGL0CqMMjw5D/ax9OSWny5ntLdkWo3Z2L
Q9eE813NlH7JnJXNSOKXZNwXGEbRg0gifjah3aU7pvP9ccJaCM4Unf9xD68pHqsXsgX6MpIbyHLm
UYnU0YKf5x94NpWve9YQgSIkhCXKTg6woquzoug0AEcoGg2FQXPQHkSdnqESSVTQOW/j7g4eVpmT
yoLYDkvR5Yp1en65dHNFFxXO77LiS3NuRGQaKXkurZsu7l7qVzRVPoprr+bU+Gu0I4WuRcWASOmw
whY9cN85HFJotlrsENeCLu+hfY3DrkL4knBr2sADvtpkPI++NZ3oBW+mlMwKfz3USfm6nOhhJhmA
/dJnmIDT55zz3OCohn6nuJt6m/4z5uTh1URmU/Bmo7hZV5dKwcMgRuk94/JbRwNKdkW6JHIWW0fY
mz8It+Uj4a/pHr8l+/N7r19CB+9E9FHv0qrkRMoFhQcnMDwsxsP3mvpwiQwjoOb34fLDSf8J1mdk
kZrJ83QiFiZOzij5aO3nWSdNKaHCwXnNZlwQsD5Xgf8LkL7FFhlxsF1/vnToGm4irkMjBCGQMbbW
Jz07i2QaXdX3hJi+MG/eqoLKrQiqLAQhEbIviVQWf9Y6ad9PlEGU8V7n+j26ywc0LI6HHuTxxFwI
Mls55089pJPwBkjkutVNz4GfRMrfcBVjGbysFYhU06h2LaI2bzAbXuKZJ9pfN7DDwJRC00TtehT/
Xr96VOhDP5/8vqAzB74Gvv6fE9wI44a09wFLfxaQzPynBdP9+UHw4cLwjLkW56QawZ+RtUfT7ajk
CUoYTlQqRghX4ce2HRSHGFz5aAS9GlHnNWR3x8hZUueHRXbe3DGnWY3IZCXmExqORre0daTUDn29
vW6dd1F886ZtXquAYnwQqlFgMMyz/ceAuXQuzWosBKguR2fwC5LQMQMt7C1jNmgjsozbU897KMP7
sTVKyH79uKAMtegsgK+HTgObS2rVGH5+rNE2l/lupE51Lzo8DGF8uewZuuGM4yxdbmTX6Sdq+csI
cQ4jB5CcC59oTjbyS85c2/bXVQyt4rzC63faLLCxV7t1xsvTqqRN391je+2uhblNo4bb2UP28mCK
bstQcqOSI3J7r6aAlbpWFPH9I/o8fk3vUqi0xVjNyfx4urGTBhyTuEF4nOzj4Am45/MeHrHlQtxD
dZ1Uzobuh7L/KFnkluSoG3PLlm1vFiUA0aAtOQ+5E41ZXjz3irX5ZxF4E2q/EnKliIooeCRd7Phh
uf5rEmXBw1BqHedkcCFo8sTFeBfkX0vCvXYzv6EnrTawgNW35TCIhl6r74OWE1nlBFE+OQiOVCB1
3iE0BwOi6EwG781qiISWpaR5FkGlnWtx2nTePQ51036jsHqE4ADt5vVGWp5vI8Omlg9jngn7ASCN
7T3/IBRkGpJ+QaeRFnIYivux3NDoFtA7IAyj1C2XowFL1UOlOlxy5aq2ylPEMPNJcsvhlEv2ekCN
sLnrRNj5x8fLrOGFun8pv1GB/eelZQcUU9ttsdnAdJanrRzqp/AtJV893swCqoNEC4usdYzW0N/j
+eAWBdvsDCEfAXycrgxkdp34QHzZOXW4Uv4k2TmPiJw3g+190lSjPNHe5MVjzTccwnt7glFLP/nL
XqECy7jAcqq1G4Qt2B91pm1MUZG1BVOrPU9eff+rVwihboNV34vzoCtxTgDRGIayoB2f75o0HHkc
cqUFmJo9ENwqGYhlKXSjCQMT3F+IPVDDqj/Yw48vQ73xBpFDov/R0HCbZK2p0VgSUF6lfLBvIasC
ebrjbMGtlLoCoy8cvzE1SRPT8Vb/l6RNiQd/YnnEb0xvpJQhWFfFupY9Y8uh7k7J9yoH4bXas5tf
HEZU0HaBD0/6X8rUpeCX6gmD+67v+oojH57bkOMYk0rRO7lWVlfCIyQdtLlj3EcHd689nsZ6l9J7
CniCHJ+eLAPObRFuJrP0gtkpcCyaAU/rixo4TKf2XVwVJFCGxYVOhQTmcl55STjkRdq58bKFikQ3
hIwqE5gKhE+XUFKA90+lERRFjxR/M2ihCFR2YLgKSedAu4cIq552LcHqDrEWe/EWFDeXRkDxRf6U
Ds30uSzEL6A186N0Pexm8B5iZ4RD9bp+cepb1aH8aBHoGjpj3HDYhQ2RUbLgYNz0OMmOMmNisaM5
w5hl9YG8vLygzn6AyY8i6W+Yb6N2wdzXQaLdEq4sBZwav4vsdejg6colGQsNYobe70yiPA5x9SuO
DviJZe/53cAZwf+zyHX21DHzqBtnDbhS1p6GPgVPrUz8MGP2BSfOS4nV5CHRW4n1SIPdk+PtRylT
z5PFdlePpJeMpw3W644jFGVjAWsLqWvLS5uNZR/MCdf70hDVAj+ynskMTBk7cPkPEvJk4xuyO9Fl
3ySdnhOUteSklLtWX5nz07OO4AlkmFm9F97SdPceQQavgsivW906cR57bdfJvk1pZKK10Cv4ecQv
uiW+6ogKJnu5K60t58VoeCBIqvktpPowbe2D2XxaNwBukL9sVBeEaeco4bnJS/d02Ipm1GZTBpOM
2T4lIgpCkYtoURUT74E1RiL7b6MXCUdfL7GdQ+PHbIpeLFqxFMJR7aMsJEBg4ZRcNmxs/vhmRvkF
y1MmB7Ppy5tlv/S/x0GJbGbG7SpmTnxe41jvyiRklq0nV38zgr6MVCLr5pxIOX+37T5kAsrOavAy
F26kdueJgTfr9j885JQGB9SI3l6ctMvxaDytbEVgsnF5e7jZzNP7r5wJMkApMYyzQdQQc01Dau92
icyi36FE36o/sbMhaneL8OZdiKLWqSGYSYQfmlQoC9rxXcSsCHKccDwmptNkHtvio83uQIevAGEw
rfwPlEUWCIGro9bg5es2OpEa/4ybfiRKPHDxkstBmsnnf05e19VmyRpmkWfXhLsFuLlOhrflKo1g
Ts7EPFXz5nO6q5YERSz+tmf0x6in0XFbiHEi95REi+0XUaMBFbreRZ0rAHSMZxIAiz8SX6TTNBpo
/xfb7T3FhHpKt9KLg5P7eiSeT8ZQKIM6z+mQ0asPXplNOetXNPRmahAmWjMQiVdu0nmJQV5HQYh/
UL+BEIdeBJee/hDIFxjATn0SohdaUfJK2wrqmlm+rGpx0RvfESYeD8INtYhcef2xp12FAj/mUv43
cepKhBv3qfFbjZKTerfvOx6/dncAEe+tyaBukGJTEtiUI/cBnvaSks2+KKHC1iNAZbcd1CcWvdsk
fAbstX0DfJ0a6PCTrI+12JMFxU2cmofzRsTKys7bNcVfETrZ23c84LNDzqXhthoqsYXiKNlohMlf
PcYOyIaXWgWHHGGxzIWWvMZdoy9Cu1p9dW1YY1a12WtN9ukQh1hN8kag7PPRsaqQnpBDuLXJ3ivf
rgPhIc32ZrwP4rzRiDGVHU4OAVQXBXEHkAhkDVq/MRvI1Z5rFYz+j9ejVNzoNug+9MibfYYl1Dlp
+LyzxOZC2TbXqycAwSvS0SAZ8f/sjGmhXMlLUjQh1/PXiH4DU2ZbVEEIuXxEaHF5nRQvjhZPLFC7
qy7jHObo016LQwx6Kay8kxAThDdCBCYmCqB6p9w8wiE5O6tGCek+ziEnd1MH0sG3SyVFiszuKmsZ
1TUjNmwW8IRJl8215ljfyc3e+uHlfG+ZqfdTEv/fSMF98oyhEff1UcSo0kqV/XNAgybLnGhR+gwE
/RKeYlhsDGsljNU4pbbJ9RGKjm3bNZFrDx/L/cJiRHcOg7aI4yXhFmsv1RBJiXD68rnt/dHUqHvy
LeLsNX+2qkRkMs4LKjMKfzLTfKCfrOkxMgxV5NNpDQMSblrc9huY+8UxTCN7PfybjaskGgriqPpc
TT/L6G7DlB0fEvVVj3fDl9WJrLCUidyHp8ftdxv6Jg3zcgxdoXreMj1P7WeQtxoIBsDvNTqFie3u
esAAHc8iRGkxNpkQiGKbK+uHOgg5uMGsXO8ZVwJp+fBZhBQmLOK5rqOWGQmAIP7/j10N4m9BiFLs
qxo5G2T/ZZdEERdfAtpXkqB5Ekpy3uZBOLL6h51leZMQtD4Tr/2NKkvi6uoYGGO8gE4I61EqRN4F
q11mUCPGKlLV5uDEtSPhNVXT1Kr/SD74rXIO8Bo5brE3lwEBvZbK/cyJb1l1EZ1iMdIo017lbq8v
XxwCwGjXlRih4Mv62P9vtrI6HJUfUI7+s6X5n8SDsJr2VmJD5PCrkXqXaBotd6vMC4Nd612IDIt0
6GQuhoZDq3T2osn2sFy8mvs6TQo/ivnBKAPYD+zyFIb//U7HuDfEUSGJA6jtymRtVpo2Rsq6kSJc
wdfbxfDLl9zalVxXVkN/dFqL82XO2QAe0Zlp6c3OLbkKp7Ox8kyUvhDP3xW2J760JQTrfu9A7iB1
Sj/oaz7/TYmMWJ91ZwqBfNAoFNTAEfk/6jkubmh1t/VECZyUbqTeSS8RhjoyAa8X8lb9YoE8Po6b
+fw1mvzlGg0VNPqHwhBRstRWVPhJDH5xDna7vokrBFc2Uu1l1HutOxn4sAL1OwFy/CWYLVW90Au2
s0Q3dyn0dw8o0CatAEoGd+1dw2odkPNW8jUO7huv5DqexLK8wW7nTXBe7k58iNJGsDDypHMbs1Ag
07FusKalgWAqiQN3+T7OwKsCI7y0Eql2sGd38wINnWH57JB5gnLurPG0QZG7mPDKQFOmharffTB/
m7wF4YDEFYf3Xw61vzsLulUfs7XRmr/gUbHWB0rb04WBm3IS4hiVNoCK3gXtjIhLMvZmO/EroECR
zbXcY+G9DAn1/gJezeu5eSs9T9vSgpoIdqFlnm8gccCFrUUnWlSGxbEH/8mRyHak6zRTBGWKqCnW
UCYiCVk36pvNy1SxJ21h/cPBDtbSeJbjvJgAyujgwjroxxu/9VZ+iPaZ43mqBGwj+8vw/nJLH3uV
oeXQLJ3OOImaYcme4h7DIc5eOSsumX+AA9Gd9eHsphSHBnLXxvwMuVQe/fDwCo/fd5U+TeKt1lsK
lKcTFXj2JZYnrMXcbW8KLuKSZwWeUKyWlgKJDMFBEvuYGUsrBB+Ejn3cQUXlN62mv2CdwJdt9zBX
mMjFDBlgmjUYyuqF6qw1If3F3VHFnTlCrceIinr41/ZipFhFhikdaG83m7T6TiVLlDKk0r6y1kNj
1ysObC2fgHN5uioEi/YPG05h7cwrUUFhIlId3vTFkUaJZVFzTwTMDVsMT9CenoaRgfQT1bX/Bfc8
QfqfPcabMIyW6ACh+JtMtfzQQe+sjUUJoFhL4Y5YJQUoXCiHXhoatltyekexleXG+ZdfUJs63j5k
cleRTz2mR4P6pzGPcCFdcCe2qNLUGaUMt0pivo59NCxZuVj/LBd2fLG72xtposayZ0yLuTNaUAjw
vDNJflLCz4+EtXoiG9j/eO0kNwYgx+HD5F7oxkhx8YaTO5TjzETpAN0HiAES8aeMNhQF/kIaNZOT
rk9nCEaQGITLhMPgiKfNRLMXwqh6TwZP/Ik8f6zOlphP/BAyh3PSrUM0R0TEnup4+SjTPOG49wgV
+pyUvpP4TqZM77KbTzrDfta+LjTYQgZ7Qgq1vRkwQ4ZntmlYIiM8rMI9DjU2cx/DdMGH4owXoXoh
/tIdS/ZW9aHjk7Cryh3CzvwjUR+i4eUV+L1gHvdUPkpnj+KaLkUjrUiqZP8WKwpQddo4WHsdHvKH
HXyNT7m6M2RZeXTt4us2RLZ3jgAlNITrIpCMDnFF062AVzUtUqM6GD66727fObM1qR1GFB/TlMff
tzmMiwxD4vVJVjR3NhwIIVVNqXpOPFlGBuWY842qaTmiqImHj2JnPVKw6azIzXDvWD95fNJeq52I
50pxeU7aj6T1do9aQ1g4ABnNXtU6QiVlvAas04F2AO8Wx/oN6Id4qvv/BWMEWTcqa9G7+7CRiWBY
CkjPLEmUXAlDs8H8/TJJZz5JxikE3QGxwEvmxL+5+L249cL6QLw8Rai3QT6zJu7018TV0L484lr6
1X5A4Pdp5JY42aHQZisdrRYD20AIePm5VG/fGmpzk69KX1G4Iv99MgGnQ/6YpCo0zaKt0pSrZnRq
9t9Bx96g9Erutwp063UOYfeEAEjSovRkWVbYhO5iiRqLUl7jPqyUg1WIwurPgQYQbpHsyQT6zbfw
HU6DvbbcU2gL8nS1flsoQd8nEhFkC6NGESomgRAwsuPJZx5VYKqh4k6HBMzxDAjvauYvwvnFHh0r
zsH9sk0j/7WrM0z18p1duANBt4BFokC3hOzrw/UbnTJ1rewSxn0Q7VKzL+niNCfjkhU7O7Xn4O7S
oIUtYkGnU7Tg8MB9NTAGSBKvaaMHIAzPvPA8piOeJtTdtDXW1txV6qjZZut+W4Ey60RoEUSWYJPU
rNC+Uh+IPTCd3nldWWlpXTflpvuxIWZAL9MU+PZ6EAFNlL9kaPWyrCGSq1w8twvNfy1Mr5I0azKQ
5bTSiqAumQoy+JSRB96f4JX7++ZPuN2znASB5OFOQN3krGjqIepVhr2VsHjnyHSWjHhNhWGX/nGh
wsq6+BkWNCaFfyq143g5PYQ1NAIaVTaA7XuLCeM2TcY7MCeuiuAwE0NMoFgJhJxWGQtxYx7cveTu
MCvQNE5coWGWcq5jsQUCkTSyUKIZ60MFxdWxxCrQEbPHKMkYaXQiZ0JBWcljRWU5feh8I628XF8b
WXgRZuTlNq1Ta2Kc9NRAlubugXTy4NCz+rYvnOIV+AXUjJh9SE3tlaqTdwdCOVjf9V2rWCYJw7v3
y/5SpL3A03lBdPLp9ZyxtYQ4cYLpDJyPPvOVVMeLZSS9MnGRx6scYejH3/W/Rok6OXJgG3WY1DZb
KPGqpmkNcIKmvHUNTZt49WfZWrlc7UJGWqJScI/A3tIdQr5jRSUTNrx2vVhm/PFzpQFJhyqHUOgF
N1Z3Xl+9l4NE/nsv4Hd6Gqvt8AGJqYK8Zh/wXvaCLmBuoX3o8KJ1T1n8MBTfWWDHOcr4s93qOfBm
wCfQuS0jhidKKfHoLpBtp/jireAsV2oXd2fZ0ynIadFZdjFO2PF+GTqw9ZCLYzt/mD1ZlUMBtO/A
HpZzEmkCY+WwMyrZ1FblnWgVEiH24LCDTPbGgAe/GgTtiPQ3ODeTZ37vWhXWM5DFh6oQ/8YF7kdJ
4UeC0VSH1t7B8OGJJTg67vDz7AITDH3dTYP8ifyX+sWIT0ODBJx72nfgJdTga57d6Ouhzl6YZfxZ
mAwJwttoYur3XDipR7qDxcNN9Vppu91rJGSvINY3RRFs4jNn4kQiQmI3qQk3Kow9JG170lfqSt60
pJykblDU1hQ2MacekhaGgYkqm2sEXUWgCe/0mN9TuJfYRoUVfCm/Agvs8z7CcjedhjszIvNclMxs
i6LnXmfG6zA3kQDQ4wAO6HSBjp0MV6XkRLX9UMdf0C9SjQrYLv5HlbsoV7JBBSg9rGW5opVRA1Nh
jXB3rxOk9Opqv/ADQHOoRXVgFzxOrUhcvTLQeostWPy74E0Thb5AvoRzsOK62H60caVpHUsyysf6
h6guKkjMX34wEmQFahbWDzgIw02d56C1DAGqMOJNsHY/Fj4MjG5EUx/HtR+0YnLjUPGGQa5Y4Qne
WvU/OAS1EClkBvSXF/yuq1dZOnvTwztuqJJqRF0ZOiDb3BFjNXkiLLK+bicIgxXkhlurwcDodNZ9
iQS+KR+rnZmSVz56WkgK5cm19S1T8p8BZRmFE+OixD3YVAJ5ojipEqc8uAlzBkiti6r0wl/cAO00
BKEyZH8ZE1pF8jtOzvbCNltoURPG/oEAkRP93/IOT3T62/r9iLdp3DXEnEa/72l+QvAppdVAX0D/
tM+oqWDGk7weyKcQdXsVsuhbwiPK5yHxnnLF6jq0D04t5ZzfNhzaK2ismA09pNL+WR3ve0oriRbE
hbkoXQjnojq+ev0DUlkpmoqJJRMcOUHAXTZNTXq3eU1vXs1HYSVDJhsW5kFZ4Tji7kBu0cTM8cgk
CiJJoc2A9g7WBHbbrdLWxkH8vLU1boQ21Nt+ppRmwiBt2eVqGSHO5/WJT4nrfu69OB6DtSNLNwZx
Ie16TcQwzrodndcjzAz4EjOMon3LqthSUrMx6P4eJNPSrEVP2Eu5wWlTUya38GcnHXgDR7yotCo+
NDS6sPlSzXaqjbUVB22AxSzOjT+ze01Ix8FbOf3GhrpSlImJ6CbQtwvGB4kc4owtJXWQiqQu0qSP
FPdxAkCeNdJPrF7y8Q0Ld2WA7MWtLZjO3PQC5ePijwBzuF9SWB/dMISeiEDKzobK9sBoO8eiIIhH
01uohdgve3c1QE6EaHdGHSUxiENs3V1QGXVCfoj1MOPuj7m5PSQvJl84YSL9sbvUqFY8Xjb0Zck4
2bhlHJx4ErcbvZ55hX0o5NtSJsBy+XlP/Pfpcd0u8xWFvAKjP5LE2MD5sOcfVRrmj6c1d8EA6rMl
zXTOTBzbfZpBR6ENr11LyuWyLBmicIwrLN/CLK+7ALz8dJ5EcuY1d4RJtl2KEvNuG8FdRRx6uqM7
P7h5a4+U2SYLz+Mq/3DCuGC7+HKFLQi3AJJ9BoSZZbTBQY+tZJq0qpeZHcI1i1ldw0VFw8apdyyU
prnXUCX6AwoSkRJhLiyFzqMuRXvRZruVM0TMF8+VdlI3sdx7PASmIpnMzsjsjveHYiltYSALpIdF
JuGy4Vk/qNmnFJDnqCAmGCkxdJHaIm6Hx1XMP2o9hJpnGf2cUzV2m1YOwK9kebJ0mTjUGiBJt/zs
g3P77QGgZZ0pg1EFLT65/p+ID/DmzrmOEX8oVYdQ2WwO/b64vjRWMDJCfRqaGLFWRbLUZRYrkCEa
O5U4V9hNniI+MkT0kjLideUhsC/iXHmakeOi/pIgQ8oYvubH62AMoxMJpEKJiwNeuxd94pHL3LSz
ZGw2OUGoIMERe0cm3dK8gSkcHS6EgTgvI/dMkAEpcU4+GSdY+8ZyswWv5WYAWVlgIU8HupWg4aKM
Z+4L9/sEjrbvMYCNhUCDxlPYJmS3LpmX2ifgT2Ht3UaQoOaU7R9CUwEFU6QDckoJl8n13sNjA0Uj
xtj0hqmHQuDBJxtjAspxtAlEn8TofHQ18ujHz/iw3hZKG9OzmPI5jK/nXtXyhMBrSQV6/qc314hT
1toU/j7kbFfUhxdgiauT2YL/bFsafYblWCQ45U7BBJHioliVGyd/+UF+wrdD6WRTp5YfcfVdVmEs
fA5leu4WfqIbHNs6l11gTH0RYyrf71+Y5A8U28kIzjGASLC3C/VwTDQ9QlF67RyzHOuWEmCbPbzu
j/jVoZ08pVbgeYG3qo46ITh+rNec+ensWKYq+pqwcFq1TF+P6nDaV90Si5aMB05io55QeRkzcYNQ
KxQZsBWYZRwnCH+DiH5yV8LGSdO+Tn1LPHfPscKIoDV63RmI9BSA69itvTUYULHFmJjOTP9AXb1i
PoFZrz1MQayehezmjiavgO7o7l4cNxyyOBlafU7oPoIhAORt6YnEXw+8ivNCSVnoesz6Fo6leb1R
KQlw0gGqx3zIlTQbzUlNL3G+6fMZdXpoMvXjfw1NGWbbQ/jOZKTJ4PaczFk5v7tf/8kbLXYv0af4
F52O1+Kdg9GH32qBI3YcphPVLQ5pxqtzDsa7bVBZcct3nn3HoucREPDNzUXC32VYpLl9ifoZB41o
q29B0iG4LClzc+xdssoP5z704RSQLtnrw1aCmYzvk9DkPQjN4bNVwh+8+RIFUa3HNd8SIldgkSFh
2ko8kHkc1GbT+GfyAGWoVkDqkyurbROxxk1u0TdNZ8BwXTCVvzleJZJmlEi7bLtAFM0sbVOwdT4m
f/FXcqORxKwFUBzx59iNitzZIBecl7+NR3hzwqmJItxysbGIdPkKcdR9lyb/8q+HEADdl0M3DoAI
ngH3PxltQKEq19Cmvgvxhy9ZVpmrFFmtMZYlWLXWRUy0r7wRZhATZQTCNqiRebmKbmTq3y8d8gAk
lK4t+jsKCjHlYjJJxJUdhibGLktFxkdQsG9tH7uE4LEuKlZCuNL2tEEaJf8BK+x1p2LViCyVwF7/
dXjZ2ExL2nSXRgXIvDTBRRwuGEqyrF+EKCEjM89UIhN/8OxQZhnN7l4yBBjwPcYA56Ovje8yd+i+
Sj630NCIm6JOKCmjPYMzUfzpznQe3f7fOxCb6joBfvJzq+E00XDnLtaAq7od/vLfAGIZkJ/vyVZn
b+0G+dRVJcy8ENP9lcIW2pR173kxILFJ3MW4LVA1PxOUsSndysXY+hdMRNS3BXm7HBak10CnkWMe
/giHBbif+XNYnnVi4ol0zarJZWtf61nAS4YMC/xRB0mTHm1+18bLYKcdcZyMDtikLJc4RwZ7J93a
CdPFauGMZUgQPaUsTSxoxVwu1FgTJEkOB3KcGdVc6ExTG3dOU0Gah726uIMmnsAztCPGnKhfEgbh
jH/gRoTxp3dWv0/ukxocUtz8a+8SIhGvhvuwVrdrJUYFECschf8LK3F70wGkj8JnJNQq0wm0gw13
2S0Wyqp5PU6VkVCtn1DglM7tXNPtVI8PJ6NaDBMWSWXbjeW394brl7G5N2pZT6yugrX58/J1slpo
wYd8geS5iEk5/DRzIxdRerid5uG6O57eGY+p1mmP3dTW+xXrzwBr6qmBrgPAk+Edzm78yeMSymbD
NQF8/iLe4ADGmU6Vw+5nfl9kBkx1WK244DJ3zbxtUlaFFoanaXJwkpIZxszDMZIFyONIpFblweRk
5HhTeYX80AZKNbPt6qJmFWMZaRabW/u0dDvE1yjS3bCnqyEONYc6E2cPaSF80qp9pK9Vi/B2SyjF
kt8dW6NAwiB8QYVk5cwLJxhe4pQfzM2NzOqbmBKA2KMSNv4EtAj6I0oAyg2n9klR6IF+I5RUGBwD
xaoA/mvuhn49+YOoTbGHn8fD044e7QhNhb+vwjn5dtfUlm2KisBlD1eO6qEyZuqTkajja4m+eQMq
upBfY/BcIL7TQ/znzjn16nRtyKZYYZSSZc76oLz0CABJDHGYAMiL2gbpq4IMgpDhOkX5eYmUYNAI
irSGMwvILQSVxSZjz7cQbiPxASXI3QCoDK9WkMHCHzfaUTtoZ9jRmUhx5J0yZy3sDyFmrzSlBBZ6
c02jCy/JAe0wnekFy7mkWEzj+1wmkwMg9JsPyDu7ClETr8CK/7nNAUqA3fhGU+++nnBS5PIEvEnd
GQb/GJl67l4WGhgSGx4rbFOo5of812xn9NNxmEMjyOzuYODgmjPbjADdjepzqo96Ny3nAAg/H6SM
bb+QnxfrfDGSoOPoSafR8kZydE3AZca/ngRHT9TnGRe/u7hjeV+WvLHJN1W84Bk5jrOM4FKWNgih
wfgIy9A0bRkOG79sYL0+pvmku/vlcXyEeaRMlbRcI5pI0PVqNUtPH7swsQBpq+/BHJnHs95tvOhU
Bg1knCKFQs9BH+xzVb+ixz0lfrdVhrfL0xeBt6YrhFrzCP9CIGhVGkCAw6Yn30/FdlFOSyoRhWpJ
WkxV7Dqkia9g7KMtB5XdTBBs9CeL+17ml/EZrHcMv4vCsociAzff+XpDMjJPx8pTZjuVOQbO3HEl
xOhaeSFaU0rL7WsOmoYQlSYoAUDuzwNah1d15S71nYeT3Z8nrI99Veelz5W+M5HkQT/qh5+IaiNm
qQiT1QfBfsSCAKaUs75HbvrcZADxRDy/ZnGbL36ycB9be/t3tP1RBLCab0CziQ9K+vK0LYIYzv7l
8Qjz9bOU9pthsxh2AoGRo2xNKxR5OO9VQxswHq9B/Oag7LchBUK9Dl1nZjQ2vxZIyah0iCUa7AOj
bSyqG7nhOdTJgBdQzKkIcvUwpkorvyR44eVCgsCsZKbpM6n2QOtnCVkxRtU0uSqnRwIFREZ02Xwf
Bvx1WVHCIxPJuuepqfJy3+kj292LTEktpIVKosc96YKrm6RfSpVFohQTBm4XsGnBKHMESP7+2Yca
j/9daKeqUY/pVZqgVapt0b/BwoXlofAdC25/Vtxq1gOD0m0J5M288xijcZSfYTQH/EbBu/FBLsr3
ZfFOYcZwvN7IAcJfvjPm6tOPZ8JTKC1oOpzvls/YjWchGMkXkdY6smVZWDYQ+jVCuEP0haFtLnDV
TZSi9SyKU8Xgg359A/SNZX+X4ITU2ye5Wp3FC7ceaEEmteFLfqiYEH4DUewEMdpPBkwyUQx4d7HK
Hf+BPAv5rEoLKmn93zSR8w29GfBBrL4qaRtRyQtGYAqcZtDAso9Sc7/RvNnj1zbNBKhCu23qW9n5
76OzmDelne62YfYD60ji++vTLQYYIreJzeJ7+wMWAuiKs9IxnS2YXU97lcZPDwDJNjoDf1DTLefE
4p5uA4OVbKeZfIiitPz58sfDUfyoGBV2AsLEEhNeZli4JRk7BboU2Rdrxz0EsiW9Glcvjjt6foEw
69ltSXgNV448I1nRTed7p5iuZBPZfZ8ysd+VLj/hKmC1LkhJL/efbzBjSBj3N5VI796A+sdTFgj6
Srf6xMPkes7UOBsojZ2Ck8RiZ+VhsYCb+7nOXzIhAxcM/iCWsaKW86E3Stbugl5jBJCoNitNmgqh
WMH2yEVArBIFjbRvB8X8NZutFd3jNVzTxG2Ldo1euEJXTdMn8oLIH20NVOlAX2iPGymXuk1851lq
GOaKYGRE0vOzP93nSPsnX61EZ+vOR/kOUeCFNASQABSM3f7oEVvdj6Mr7NF5nS7JosvTUKQtHZrk
HsCdwkLhgpoWq+nt2DBQT6BVvOY7ARgxbdKx7RjFirCScUQx4spNlw1we3C7Utdk+P1HKCYlMlWX
ZhK47vWXSMbtAsxQEo+Rb2laFJZbGpi1gyYKpdxOl1xllQX1r1igh0njvgGB3K7sdArctRkIHI9E
2DHBWoqiTb469DntGFyUT9QCc2FXvPAVs70EVPK3jz7ufZKyE5sCLzyYiN2A6mhWDbIrOwWggtOG
g4XhHHF1kOo5njhnk9Q66pWSDHbezBeAtU3eSjkxXfJ7yihvmV80kJgdeo20T8L7lbxYiHg2aKZs
qbKKPtD1i+ytnaZhNxO3vZOmk3zVtMt9J0+xgCVDHURrd6vXbg+62yiTbQzBFm0WjZKnOcNVgF1g
c96Npl1uyySW2Zv1yrwlh7WgwTpOS3f1tZrlh8NcU+f9/vGPbxl8zrBT3D9qKqigUo+O5+Gtrrfd
we0IrqlrK2VmD9EydY3ZJvQbETMZqmYyeZ/NHBs3oNmvoPXSZFldZBKiFyOLrAELwZ6HWd7eGlvN
qJtNkHIIwmi9omAxhqD4lS/9T+tLy61FKhCF6lPN2hfVxLJejekNM98mFDPDsx+gu2ukOB7RkMw2
5+/NsRBEuI+Epn+oUUAZFMupSPY18wdKS0MG1HWWL/yeKYbmGlD+Rgc6OXwmnEXIQUY3uTbPbZ7M
GoOJwY6qoXf2WlT4ROr2aVKUkgGL4MY3gAeBtERrgfrke3GTeBYsQuWG0I6yPTPLsEbSuK8CgqDp
hAEynUhkDBcwQ5WaEwbBzDAlYk3+AWH5G5nSJwkSMVFkr5OjDC/9t9LooB6bYmKY7/3uStaAbKGQ
LiHEuXd+9K0GiaJFp+LTUdfUvmLGfafuwXqijV09t/8EcFmDjmApYXMIhFSogBZNR9xt6dRrlb6A
BpNUIsZUjTV1RKEOUfqowezqKj/BFluFqvE9rUFuUpEtG0IcuRXU7NITOAmzuabH3KP2qnScDjrd
xGREXQZuOFvTMZvBiIbbKOpIOu35cOFbf3Z7KSrQLqT/o6qwttfKgoPWcd8RNrafiORoqL+EA7HB
QihLyZnc76FgT1XiXF7o3jejRNpGU70aIL809hIDMlPw9HA7NULYFmVPKSiNnA6ey88PvUNfJWsZ
vx2cdyN1dUyWIgMTbXe83RqTeaXAZ8mq2fWyOYRnExdWNpuoXRKuwOhB1pPKhZbsaLYe8kgoSJ+e
UT80m46yEpyZBO7f8QwcvrHpF3i1kPsiB+1YEpSW5vMU24yqP5rbDf6KyhzA1EHGYi+8diwabmPF
PQVpbF7Ieodm7nGfCAqLPGCwofGM5bb4/1LekQIsfZtlQpF1DYuDQVfJu+QMnHIyVmIj3n+oyucT
HXi3bHQOEcOrzV68uTGBjPfcLkaXyUMVR4qKw0wkst5uj0zqXzW0xFn9CZxapudyq9WxDa6sUQQq
kaWTaWt3L0jQBESPohvaQfLxTc/xleX/mwDkdhPSxCEl26OHSHayL3WlfyMo3KmCwp3eb7+klG9t
7nfSOjbTlgIUcXUUzZb1Kjkx+9wRWX8RoxWA36nTKLFfHvklX9HXRUiXCNC9JTjYRgg1Lr9vZEDc
JT313OL64eDxgGyyBiFM/DYrUewrjfnG9jxFMPmjyhFTumrjQ6Le7JsXwCtELSYHDie7HQmhRa6Q
IVgm5uh3kDtmH/ML2TfXO8MDxPJb7wBbSl4R5RYy4Y+rsIqymjq4br1FjjvnJlqWJpPdXaXGvGMc
hpg6MMlE91P3POvflywh12J4qm/ISUKU78F5aHAI5aUAVHf7gCXiw5Et7+9szIvORIUKueb5pbsQ
D4HSEVlxlfVZtFcqDGCI6SOvsM1m2v1oNJEtwFfa6xtIoC1BYKCeIvvyGzLqqeX7TV0DuuFZgb0g
jx1svZ71vC00UdilA3W9hbcwqeNdO/94tubJKMwFiPCVqO69yt4vThyoUZM7Z8Tdw8VNHsLDD18I
GZaC/NqVjc+lmk9yB8K97Gk4oCnM+Uj1S0tVEZTpDcKybA/d8098m/6/9lOYpd/yAer4zeWplxmu
Z4g7i/iqdaGCejRWnnqbn5WXVytx3HPKs2SCpk1MTq2dSMKXt1KvmueuGF0bc38cnfWFSsefukm9
yUAGETxF2TOjkP/ySBSC4K9s3p1miEHWtpeAWO9TmXs75Pe+an5GLE7VVFZ4imF9LzW8T1vXKyZA
tKrgSuIggkL2/DcxPwH3FLyRU/ksve6f7hqImtlJLQ25Ae78mIBh0/E0Uw6u2EBNdaBwULKLfvWQ
Ubb+Pz5XkE9ord2GxbXaSRp5C6xpo4UAKN7Wxh/WkTuehLHu2YdubcCXSqCoXF64k/8zStg/DALL
tFOk1Sdm2tBOFLWSqMCetYg0Gu6LS+pBkK41BzfxF/+9be2xCbqKVNvPfaqu1fUXjbK/hKbEt9VR
HIZ6SyBZmwoZ/qL9X6/Bysfk3KrHcR5osV6/I8ToLozwHgMVg2+6aLFIHGFTaoTuP1eWdMjN7Ck+
ySGJ8fnB4Wr3nnV9kwK7TziEy2MYpErk0NORHf8y7LwJYuLfFjjtiWb86CyczK3vpl+lJ3OdHRrR
s6HXIycfrHTEUvL3UFG4UudkEPSkxis9pSAcY4BYeruWpvzsR0wGA2ODOte/MqFU7V/FeRRe4wEp
NhQdDRr662J5kYBMUPWqDYB84g7OC+ckTWiAuyxeHSoUcuNfO+ZvCKjE/VLg51vQkgVBXA0nfb+P
3ToRs9xywE1eEJnhiiZTttgvja5exwYXZY8lyuvnXz6WN5tHFAIukkkFaxL191Mq70Kq6FEw4avA
K31KsAaUger7uZoB+0+KYUV1M6hP8VLy/kahBfk/yv19g2wozlCb/zb4LdZ24jU8QXO/2Y4Q6ZhZ
bziHkgtItwvCUpDcuNh5t3sW2uVTvD8VL0GCTJ9L5MqsiYGcJdk6sZSroSX6S+c8vssTcqCn8aRC
Gr3wOWg5ZCVFwP2AymP8w30tucKNemilQh1/b2RF2gVv2KBaelby49y0idyj1J3j7hMdxknnsOGm
Mx90S8Qba5icKPx0uVUZIEOglHEyK1EdBuFQp0wBDV9gYACbwA9s+HsOhIUlJVtbvOFePCCfhCPU
Ffun/AaihHJpr6RP7eWrUwpf9gVOCVFZzBuYBc4Acq/0IQ7RsqEkxPqkCC7esD3FWpR4lz0Hwm2e
JQm3s8IwQxRv50PntU0Pqga6ksSLYgnNAaE+GFqkhvqCLAZJ1mFbox5GQjcf5H+5Si0BI6qzNlyG
GCC0XYp3fCEHktIDG5S3fOGTVEFECb9Wg/newMB74DyP5seDwjaNPY8EAvsJ/voy4tVlze/TKR3F
zs9VIb9QKgkxHuvdEbRz0sGxqtcr5cWZHzstAttX2A/2U4b/g7G1wIFb9cLgAheW4+21mh2GyU1S
wXFDBnIY+3bbmzKrQwNJcDfwww8d+jaMDoPCjSG7EEZWSaHmwpE9GYI5+b0Mx8YW77N7JiSUZnzj
ZGOFuLrZOpxEkCVvbmPLgET0X6MdmuIEiGX3ykLa2PxLJNG//sPiNBQu0vOPz4cOgr8M1QexdH/C
dI4HhsH6bH/wCixChWO6iAIx5g7RPEMJ37WZ08QVWfteU2GHtzhea6pevQ/cmjElsPuGnMXcp+3c
9Pj4E1MQDJAf3KzeH3Lbm0trd7S6Y3ranuUf1MG+HswDZf4LlGYXjhTpIGCiahNIZrfinX04jhiO
UzgB5iVySLOi2ACeECX6p9eCj9E4kbmvSkrjxlmNo7ghiRBdmNExXKiXL62E4RpakbJPxijL+L4s
Zpn2VKQeHXqjbz2AkqCkINzl2kOGNcDBB9VdrzbgIl8H00fhPMPzI3y5GdFxdMl66+uDmOM4VLA2
e3FjIr5fvL9gr0sTWJX+ycn6RxGFVPn6odmAgl4LWpiV0lWFh637jU7ngcsfnrSz2bO8iqStxOpE
73X53VuhxXJgo07ky1GbaYsnnavgxmqh1flAXDSnnSm+SApGq74QYzXsMpuhRALrM9iWxGbphUdq
Fx4yJyo/UreYIhnfFwZXc/ReSeiJYMhrwnNH3x3BxMsvw0R3F0nZQ/FEbTJoXfxw2J2mPsPUn0KT
SzXCrjfq04xM8JBZyw+jktDufcnvrzjje8NSAEUK9Aqyc7vhBsPy46yCiXCvQqfJPnxrprWFI6RC
nWH/FElkv4Lx55Ei1P8IMxqlwqLa9QG36RD9Pn7rtxRjslrndiOx8H14uNWsoXL3k0rguvU0bP1s
bn79aKuVQ8ClaEljS+iYUI2Jz2/cJkweeekLGYDfmVGOGHsVBdIYUyIABqcxAnEqhTtoW96WWQeG
Z3fnLjFdwZ9bqdtD+zvc8uYpX+P1cmXrZnfFVuIBVvS7V21k+jQ4PiitS/WsBdf2U/mJOUOd+MKB
eBN9zJ2PQXEBMwcrym+q78g7jKJUVDodoMFFl1poJICU1hGnT4LgnFuOTsVxdrjcN2EJ/XeqgaRf
nWa5+mCple9Le+m1N952Hoa0zlAAzMP0qYXdCCljPjftypYLbjj/f30kA2Fp2pyuPBQsVDORJ861
4B75ajPkm4ohxojo95b84RSuumm+ee0D96ZcUscNVa5sl6vNWgkqZYn9XBr5efnv4RooQr2G1Aps
bE4nqMeivqaQ7Pdi4TBcVQXhCRbVvXwblrXTMJwgg3BEnUhMJPcOXLWSLmmeVvVjqFDo2WfdoZH+
xUwBy8LP3VClMFNnZJvhXejlLsLYTf5H7Pk02TArKiGv5AnaloL4S390V5N0RvnZPq9mrVn0JRNd
mQ9zHtxGCFmco94IjpfY2UgNZ/AscoiRzYfJQtgUjJm7hcH17yGI6DeqUoOJZ4pR2vHmbyBXvo+M
kVrUHbGVlwHPMOhqNnGJ3aERWJ2WvuDpGjmu9d+6ZlY2XTJQtfiEdXTTowdv1LxgJ7+26XcDB/Jm
/gi7mVKXjr6ML1lPklDtJqOAXYUe1leEGUTMd8mwCYWowYa2GWrVN18eW44WM4Of0q0o1aCcVBW8
yzS7sarsP4IDUbzuYRixZ1mbJFdUrtY6Wr05VOlgR9BEFEedsGPn4DlEa6AIu5MvoDVGTjzgfdK6
tHvDTJGeB81gq9gQufNGc1NptgXaHhTA2SS1cT44xNEOZ8tP8O4Qs1i9UYcP3asp+2vSaC/wP6s/
7qpBohelfLYmceXcm1Qxr6ZlqcmMPq5Z25GehN/MBbRGfbzYVmIGqNNwhk75r8sqTkuvcYJ0oye9
SdOyFrj/xHc8H59as5cToTOMJrYpnuz3bzksEfQXyyYKMG2akMaNEhbT1GIxemBR4RRtxiYwtXLg
dRxNikE20IkpbrKAd26MSQUrduJBZnLGip3LeOXuIDVFsOn6QPF7vuVOkqVDoYyXDCD7FvW4+y+B
DTTZ5yiLLPRg/TIRN4y0ybisQF4lblzuptKA/CaSC550PA0t8NXJPYQqUzvUEhXgO231XMVLL74T
lgBdFhDvF7QpSysCHWOGc6TRXjviaoQMQk1ABoaAO4T9e8OHnT5jrKbT6+44/KaZuV/AUAhNr9D8
scWXlJzO5cip84om0kSfmDEzszYoIyjuCT9dCJHaug7yI1cTZgkxY37FSzXLCqjiTnW5LLZoOtDR
acVugyVFYFpF8cX9ZWS20vwXc/JMZ6fD1/zoZWv7+oRJRCSr0uSufn57wKdcXvo3qf5QWMhO1E3F
FAsfye+E9zgpGvC2c/0ul1ONdpq2CPFNlio4JsyQoEwYuZ0e9yBMDkGyt2gREe3HlcMr7Mz85HcM
catLGncJGljTwXPFVSai3PhbXbg4lbsWUIIjpt+FSQOZO2aSa+ZUR03lJDlPiTQQMNZZam6IpGVb
nwUNCNlWaI9uO2LpHzQtOzwR813qTDkA1Mlj+qikKcWtbFPXYsCHD+aOvW0xute2Zd8mHYNBL3RB
/iC0T3EXe0WfyRvTM5t8E615IqFwsRHufdCEFCstOg+6cD2FGbAMq3PD2p6ok81P+wMPhLYHYTrm
PkgasUtjnvAtORbyWe2jzVvDJXH/EBISM0uNkwg5Fx9gEC1y/qvXFLTutVGgX6zxYaWDMzDeQqah
6mDgIWTgorZwv0myBRjP0mZmPSnHqj63awEdBgPoS5zjAumdM67sTfPHBcU77879+ztdWr9fWjJk
QM07nrFdpUbIiy2KRJw3ZEgpHGzfcGJ6Heq7OUtyK81EBEKP9JS7c82S3Y4E2JSXelfcvzv2oVM2
sWnDAtkAEggiznmWaQg5JTK1rhtYFAQwTAOFEUkoi7KenVvxhW/8OSym14P0PTocpaBwbKYHEgGa
dJbBJbyRFiLNQ3eafjrYhQLuegNGkbYbHa+gzyO8V/LoUYCUu8ZCUIBOEpvvd1TBojF0+i25KLlf
qiJ69yZgz+CvtgLV+MV/ZwsyWcNBcCSW3kR5/rdbTi2ujUitn3zhUKys59sFBOC6tIVK95m7sQ+A
zw4kFEwAIFZGOeihQqhrlgIOE6UeV3MjBowy20E+UMawVD8LLOKX/ni70o6W8RbUUNZpIQzP3VdE
9/MIKCK5tY8p01cA7dVYpGRYyCcnYNtrjMpcmTGfIMq/bfmAflKlIoeZHjS/pJIyloyvZysVu80L
IUuev+7w1/hBMKzNzHHKgdo+VFE3YT5hZyh9nYXzsDO/EwvU+Am4at4axPcK7sbkmLP2RolZILVy
tJq4evyuUHgvcHXQ9m/kMCG/aTptr85mv+xemQXiAqzRu6limf+lcYlf448KMgFCosjaEC15BIxS
+28jX7v36N2ICeoUaUzsdzuzGUqQps3BA0BeMpcbNOyKwjn4/SSqc5KT00/Oau0Qm9O1JA+/9CsP
izA6Lu/igPRZ0Y9VxVIlNJ6XEuogojfIedV+HJxy/FxVJPse155rzHHEcrYPrXH/jlDWwKwTakST
PgfQVl/+TkUv7gVhbe1Vn+8pUUMvJvz0SbnryYVyZSkAmvZEFFZViZKbx9BsZwHDuApzq2BYnLoS
+l8SARs6jPZOyxSP0FqV9APSbo6CC90dgreiRnbVbutPspd8vORw+J5bLEBWOZYcFBmYPVqxTfyx
hK37nO403IBLbHGG1oYMLJBsg0LTRMTzBNskyNcmK+SuNcBSfU4fcTpiRv3R2yl2oCidB6nesLa+
gnyf8KQOCqZNajN3UYe3RtlOv1qfCUns+74NXuFB1GMkoCBynZz9K1y9URNn5DmhOYfMktSWogLQ
tWWpZCfvVy4IdVbpkjueutN+pCpSVCDKTlnJFxBdYL9fx4p2lZ0AxKexplYMucRz3jY/gRfsu6zp
oShygFayZm/2PVEbdHvIA4gQuFO7EGawLlUgejbGYTgnojgMlJ94klb69hMDoYK0cluc8GkhYJz5
7NHD/QTpU1mY5mpiZvMNDMGMlCjkI1JA5osUj8HZWJUIlNJwP+PqGOsHmgMtvVTOArKkRzi7haYC
mtboCxEtyh3BA85rN6PlhAt0+bQsmplYXcK3483Npg+XlyfCsGuAKM7rcWpkyhz2pY9BHl+2vT8y
+hQZxmw3dHEBV8L9RGKMpRxb/eplVRjE/cLKRNy7N/Bp2E9xM8FAqQtZq+1oU0l2smIYAw4FkMyI
8F/Ca8lY/kTb6VFlWFUaEYZUVhHygsvne5RtVwSSLdKXAgg+jQhBBaUeQvd0EHtfgbdmrtMgaJAr
usfX8xnDgpCPsW7oUEicA7LXCgHYZMWVksKExIS4e/DymT6XCdNSgokHQhSzSbif0H/4mwQG5f89
XZTE8WLFo5tO9lYDONIEh9MB2109FiCmkvvLkGy9oL7ivZOSe6+Qwa+xxKbHFu+onxUn1bxbLhde
Rr5DkA7pVXYFCqKk3OE6xXQUo56s+48s5A3GHcS9psQZWiUZITONLTsMJxkxmpEncb7pEmoORF/5
gyMU7mT/TL4kJGVsSnZahtdLI6wxv4PsaPiMktjEOKtUQ+h6gbTSdthx2PptGVPWfgjVAbic02EW
RCptBSVIYNnmkQT2yFwdbBUC/goVbssgYQWbtoSOAG7BjAx6lW/oWDEXzMmPb3Pmzz1kkRL0M9Zi
Moj4vT08wZKjfk/CGIXjMOKszXInFF4/xyMfkGLHSR77Kv4Z/w/3NbcDXnsOvlAWzyTnH5XNh4zE
PrH0PNhOCot700K/U0+XvPzeCmy8t6SXZx9A+qOZcI4u1UfofU71c853o+qUhCkerQ85LBctwhUC
9CUYJJqTfb/U8BUMe+kb0/3lukjf7RMVRzKpZbvfl9ww7zeOx/HUVXt6Y//SkGjY//Cs7zEZAqnn
zvunQbB9s14kA/9mnkgozHB+h2Fmui2Md6DcEdPp3T4HgyIP6k9n75qhNAWU0t94/H7p/IChmFf1
4VwofsZCkXXLxktwMmcSrRdoINEWbUoDph1/wSE+pv/D/GkM6gM4dGI9qzMZxJDoWCFk3Etaqofk
bzGRPN9z0SYRPjS6KZ+xqPy6PWa1e3+RbE+aFQ2aAXk3a7+IVJ+fypfhBkzZBEo0mfcxaq2x1TaZ
s/H88WaST9py82jS2awGTxckTR4uYfKolb0qR/gUZzfd9KiKShW0L2KhzoHbQtK8VThCv5d92D3T
E090vvd6ls8tmcu/Zs4+gmx8GvqqLQfyjbLKWQiUXOqQhzCdwl4dfjWODadLO4v+aJ4kDnF2AUal
p/ofe66Q3KoESeTLpbtlCfevAQQQiBHNx/y5EDys5AlergKDsFtui2TAufpAgKv+Lo7a3qT84uoT
uiZ8+OS0OO/meIoeEEjr8zP8mEjhNZTUJdeYT93aVNsSTJzQZY9Alhb4BJ8/LQpl7KePmzpRfecG
KiGUtBUkFeoNRKrkT/O0HU5I6oeTT924rjSMAEaRQv1mcyRa5LmWzIhowlGoJXOHW3+puStBWfgl
iO7QJRX346VLxLuV2fCSyW0g88kGMU/0eFQrWb7XAu7qBoVkBotMTfQpyOn5yRgJlkMyxgmhgjYm
Sgjse+MI7mIq3jlJVltCEoOuyd+ZHa3aV3IqdUSe8PBfR7S/xYotf2qI8CHoEHQ0s0e+FWlFHQoJ
feoQilHNk2EY39NNXvKSrpIRFpnmHnjXpJF/k4mkhOYIuoX6P6kPXS6hofuyhqeFo4Qb1GiouuAF
bkVSOKvWSCsCxvpawoqDVy6ePc7effF1/Yo9AL3De8NxqSSFowTwjRFuL3IPvSv9DwTBqOiD6xeA
V+q7WchZTDmvFSN13pIE0PHnF1MJYf4P8l4302uA0SDZ2GDOFqCvxKIVSYy/fUNdGrFlT5cg0+ew
lfOlYeMKZLket6MUaeMnvf6NNY73HTeWmX1ZDvn/Gb4dF1CxUnwl/Sh/0EK0FH2AIBy9xyPXPZ3U
AMWy9wOeGK5jP5Dy1XTOdMbU3wFEbNmIG2JyAzUCD9L3yaROvgkknVxpVv6pnArA/rkfxxhCmdco
JPOsrHTukgHhdrl+oaZc/tIPS1gJlql/xjDxOVPUgjhEa7MWsFkHZ6M9lC4Zgbx77azwyV3MpJ0H
/i5pxAoCtI354LKyDzuzr3ovoi38PJ1OedoWQ+ySMVDVBVS0I+/pZl+YPQwY5WCrmRo1ZZ1EhNHc
iSjFUUY60sWJuZG7FLr6ZB/veNSJpI/xhL4pC35Uj8xEXL8lPeJjBkdWq7VPKqHFuDuD6IOUC2Km
euoEPW/VOmxRg+yj7XQhWqRLcZC3mMwjZnO1GbV/b8P0pxB90PDKB80+IhoMI0vmW7tNcnPEcjLi
bZLwAa9Th1DuTCNi8Z6fKtNedjv0LLuNP6Obp19qK8rt/oyTkuURBac8JfnDdOP4CAnhfRymZzeM
P25CdjG9EyhkKIa3GFXTNViSgN02ZIdUF+9Yps9t04RF3ZDXOuCpB3A1v1nDGMLw3ivnb0xyD64N
k0Eu9VymnvS15jAC5e5c3EE8vBs6GiWPLhOCZf0a7VeWqhzmNXi0LEHwr8zi9shZIyC+szjk4ZWt
m1VOXIW3XCFZAbgwXfBqJg8aDIaqgHPNXgeua2VCWbMK4iCehSfBxxJpivu2xjZMlI9HGPmA9nDC
Z1mUtewxX8jiXXWgQ5+oncE6LMxCz2kuDzO2I0ejJTazma+NsYLJV2qe1lvXyZZo4AnvyiIg9Mfn
E5MzI7gNLAPt9mK5Wv5mBhQzWbE/t/LS/WcqNSVqi9wJNQ3XXPAuFbyYHoR/flzElc9JVpQZ0diS
WeGe0VB0aZZn2UtfR3+6hliU6QBbadiLGduC5NZ3y98BrvIxPQykaKBHva5ifWAJP2xF8zeR/D6X
3ve3WeI3pQNazZPNCo751Cw1ey5kWgf3HmjMdqqmV1LfBXZ1Y8boqov5RQsD7aRICsSU9YUWRTBH
UDuHz8SgaezZgRWr9Ng+ArJmjOB2ttrxYCaMkr39ChtYFQaelYwKDzPVWKwhoD4So5oFCvJhaLx3
3izXEeoV5uWLg+S7NRoo9Hip3jnos7KcF/P3spO57HK0gkYILSEMkqS8xt1dUlobOnq98hJWun1y
BvKBS/WpPVeRZiohQXdlC1FvnUnBS5mlxFrL1vP6pxJfu23FNAd7+p3db9huNTXcO2TztOY53tUX
QZ1eUdVxaZWdpIuboMfWz7RpOjeofCM9tP0QQYL/huWDiSlLSXBUCk4rIxqZW+mtANNxvQB5VTcO
mUp0wPv8WpIzhHoKSagH9+vqDtIiP3gXLdWxG3ERHEwMbjLxnK2GQ6ZZoaFZ9UJibX9BiShs2Q9N
ZTxh9ZE3CbNpRVWAO7LSi072LhnXST3L9neyf0Sf7yZZCV+kYt3a5Pjl0dHGnn9luzSR0m3e1SeU
JaBME8yeseIqfVQ0N7EOe4qqZMPYlU4Dny3RwQbvBnNMSuHQXK8x+/thkLEPqSLS1xsez5er7GJ6
CCy/6W160PcfTyW2vc5GLdjSneGyVkJiRSIWMih/GNfpraDiuMYnvzMUQCW9RuooyVNVETPYJ3aJ
EKt2bvIECn+KZDCerEBjJHH1AbZatdMWiaZ8/lm7TNxvoxSyrpVFeaAbCUGRWX0H6oJtqwrk7fvF
4+r529F7IyNsINEXJpEClmzCD34Bj2O0TvYQ1NlRuYced2NgTsG0XYly/5wRVkcpVdIPC1VFmCtG
PNsC1mI2WaF2C4yzRr8S3wqiAWWK0lns82aG+qtvdf0FcJcidqVqB3sJ8PeVRgiIzrX4UwsQjVzr
D2/PC/EZU98VJxXgvG5lYSAksOfEU1wjWXbR5rOSQrR38iXkMluWLFKlrw95LJtJqKSK/D4DtW7X
BeAn7SSTG+LZlMMWoKFveXbjnAfAykSVe699Zn/w7ioNxnQCRGEXE2R70Pw7IRNgVFiNu5+lQx5l
ItEJtPtINTtQ3uO/ahfkYS+Ca/UwYvn1V/V9MyQYXIJ7+NBV/qmTKp+o8yu+bpN3szItcXZP95nh
fizytSuviMZSYRwXC+BkeqNXvlg+5MBWYkV20OtXsSJ2nBuv+b0B3QekUSuzwjHuZ0om0BJwX1o9
yW3Ui6d3U8j9iLKcA8ibG6v190wgoipu5HcQGsmxNZdYdvoNdXomPPgVbVucoUgCk0t/3BiL4bya
GXm4JLcE3nUW1vz0O+p1CVIdiCRYN02Crzjqn86rGyuwh9VNPYVFxtF/T4MbR5P8+qay+GUqPyes
DTimMe+GhIZMZea/n49x7INjMCRUMkEqaS/6Y3xnyF2R+jOjVghimx1qhCdzWMPAbteC9Uxtiyj3
x5bFFiK363llf3M4cYb1oeMuAoxv+N0giLbe3I8xJUrrMqUBJG8eGuAf0u1SYnA9H59qGbwsBfyF
YTTbqmmGyPMse1R9IEgFgSGwvYXjI//JccYXpM2qZBv4dYkGF51ufdE80C9Ci0RQ/hWZKL5Ge19T
BvlHxQPNqBu134FFCJAzF0bpDqGSH4ro3rqDQ689KptCxI5XvomFbS2hmGq2RbDZJQ8d1dzFf+HQ
9YPIa69arFIpNqN78ewYCdf9fQH8uWKifBC3vup2Ky8xH5ADXyUJwT6qE2uCSxN3Q2UnFDVcLydJ
RBk7mDbzbY6zbdS7KGegsQG/snzsSu0fh0zOm2H4vDdhuCNNMmnOT7TPK22YrX9DsWDzxgGBZ9MB
NwkLn4kkQS6U6nM6a1AGEeP42cz72t+XVOJ0sFtqAkqo/TZEQEHVB/r36yBHmDnT65yLjSl2/Dzm
MPizOH8Q1EL4ePAaOcy2hFyqlTzhEy2CCEsI4OqCs+I04NoDmiZ2MdFXju11NwPvwagFEXtDE2qP
xa49qzObvWIJbbYSBJHvW+caOBaLrwjC6jM2MuYopT0tXRwWBUz9nC/uvigKuzdSD8WnFHxEHXyd
6qiitkapvHCZBUY+PvAequyGwt96atUMVi6ZCqQOki5z39HORZ8KaiH0bQ73W+pAq5aaLCdmgDZr
sZRlKwti5oBLy91Dybd7efId40W6G9lMnarn5aNMtZawfGrVdf8TgiEXDyT3XcN2HwvY4U5mSor6
OpCZPWsKQlPGXhk7QMmNV7QWUx5cQfByJUFkddwIDSklPgVO+ePWIFsz0IFoJqrpkM7CfOh64VhA
rcrZt6n3EpLBDDobOoTMpWeC5PFpctKIX2+RpAJEtQQGDd4v9U12VuGrDrkLBYXEXJSEN+xNxRKX
NGf6K9RFmDAUrKBmuPPtUur4llZ8p29uVhXetPsElaRtYH7SVPjkY8gmNADAAzCfFFn0FIXAkVx0
I4q4eqfItAl+uZbhxyVJNVsBY43TIonkjXaExxlMIx0GG9MCZMR/IBe5h7QQ2slJQZXgSL64i29t
LH3K59b4ONhaqWH9MzK+GRNkahWroHGUnwBJd/muSfDXtkvIlBL4iY1cQLTx4Hic/EB2i4U2uYmy
/sFSQZhp7GSjSp74qGnI/NkmLO35VAiFgdTBNO8woYNjica8I7Td2w0AKmkdldT/14I4dHZTuxfu
3xigOOUcZWeKHTEuac94oSNlkIyiyxO3VwxWH+vDv/R4YZiQ77mfgIZWy7ay3e/ZaDJI/atDqsRt
HbACTeNFHp4zkT+yU9ZTmLUCxc064xIdRCQp/iFodCbNyGmaEjuCuItQnUc1+F7b2uHM17KuTgkC
oBnRXC0cd6SKkl8pshN0pcnphRsWM7GuQE1/OQVHUcif69eYC7TurmAnB5IOSXjbXltb1ZmR8Meb
A7gItscV7EkR+6ieMdxfJo6sCx26EHhaReuxBX4/ZKIq/rZ8wU1wET552Wstgqq8SOZ3TODP7c40
dmPmssFDMrB6ok3ZUX9KNijDJrksukHhufd3imGW4aWsHYcOGaS4SzfcID7HVtF2oTofNw6NiSd9
VOJvfiohGCHgwjnsjFjrHK7n3h3CAfjcCNcPTvv2bWhWgrAbYnX9xFfUgMn5/mspAY/NszRnQii/
fublseSiFZZWOM3721eADef5x4ZBZboIAN85G4nFVT6C+3rWpLJQPm2ziFFUquFV4W0fpayZOG+e
dxBYShjyi3/HlRO+o1m1vCeVzsPQm7/GlMlKxLoU1A9s8sDhkNTAIXrSYvgbmzbxAUEasauMH3sx
TafkU8ph5pQGV9Cc+14a3oHNr9qJgOh2EtP7gJ7EDqL3fwbbqqV52nXitR5Kfm2RjExulH0SKYl+
Zw48FCs4CsI9k9IKTKAtAAwDrvbH42xmURB7sBW3l1Lbk3GfnyCZuwwug+ZhN2y1T3767+vL9E22
CoUtNlKGZThryUXOb8gAzpMhdWN13dzlMIJGGRNXGVKf8vKNcyG/VxWtVYmbuEEpfVeuLQ+uwFn2
ZhAC2XfiWGt8sB0Fml/+DfU7wYVgQB7/1CI4tCV/CjB0GypXhF+WdjR0h0tUgb6JA1dSxXvY7TAX
E2TAeNFqjr1rr5Hc/MZ2dm/BiWcOytU6eadI9PybZ9qP5038zKDCJsgEoUI2Yu1vFoPoh3fPepCT
OHU+X4aiJ5BBB5sNNkZAm+1fDFuXRxyymFKkvUiR/ZT6zIT9+je9vkJkRJW+wGDdOLQu+mnnoCIY
QmhdJMX3g7v7cV4LNB+IYmXX6Qwqn98pDyeGpH5B6eyOFYGZCAaLKvsWclnP5qhOVFBYo3sUYMpZ
w8Sl7fRcDlcvKnh5PCL6qra9O/GXNJGDQWRd9nSVoJCGz9owqpuY7CxLx+VIhQRz6HrLYKTG87Ro
PTOtf8M7UdfoSOQqj3ZN9qsf2g9c5mS5JrgxCK21mn6/BQdDaaaVlUfdVbwut7IlOb+TnUAvWAQK
cZE/XBFIPKgTAjmLwqfWuiPtDjo5inJu5Pnrm2+Oh/VtLriAxfBnWA9JTWhPjhjCTeKazdoLXosn
aRvgKLs9YcHylJ2aG9GDLx8Mdc5Y9LPnIwgXD1r4R2+1h6ck8PL1veqvzFirda8TtU3XmRt3Wrmd
pjx3wnA9/a64R1UrQQjmRJilxcFRL4CVqIJ7+aULOdkiaEyEMtKZ8CGJAWEHuHELicykuOVL0nvV
0k96kzz5ygmBOSzlfI+HKAwm20/6j+t38XGF90DCn0bVT/qyuL5jn5q8GYD4GAhjA5ws0mImblDJ
PwSBZcSlBOVUR9JscjWbQrpubd5sFkiuGgUXqnNBXGO0FZUxz/xmd4ejg+VZgpnlLeYDzw2/7Tdv
srV4JIAdtX5hXjDJOVLSoJIZtd5SNYvQhQKdMLcrmczltC6PA3DREWewVTCVQ+mCvBDBRsxrle2x
nAypFVnse0Up+fH4Pcd2SEZT2aK7pClq8NE4akbbDj6Ou8aeGNSQ8QkrrrM1SAGnkqbLEiT/pgaz
XssraSX5XYTBXNDaqH4egrA3NwFAf9P1lrzb6Jct7r5mqZcdrzU6gFm2e3ZnXsJz3GbzKm/3ZCYS
hR3J3NLRiBbjO0Gd9jm3k/QNnCgQ/yXtn5tNCe1hRpjZlHMWjNBXlaIhRz7krVaoOcUdmj2y7fhc
IrHMTqCU6T3aXyGAI3pe/GlbUWmePXPS1tSvhZkDFRdaQlcEVvhQDXPL2xdrFkjDN84sihg00OC4
zkXogWTUf1iO8jMBHR4s90lu7hEq6IP1zOMFkvW2o/JbkpiXjlyEP3LuYFhObNxXrm0NTdSxz9EI
Yzm2mjHxNk6KCpWW4r96y/3w07gfxNCsdFv3SfdhlX42++OmlvphzApqEEJtbD8scH+oey+FUZft
SGR85cwgynWQSm3lg3cMikadrwhLxhRr1z5XvuaPc99r4NbtA6BolJ34hqKOBMfZOMu99TJ8T4M7
T56Xf6v5OZlLM0iZ4TanaIp4An8/ds8tzHcz4gB/upNymiqahjwgH0ldXfFD0HW110YKxs/Uv7wi
vN6N5YkCLFFpADd0RkAKCHpWrCK63c77916ijMYEIPq1aN62VbZfm0C5+vfSquuSVjNRjvlePhgn
tDiOasZ7La0WImPYIlcMJ7T6w6AV5TdjcQZR8pdZGtCEcc3uiCOhBXHgalwa3pzhOR8N4S1W0KDh
bzz1uN8ao10/Y+qPRryhlVODYhI/TIFybEorCf0B1KxPj2OjCQRlUbYNQmR/rcx5+Q2dHQ/zizn6
uLEQ4S1MFCS2HEE87Nyr/4Z086hkL1oGHx8fvDiGwKSDaRYNAa7E1RiJLCQYoXd8r84grGw8nXdj
rHpwnGjTtXsEHT93nG+wqKtCxLSANdlCqueWVgdEiqWWrgwamM2ekuPxRc+vZ4ulnw/u2nD4ejma
hpPvxQ/BkT49J8ICAKrs8q+5622sHzohCzUgbBRs7fXmZoyF35LFCqYoQDxindyr7tK01cfHsEsW
VhEyrTI0Nb5/ru8GwX6SS7eIPa/JEPE2ZUEdHCbp+sVSPCtg+fgsmcaMEIb8fSlSoYvqFNhrLiCF
EJ9gUy9/b2BIEHZllukROIytx6dvZrI8GQutlVEts7ldCeHgeb/7mCWW6TRBsmmtzwgpoi38dvX/
ie5dQL3LGoMeq5ERyCUVjkMcjxbq1MywMwtvy3UjY47uRNgFaSkVIXLUKxUfnTepLQCzXTsWm5er
jGaeitga/fuae2YW3U1MN9VPPQ3bCur85hCCsV+Q0koR+00szlhWNucbG2lQdWVGCnX7hhcW/lo0
TPkTiPKpn85ACei4l73inbNd+SfPNFeg1nSzTdMK9+Mjt+tukMPt4yHhDUo6krd9rzMDXuO+Oash
aMLRsZMLEhFNWoZSkISDwJwhANIcy/P3myfbb+QOeR8rawq/NE1Rd42g8mXwvIqK9mF/aMApcKM7
sw7ALII6QacqLOhud5+W1kohu/kIgoNmpSaYZ8ULNW0ZNltVz2us4tWyTVyJPvGuciHZ+qWtRD6A
7YQWKP6x/x7wTihF0jaC1mKie0lyWpA0VGfh38S1vrX/8Jape3haEXMz82EVpZppTo9BQyxioFD8
TLh8IEdnhiTG4B1XmF8fxOSqTe8SHJHJUoRmJoM8hcvjIFWJebPUJjzzFug2VbW0Dh7NydrnaV4i
e1EY25IgsagHDZxtXub5NLs9hnAREOLm6oFew6Js4SOyypzKbd9Qc63s8Ks/4NnUMd/VY+AcvKuF
U48ykm/06VRt7qge2K8uQASbEMb735OsC89MpEP5Sz0kM5nKT9MhVXYkE3qYmPaKhSkDBXjNjXVo
fq2QhEAhD44Xt8szt8F5NCGOI6BI/5jyxn4sGzSPkW2ESwZ2pUSUoiKqWnUNmQwTQMyktztaEs40
6FpnIznxMjasH9ObUr299fYLZHhGIm2BBCcgYvMiO63a+DKKNkl5UK0qg3ZA5hzIJsnCwsNl5jwZ
iw2YYNA3CtlpaD7tdoT7MQZj1uTd4g0w7Z6JBNaYC9Yt7MXPTAyw5V4P3IprHIhqn7VPqwCP4KVg
m2dJ4BTVoxBxWHqWdtLwPZU8LLOq1ORdEhO+v1nBYwcYPMpOecnZGgBW0ViBh4Q2VlEiYlulwjJ4
yNCJfK6Ja8LfpcakniHdLoLi/g8EXPZN+YxXC3Q4xAykC9+pz2bH/H9tIR/qYiOZXDaaZ91QjU3f
ZKNzsE+AVern0hUDAEjT+paatgnrkUJZp55puyZbOGktVXXCxxEuU2G/TLCtfJocxWOAO34BMgFz
1Np6xEOB7sPBW58wMV8kNQltk/T2kJ2amIg4ZniGhMzDUY2qaCu9dxAaOFAPh20uL1zPMgA7HHc9
yTK9MmeIhZcPpm8l0AmX3jcCXDL/b0xDbx5bUe8ICAs3NjhlrKABprp1U73u4emWWl4ojK9NhTNa
yPHp5Ov29bFP9uNYLVC4kipwDMIzKl53MuXlE2psekFnIG3pcdw22zAxTZDf9xYsJUGaOX3dNoFc
ZH7tVIjQuNyhGnyTiHZuuFFoMhEzq4CwV2N/LsaYrHju+IybUxid0zzYOIFlIT/rzi/BIo8LxVpp
4FtqdncYzJKd2vORJ6UZj9pcyW9AZ7c8dIG8qtSnvQmvElm2+ze5dWSRv8QJeBsa1P7GZDZRe6iD
diJRhAsaEdZhDPXdDu52I4KZGNmbv0QXHAF9gkSABrxLOl5UC8dUoIkzWduzbG+mcyZ+vo1ADNFg
L3MdeFbk+QJhIuuBZtTwZj0VJ4Oa74RkF2wC68HJ1F9KDL2wc4hBdMOWg7p2TH2uUML/LK384N1/
6DNDloVEll7N/66xWkOpTih6gkFLMOdSRi3IoZRNVZROZMgeQT4fK62LlSab0CA+5LnSil5S0oMt
WyrAQ3RMrlMo1cDbiBOtI117r/ws3h9nN+kY9+B2RPub7Ig8SvclUwZ2QOLLAykiN5GOMk7mjNIx
+AKSnJxI3YG6LAyAF8WW7xCtUV+rZfSnRSdy3BNR+WBe+XPgZzd1AHiPpfnTaS8Cu38qn2u10jgi
VGZ781uGWz0tfk9sWbsUL4jXtQyda25mOAuvlJrYaFxk8S4OBZx/kx8THDHqT83xUYiTtzpiAPwD
nd6q+DFsiBMOVpGRJKvk0BCd6L8eY1xQOqsr3tH+WpHhKXcjccYKCJKLrZzTxRTfR39+HTjPwc0M
/lL31npwfy/yRA3Fn2ocDauRQblOpvWGt1ZEEdNXoB3+a9Yry5VOLdLjI2dAaXL3hTXZM0Kskbi1
qjkynCvqkX4BmDQEbjcmoSfI1xipDLhMX0lzWmLl1/p2HBL0QlrCqwfbnZJZSrYKPYi700uk2XRN
0rLplKpPCSSWO0Fy6bjbczxhDyuF7GkojUzwttD4L1kzWw7k06cep4ZUkRyuCziorQHoSXNQZuEk
oXDA8JK5mrN+LR+SpBVquDXqdlHf59g2h5+q7nWNrScQRb3qAtgEgoQT3MGMVWSKqAsvTrv8vrKe
9QgLK5khDQwOMAei3vEJCo9QSTZFwu8dw1ykeQS/5+rlwSaJ7FmD+pGjqLQsx7Ey+ubJZKOr706X
6uGggHWlLOGgXRSPnKOpXJ3OWv1N7wkyVQjnlBXtvxMY79mpsJbl4xr+ym0YgUvezxtHl87xVREv
c4DsCUipI+enW87foFBVRITb8H6hpj28rIDO6yOS0xAYxzBqHzzVE0YBAsoUO0mjqyMCB00l0lJL
coRDHoIeMxnqHc63Sb/E2729gM5h8d3UDZTRFtUwpFn0FLEj2RDRCjPQgvWt1VHwe3PvSnchz/N9
EX81/8R9DCRBax34VE30AdVK4x+dXAUsTprJqmAnFFgxGvRHGCgVj8gBUHv8VYv0WDUpbZcEZge2
PYEU6lTnSLqfq5256rtuMNLx6k+ZesW7mZcbeuJm1CYZNktbGNP+WLGa9lahg7/S+qvNj77ZSL3k
05Fu61k4y8Y8qRf3G/hcOtHVLSkBePeyjcubWO1J3FD6k90kBa+IPwvB4R+gOko22PS8obeL+aqA
sBwD2DF/NiK/SnxNOxUb1FYEK8Si82Jrb7sYpINfrdhdqG+I89s799cwNce1g4op9UV7RjJvS/Gi
h1TMqKGZw7dIdfaUtdJsHSQC8vcpyLGeEDaSq6R4dTpYbc3ZEUAUO6mXogWSoHm+Y0Ihztri5T2W
5zSLBr9fItVwpKDHbYXDUn7XGlBByW/pMxNCpDMgKdEL7PbJuI6L3kX2gVSOhdyyVXHaKxQ5yDs8
4kvL4zVCTjEQ6QcS44VOb5rxIZZBVmGP2NsbeuU7kLuYFRfVGUBjypZJmCzRq1SYNO523Qkv3f2I
nbrrIDwjhJZRLeksyvF7rzJ7wR2JHLIVka4LbaORGIgMpNJ7SAkdImFNEM6VDcmg67tK9ON110P4
awKnSxjsqz4z57cYpJm2NUWYwrQTB8PN80946JDPU6Anr9LpwVLxHKiqUm5lGnnNScKOv7RC1s+k
wuJkgoCOC+q/esOOYq4o+pvHBDjgxVExgUcOX3J1TJJDc+AzB8JhRqTGmB+jRy6cjTB4AsxfSCQ6
bzm4Kn68l3WF/Q2jsVw6V9Zq6GDZg0HZUABUJIYULb4yf50jwZp/IDZa9FfkI1Wl216Qf8JaidSQ
kC9+iuy1AxTbgaykPsfooqobbgV+eO1KjDxCpQIBgItOGtGGPbTATKwqMVSGBybrpyIqsXUDECux
gLIxtgSxXH8M4K8Gtbws+parHnsd40Sz5JJxdwe6fV411kP/FdzM5w6T8wYjMmuvGRndZIDqq+RT
Ebp1pTeoIUrQMi9ir2b5+uWP3lw9RAM+aSaUCqsEJYcUp/KOTcZHPNCyAv1XJtNx9y685WQYOaHn
W/VPQXNlE+0DvPi8glEhWBZFk8OA2bZc+V7U3YsbCVG9NxVQLpebPUtSVQ/ESQN5F+RXtt4VyHFY
7kDM1f7A89Yp0bHvuWCXiquoXIvBAwBQTGjEArDSsQM/ujSNCDFA0mSZwAqkuMcRiSy9tCswZyJ4
UjC/UH9vHcQo5mNDbMAUs1Yk3TK4pcd8SeeosxzL4yJx0y+v3NPFSDtgfdbnB4WCRD1m3lA4Onq3
bYD0LOplD2oDVIncfUvy5VjrdQZJTn/TEeKYlX5+wvuR6mh8HGk6jCIt5/ZdSPXMFec1NCgCqgvs
rJt2j//d3SNvDLSCbAZ7O9Bck644rrsKRcYqQCchipxMr3q05C09MBSfoQL7M23TwuMY9qK2C4Nn
9aGQP3hfYwHr/M6HhC/eedGCkG/JUNQ8Kj1S7mVr6v3kWOIshNBqoeMPqXyvwAJYifmUhm0/nE/n
1O+nmb7qiMOmiQrA3YTDTjd1z1juBoUFgXi4/LUOtOcRfARR2fKyo1JyK1zyeuDxrctdnvBjHHXs
keAlE72nr1ILlOIs9j4s0nqdvNVjg890R2M3JJ9VbzAUvzC5LLGUgT85ZAZU/9hFvp2csL/UVmQU
HMdDr/4ufY2UV6FNvrjjA25UzlJBxqKVQKiV4BlfzVqzpR+WiJOESxairulYYX0l5I+KRS5vv7w4
psfOuHv9db8fcMfLqesQKbIKl00qDrLsiE3nRe8tD097g90isfhiGx8cqoGYPboylaGLfD+A2f8m
N/BfMtGBBEPA09sPToWaKGdy8PDn3tvNRJM7Xo/FFH2NJdTCmaCHGmJd+kRnHNR5PfKRvr3j1JkZ
Y/nDWlufEdAtIFxioH45Blqf5qNPJX6fAD2KlgVs1Hw3JUVGDNBAXLqlyiJgISn0VCnGJrxPdDuO
NlqkDmFW57ipbT1A5I+NQes2naCR0aaWsXBg5KElVCpbSQbLUmNZ5OTL0wYa49OoUh0ynbxzKrgE
qirC2RVXB8QzItHFcigXcgpv60ewG3pvcg+dv0ZxBvanB1JEU63X/JU4Y4vRLWwNhJ9u4qZpZq5q
qMaBkNDTQ9HWL61A4s7ykAUmQEeBFw6o72/xGeTtxkkX4gnLbuxLOGti+SlcWpFicVfglVgPmA8B
xUcZ9l5NxiOZibUuP40+8MiBwlYn88EOVY9j/DVrqd0Xi/9JlP1I8X3DUwb7VxCBeRZc8pgg9Wk7
ztijABtKqdax4383CMtnqlfgvz2rpNflqXb2OjOsUqsChWCTEqnezVqpEkyWp8lqzZBw8soJKGEi
3NwOKyf28yijifQUJH2FWpt3Zyqn8chvKmqn0lyQOFNQ3WscpaQ24u4Bye17amNYBe48DmmvMnVJ
zbFvmBmuF2LpE4HQi4JgnYwnMHUokWe5QTQhH6lLO78NXjGBoNUfEzUr55cWlHDFuLxaSwiw84DC
l3nqpvK5peiMA3VuBYgTRN2pLTOflpuBB6yybIZBZD2GrmKEIHKXoT0/8Ou7wmWiWQBnC7rgFA7r
eXV+2kIv7zgSI+tLtNJpK1+T5EIthta9t5OV1nX04dXhKDeLeRIIML8RjB1Mk/4fxnPXqMJiRoX5
s+QGZpz81Ti2EWoO3eW3Bf/SF7WTDuxc8aTWA2Bg8Pg/LVv3splQFdXt4M/h/u1iFzGTG/QacV+v
MiytfgeI7JxzFuYpJlc7iJRN5G74PiTn7lBJMX9khK682uwzndn37bYYm9y/8GXRGCxE+gb/iT8p
EZDsiH3Y76Qx42efWB/PQWjJXEvxSrGgw00JFj1gjTY2qFsoMgxnWM9bJG+7xNpExXPmeUtXQGOV
FHTqTFAdplQREnSfAyiETAdulUim7pF+SJmKYK3Yr5RCWWDS5VrIpAIJDdsUBjGMET2NpCHoMfoR
K6AR5XFHDeJ4JXxLoWcUwpraWYL3TGTVL0KunhzDJgc1T2ZSG4IsIgx1A53mRbjH8zsgv6hiZgor
VEzmSpa9Uv1Yb4s8K+0o2yKn3l/vTYgvaPv2JRhD1qjHgY5NRbr5zoP0Te7nASM7u9Mlr/6rQ7Rj
3hCIzeiJTwez15Q6Ujkkm7kdVuxu9UPUTzTSasFurdIOi2i+y8v0MsbO+LhgVZ8txUNwmrr49lLe
veg/0V9J4GOmNmc7mmmScVC1LWVfY0YKfSa42opR2xzNmmfEhFUcG1L/BCIJe6StZXpfAkJWDJwO
s6VADPkTxga3vP3sb/qmbIHbdAiHh5eOPXkAvs+n7c9KfvKleLt7ImLYmrAh0LnXDsFiDfjYLW9a
PGp21wldgbjS2Fh/gbdQ4Jup10SCHL3b0TYMe4mA9PnxsfPIWmeEG5rowJ9rPDXIsw0ZQ9D3zir8
qx7XTsCBCslTIMvJaWKtrAFXKy7Jx7h/FmrXj/oxbEbjIItE0rxYprAK0F/rLg12IFP3gk/oWjqn
OLQuC20RNUTz0vAbefzyUr0h5OCRA4/u2ldRIXHxdFnr/dp7cmgIj74zN/bwtucA/kiiyx1c0Wrj
Bwr5iQet6b22aWzu6Bq6pHswAioTL5aFPoyF3WnVHpyg/eq2ugW4mHq3Y6aqrYuJ8IsD/gWmQL1n
K0CK5058dg2QcmmqdOxhuRwACLpb20MSY62h02i5vINEF3/npNf5+WmRR3YafIHMy7kw12SMZYO8
1zU2ljKtU3/9fUolBr5VYDlKPNOoCh3wtwoQ21Nfzi/nKjIv7m/kXypikV14Dy348eoiOnbGePzh
1JqWItumzCKzQmJXFGUxdp7LJ3A1hfYH7CtzwWCrE7AxDKj2NWIpoTUgVIzo2cAD2J9GBbRDrcFG
5e+bp4N92WUB5vXkX0J9WP/2o4sqIyCK9EdyhSw/fd1BJd0h58MMk3YIo+C3aypqP3iyKcQfiSxR
hidZl6UI8DxIj2Ml7H00lNL0m1CDthBuV4uMntGC0OCpE7q0RA5cMmmiLf0lKrd9W7A2XHkgVZ9F
saqNsu7+Eg82+iaEJ6bhw8iTROxoHcrEcc/9pOxOQTfdT/8SZeoUtrOlPIH/uxdUhjaTBPM7gu7K
Gchm2zTydgWmjQiEA1Av1qFQdrjn8HusyANYLZYyre7LxQf5w4mih/Zb1Ib/xXSSidT7T0utA6Ti
6Pq0uhuIN+CBxwk1nSVl25RR3ViyYFTl/cjQ5GCArtlm1knBD8luwi8Ky4abefnyM9hXTuGSoljg
XEIovhrc7sk0WFlBhGxBu78QPBCTlTKKnpe/tBh4LyZTzfNWyMEeXBXKLLI5PvbhpnVIYHtQsZbz
qzWY7PDBZpT89X9/gQ/61E4yiVlYWe+pnul6/9GFB+olDWx6VFUYQv+lz59D9JolPUs5lS9vgJX3
Gq+ZMRLRJfoRCyeKl4UvVncx2R0YsP9V7/k4eF/Uy4Bu1u4tgQUghxTEGnZfEW0EKyL5kETHvo2h
P9H+EvP6jGjRnIXNU33Y9MXSXRnKHLs5VG7NuyUj0MScymcnyvAivuZncCJFzX5KNR8jNIJAlpXR
UWZr6kFRNYweOKZP5nnbvtn17t5KVUumDktUYBMVFosCLx/d41lwdnuhoUOoFHCVaMBQ8/DmDp05
gMySXpGWu2g1pqbJ6RLjGBvAuaTgf3U61M9jU5qJJKVIbWcN1vKb0xmSKuHwVeE1a7nkCl37uVJQ
4MfFtye1YD6uA5jbMAWdX+Bw4MA4LfrC9deZFFYhsiZbKa4ii6ejzh4eC58pqM0w+U+lxaZIQd2R
bmE5abhrGJCT7hL0wY0OE4pTyAyLv3MIwaVFqEHqxX3QMiWZbC3spyIiqq+R0154XSnc9HvX8QPF
wuiGp2+G6kKqPyD50NmWRiCqccW9XeC/yL1KAW7glrKfomoyq9nM309BwHhTGpl591nmwL6fgVeI
25WmATu1+Eb7uamsBYV+7WjnYZH+1RE1aST8QMeAmZCji+LHEGdYb8us+bfUyvbAgwW6yVHshpKU
QDuFuSUWMsAdL77kXe9PjFQP/nUY9AKta6ZAqeFr7ZJR2dx1upgBdtglbiWWWTYy1yPdNK70+zbG
6Bm2iDfzZUvUn1b80PKlZVDpJ+9Kzz+D3C+kGAbBnb4TvSoMmTVErGrzMEEAbE8mlZL6WqCnhuzj
adsXjlCCUlM6HxRnq7hfuk4cRiarIvOsfO/Dr0wWNkxfIftF2KZX2wuYNBaMoM3nHXvgzLKlv3uC
160yYW2+S0RWddeHnzyEBDIvDxRK+xp1iII4LKWolgbnHNcSMXdTGSut5+/WvJ3r926I7sOVu9HD
u52p+nVf7R+zJ3inqh6wNHoyjXWgAZS9ZCwkNNIs4LTxhsj4cj0DdmH9GsAD7aeP+v7qJqlPmnMA
rAKNLEan0KaYsnU289tICHSIRAjINcvU0NduTOvCane3FbNbGyi6xlFpxQvYJWIhR5R8a5sH/j0O
ALeuw8FE1fx3HkI6s4zQ6t7H2m04t7Lha8PntnWs5AmyLZMQ04XEYDlY2e1JNCmjnkMVGG7O4yct
bQgyFWgQ2sAergdvkQjNk9S/52OyllicK31inlJyLLXx6vZL1FzYCJu0khUpWqGvGHTfnp3qncun
quAc15SneQeKwK99uJLvDH39fE2uvKw1qijknzM5b0xtjZTRGUw4kRPwv9UcWDf5f5Ni/W3g0kp8
xU+3S2Ja0083tAfSa9LTF+XVhujA0man0Wp2rR8GMIeRpmJgqrFCCIpQfCzk76vNuc1WI7zKf+sl
SOvgjx7s6YKu3wVBANnc3IvYbl5bs/BY43QwjIER3gPtv/AtEV/v8uvjE4oXpc9B8vuSodw0r0F7
PRZU7XhMpvWbpsT5cZHpDx7UZrDxSDwwQLzfIk9CumNkgE9wV6YuNUVFACdOEOF5ik9QetfCkNts
ckDRtiPJHW/azW29MqWx1v+pFL44+EDuADJWAo5/fkH2DuXxUsPcIpJ/p5nQMY/Pj8fb1X+atQMH
XtZNfG+HXHx89yuVCtL1BFlr/DhPDXkDdHRPFbD5FpoFVmLzwP1Jue11UsD1bB1lPf4BoVf22DE2
YXKVUscLK2b1ZZMYvjgotOIm2bImwIWEwJHza+vorKOrfcFtmcRwQOGYtG9G31Z8pZeUS9HLhlPQ
boKVVe29/i/EjjDFdb3AMzkbYrNacFXewJYMfPRLA+I6IuuiwrB7Ck/0c7WXCeT4wC1pUWS9SlE8
I6dU8BBUmiiTYRrq8f/h+1UiplTnd0CBXmQgoEBkWMYmRAqbo0775HkQXZ+sSZ9pY1aA+UdsbzqZ
wnHGTD7pkW/OkJDWZO6MzbypniUGS7ztdiCER4h0qFjmXX+uM9ftdZ540HOzhJzrq0Du8uAN5H80
dVLiHfCsDsQdJwMJ5mut6AVAIWMrb6yMEjXUV/jc11DAxO1KsF1HitBCHKOWFfC2HdZDnlagO5A+
mR3NULUtDFhHwNIlxNzK05X9WxSoFshyw23wZpR41Ob4qXWZL9NY3xiOmOdnpw7URm14ZQ+DkW/6
6gAVFLEC3xAnGnVtgEw1aXHqdh7m9C6HkERn1zqlO5iuZdV9GFswtWiqxx2U1H+6vQaFK75GCMyv
/+XWgHHb95z6teZsPvc62IYncRdYv5mgZFtnPr1RlWYqxMxkF/uAYNjYRPoHJz3Ih/DsYXkt+aN9
A7kKHGJlEvs0ZqBXIb4KJzj72VWJbeK3W3Y0uV2iH1l/aOiBIlf5i9tuti6wOZ8vv8w4UsH78IET
2WKhT35G7b2rvdcE/u63zkaAZKTjJyLGWlfZ7h76URjVUavVEYn8OLmE6XlTfk7X/rKtveI3/075
tNLA0y3zX6O8HWtqie2sqnH6FWjT6XYHH1nROdDuYZSZ7WLMXDQvsmXrJlD0cU/oDi7RlF6s8xmP
rGwg/N+nNaW57a1x2GsarSNZCuHsUTQQYyDODPQDc7CyVXVy8kXzZug9NeN8Y1tgAwH4oXU50OQ3
7Es2SQq4JKNoD3aQ4HMyhtXu5+jMAPBMVEzkuVs6eNHiA8REavW4lT0fhBfY4uOQjJjH1vSIFFbx
HJsIQ1uvkkWtXO374cACaEuZhjCMH77vr2FeabWXWI1roSeBBzTN63XDwHAUa6bHJZ7DpB59hPmY
nkJFcfDB9+1B6JlOM9dNmbNnqm3MeeY8x6agSdG5nbOrnFGZJh5s7Q/0NOS33RwQnKzE4aWaoQuq
XbJ2tQcE3EvqiwedHRdBQ9V+kNT5EOUIxIcid03DabGYEwaj5DjUEa9e2D8WcabNGoXdP3j/1WkB
6OVS+4mtCbocFwldbKxwSvnmBcnWNa51qio9+nOm2KnlkSqLbiBgu6iY/QFYWHFXzm8S9FjBKAB6
PCrgIdJBPsttR8ACBb9lUshrk7qDkYXpFCUve1nvlWK33ZcOvasZwIa62dSnBHfdA2gv+dfj8JvD
fPexoG3du+dq4+q+oC8YXSKZ0UFgCtRHK10asSA7+hCwIplj7sxrbN76xzQCHrxV9FJ/4MYH1Wcj
fB5CMW7w727uKrpgrEQl09EebXgoPl73QlmgBzPQ5i5X7qNlUhLqYxX3jyTHkQrTQ6aiTSwPxg4b
UR2flAoDmR1ENnrAiB4jNnSU9HWKcPmRGFnNRoSZbzurdC1rcpsLZAo7nwQS6dccJX2flTZB8T6H
h32V+nYgHT7ZAzGlV4ubG62MDmnjZi4NxQyc3rNf7H6jMDhis9ICSI6VnPmXQ2OJStXyVSN/xhgO
d2KseLzXw/v1yha160ffikPvtyjUn7nOirX5fNnenZp5icnNRzO+RTIzloOdJDIBjRy2k7ZboJT8
elGolWs7bz17Qex69v0VOfIlVOctmvK4Ivlj8v7w4Ns+9Z8DC7EOod2a+j0Kl031E+ekqz87hrpF
6xksdpiVAYredFGwJfcs3QrOTl4r+hwi3ZlEzN2HLn1bA3n5/mcQGXveJAUCwcWGRNfv4/wLp98/
MgnclwQE4+5zG4ZS9SUnLDS9eaFtTk0YVRtNwthQFMI1w4lrYf2vqXMFVSir9aqmuyqREfMV53wN
n9jq/r+u4fTwDU9aGOvpxwFqJxFdYbTBcb0ThtflBm4OCdRmZ84P/ZxN0K8WPgjtNR9OFQIOLy9c
naQh3lTg8kUr0du4ACJb3XVAn2vPVCgCC2qPER+VkgvQZ7KiaXPo5aRoLJ+eckMq/yCzPXdP7KaP
M8HmIo1dpsZx/4yafcD2XsAYtU4Xvc7Ak4Nl6M9VZcL1+JZBvc6VuSMa6829Byzy2MoWPt+k1tK+
ifeaaKDLm7zxHi5DtRwDAZXnJ9RqJEwnVPRCbQDj+q04tZpwhxY9vcs/xr9udX3wNez4oJBo3res
AD4C+zMivaL6Op7UMPW8ZfPobopWXJI+pk7fokEB8cqUHZMHi4YUK+3/zHWRAb2A+d4IX0ue4wB+
gvsN8AzdLGYQ3JBFSU/N6A4GIE3O2jMzttkNb4qyd18KUbChhzacibFbTkPzPbHprvUioC14gHzr
JolMP1iB3S+RzT0DL4yXtRCh8JS9zOqztJmoGQny1CF4N3Ns0pRZkT+Wk9yg2+TiO8KCVUYVsppD
sc8Of29P/FoBIfUfL0V5DR0FNbEEu/9TbLcJ+gqe6hlHTimMmz4hNPT+2ORvFHLu58pWd3S72RQI
hzch1VZ3fPtHCY5xZcNccbuMFvA1rpXIsOsF67/++gjUytrrsh8riTqHg5tN8hy9qk2xGDfCkpvs
pANv02r6DaiML9eOVRljwNhoiuW/552SsG8jWdZieM0SgLXgCWM3TC1Oy4X2QAADpnw+YbEzeQLq
x8Jl3Ho3mOBSq2M62yFVMpWr04ThofWIDD2ZTBN/5ONsD0ru4Hnc1b5uUX+0U+xYtw3HqPvCAyst
OIbLdYSkh+budokbzowq/CraVUsQMiNgoRdPf/qfqfmy84BkziwQWa64tRDnh8C3G6h3sU0rKzUj
GH83zwZorbRzg8uqMRV8FYRmewYJtFApsKLbBV8JNG0GYXfkkNT0m1YCLnVbNN5vhTgHIy36F5PS
P+64bLZG9M9c1nmkyZuxNTgB849gWxHpu8s4KluYfCInGXUiSyfT+BrS7zlzPnyhyH/umMLvRFt8
LoowBCN64HAhWFhupOBM+atMNNxptr2SzljOdV5CqK6EpdJhroL1vkTRzYLmCWMjIqhpBh9zYq64
WQV0KW0XcoNYCbkiDHZmhoWtECNF+F8T2aT5Hh3n7L0OcwiRTar38XtKUf6A0jJSHEAd0j2HgeVT
+o5AwXWojlsEe54N+5K3WhU/XMy6L8cqwIxgHx6jc8hpZ7wAUkorpRITH7shEAuLeIi6tViJUsjG
IdooG0KaMuOkzKeK69nZut+J/GFQCFHHDhqe24zUuThV3mvipY86fvjj2A7FVKeupMqi0KV6swTf
AASD+jhd7ZlQo01bH1PHs94q2odty6shMnfm9ouaQFSUay2oo4qqs1r9kArto02SvZmB6RDkOLAC
BPFloCg4vwnfatCXAT8KgnrKpnfG637wtiVAS46omdu7Y/FmaOseAY/vcMy8+eFKy2zkaCje6k81
2T4+gJb3T5Ez9XOxBcUgiIiQWh30OOWnfo34dGlriYX9+/O6I8+VYHBZtdksTeze3GSY1GSuBlLZ
kFGR17TEyx6+PPL2But8AjnWB9pS6W3ShXMR/ZWAmvoxO4fZ4qQ7chDSxOrFlnA7QSZYZL54geRt
c+Z42d5BY2QjiYVCDX8QUpPQAuOAWl9vMSVduquQk/z+jL2lMj14jkyZNNjqTeWqJQ5d0pzEkIdx
73XJUWXEXZ2F8Jeuo+EG/n9g/euJnsmm/xs2XFkAnyAJgkYT7lGYamPxdwOCSuWpPAshQtmLT0iP
G2BGB8dvF38ryqf6AYpSVSG0yCgoT6IXlqBFM4/m2vp70rz/SBoITLOuXuh8xt+d+p8PYNPgqA6Z
xSRgzul0zROXxWH4K1zb211B7KHQDWuU2EyU9bv3EgfdhV8214H13D3sD6euBpYLE1WDcelfADgQ
1r8FqUc0sxnWZPkTWTBrIsfgM8iFHwtCOIptuPUiGCefQesvLM5J+1nA3cqGQKVORUpBViGQTRSw
KLHfxPx5MRREIBvrQIpMAFDjj0Ncuxl0DGZR5pWGSKaRPUw+kkfAISha26QkwO+f4qEAmjES0ZKc
YzxqjMW1ckgmIUMYxFFmK3eI+yLUo4dDUIrw5fdjttppWILmyvgs4caL43sZETsaIrTt1LivUH13
sdTdNHSeFWbwSVFqlKtzEm4Bju9jd0mOocVkLpXWyc4Ot5bzA1OLW5p5PXLMoMYWY9Am0p0NjrjS
Hnwb1IszuduspzQBir905Vx82MK89Xh2bGnUjyR2ZG/uoMJvGNIisXSqlJH45LIfm2zTONL/8N4w
tY91HpqG0vOMvbTJ4Rfl2J2MBQ1zXoADiJ3hopJmvO+Rn3eeVK+H4XxZdwG+Fbwdp5wSTMmlEbio
lEYdKpa6riiK2SBoJZnKNBAguiHKfDTsf8+At/Fk0BCVoH8C5ic8V1lpQCdZdYubN6ylVuOTeAO8
kcHCi8Hau2G2cFH/U61plykm3/TyJ+AA4bvWyy+9Npr5KOKrsMG+G85gN3RwF6XlZtXC66Y7sBTj
8RYtCxBheiYVBi67iGauXWmb4XimiLpl4hZYjn9cWUocr4V/WW7wcewPhCMeohuhc2kO1fDKj38U
61bJkMaNz3UHzxJokf7G/mJPIgaKJBWQDEfh3NvppxJLUWZcNGPiauRNRPtMpmmwoix6ddaHOQh8
aAJeFk/ZoJXqQY1+Qk5LhvQJDZiuW35vfKz70wEUnPIwDdLRRkm5ueEDvzHQUmdm1ZCFYfvhczV6
fB4KIT3PCHSTlxMqJyiYOAuXLyeL0cgfjDSUe7CAzPxPHg9BOcaWQzpp5Qfra9xJ/XXddYXEA6W/
cXptZuLaVnNtHcchru0JqCUhQt9/wzcA+l6SsArw4Y2W84CXqvJonsJTovYpk7szysV9UIfasG4H
OITy/yAhYNHuqC9B/yHixEr7IXbR8cMX1HqyEWNt7Em0KsAMAswa62eyzhJw8KkM7SQ+fXCXLZnX
3GotAjVN1AhOaiSBVDDPaTdRchHU4+uHpu4f7cgk0nviUeWtQ0gcf77qhULvDjX2hBmd97i6RUMm
1fzk+jZv1so6MFky94svyyNjOeQCO/1Fy2WZKeDNq4cPunFRV2Ti6b17LGSeIZuez0Vu2zKPWxsv
3oNRmiFgQeDp+fV4cJ13TTrpVI09SgXC5MweIcbXA8knHTDW2Y5G7gS5MxK4PmkSeMIDjI8SzgC/
Iu/mbgEHcnEIn6nzcaOqQ0l9pn0evgIAMZGmn+tZVnmoemeHI5++kDMEKd0d+GF0StV09GZ16cj7
4wK3TnPrdW6YrennAH+IQdgfQlpj0XTXD/OWTEYm7lXsrvp8WHswwVpBP7lN1VY4ayqgNQfvDvJh
2zccAKm3EQVGrSCahd44IGvYrryQwV+36q5EnY4zdmt0wYQWtBbGOM7hnm10dxKblDnUa2jfo+1k
I4/xTn3NWhZrfaRQTsch1sfIXFeGZR8iANACBI2YnIow7p/6Gdj5Y7ZzxJcW8QwFApGMScZToAQv
9vXWo+eRltxgAt6oNj5bruicwc/kfjGE3+CD3uCljzm8HZHGlpIX5HjyiMht2gHtyzExi4LW/aIO
z62nI/BqzLCRpUTbVSW4XBPQzL5B7ip+U7dL5AB7wyGtg3qFCzSqdDOGFZ73Y5a4WTsDGDCbwS2O
OyOHU2+i6S5uv4OW4pUodZotgCPa+jnVug9YK5Q+i3Z1li60tMdSgGQv4BY72bkiLtLQjRudStpV
NiEMhlQLCJTrt8qVPKB5QwlopTG8l3f7eNwlsjNGjW5Wdo6qsFn3fLnU2N+6XJeorpKTbv3TN6Lh
M+XqDkreiWuPMxysgSuK5FSiWEih+kYDS11k9S17mcgHT/cqeXD2JF9KTb7nSBsb9UI4w4Ygqkne
boje047ljJ7d8hlVYJeMUV6ftz+buUyjUY42SiVlR8ZQGtf97fXQoCzcKbrV6EVjnrhvMbCGX53C
PKWMwCFjm3M3mjRVwItBxy0VaQsWLZ/RB6Z0ygTTPC7bvMjR7Xb9Js0VvnizClS6Pd+YeaiyZKV4
yuXj5mLePzs/xp0HZn06nUlbVWrw5iQj9UKoleSrO84yfzmznjODA1G6EzefEMr7xzBjj7eboz9l
Cab7ahKn1jyjOHZ6cn1OEghAgn2qLKZ05848Mr/+8VPtHEdhTF+3YsKiAxKLrDonmLiz+7V5glfD
LTlVhI+ZZroOteD8582tFNFsQqA1tI4TlpH3wDpxPAZ62caowBgWeKR2NC7kwtmov+kYW/b1e5o4
STxQKuLKiCNq8zG7w04/HYLemz7Kg6dqTeaNgdKtW88d84BIYJbez6qK0B0tTNzPyFPUrYRvFO6b
kwst9gYhhwGuMa8INb5dkSfNU6GoLbtncyx//QKHDujIX2pPG7ci/exaLjJFm7PrDo/iAmW1eODC
We0pjtwK5yHkRYNXhK09Wj1DgTApV7QM+gy80rQZYSUOEJrSORBa28zxtzQwoHayeC078tmzbUAM
ciosUVHfN/0PJpvRccCZRyQXD+AV2f2pAETsZDKqH8aCJzexZ3CkK3zZlVGWvqAW+JpFKpTwyQkA
Z+hYrlNU2Tg3nk7Ug8egQN3pY7YPZAOtiDM+A9L6PzPMrm/7z70McV/hceNlA10BuGbzmoTNfFON
XKeEfniQ+v8RWix15cOmZM6w4rBRTslpJNMXy5pQIUiJaO9BvgU/FJEhA0sfIGXN++ZNy07YCANS
ZnyF/SgsusPlSgOIDHaXendihyT9uOCXG+P/LaUyE4mjy4JbbuNOZRzTSoiHMqCIOxxC19SO2use
cqF/gdV2D6sh4wqUwhF1hTYDSopTLVt7FrtMWXQSnzeyY1EEntAdvuu235NI+XU3hFUEZWXQZYXQ
8gIWcIMGVMl3p3JUGbLeqWYqzrzUXitXYonP4VwmlCMJ3DCXW89OyH6VOrMy5GqQYZODMZM365PG
xSMFNpVjqYOhPAmXc4cNCoAZRHW8P5knB4B2DyTXuXoiTz0cVEFGM/byZOKAtM3Pxxw117+Ve2DY
m9jrqZxmx+5gyRG3MAyJVpOeCe6zNBzBYh8w+lzHkCKQ0Fx6tMvYGnuaM9DBDXAWoM2GYErLs7dS
aXK9FgxXbmxlPuSd9PKoef4uIKhyGbF/zNVMGmYEujo0usWs/XdmEi+D/ce9p6WF29IGX7ZSNdtK
zAx4mH18zjjscaCmwzOIa6nWwENgiy0pUc4EtHw0a/iJ1KD0AJeMDprhNh1W3GWqh1KduTYSFxYF
LRDlJR7tfJ7SAP4zZXu7B0wkMbbrpEjfQKp1bkCFvxuw2nkZZPVnCNMzROeOr6jL02FUIP7IqoaV
/M4c9F42gR6FXrpE1tCt5/rdJ0+4+mrK+n8lNMwQTVjSeCCTV57E4dMbhB30NvAlkK/CVq1K0Gjq
mXw/1EM7/+GEyZoDbgL3MmGTWwhL1GNawsFPbK0kiqz4SU4qHEucXBbvWJN4LeSM+Qd56PjsWo7T
SntDsEL8eG8C2aNnJWlbc8xexnt4aG0ZKwtLS541gbIvqGOpbSCl5SoLGGTsOW07yjY5jAE+eYX7
s6RCDnrTh//Kchn+rq6BL8N7j0CtaXcFFVy9cYbiI4rz6EV8xog+L7fjHFrkpYskmQlo/H0g/u+k
nhjGsVNexXZcnliftRG2ShcguziUAxTXRWLGuLxvVtNp6qLjtQeGWu7qR19NgcWVMnGxe5suI+Fr
4i5//QMQcFLSUNk8qNx26s0kdSzh5gisrdwIl09zZ8dOqv6H7No7Nd7b7Za5D6xA8TMKaYf9JMPb
9zJbKPx72LqepnLdmLUg9y2HEjfrkUSv/8gQ44MR6qTOLeN3lIvNZI8H/veWG7yuoG1auV5dWADi
VLUm4bnFKIN2DnuSD0N01/uPcZOPij51t/ly7aoehXxWf2mgFW5fW8QDdsLJOBZXJYtCKTNOcB3C
ASPna7BZ2nGXEXim1YR91+5VvZYaoS/Z9lmfC1dw7aMSZXCZIxbCv06bqosTNvcfSc+DVyAPu0pu
WwBsSLhslAtUbecCII1al+FWCMteEgf4CFM7i5Sv3tbiZDsN+Mu99EHQzwlilWwwfccrxTnQwZ5i
aSe6m2Q4SDCO1OmVCZ65wzzJAJdNiUbGzqxcN4Zj4VwWLeOTKk7rkT2/FTdzxbS2UpavFiYh5ohw
lO95fBMXLB4Ql0ra9p8Vhx547Lvqyh858FDT+KewRFJtjwHLeOrMulzGUOYht0qH+QBONADW2JmQ
yZegfcPb+KmHzptKrbiLG8XOVoD55vW/8cOGybikouSNbkgvEqK+Y8y+77ucVWKIP3Dsbr+76/Fk
ek2cdNVSnX/YL2d6I5zsa0rYZzJo3+FZegILa0U8ZZopaPnpg2ePjAo+dDyy+wbhvBduujz1jvG3
2wbqto15U1HI0Q6mLeqtwnrdKatTP7OzJC53ntZY/MJIKDkWPoYsLUcMw1SK10REZzxhXxWxX/sl
nFcwbLgkLWRCTX+nU1SprC9CNoSteIdofg6E0jZDb5NBMn1iYT0nI90BF5scm6eXlxCoEilw0HuK
FLQKOcY7aomxF6YYV49WlnGGvkbXE2uU+JucjD8IF3CzAl5y9nlagxwiQ+F8iBFedIYxqJ5bvO+m
iAHRKWZzZdUXc9G4mB/T3XL0MJNfQkGyIldiU60USqr6sToW0XHR9YAjCreAKs6erYin+6UlMmMw
fgjYBa64P2t1IZN37H8kNIjFcTaFvyVE81OsdAXr3qwrPBeZ9xawMbuIW6ZW/NsN4jcXkaRp/Fjt
qNpuKnzrxNBquW0cC2EYbUbJp2kVzG+nlx7RGWkpDMBJNEwKBk4QR2uqcW13YSpdgyLuXEmhN4J+
R7QeabJUavAsuxv3qXBAzbMeryvVoCp/EdZ5zQAs52olBmpwZxl/U5mk4N38QUvvEALT10x5x/nD
Li3NlboH42Xrfyz5HMwxgNc6McRjaP8Cc+LwRpbf62PB4kG6zcBGWlr4PHSVvIs5+oNnkbTuDZve
ppUeQbkSpsuGq/IWmkqcXTxARI7W9xKTVBURd1OmewmpOxltt099HI3CHPFnAhP28KVagmqCGVmD
IKPAIEyOHYreflohHTKaZyppha763mVf13Bigi7wHhJoLxfxbYLcHquGfd+JrTNsURdHuIhz2R6Y
ZDf/Kfqo7FHnVQjPSbeZs2jcofPoGpsrqwalE57pP1MLqmN7Ub//TOSKJ1DjejgN413TGY5TBsrU
v9JH8EgySMbsV0CmQoWc74FCUHv/TQzvKF2NtN2cymmhigKwTkmU6qHvMJpUX7TOFJWPVMT9obsm
aFd1tK4dbWMxZUqK13ET3xOjIOy1jtvr5WQiW5m9YAcUwh7P/aIy/g4Ex9I6BznJOMW+Yjkjb3En
KMiBvdOWxLj+xHRbe+CCbkau4TMvFgeg0u1oyWscDjfpOMvUxCSP4c2+FtS+EwaEiYIaldBKhSMn
ocrH+RC4qoijNmXZ4a0YbrUYqUXQKdnhcf/ksNXuPkBg/KvhUFo5w2MR7P5hWc3NLKASBVflt3hC
3NW6ZgrKY+ujkcrk5hARVdbFF3dGe2aaE7h3Um+uHwiouBiEPvv+O5NVicr92cfxOKZnabyn5G9p
WYZ0YAvh5qMCdNJ9K5RvqH73dKqZpzTIbxwyLEv/PpknLGaLQ+RsBRpd3DL25Jfo6V1EUTwawJs8
CfuA0CpEQxJzFwMr8qPUIv4dQ3jNeglyH6pOs5If6XMQa2nZ7OK4a6aen+knTfOtO99LBReJCs/x
v2LLsJzvE4sbt+HiE/I/YmxBkBxzDIiPyYDCvxlTwL0aLNnziZ5EOlkkjcXOMGrhbTwSjufSchor
R4QVoSthEYVBxWoyVrNGx2qEdfs6xOfX4EY3UCjlRNyorg4q1hli4otFJrvarowW9hIq9rxIkwiL
OPoe7YbSZIoq9NnZoBLA/+S+HHgGT0itQjTnnRKsK6z6ZGjMh3yqLQuFuOJOvLXz5Fh5e5EEnF9G
MGM/cjPuSbhhre/Imxkf1QjYEGMOraiR1sEjR9E1sTY2PmsMrlPJHDnvFCeIOuVsFU9A250Ib6ZD
rGo8X1uGRelooo9aWphwHB11QzqVXx14x9GxHynDp1UHO4CviBsTjKUAppixXop1RQtrucClh+Jk
nv/o6e8nese+Evd7tGhWelxssH+tAUJZWNpjDKiOch+RgphjMFTpzMpS06DKUdFmuIUr6nc6WV1A
iZb68U3zh5GQaD4aKsI7oId7iw/Cl6D66NAxQkRJ8aZcKuBebgg0XmfJkXBCJfB8f5M5shC1musX
3VfB+2XhWSfwT4jkVZvtAS64FNBq+L0BgflmD76ioS4cwWwMXyP9wueQO4XAW3bX9tUmloqlJlA6
Ml332PplXhJ/Oisf3oDcEdR+w7QELbmc4EGHfCxmHRTKTIGgs5cm4kF1D52idNm2LRlmQZXyIcor
OPxHIBmX1lkslIBz/P00qAhw8uEBfOZwohi8uh5liZnairJOcwpFp6WHWVQwFd9aknN4x1P4WUB3
rtARZnlSIfedkciv5UgZFbPYamy3+1taiPYAyQqtOdEH7ksxCSoOPR58GITzXyDiH1V8creszzdj
YTbx1A9H45fMD3nPk/6cw+oa4dxZINL7SKNesVaF108QL/SE8vz4diEUVtnzpK818LoSfI5RmHGL
NGHC6zYX2UTAxqs5ZbGKhrq/AoDks0oHCjYj88DmjJNTOl4VCKE6sNQsG4NBS3U/U4lYlca6ITnh
KzFPYM05hKQzoC54/iC0kYlbcTrmKXCQyWhiom4v9KEzTGiZ+eRhqYg4WqHJuCEgo3m0ycJogEFX
haR0u4+QyvJR2e6jeo6pb3b2gRlIKbTlyx4BcOMllz4YAKLkdYcqAtuL4od1jvGnz6yanYrlpcqP
Fqfw0lpwp99ehSlBIX7bSej7WWuoHLg9f/2/2FXfQ6zo3QSVXKcDBfMGLDilhV0Xxqb0Ci4AuSmk
Jfwks128ev1bQQ5sATBk/h3YU7QY9YhbY/cEDEmHwZRPChPR5BOvBQYHB11Q1cs3db9AIC8FSdwE
ZdlhJdAqlT7xssJ6YCy0CCotMwqBFP5tjZbzpowRNpWees6m+AxDgqirQdnADfo/RGdk6m1qOmCt
gcsGl+zEUBez0aAPhAjqQS9BqTeAZLnvXCJxrnYPRAAJDqNrrbuOiN9M/jqM93AE4166HU0tQaWV
iOlM80bD8AGczsngRKBxj7I8+4BH715H1xviykb7kDIUCPWYyoSCGk5boJKyxADMR6WJCSS3xmB2
mu4ByYOnvHu1zN2r7CA5v/dxvVq1TeT9YPXCbbzJP7fV7037k3Si4kmxvlIpzJtRb/ub+iY/OWQ7
VboJ/cxQHgoyXYwRzPrqRyrARiHBnnkdhRHlSQf6Hpa61/uFfTUxNTg4WxSUwVHBH0y9SbhiKO6F
16btwhvamSaxf10toxVElh5mJlaoEYwqCMjmSMIGnY0V8tMw0UeVM4LkScL6kPx1/oBZhCOJ9sIK
YjAmI4NBMidgWzeK9y9kiu0YbPvmKcf+/1S0nrHl95VeQpT6Fs1hONa07eqLYWGOPWZTDykor7ZA
xCXIMa/qUdP4c2yellXkVjKEOHUBLaGJnt81sPMh+0A5OFgeLSHy4y9zgTTHgxepJL1jaARW3kGb
U1eoVj0lGbG7vz9MjjbVLnC+YvWzeTHGB7vpyf5OqdaGv5K3aPZtXbsSAhNVInH1HbxWupORdBAN
3oradK5t4/4qguWm5/kkQTWGBZ14sy21ofyhVDQjpchV+KXhiSUL9h0uMPLkQ8829GayLSdx0LXk
LiH1ldR/3FHLGuNtk0OQWmMC1ZcCdH4B0m1rZsH+JmB3IS2+/AsABEMmtYf4YD8rTMSwNqVt7Rif
kGor5C10yeCeHHBlo2CcA4XPacqEcigzNds5obK+BP0SjRvIniImdOqdh7eZkl7KcEgwRT2WvM38
2z2bU+gdpfdNgMwmJp/qVF/V88vjXwYVQx8w1w6ZCivNkMmtt3+gLF0Rq9Nxv40rdxIXEjUAkhIE
xmfeHA2/nXPCN6I70/W+p2qzGe00W3L1cxK7c5Mv1LBAeudl52UPQMAn9nRV8HQZXBCe9qI0Jqn9
FTABHOZ/iN6vJhaIPQdc7GJLkSz0kmi4GhcRgvRqOkADtPsKO15dKR7nmYjYOVGrXfikx70GYaMY
ZVqwRkmsMNh+xKd+by38FdssFsVnaSSdp6XkO5phMD3WBMpQqm1pBH5m6BCjJjaAza0vkNZBUsr5
4qUE9jB0Hg/z6v/yqBYkRvFBz2xsbEy6PMDFSfe6vu5iVVEbOZKQTG7mJ0PyuRizIrNRwBstjf/K
MCxAmexM4GLavLd34EJAzOjTLAk4dLJTDYI/VWBxCcdDMFC9E53+5VB62i546FZtF8qAq01NXW6e
tUV6yZ/e/rQ9u28GNGKkgSMhXQ9g0yxVB0oRvLcaoMCLrLotn+HdS64kAHuaW1inrpmGq1dZScS5
wIL/HWffTSWnPwNVL1aS+LndvuMX8XNf+QPhMwtOlYQJjEayC1wUhSO/gLdtZdSxCRDX3Fk0ho+n
iOSVf9u87l/4UZ+m+daud+26MgmcX+udXTVxcdrwIEPCER1ZZYiLs3wjs0YrpbnuO1BuxcCtaPLu
1fZSz6kCMMjOBQcSR4NFYE2BSHWiOG1torzIL+TztT5YnSvW9HHMj3Jj1H/7zH0zaawSgS7aMjxO
gbc74aoWwAFllC4eIA6kwZ9i7XGDKNKRn5FOVIW5+ElwVLy+oDDiRQ0W+FlckUJCAAhrMvYKzWOW
ta8kl2p+OTNCJUASp0ZGgMcHtoUVmzPkHAKe+NcJPL/aTbKru+tHcKzNzkeWdXzO6It0VIk4AFzL
8VjEe1nU24jJHUEXj9CgbiKNWPDwNsz+Vp1P/PW/oAaacjgPYvPsYDPg30Q2zHjBq8Mw6htWh9BY
/PmI5rvhMe9WzndKogsEVXp/hx+y9L+MBqGDBJ9fKkK3LEiK3vG/0wrzQd3T9Z6wkNm8Y24oayn7
qNZ9PzzpwjP2s4N6nL9OYIDl7TwEwwkspIt2sSTo1GUAiNvtq96l+G3YL4SzxopGjUCNXxSn5/Nl
ml9lKAg0Ls3EpPtKIC8Nim9rEPYYRhcmj7ZqXqAq9ORnqTFglyPdtdqLjcbE/MfAtaGs9Zc/4CQA
P3waHTGZs23+euML0OSrW8lhz5DAwE9/3IGYs/Jo0NSGeQoqPL8RN8nf0pshO206QpupBA6Bejae
zI2xGzLGkGtkLDo7A8FPtJ7IEh1vzjlur0vJRrp8AdFBeFsOwQPAlr2JQrkG3iSn1HBMoCn5bAba
EFSVM+TVXMd/OyTlZ7rxRFigCqDiHvJPr4Ti3ka9p08qWcLd7GKoR6ObdZ3XpwsD5iD0iLzh+M7+
Dyec6FTLnMMDRPSCI69DkZsjF33vchh/f2AEefLDPoRvhGH+xDhx6KXhjzTfLce9m8FaH9SEw6WD
TnBM4V35GfMhcamig+Dh3VCMlshiVhEC9NAO/2e9UlnDI4VyXQ4DMm+jwNRq+kC+5hIhf9PDiEPy
986RinTMTRB0lFZW3W4w6A1JlK/fy2MMkK+hoLKUCvQjjn/lxyDNZj00VH143ZFAIZOS4JR4T2Ml
JsN1/vfoSzt2W+0Rh9L0WslF5Xs7yyix4PZ26hgrEG1MJH4Ctz05J6jONHLB0bSaCfAqMv0/f/m8
GyVJGClNjG7UhwaKwuG6WstBdv+YVm6b/9gqbmNMbm/nkzg9Bh+tJe4CGzigfa0RAvuvnr6VVCvM
SMNYdAejy9q6my79zPNLbs+HsoGPBzC0CQf4My9YppG4rmaAjyeKKxL2XiJqGduxAscrCP4omlwo
bKlNR3iml7hSnqMQ8tI66kDSXd0nr+DC2Lllmn0bJRAleLmRUI74MSBom1oyezu0ohpnMUsKWeoJ
rkqaVTTGxRMFQw7F8nT5hlTfviO5ruqR0K952d27yDncBIonf2qKInxkOKEp9Ln4wswljzGLcsmK
ZbGVs99wIobwAW30H7mFGR2u/eyU+mBIW4Za7KocJeD4hdid7T3YrngvdqFAj7SSYL/QE3hUGkPB
75h8aiafnVQgYYTQCCzbXjZNZsikn/7ikNiYFO0DGd+D+99Gm8iqDu0HgNEvf60jYi5F4BpGRmk+
WG6ll2HZYyKgWtkreVls6/IbNMRCTvFGqaXIvQs4AR7TgbH8NY1pGLwhDFs/Yv6Uk6s9FVhLMzlb
AjmrXnRnJgNH4PfeCPZ+PqFpSoenoNuWbh7WQYRihu7Aj7dO5p6b6QOrwnW41E3xB/hRnut1yun4
pgecT04ipHNRE/T7ZG7bOUdJ+KtH8hXIC7mte9cik+pxH4ee8KelQ0ZLqXAPkuVP3vzJgJw+9m5C
XtEtMbJ9+ZPsJsV9nNucOK9OiwdRTUh+ALGen4Rlspd6znIMxZYeaV5Nnt0UF1WTN7HGeE0iknvY
UAikJ5GlgnFekQj4u/c3nAa60xBzwFAHyA1HnZuuypvMI/qBqp3Us6VjheZMHPUX5AhwU5qY5jwb
/K+20Aggtgfhytj6dba/Qp52z/fISIfAzsTkzhsVy9n/SabKDTyR5z0dFG8OOp2D8fdaie2gqHBl
9clL6fDt9JGKFSyzf+4/UJJ6zLulGQsw6999I5xj9/ypqYCUdQgywMX7RTTgOf7Gn1PB6S8Ivn3m
ckyEtjM17m7Zmea2UVMTJai0Yqu9aO6sWcFAOXz3ab00CKOEB92oYuc7J+I6y3L9+r2AU4XAStqm
zqO4lMZFlNNu2Wfon7SgMAaGM14YflAHuHvhs1R7VVYZ7fx497eEml1iEr3mqh/orw9aqJMWCWR0
PSrkB7uzY52a0DVzcCmfYJ3ZWUJKgj5l+zhB9flEd6rRCsnN9BWrhuuXCTiVwVHI2CjBJRIEdOXl
5464HxZnYAFAJak2T1geeuzNsKN8FZnZhVYa4IL9hakBtSeDi/jN1e5wiB9zSpOEnQZQo5JPv59p
HXhAGEBo/+xb9Xm/EZl351B2WZW6aZKR/qQSArcUA6jMmhN4BWYqCUcgHoBu9Ga61QECOTqs8S9B
mg1OR0XMS8pNp0xN5AkgPyIxHewZSF1WcUhXbbATobodAvoSHJdum7UD9tGyMpbUIIYtqn1iqfC+
quXdfe+JBwSy1NZ/Zbm9aBbNbdcG4f4gjc5rwu6qhkd17Sa9R+w5ASxLrym50nXf5Y/fRtyN3GAG
5vMmaiate6sv3fCKp2J4oCy0PtkqbMAXdLZVIXE0MZQTEa7EIRnysv8zxBG7oQ0tiTxazeMI+Avk
3k81aB2dJITPTla/PaUVuhBaKCzWCloxxJriP7+LQL4hYrYDhCRNtmgOslymrdHD5wSD60TJAEV4
pmDj5jL6KV5wR6rLUH4OdgnGy8+jfzrlLuayZLTGcuZDjhPazhFj3CWAs05WlRbG61v0jiaAFvbm
OJm8dlych5pCsxiQl+BYTmBibfGNohh2gbpYAcbxHWTL6J+IBhY0jTcScFTwWR3Y0ED2pj4/5DFv
p3K6wssWiK0t1Iw8SYwcqj4/DUQ6gIVHWJPGG9z1hiHr+amOWNE9II4gskBHTeCwI/dV7OpMXKWL
6x80zS6vtDiE1O7+j/IT9ooUoprZEpBVE42QOeOOAFgmxzhFjvQ0+CLHUuppUzeDO6TTk64rgRCG
Ny+G4g4DHtPjjYEWV/Og39mUrULPV9jZkRSKcBLAc+FhcKaxpV23MFeoYq0Y9Gbjs4TSnqr7IeIh
A5LYNFqlqcgjVxR34wCLfWl9OWWpv/Z8Q3mfRrkhtQUtxx+hJvHxi4zzOIGCme199oYsy8JF9WFk
vkoaiMI/B4swSC/ZXGOe1SmA0z1cTX3fKPGAxyybAq4GuykeZpX4hA9K+Vsxnwz4C+LbtpU2VnHo
7+JmaGKWsWlGj0J2wbnh74Fa4fW1nlADG88jk+ZIEaDAIfXY6IJOgGPhrDwhxJh0Ku4z5EtAMpAM
zLvZ0IN33WxdKw+kAdPuOPkpDV2sMDLETOLBYECdKByzQECvGRcrHiPR+gE8AUQPE3lN30MfuQWB
QBTaG9LMpaAPjmmgVxYTvI0BKmdh7IrjsT9NI0AVZyYDkEj31jOIhc+36lseQmXC3CYp5G6IEnVE
o1/ksmJ/BZFKNG2u2p0wZGzg3/Eq1XxXxzjEXO3wm1N+XxFLq25Yy7uKnnUxokTMUmA06KvLuEdl
9MVz7VK8awwrNw8iwe3IlmA4kHP49dZw2Bl4rNs44RlfmoBiDVSvAtHTg0Z3wxX3aXtO8kf0oDbr
SVIJz9VmBR//OXydbbvSLjximVHJSNfW2BfIN/MzRtWFJVuXOW9CiBWuI1zokassVB8i08Sbfw2K
mbCXWfpL/S/2phhpSr7whSCMaX02AwU4H/9RwOvgWkMbM7uMfV4b6GxJoAIZWTtpARomcBEPlhh9
sM1BMUt3V9dZ3QB0u2XRLKBtOCq5GeJXuX0kwMPNNl8m5qgKH5CDbJk4HqJermzTGT3rODbixSgx
/wwkTutZ1KPU8z5l49PL2mohzJ5R41jzsXNmQQQBR+sKdLp7FZAdBMw+mvXNaCtTv3C5wAsckFp1
Bc1neF+Riwn9h1aTdgIUsZukOJt711hz24/oLvvnMYEfSeDbEwdKrxxbpHmn7L5L2WFWNgwEIO0E
7C4uam8ZC+fdu6n2J4Hj3sNqKmoGgxlfsXK/j8wNZG+WP661x7JKHnNYwYpllPf7+rDp1RqXaqQv
0ztXMNC4gebJU9IRwSISfn40fhj5DTaCV55wwYlprNMAEuBdEDhTVnTMwuh9xOXcENUm2ofrfXYa
YnnhR0fwCbfpZJQp6fiwLD/ow+f4fYatd4kTSf0iwev96H5nATqeKxclJH3lLQq0QTLRMAbeDDaL
t+rrPSdKmX1gicE2yDU9DenDjdZdxXGWKEKRdGmEYC64aKy7lPjydyCErXZxlLqROpgEObqEOZv2
CPaN8tgd7SuiQzQ9868ve/oa+fIfT9hkBll2lB+Gmtpap8Ad6J3xHwlDyXUR7Ha9GUC7VGqpBzMs
0MRIwroWMuokAINJ7dqyz6WKimILUuHKi88L2p4RrAA6YhGQPlYfeNXB/M38tvXEpoHzE7yglaYN
TqSQBI27KcdIMdvCCOmbz0VnJq+8+Uh6UMqKNNjI++MJxlN6aufNvDYDACIrSI6euicSAUNdwNox
U9WeXMfObOK5NYAz3zZdwbDcmjOwkzzuLaLEEl6DXVgr/e8KJgiAORTFN7vKrakGzC+ABt4kV+kS
3NcxkCnJneXJkQRgmCfTps35QgrpqZTpYKICkcYRf7OsJol5VpyvVlAIG16/9M3UU6y7+yiq5M4M
dBhOm9/ihN6tPYKwmV69QthQDvGJGDuIeUNd0IYnUk3asrvpjvarngzHcItC0JJ5cyvnZNUgw/g3
Ir1wi0lPXDUEg4C4jCU1v9J33RM4BzJ1zz+8Re47Hg2AD1gfq6OnDKlVSkVizjfJ+7iXtijmvd8g
H/0Z7fELta7WfVfyC7rwxnIlZmQf//pLgjmHuXa8i31eJTj9mMso5rbjIYJIDQCOmX7BWSaQAi+J
6yOTe+Y9rlBciUzLAE5H0P9OLk9TMTgNUef6aIzyLuBZuQ0CYjEUDpYalzaMgFLZeIhrlG+rGwCp
rYdAyktSC+P4RVJWwnF4Wn2nnfXW1lJpYOXoF7RLiN5WAc9jeSud7PfX6ewfK5rONuT0A0AHwOBY
fplwKzMvtk/28ZGM3vXCnMEGILLpJtZeAq0hds4V2HoOQcJTTXViGLGg6ykcO+sG2MrveXwfgdVG
OCeFO+Y3yl1Qk02AH71w1RR1tHKQJWoSjOCI4GEEjV4LMGAg8ewdwKNVYp6ZO1QG2sYkWP7iQbAF
VTeV5eOpwWKUsa/MwM91IhPlyEygnJPXS3STYZMfzZIWWXs7iBmXrPrck5gEiVYXhyJM1nqluDY3
3L0vURUfdBnQh2RyyCRTGDp3BIAzJaeVPH4EyLow1nWMVJd1z0kQUXRJw66tZB5SCiGsvlPhmDd+
xy20tF51NQLuOYWr93KKIfZimBAajaV8i81s46+4biNTOBxlNMVXzVTsClDVbTASBfgRsHe1pNL4
20nuqNTvilX4paQmki8MSzlF7zlQvY3GtL3cp7pyx7DsFpeL5nT0yokX5RsRbm4N3zIRTQRByUhR
e5BW8H/WoCfC3SOTmuiYmTsqJygQHXChlPM8EBLPetspiUb/nVGPyaOeUUfWe/YWodVIspR4Zufw
VR6Uy8AaRcZvitRI/Ztu/xoeJqj1rh/iIle26mkLg4Us6dE1MGUQ6GCVJwcC991tletfgW0ZAKH8
56G5mb6SOmAhQFuU6btQ6+2U5bIfBIkR1cl+DMddsh+mFUiQBz+geeZm5awbJFxfpwXWbtnvOGN/
2ao7Yq8BrvrnG/Mb7tiCAwZB8psuwKhH/nfZBpkwPdkE7phHXoTNruXbWrtr+1ggx0Kuea7AASWk
4nrukBUzPmC6KGUwzsSOzVIx6/3/o/brWv9uDPewJTvv+GVgbBI8SqVldaSJVo8D+BMcmOtP88Vh
3nGMpWGDzpo78pbMZfm1HgbEjMJAcMFWA9G2KpT5ApPe7orECtR4PqZrwX+T+oTJ+7iRQG9aiMcn
Ud5M3CpHHv9/UiToPJx/yXdVKjvbY4zbQPFH+BRb57aeJ9PSG+2NYFfYF3mEPuLXqHsa1mIKEuxM
mSv17hwZDEjHoHHmibLN7QZYqYTAuGzCkhh/EWBdEa8M2K/dpbCNmVuCjtqgI7lugs0Lm89+coot
o17ZSVr9jOv9brLoNyODS7qdUdq/wzZOBDHFfSAvS3CG1+SpXnPHm0d4AVO9TOEmMaU31ZZJgPud
YQih758viml/b+bCEuwHhKYYTtHeeULzJ8madwwpI8hbevBs5RZCJ2vNYjTa6/YV1q4MYjxMwHnG
WIJ0p4IF6f7KSr0mJC6/SSPcYL5CpagYy9qSTHwmpj2rwf7t/Y7BYgU6pWpHIKoMeIA92VtA8OAf
RSDQ3TqsTIdv7OUxuual5yCx/AamzDBbGz19m2A3LPR3bQtrByYG3n0M16pwEPXhTF8CnOZxxpkZ
41C9tRA0onPATNdGGTV0qvacPBs0k2/3k/rb6HMXEcLve9rwK8ab5nU6wmL6SlKZJpYKDelmxgDY
Kor3QGqRnOP4jNL4sE+pPHjhFHFRqnn6I0U8OQvBuSB201auKN3lbhElkRtOb6qX6FdJx10bH8Y9
sYBJrKccJOJvtQohGuzWIp2drk06il3E00aMcBemtQnaemYtjOAra0nGIqb22SMRZ622PT83l0Qa
29euIXQLOZJiAt7A8duiHEaUEsGmgtBatV8n0H9i0T5Jby1NXDIQHsjhweB/bgYj0V+m1LBK1Eyy
1lFyukOr/kLz5ArAHMwYt9fF8WCxjxBRUvpWfA5q/1XUSbEDiOhbdOTWQ2drktx27bcb+ezfVZXs
AQWd6LfmFM3+H48j3KoBnwOAiNyGosVJHhewBr9a0NeB/yyrWQrhk04nbXtbnSbFwLqrzB8dY0KP
c1pGkifcJOCHMWrEFTRvUZn2sjIOTkvMFJ582zpXQbbAmwbrQgWvRDaRuFtnLRTNKE4iPbVz2BaC
0Tmz0HW40zUvLNO54ZgXD8XekhDsEFpMjS3UOPxaFARefnzYQ8Y5Fhe8UVF4TYu+nvPlmuMKVq/F
kuBgbV1xmlh0Ws00F2WjH6kln6Z6vdQ6uSQb1xodMnc9vyYqODwQMJlOMZxGDvMU0NJVfbLY/Ty4
iv1I97i87yp+y3rF/c3fTyK5cCsSsk4aHOVzGLUubatLPj+9vqlBrdtgNpMWUN5erLkH++ytKyxD
lmC1Yshw1MW78EedrfZDtesT4mwolJMayx6sg2Ord4o2HTnTdHawuLdtSEBW3Mfiwgqg7NmjvGno
gl0Z/PDCe2lcNispwstfkL5ZnVrVgCXMTL7jwibBQwlifYHA4uOOW3v91x3XdkVHS6Nag2PyuQJS
QcPdese9yXqpUc2lF4X4J2kSJu4Ad4b4gUxZRA2uaZeLwYSsX9WxoOaO4XXrmU1DggAfFgsOAWPx
XdwObLg3qDUwF9023ItRBRqyUAW+ElKSqcdfx2Rkc4Zp6YQIidHOc7utGjwQHgadyOKU6NeVZsp7
4P+VWlxRx6z11Rgg++gf187Nl1o0igmN5/5XYkaOdTET3rxGE2zLLwMzJI/vmh1GARH66i6E4jq9
mm+DWhZiOBQmAusn6AVGfvg8Hah9D55Au/nf+/TDPllqeqal/PdjgM+5stRIizmYeB1GCgaz+hzW
MpsoAm3jTc1lGAnJXoxfCT7kZPrXRMdW9nuvy4WC8DZpOe4xhWAjosjVhpL06qBEq/o6laed8N4x
IAqctFLXW0LG5ivmcYIoN/JTW6W/gSx1SHiyjyCh8WnCU05EpdYobijFhGQgmUq1naqrSmgQClLQ
IwZP6fDRkXBy1B8Lb4pCmrQwnTaRW36jGjMfUs/IQvmd1hU8pnFUitw945e5J1Rd6pxFqM/v73+N
yZvWo3zbHTFg0szwSsy14+rn36hQHBa136lwlQfvCMS41PD/mWViQcCtl/QxiN4L7Z9pbzEkx1fl
8kYAmF8G2rdqe86LwmWXDzf6oVQfLO8+AcDcAnOtSg7JNYFk9asqJimA84IS1akucovAN8I5iGlE
TruWmJ9mxpGsBSAJTbtFhPj/Ob+5eK2wOWCVRa/5tHSKOtKj9c9gZtpB+2K6V/TnASfm5MPt6j/8
HZ5c0Lm2Bo9hnLWWMdOYW46Gc8fmPF+y/8mvW3stBM8M0T0q/UlCBzh2IHoFwYNA8PQSYIRO3yiP
Zoc7TBNFRI6qUFwEdnLEH+UoXn7SytTpR3PbCGVbzoXEtuTHbezaVERMWl7rMtVH5ENmKfftbeF+
5vnDPYRPK6owo2xlNak3IvE4lmdmOe2P1FFKttf/GnACQ/d4rcy+Yv8KvHcKxwtMERzuk3B1kdkn
3/4D69FntLCwVnGkB+r8Fd73v8Gny8dOWxgAzEr8n1h8xF08PF/gPA1Df6pBlBTiZtItqesm5YqP
VQ7R2oDnC4G8wipGLKBydFlNSv/mVuOcHABv5V9i4txM2+udUeIwI+QgMUGInvshP+RIzu1xndjq
emqLoGXK67quqMiWrxrGLrTv48ewgORRO2sgWZkOvqYHOYAxsLzzh66jczncdqdMC3WDr6ZmnYN2
NpsoLMiqIqrEz0HMy+RLKFWyXdr0qUoKynTEZueAIz3zMKykf/nfyWHyNUyZos7XPxgDaTtHBRym
+zHgDOkcHq5ofMxy0zPZidnrwBj42YQhlgTkOoTRi2Idzf/BBoDoTD7OEyS/XuvuYUiKaGhUfCj8
SySffhqskLCKEGjBaHkbbXfO2w0QeTFIEOooHV4zFWDvaMNQpz4jL6v90Bbd0oDSWHbrpsY9gj5p
2GVjujVzrKfFFq3ZgJcF86eVeP/0lpdOqvPEiGMA7xw9WF/3yA2s2iPToswxnvS6eOuaMfsYNSsg
tfZDeETC2zOilfFYMupmiX7jsDzWf/ZtDKU1I7xzMCh1A4V0ivHLrozcagjB+KWsaonckQwQ1/QT
Rp29TLOQ8aaxUvdR/wj5EMj8L/cog0bK9d9hCBJfF7TUg6JQf+J602d+oXkbvdyXKtXXVYUgr1wW
pSQWr1JA0pBocvET1ivzU5F/mXfrNEJI0BmBFz57KwPgVA/uSgyFlK15rZBp/AmQnTaH2SXt95zk
dYjcIFpF4fJF+ONJi6IkMavJ28X30w7Ibx9up4MWTQGcNcMuPPgMURla7Z5oCcKZ7QQzIGnIAIy7
y9b7AAQDevyrBn3tgnRaXbdCfitVmPpRhx9PkIeRNBJdTng+RSIuI/OXiNn1Ez94EJzggICTHjA4
YMmGF7TyKs730Q/eZARJ6pzAR+VvPlFETOscrStBFrZ/30sS9N2JY+mVwGfZeoleKe3g3z+j+cRT
HReg5GJ3nRo1u6f81NmjqK8Z8s3gc2V2sZtKz3DlaHGnAlMvzyYAI21+ejKqvL7Jf6SMcz+mJXWY
nPQEsWLj8naHU72YC1WgjZW0QPAUWeu//0vGBl0E+pjO+HiShGsmQjzy0+CqIh2RBoqmzzvAmcsm
Uc0AOFto+sidXc8O2Ow+8Y0N3Jh7fljZDPhuYbve5aGbgmhHuEPvcmtU5Va5pPy/weBxwsK4bFKU
1yRzGZhTNtVY4UVRLL8AAr4WHycnBjGdDpESCgZwoxxsMJiaEUFdl39d19KqKo7QXENrbhZZW2bW
kEpzgV+LXpVdYGObHnOzxCs7cs1cY3cwWOMRw6HAelItRABlL3wgizPBkz7JxAel3NQhKR3YPmOs
rEGTKECR5JCvZXiQyD8Xrss2IIoy2kfguWJwRJhhuQQrlCT3prMbJzFbJmR02OVdRjv0WlaS4K+l
DmYfz3zurZoQ1dpnFocQuYP2EB7SZ7u11eBYdZ8T1ubBjXlF+CQjqvel9RP56yXuTa9KNITNYW0D
X8L1i/fAoFb/+gxeEuDW+tW5ZduksTWb0KgTGZF9Y/WKNTD3wuNMnulwCWDLbOaWsSdNvL3B+tAc
+mEjSxs+6v0ER88NEgQTZrM5f/e1f2/iuhCfswPx0AfRuP7plaoEDtVut6zmRl6fI/wD0fIq38nB
E0KD9GKJWeGQePfvWmAjjoeTDRX0UGVVojBkrR2tte7gpeiQMUX7GSJLZqen+KzaubayHxjHlqUP
54moHtUWnff+ttQ/tMDW+CfcsS/O5P8jDrXeBdcwsHw6FO3N6NSnFmFNMe5m0iHjERs8oV7MJLHs
7thA/h9giUqNWxR3vTHIfDCetg5ar6vQDvHIs2WbZ2pBtEcIOzPnbjywtlvSqdGjE9S8oNaO5nEi
svDpMQCNkgGYPa3kWH6Rn7w8d293L5+G2QQ1qB4YMjN+g76uEJedZf2149IFjtuP2awBl1hHmAfW
+OcCbSS5g00141a5TGMqLLMZTFPiU1BD+xcxK/SX0xBtyZM1MPzjNuBFUYs+WREMqoF2Cfu2u/41
CLctRkP2fA+BFunt1+YSNzb4xJmFr7kHvBBvUFrEQ53eCHbUHRsl5hX6u/nKgN5HS5s9vfviixTe
pB+cxGVi2us04h76IOhmcXVQlvA50aREEsRnelFsPKld2t7bT5bDGYQLKcYTrxICBnAAvTi6yS0E
t5GTsGvGIFHZcko8Rq/FjgcyHwDHFEYixGs4oYYcgORdQ418NbGy/O5stRw9mfaE9O9QfUzZtDsB
oF5fEdv+BBLqIYgkXG8aiipQK7G+pwTxejj1rMmSIArA1xfjb6TfBVdE+b2HbZa/e1cdpu9vS6Q5
Bp6hloyD1wfFS7m2HQvR8reRHNhOg63Vpn43A3chsgSL+lXR3y7cyFqN7is1r4/PGU0q4QnDcQtM
219QDx6mTCMsAiFo8GBWc52QLJvCa5mb6yKi41XoPrjLvZ+CaH3BYOaZFIYXr720FXgg3kVcxk28
TFaRVZVw0yBKz9VJt1ZHZbOXpoDKbiSuQWTZou8deZF8P1a2LUaoeNW9DvA9PRAI1KigL2tZUcgW
hT2ZYxhTs5tIcxYFPDg4ppJ2dTs+8IsDWOe7LNbGXf4Sbve/HUPOx1Ju+xO8M1eIDPcscBGRlRxb
KpFy6GsadSPCi4/tEfLMPWFXmWl2IfBGGAQu8H6nJTmlpbdqD2pF2bbS0iIS54mQb58OYmwqyCAw
S9mIkT2CiFQgcLE5Hi2keM4EKmBwkveDeRYt3ECUk/ARUFyW8Mep7cW8QY3WO9K2eJdeosaPNF4R
JtUZfI5iFweidG9AHQCCi6yhsyX6RwXROg24C8LKLiYedds4Z7wabPp5sZDvk9MZUr8RPnAaXopS
R1oA3xYgWgYj2tKoShvT1JPaMYaFFaUFI/g7cod2Z+mKk740dTCF0X1DzCS6mKctHKar6yFssunS
7XciH+0xNerzQq2BwD+J1GKnvDN+wZWXVrFr8k8vQ/6vgR6oUHR48x8mkUbI56psGPNbrNTC9TAj
XkKwZmUuJPvllOmrv5UgJF35olxuel10qqrjEXmJZRXr3aMZe5YIVQEEG/vOjCV1c3vx6xAn5Bhl
oaDL4KY8ERqzSE08Q+K6w1reLJY0uhEutM84XryqpVPr6hqyzgEqBVr13HT4ckmoW8Ayc1pX2DYy
8dCOZfMF8JFqLTDM0/1Zf18CF3xXRnZ+uwG4eRehBRouXKQkkUEJgKYL/2DZckFR+P+tNtFl1QMZ
DIH6agDgaHXD6onQ0ImI5tomtueisdKcuoSSOL+iVHXLQbHT48bO7bortDPUUsN9vU8s6iCJz1+t
N1EFvae5+GwtqFaAXxnA9AD2YCi0pYntxPCN8kiuo0lnIngzlBb+OwaIQYToVIWWKGOZh10LII2U
xlQgwaL0kcFOBJ56zz5XiSu6TiFyif9VGPKXwb2xNifwVrXLaBKQ9nWpNB78YDFSfYtZOoc3w9V7
auB8yl4yAgYr1WWHZJfic9F2OUQeZ7pB8pJ8RJ+sl4THaL63SKBDASiQSyiAuOHB32K0p6moS6xt
wU5qJgYfq8wcyEZdXYRw0dsz7X5Sn/PW/maDSuJL/xwSSUvRpEkcqJtWWn8qZQFBNU8h51c57huA
3U6O59rzBk6z9YGQsL7J7INbe3KEgoOTStEhHIBZA0vIjl/C0BVqPJtK6XtFwIbieysaa6Rr6Ter
eXmr2Fm0pH520M5Z3/UiLaQj3+keDLK650NSxeGP6dAa+3sMZWgFg21323/QFK+G4xrZrrkXCUpK
LDDd/uyDXJuGdCFQv4c+DtPFQ1zAIqFXBG/IqminmvwH3XL7xHqVllcOkNxcX1JDhIdeIdCwapTz
J5bZ/tSOB5SLuzshH71XOdlwZxmS0rgVBzzFMWT86Oe5HCdD096qC2ki8Pcue59ZQPdnchHZKK50
QXqRFgbjAy+DUeqWVDDrM88+fTbwUpNWhc19EQIv1W2QSdAC34X4wWhDhJEws2wUP/qKagScllFM
X6/+6dsHIS4f3df3ar16pfPDzTW8MZsNjH7aMw5/eDVZTu3YcPg9tXwybL3h/7kyITcXLrt+Z1dx
jJZU/48hToJctEgjW8gd/o4CFxcj8rt8mzD94KNbZVKmWBcOzVUjyVBPX/1ELfTYRELpDwxFG9z7
wzVA9Z2ZzGJopmM5SrOudbXFmt5GGXJuFfAYGmU9hOqn4WkdmdFWNQbvZ0SiK7IC2It5SBR+gYns
Z5O8BULPAag6Yehaflj2qdr89EWZZ89yeZnlWRIQGspmbvPDCpDj7DR66j83m91Jb2Tk2ZplyOKi
FtykXD06z85iRO3VD+KTsRA/BBtiSCte8P38mb5v4rwNgMGfA/B5z+/sCL/mHK3Q3gXcaFZdtmQ/
DxVwk4ASIg82VAEDbOj5P356eUy8Nme6gpF0pG/XrhEX6NSWuMw6OYZDAHvzaZxYiITIjdBQFx1B
Acf1ll0XzlZaF8UOVp5kLARYCcthMYby1CdlKYciAMeGmzHkW0CjZ3CveaBVy1xhzcbVMJWDb7WJ
SqrnXFVNtRM6FWP+e9QfxBA3S1lL25slnfj/tJkUz24f6g+AYpQFV6j5lJGxYti1pG+CbUd45mLW
1i6gdXTHXT+otP8AsYvcSHqYwVsFK/Dpf8mtvFzdf5Ty1WbQekpwmxeLwbEDMp0Yxhc/+ZnPBASr
XjRTpL263sNX78axNQxUtwKtAaRd80hla1MqEyNYEvbmgOWZk4tf1PpVrh4JpGZF4pwRf+H1mF8w
t6im0A0CXeCI035NkKOaIyI9Ztn+9a9GGhbdisfswLpdswwyliXtwS0YeL4xeGW9AYLS1v1LmaKn
V5nYn+Rs1JSJPJy/3F29r2pf6HTgdHPghhfyEKl2bxSa17Rq9Ud++U1ATI760wzRC0/DOPcegFr4
iT3My7EqKwXYY3lyXaFUfXu2ojNLg1TLxVArbYRVs06nWLXr7apDTz0IzxMdnIOtJHDyL8XdSie9
dJHoisfw/grbf9664j+uqeEGEYiY3AHBO0W8dDaVCPVW92xQc8ItlE0aWMaAT1jZBEMWrCKJ/cF0
VZ52yPpKDbcXhPrAZtV/VuvTHwjZC769aA4phytdLhQfe9U+vmv4QqDgZynIE+EOf6cUw35NCkAP
YTYE2J2zzomuR/HDJ4xvjBtJ+E7gyspLnJNepNYwIql5YwUF1Jb8FcrYAW9RI7BAfx6cbd0Qngk6
MmIGjEULDbzWebEhgvBZ4JehAitHyM7sY6N+mIf4lwipYVtMpyprn/35jhN+J04EBgzKHII1KI4G
QRCCWPLqvHYBn71SOnqYvk7EFCBaDG3/xecjMpgQCQhUpayxs3gnNupooAi+NfJIxePTAxNECiqa
+XWUmk7jYHTSWEMxXEm4DYJ2KbRNBUm4+tVgo1CmAlUFZmEdo3Vy0zUJ7j3UQDXbglNTYlSXfHNk
mXdhi20ydGAC18x2FOT60C/h31hYdp+mWZU/MvO3GNLYL3+Bc9wCrVsHBSgmINxsBdk4RBZBWK0s
ZDfNpbn40jpYybmQKWXvxZrtdoM6oliddVVWno+yxx+5wdfTUyCRR+yPBmH4d3PqfYyAnwvmbBld
MVkNZwLOn20VLfTUy+vU85h0ZV8ge5O4YnOGArgDE+7o0FZMbxqVemBTzHTmF7/Xd/508avITrvO
6yxB2OpP+HA2Y+IiocOeE/pZDR78NzRtSYjyFwuqQggzRpu0SLOd8saqyGQhkqMYjke4NWa20NXY
ubj5bGVt83PmKmOCTZmCXOwZILBenUP/XwFIiuOSXVgLjQK5nzCQYh4FJnNyXOvFbZAdZq1TzAXk
83X5arjYIU/0yDvXyPrKE2Xz8cCh/76e5XHEQt1CVlEdJwgHWMOI1ewj2FwQRGWnm54MyTf26O/5
XwFLag81uYb4k6aA2mG2h6AUZstxZbK6P+HhVMhydFkYrrQ2EFQ1iPJa6d5/qV3YAygJd5m1O6YA
9XcasRqgeAZzc+4by1ZpGbsB6byhKrcdwLhusb/hLYDWLgxqvVikwD1mmVZxuxIhydx9dIigdiSn
9DI0I3BtRGzD2bpAtsoxG/HdAbfeu4rf1QwzR0y6W/GK/C2AOtAD3SEzwUL7PZMHfj3M6JC3+EnH
BiI3MLBgV3kiusvu7ED7dsuYAEdPMYR1o/5O9A4eym/9SmgWmRXzx2vQsHYOn7uiGJUQD+dK5pLQ
U7TdzKQfNkrBBguqPbOMggntwP2UpReSDjGsB4vBD6lKhRR5Alf2ukeaGyaWhkrG6EYHmTGL3b5I
Rxvr45njO4N6/0GUichAfHExBrZQ+GtJ76DyrrUYRfIrK5PcZiUeVwMomRRYQBmHGQDsJHm5aTG4
51mpA/lYZkTWZSC1N3WhWFWG5aRNGzx1sfEu2tSp6zWLLwAWJiCulnWxyM5mG4NVZPYPtKHuqwCk
ryYLlG/66NV3BCGsRufS/dQEhcLZW6BGSNz+U9Y6DeKzXISHRb4lkdjl1yar0InYCp3zKM8ROEME
cA7AyBhHmxQysEAqRmyMJxhdfzc0zXGTdcVN/96Qv/4jRb0FkF8NmC9X5Myxipe8VcY03XUgiVl9
v3jgamgL/iuyG5qQ+ITz4Iw5cv5KvjjimcoxvVTNO2BdH/EgakdgiWFo+bNCz3Haxq+DKBq5yCEJ
w9t0fhFgOTPiiy0q/TIOMXkB+XsmCyqLS4ZMhnHLrqLpq2DNm0aAH4zIfyRdu/7xpxdL4WR8sT+T
R0mopxKeVEaYzOIfbiZl5S9x1FjCTS6eQixWML6I3Aw6Mr57Oue8hzQsoBZsL4pnojXI2ykGhMdL
DQxgZZ+7snwNazX0TCTi4ssTJ/4cxEiOLed3evhCMYmKeQCOYDs2xmWRuqR91lxVYZbQxN3tQbqT
FSsLTCpWE3XoTWzTd3seWfRA/9Xl9ho4lOlRmFFpoM1B/vgTVPmxBhqpYMcH1y3hWMIIWHmKyprg
/zOhD0hqJNaarrdZ3eu1ylzm1YQMyCQ0NoT9B3MIvKLgnkCUrAEpxMtBZ2lCWmg8xeapeTdR0L4H
k0MMDH05wdo2/L8MK7HEDEdmZuPmLbf5U4FN9nS6PxiwyXKSQeY2qbZn9ikdXb7vsyTYiJXu+0yU
kMGW2EK+7xlZNLAH9kq0HXCbVjAzxXjjEcp1PoM4T200krLax9PqXncK+3+eXcngOuHzjRwUDOus
HEtl/COcFVhVX2Fem1CNfOOGwPo546IDLbe9gOyx6GFHuKh41g3klwZm7f21DwJ8chrXl360Xi3R
WrZ9bIRcZ9JOJjS4GMPRD7NKSzVYNrMtz23LdHhVyMxmh3CTRcr5qVMCaxZpfZuAur7OCAhM2LYP
SEcdQlsWfd+GgsyEkBTQExlRqvIiQij7aB9PZL/13J0i33q+krN9HyLC1wKXUwSmAbyglBKGXX2h
cmGAfaVgqfh9rU92VqLK82W/UEcrSCE+LTaIV0Sq1EntiNK7isW5Tphl6rFZXsHstFn/FZLP77U5
mXFth/IanVLXvGpB6aM/JrA+wfCvPDKcGFFmOPmuKFHcnfTQZehOTII71tCXc6Oh7YL6IiBXN/UL
GVXsDDc7XnnTd4ivBRjnZeLJdH3pnOCxZMhGee+hGEVmJ41U5ghlrEK7YP13DfVOz8DDvKh74tj/
y7w43uvWGuvePhCweoYi6slevvSHRWwM/9oJ9qWJyj5swE5/sZOkWhH3vorOJ/pJKUsYg7CKtUsi
jMuTcSXKL3kzCxEUfiWZ8H9pQT7wxODjRupfxUswLPJZZ0RJA0T94PFVw0mlLuYK80OVkH/OOoC5
KNcaU0YR6Ru/DkawBP3cBCfhAmALQ7a7jl40f1IUcqbYWmj97cP5oPuISTfyYvMG0PHWMPY6JUGc
Al3rXVQMJjcBPGz3alC/oY82jiPLkVqdF+kiyeNUb6aQha8lOu0sHkm3bHo9hGRYEXzTTLuMLyR4
po6xKDKuYU3U+jZ348fi9vMf8M/A2HfZuxpMN5yeHg7krbrxCGSlYAnnVQCOXQf29hXaiYZXvrmB
+d+d8rX0iPtgGKSMWz7FseWrsVY1qrJ3BxgYF8Je9mXSC/6WU1ZrA5nayBeAXCJi4vDF0CPdDR47
d5KYjSqhaWPTB6NKhKrZ2fsLbhhkw49gLHzlR1FWQP3mleQyMiCa94wjwBiqSCNXFLOE5FBs07tr
aTayP1oVPo3rhZeaIZsQx4m7n0wVCo/LRh4jiLTXqsSYIE4vKUoIU5iuvzmiq2lUVUiE/AhQA5Rt
nuqOnCKN7Tz7aF98qOIvyOuPq3Lg7uN1yCDcerV94hmfvxz+33JmoabxaYnGvOnkKIk3GivGx3dG
TW/efS39rTbTNCztr2h7K9bqNwfdeN52KgiU1KyUMJoWk470s/645d2A6XHnF55DAFdeFfXRNN2G
O+wiIJ8jszlb6LzvXtBct/5+ptrQM8aWE/q1YsEx0T8rG1iO4VNW7n3iZhO63LTKzgrjxgY5uOwF
TUQWcAPZ0dm8SDlM8pJxVLBDZTxFGWiM1d0mKaLLeicGzwAsGZDe/F+nu7lpY/Hbl5jGIPObbDyX
KrhQEz+oK8xVV3dSaprpM0iA6xc81XdNDC9KmAPrzYqpjn7sBFRA7E8lhywNsHUc0UxI6hkOEdM+
K19BsoE7xLDPNO5iey6GppVJy8YqZSEJ8/VJLC4coQ3BjN+6DRyWBiGGOB383dC74DX3sRmqudf1
/Vi1yFjndfnU5wI1Zt/AXykRbzsHSLqzEAds89KBdva8q/9Rmql2FAI9pXqhaqKRaGH6KxLW20Ij
vbB5pKLlYABmL8qWpxRrgcIWz6MVbJm3HeYi+x/U87l9oRh5lQe6UxGGcveM29gEg7cl0udsiZNr
5jVSR0hXQEXB1sv1nXJvnhJw2SEhh1fVEowDCCbq4K8qYsCBCz4j+hYr5ZcT190Gv4qygK9n4Qmm
xklXzPdv+T4WxhgcCiZCGFcPIgvQf7iYMHp7H4mmZTSBehaGWdROHBDk/TC+xL6vbxEYFLP1kyJX
jUeYYuzEeTVhEQzliT0xxD6E96HrHrScBDZ7xoidI4YIfI8YCzT7T41HvpqhkHSo97wIyEUlvcps
+hqY7s21p56W4ZtD7iuDY0bvC7Cnh5dlQc25Qjd4maGyB62q7iWiz7qyxjYvKVjWzXxgvxEwC6mC
x8kT2Cz4vRJYfnFJlfrKB9rAAzaBtrvzXlAV50GfxLy1ON/Yd62fD6lnulMGfx3oP10N27D+MBGa
AzYX2FiqDa8p2SiLeCQDf95WNhagG4mZZyT5Zptzv6dsdVYtxmM2AR36BMcjyjpOhBPESllTsNBB
D6PXDxsgCjKJA9PWrYc3V0JzlkKsqZy/k/liGMCyzh5BA3+zNlBKA0/ajBVCFCSj9ufbU7nCkJz/
VL/nQ4H0ykDWY5LQ1WrKR8nS1rrG/JUA6xt4QG79I01T9GgMrrQa5S+1IFk1+yeZ8SOD8fDbuqBq
OR8blRObsVQ1673Prv8CW5L/IP9lHTSEuxzm9V5tQr69Z6kh1mgEfe5OASjOcDW23aH3MmgAiVRA
itjq7J0fcYUGr2Fl324n3oyTT/0rbIVO27EmOFvGTTA29QVyVEeRVB3M+ZOEdy7zxcipvWwOqjZp
Ddd4PwCEMqxgoLjp6qJhyXG+ZlYzY9CSkcIO+9KgJmRarNvwVa8AdImiyXlbaiUWwN5RdlwCzbmn
ppW5kijr4hUOFgeY1/9ZxVTd4IJCfvfTe11J5kFIsGyMwum12KPhUBP54aau3Dj4cf8CpASa1PlS
2RAwrWUxIDocGOtpYFOU8CWGo2Ugc2RhCaMUz2Utk6OiOqJirOf7ZDl405llil1gsGmOscBGhXyq
E3iLZexEEpa6hjCdj1E05h3E+Ewf2qjyDLBFL2NL6xtb0YUfbhuGmDuNxZBevokLearND/E4VCfI
EOueG6eHupRb6F0rAFfOhBNx19Abi9T33ovu3nm12CyLKLjmS3TK3BZTyzff/ulTeMS+abUhnSPi
4/cjobmOm3O9Rp9U0gEONwaB1TcMweTynwjkYn6XJngBI34UVRugumn+SpYgj55v/mWu1LyKJqHL
UFhTHzcylhrny1Cu7vkP2zIGcPstPoLeP37ohFS87yCt+TFn2xX73JR2DnbVX4UUmALCBbeespto
fAtxqc/wh8CnaTjFm3/X1rtjNC4flnV9UIamvwFAOki+i45syXVxlpGooc4yBhfoMC+CBL95zUj+
H8G3cOQBNlck4b/zc5XWZIlmKZuh34sVV11AuZOHg+iPKVkdUFN1LQqR8jA/8K/1KZX1kZRjcdDM
fcJZdyEL8fdsSFGaPMqwNVXoBEJmPdOEKmx5IwX9KlCPg5MWaVbigdecMgylt+GLEg3lzjxRAAiY
ZI/Z+/wZArJWlyDudx1KChGAtDFkZCpXYgIF9dVXNThgFu9Ur4inVDJT4S8no8oxgNru8gUzft+5
0GeW0wQ/THCbV8ZKPBWBMA1kSMqegwN6VmreN0HhactAdg/qrjMJEiWpTinTg4zK54DRRaqKrV+T
qcPL3at5zkpEAxodmowIleunEw5WaOd+EEXLPRpm7WNiRlWPsmFZIZa5cP11MOTbVXiXaRNEsBSx
UupZ3wz4uuZo4hfabuU2UcvIv5sHm4vbWyNSe9m8NFMPu1/dLvTRXbKoe0pOIyICfhg4VH2mILfX
0mn+63FX8lx6q6wTMv4uttk0IqPzZcztU2lqQ7UyGB6BNlsZ0VUtj62Pv72ggfCxCxmjF0MvP43l
MeZ+jtL1yqeRTAyK4+w8XYt/EOaZ+A6D4ZF0RUB8ANcCzGhfZZRrzkHRhwvylJGxpr8IUehEU9l8
qUshSj1x8arVQIwd+YKrs4PbFf+N0fegKmwCoHBI1g9hrFo6wGj292jFAtsBw7VU8Ah/pdUyAqZ8
fTl22jhLd+VYxACQEsn/9X1WKEflUDstSJmr7rzl0bwjqpPpHgnlaO9B70YYGunmb3EZxkcEYyEQ
6rMfuTMJ4SGgvSRYa9WZXC5/FTac/fX60DN7XWSziTzUuZtvYYWK0qcY+B7elvbL0nsu09KYhjJy
lHrazBHBJ7IB8/NVfiFklccAaTPIP5A/Sm0krncWNjGfLbVlsDSc3Uk7vf3SppfMBv9kISd+ejRT
Sl+TP9OZ9g4hDbasA7Y2peiQIUwfeZf/iaSHGTnRlnc9r+egIQGsdGr/M90rPzLOEfxk7lcux9Rf
JR3X4Jw55YsTcBKC8nU8DB1inQauFmLbTDsCsNwVmiqJfppvu/5ZDpttF8Cr7sdV9gqfmECYLr2i
M10hOxAXXyOWZ4yIzjnJv8zuaZbtCclEOEUZ5Sn35ooIdGTFXd+Fo1mD1zq438ygyfk5f9nrirwm
3e3zg9raH0RU02cD89sPk3246ysY/5ACKajNcADGRwVae+6wiXOdqwusQ0gbxXBWYLSwFoDrwpk7
1faLWcdN53QSQckB9OdX4H8tiRZAOZZvXyZjH1fVE6SLVjTsTWhJyQiKb5d7Ne9ffdQR2lt+LeOA
aQVkhumfNi7MSIYrjnqrdc1gZtZXo6T0uycUx7aYWECNfw0TVYCtCDH7XX9EnoWpd+QoatV2hmYJ
bm7HNNoZz9iKYbbb1oLUm/BoOzCriSw3ZZsG4fHsoK5Lqkt+zJ9vnn0fLqq5Yfg40zBPfARywrw+
bqxSngNfux5ZjRbU674VEVftSQX9azsQxfEEEh9YLldzraom4kY4eWRSqDEssCZ9q62ITjM3ohuR
AOj70mbVeV6lYRR4WzKi9BuY3C2KANlpoqtdJ6n5iq9Lg/RZBVdVawOeB7ZG1KZmbVn56z11FuOy
oR9M+ZnmO7FUH+/t1QTQjYiDrOL1Fbpq5d9o+0CcZP2aLd4vMRor5hmrfJEnm60esSCfyVyJiJEf
FdMNvlWsv0I5mbJcYinCXUU/T9p5dB/9JJi7YhkqM5OZqo+1NoIkIKQ7s5IB6NOXen4EL+Qj/0Tt
+AaGZUIHFtRcCmIleRDyEmHnafkkEj7QmJUz//2bhtY8gYdArmu5G8vTuIb1DQGKOpOnIsU3UTK0
OJKEbNlErEySuJLcH7pYLGMS2U8VD75MtTaGjeqOnju9dUJO1WgndqwtQ8/9CRjNwCTm/yAfZwNo
l5+1AUq9cbFIuPceqddf8w4It0fqZ2rGR1g4VJ6iSHPpgCvqlnxA7Ee6sSyK7u3dktOCR8w2LP6/
W0c4uGvQLWiuw5VxoF+B4ukwQUm0urON5QmZtCHJAAcUj0+5AGKwJlzlPjog2Z83+Lsi7ksyKxnj
ke8Qdo/LVzVKE/ZHZ2BuMrObs0KMsvh42JIum3r3rTWgHkSTqez6WtaOwr/fKxXjfMCLzhwJ23oy
7ujLjoc7gmCjTGH9a9E6GkoOWeRoVWxrYoAuOhWRhnDh/XrKqc/94lVtYMyOuhSieoxO4RYYdNx5
3++7LcwcHFf5DzX279hlpBBnrZDBmv52oHaNaROeO91F9PlMlXWejfsL3KcVP9GEYVdgwkM8elnv
w5Rg2Tlb7/Mtahy3GM/sC+3EWl4P7TN+uJMoIhkVwBGVxxK9d3v5uhfBmbudZG/fjpj+trTKGqSw
RRE0MZ1a4R4bPoBDYXSXrZlNmPZZQZDGayIBJT/t42Jcq4GYk2extlEcvG2XdEvgY4cAdkkAk+vh
JUa66TyI5kM6iGMWsNYJvMXzObJ1/US7dnnAItlRyb6+vDDFLl01BjBq9n5kZkfBS8GEPw0nmXBm
oU0MKpSMH/wmALV8l/KJt23y/ey/M7S3CDUHr1dH3e/w72WE6r7vosSr53oBAsA/ovcZgStq6i0P
VFuQzx0YUoA7jNIWA1icwEaAWuNZGgraTATpsFL5OOlVtN1goGXGdHNeqX2pP+W/kWwBxDX9PCXe
G08hyLF7rnnyXARfyX7/F0IhkegIswX69quSw2qdl+I1QGwpLj1eExf2gS/ygGkrTzTVGil/kp3H
rFsdFsRQ8wBt6OIznyOyfQx0B1Ah5fWEhNIyJ0Eak9++P++d7LnpLFr0zxWK4/Zk2pr3WCw6pyWO
YjEINviviSZWbjoolMcK9GAn4V8m4v6iiXCPd9+LrLNE1AAFVNEImoMRjczGG71qOykRLKCkmpt9
3HsFTsnDUL3c7FbHc9A0xHIm0YtbIb2eo8MdTExvxdNd2j5dssK19tn5QH/8WeDJO86qpFjiFQiP
LghjBFr5XJTBW+5wFMkbDEjdhlgv8eJLpOBN4Oz+9qTLxINu3sBrL+bxPl0QrtiCzrDXujp6iSjP
Vq+2XzbWbwMDRsFv3v9pYNBcGiE828fTyxa86KL1zeiRRF9s4TELsZH/SBLMGCFdwUOtAvvsSabZ
YFb7FFSTVvahC57awPYF56GBSJjS6P/qLg756fCNtCoxwP9PbL/LD+HUEVBnLgdVDqWhEXlM1yc+
rlfUWK6cbtdhlpw4TSljA33Am9vSzoS3lgg4bJZMLbZfuhnZRFu36iHE5azA08H/W9wEf335BQOJ
Ia+RLSfno6tW3mANy2VUfFr9jgHI5cBTRqsyrBXxTXLbuXihb8LAx3KQrrXYfsr2hPfr89AvfrZj
47iOs0TZ7hyaifq5bR3oY60+WHe0AT0UNFfKudhW2Ql0ggwILB10HFt7iqj4X//ZWRNPGDaIaFgz
S/z5+bGGVbTRI8zwcZfw8o7pD5JWBn/2T7NwcWIAP27sBRxRPwhq493McJBF/ytnJCzur19Wl6a+
XVJV+54MtruGJIuAlALVnlKeEl0RSkEwveO6M6XuBs3Y2WtWJMtiyw8pyxsJafxOoTRQ7x/eDlX9
hpGf/wKnwwmqFUHx6ghh/ucxCYMy1yQnyj3eFemtGGU7bUJXtQere1AQtajBb6IgZQmusMMIr2hY
pOrAfHVo4mUO3Jh7ZbKV2zY3uJVnugUb2m5Be/0M5KMuYCZIyu1ozOz3CvXeIu91pYF9HdvJigYK
rz7ijN+FVro03jIlU2ItkP/kGz78G5pglbaKDoJZDNXPwj4Qe2Licfy8p8MZ48ga5AZ3UqsElkTz
Sng+o9bZ3+OizLjeF8JtEgrcqGKw7wJvTtNhhTSR0ktEyVll/Q/aXHuvQJWQccLlUccJXfNsnGbc
i71RBITfwmDmWZXxAFntaGyJc6vyOWrHQUWKinaldlxaG460iJJOnB1P71djZcrc/ZTeiZUrotLW
hMXBuGUYDP6c2GaaDn9TiqVXQHvmXYo0eGZ5Gfb0WxYhsbc/F5MgNKScLvbeZlQ0PRlbBU2xFKbB
uuCEKs4X1/MQUyJ0AAKA8Expsz3o/0yBuKEokOuVHpqKf3KFZR0rRPQbfMjy9gOajJCO4DxeoOmc
0JLZmDVy04A1caZ5sWCNHdC29XsMAwiijwQ5ZucYc379+z7Skn2yzbi4VShOa4RiCzgl42frjRd8
jLUrMagoeINoO/A9IfhKEKXvwGa1DOxl3Xo+dQkavNKiFMrplg+nxfASNlbTNbmVe8mzRjG3MyF4
Qm+hPoSPOn9Xh7ZoSc9vx1Y8pZbHxgewQF6sBbfrcVj8rbcLP+pccN1mM67FasXsdazRzutZlCu2
mYjNl4sukpxUrQN+QzyNfRpibfxNI9LOgGd61G+2tTKBDcoX3dRi5VHTGPojXH1E9fHAgtRtmDNy
g8TmlBSy8zb3zQmMTHg634T+9b1wcK8HZ07LJN4DGH3YwiloXWVMhxzFDSptf4j26Fl9Fk4MePJs
4bzh6HErH7g93RsAJSMu74y6nv+632Bwcg2R7EMx6maopFQqQW9mAkWl3sDRY4HmIhgqx06om84b
T9i8SljycguFYhe3sZsMefSqk5uiGQbNycXHPdKwvSR6JqMn79OOpHPOGAOhI+7wviRtGsBbZzND
uc52xPkxERbeHP/+2IDrpbriNxjIHUiXYaZ0Q0RmpCfHNZhTfO5Xcjx9EznOE3+nSwzGBpAUZNW4
GQTNBCUoTcMRiZ/iEQLDqES2MdxkqjCzn+1dDi35jhdfNoSoU0wWH9jGzocjajEC/uKn6222QyFF
iToFYEvER2AnjagxcvE3bw39FnzlNZMpoShom07Cr2sKN2rC7u64FNFbBXQvMQlogSxkpYz0dG2U
X7s5piUB+Qv6rBrxyLnG0XBHWHOyc73c0Xad3ON0oP0bFFhkgZdHdwhSbyNYrUGb4Bm3bymzH3y6
zOMiAYkxcQPiyu/yjbKlgawqPixj9HoMG2wSUHkBiLhig4aHeIylL2SWDZPMMVv94FrrU3rNsg+p
fAEsCGlI2QkfF/yQvlkObcWiGj4QGRgBKEppp2IeapZ1Ytcv9a6N/XajDpO1IzU39b6QI71CFw2P
Vy/BkOz7M5rjjRyP0IIuBN0tg59u2R9068eIpR1rDLko/TkzjQ0g0Ler2bEcFT+hgr3555t/aw8f
YMvBewR3L+OjlFp1MeYHZEPoTx3WojvIsownt9Lfe/RPqL7Suuq8BuUVHZ5kGpu0m1KCtP39LGGq
GrBmexZpX0wE2Dnwtr3cQ95VcWsQfKD1uWt22SegvQjxmno9FIs0kOXJ9jp/fr+gc0Zr/m6F4cW4
Dr5HIYOOTqdr1+DDWX2ijHK0E6tE/zJsA6tbX4qmzFtY+RxmOiXtmwVY0A3jrewT8oGHVlh4A6K1
hoChQGsNGAiQO0FMhnXFXyocHoPme3oRm8ylqCAbMCnH9HSSCvfv86e+XOOHgM0z6DDblnIxJ7uN
mVZzwVt6LaYaBM4d25fULFXa49Yoh6XEHbZ4nR2Gmg+uHj0gUqLsllWPekkz0ZFOJZ5QCPf6D3MZ
3EkToEvP3mabU5WckvR66OIpawKDp6VnPDio8nqK6jF8fyeiP2rJ44QnL62RSTMuRmMjgCcvj+Zl
Td73QEh46fCBLtcA1ZEvzF99Jza7hX9yzwP0RuUr6jOMZOFB/dRqkkvT22wDSwPJVt+rQQ8dbEZh
t2TI1ZwSmTQ8r/7fWe9tonL2jBJbUbyH/C09kRvtXMyw5a1WK4386XpySDCXcPMyFhr58uPRwAAp
mdCzHRDnoAY0blZKOFuYQNzWaC5v04rQU0Y/fuYbeDAMfXBQrXdjvjTjYDBovTIFbABwUAyec1Pq
uZzB2Cc3ax623Af5ehSwrmjWnsdI/MNAeIOClP+WXcFdL2JjXOLn4FaqA2TNlyp2eCsX9TEak3b4
hjTl4M2CVl/BpW4z55+9ebv/PIr8rC3LQJKgkRoVKvShGqTxm4fYy0vq1LmU/9RNX3eIlUxRZLnt
aSSy3+vQ284l9yFEXNzpEqu06Lq6soFn1sr6hbFdNYQWW3GBC5UmyF/vqgQiPs6fXIfAdHEd/er2
ijFE3HB3shh0zHvovFLOenRhw3tdTHtzlDn2lh9Yi9kYYq2y5J4p0pp4eX2SKQxhooZ5D+uDOEKn
Gu7eN3/mTiRQr1X9Ah898KjLVh3z1DF98FDSMPfSZsnn23ix86duyVeqCm8ICRIMluGgdH1ccAaI
rRbZfBiFwQl20+abjM9Py1RhaoE5ihi2kHnmTPpS7fGvVcRzD5DYY0UhcmKidqfK70Vilsjr+z7H
ih2Rgv0NFNsaMHx3LOgcSImIO6Z3X6bxGxJJzspcR046mezLtV/IEnA1sho3Su+4lfbAFeNxZn0+
gN5yEp1mqnkEmxvO3JhYUWjTeGF90ZAbloaFb1FHjOYkqZLCg5H4a3H1qyUWRbRXR6XccctmFEh/
2IINNZB973AynuD7G0tr5oVjlqLcJGuGpPqVEE1l8bK+5mAckxCCU/2spvY35p3GGBSWQAdNAUDZ
2nXmnrMq9XpR9x5z6xf+HWxT9HfMxxeWhJvGfO1EoEaW2/mrq55uLt7xfOcu0LurizqjKI0Nx+sR
IulObz/4WNP38oworAdBeLdxFCQD4N917IPV329/+exuy3zEhsfvS97YnSa3/xOb+uBcqvRrc01S
BscTjY4md3k22rl+FzaE5irJzTPnCYy3HkQjuD0ih/qDsZqgWZsEeMe5jppp0ViLy9qalqphUkwF
m5jXTGuY2iQjWfNg+o4bmgeg+Lm++++9Var56zFd5nGIxAyUd+Euj+TL4PdlhRyKQaknfkM087pP
17zMuyeabDb0MqbiXjT5JscGUif4vCu4ElqVwUtHRmRfyNGRemcuB83ji3h8yHYssNwynQNPisSx
oPR45JzySF4oONc/6BJkYRybhcCi08j/qRIqC7w40QpAukn0ZtcesEi4hU1ynoYXUBYrlJHot7EF
2fsaRZDyYAexV42/ikSTAke2BCXrEoAHTb5jZuqVYPZi6sjpIRPqkO2ZLlR7uKNUWpzcPTjOSXJS
jxuPuUa7Fw2rtmQwGztMp0hcn7E2g/1GWZbQn8bNXpTqJyU0u04Ce/qF/oBYQMJ+2ZqEnGmAz2dc
48F3x2e+Zlh1b4E0x+yULEg2lQts2lO/ykLjeJFVIbckZRHn4OZTSc6kLmYT2zmrvBCJJeBWYPiC
VWPNJRGjbQojuox2VswcIm5CO1qJqrrdbnO+pYF7twdfRs6AqeKWTG3dkns2VqxOAA/ROYYmAVOV
SPt0rxxj8azr4NoUp6FKNB4WsFolz5GZ3UVTcLQIskUUqdsOJpecaesxfV6mU1yAHVZE3wWcvt5A
uC6BVYS1sb0O4KXlfQWAAA6PwVDmmnYDdR/EEvJwA1KxFpTREwzhFSPyrrmIH2v5egzfD4bX+Nhx
6NgVzUmbSIuZpoMqMphY3KbZpwOO0UskgtRFjWWXecXKXrZJeh650Mm7iekMYfiRxE9J/Gun8d1X
1hrJy4r1m9KG6ZRE8mdjCvpjA8w7Z8g6qoq3jrYtV6pp9cKCybXgGCI+6+k6SgelMmkeIsE3V7Xi
Y7cGnY6D5lJCtfRpRPBn8kCM5b59dUNJVKZDG2LcY9hQqhy5xUd2lVzsvkQZEjHEx4K0R3UAdLAt
vjWp4SvEB6OAlekmH7DCp6Ds1bDOmqS3MV64HOmlMf6U3AC0TxUqGe8/ZhQ485VnPhrcdGT+EOX6
DmeSRY8es+SCBZJUWDctoe4E1lB0U+exrhsSfHcTIpT8d4K1/Qk0fzSJH6dr5tNCsR8O39nmEJiI
W2zt7lHOQ8yjKxVyYBwQFzqC9SX327zKb2HDGMq3OFC6SNc38l8eiUpMYQt24nEoy0SWRivcJehr
e6gx6madI5rEw/TeAaBZ16G2RZPOcsMiYu7m0ji1ItKWC0SCGsYtGMARtxSvSMhrJ6E+LrOHxqsV
aNHpX811uGEe/mb2s609V9Oh/Uc2drbH5X+TAWFdv/tGQYman+U9/daXzSvZQHWuN3vSitYGW9xZ
kScEkOI7yM0IoR9omhqobEXQif1K9IrdIBLHYCHojQgVnl5tjtVPR9sltcDZTpSkv/4AFKHcvl2w
4ziMhjCpZC9hzDNTYXQocXAVzA3nDhO1RuAO+z/5keCIsGqb8anbnLRS6WYYee5f+gIvYd+DQf35
q+71fZ7UiwAUHoUT8Lp2SCc5Qs0a86D7N7i4ZHlIq0IOxDpSj3OIW/IkqpFWfYh4ZvC0GtDRac+j
YWA/j0fzRNGDmLml4+oCLPDDK4uxKS/HF6kwjU+KeeCNcMUwJNAxeG0Okyld9WcuynSD5n13oI4c
1KAOcskJDqb2K6xlCi9TSCa2QQM8stYrOBzT5jJNgGTFxtOnPRgrunjZU2rtKpcx8OQyR3p2I5Qz
LBIP7hqi7p0QRUdE8dyQsRuWdNqbvsro5g9YUwlrTdyX/ONMc7bitB+YeIj5aSr0nwlITdJYjq7T
/Rrt4QaWo7OgoS3YvZsempfO2nvq1b4vSqmJBbyVVBrMBDwca+/KsNQ7Q+6KTDuv5eQIkdnYnbKQ
HmOuliJJdsVd146PA9v+Ye6glGNzqgr/Xp9FRuPrTP9q1LM8QGAFc3wZ5jsHuYoAqGL6TeS2FW34
VgyyIzM6AFubcj4QQOhhxhvzuNm14CodZ59crmZN1wCSccqpfiwrzHVu/Z3mYCIQx9KljgSnTrAH
hPB9AfGSfVm3LPdhbbjDdgBUCQ4uXrm/l0rdrsim+IZBRpUQOi3zv/lKqeJIYLpGgkth+Xpryj7y
3y54QOHs0oQA2Xu/k1C5+6KNS1IHR/gb5FD+12pM8oXVupVXfVFGkNIozB7zN6LhYqzQfZGeeIIp
9yQSiQUezBzCblLdH+lPmx3muJEkfp0IK73hjf6LJn2PAXC/fxI3p46uSlAVnOV5dt2rG4sNOHJY
kSzND/hHzjkSWBI3ysaBAhXF5ZNOvEHc8ckJXUnqqaOyAuxcQPEHyH7cw7ZDUX6hwSBuqHtK4jMi
I2aylU4LPp7ISUzjDLqzAuy7vOnqauPLcEuYhB5Lt8wgkKAOmRPUew9Gfs1+JPXagoBPQibp0gVj
H6gb5pKwySNIOW2bMlBAVcrt6peKdN1enCA8e9gwmnvvZYJIwq6e1jaNg9aMMTgmawcFZCxL8uum
yNJo3ySIRfmWchT5SKBoFZBiD3wYL3KHsdphOzsArcrtG/EiwrtZVeN7PLbKms5Kbw89xQafOW7f
4KoSgzgkM7aKIp1lCEh3H7M9Uw0rj99uy8TrCxHtfF7rVirCii5uOdYR0SEmqWQEM/kLy5sXIBu0
6sOygK6WtD4qsQT2GsrUHGtY4EDRQ66RRNSm4PRcOAAHdD4/ov6n2xdMKwB5FT4NRSXFnfCGBViJ
+pVG0kJo8RgG6w0Qk7gP+Pj6sXX2ZmzLC+xcFPLsZAVe8DPMOmHkkCS/sdvl09O51/e6gjoYeCKt
n8WuUu7/lImaxodjCzkBU3B/PcDoKGeWRuPII43WPv2y4yimHL2HpUOVpgXT13HAKReTr5p3U/q0
Y/OHsf3AT5ET8uSILIRIT9FeCKR6LQUtepwBbkLxk7jrdeFd5rHQg1RDTKi+RbM0rL0fKcAempng
NiVVlxylKXYWm9c0nVj4eYPVosKbg2O01hbzM5EFNp83Y+UEF/JHdGt8xqFAv3ZgGA08MYVWuTN2
KbH2GDxACdrRJsT65n4XQPbpnkYXyy+2nHXlb5ldYmrqibqpgx37BBeQTTj7yP8wnwQtrwJjv9Gw
I6COG++49d3YL9h1Rp/jEh/iQYv7ZXgKfVbpNwKte3C9H7yLkko9d+tNdB7EVVkFwda3rsKkIfzI
GbZWVG/3EDVqA9SEuZY0IbnOdj13Y42AhfdX4UYi/7NAjQuP8E3htDfaFKQNwJXAWfQagKn2pI0r
sjokGqv7UzC7UEWgyOJM6Bd7OM1I8a9Gc8o+BGgSn1ZqkOXDok8CCQbhe4niIEf75vYiRpY+VWJt
CLn1dZBLPzN3QxNpD1vYAd3glNRGIDDeGgqQ3sLhO/N0FznryIN0Ctl9j7P5riCwwvrgsvHoeP6H
RHAAkaqz33MFzMqO+nFmbCJawDHZh5E1PQQo1h6152pxKhg+5NLc9q8Be6l/2vtQcDXOdHBGMbIB
c2CCLGyimGFWEiYAecnQOCntJLRIHaBtbCvWZ9qjjutAi9hzV9jnKiGOSU7T54xKHExkr2KJ5eyo
Y4R/eiYQYwoyKKZRjwisBAMFeaq+C5X8RBE84s1wZihdPgBOb/NVl6eOJg4ds5YYHMO/CuO+Z1YN
W6PvcOHIUF2NdWmdcB8VmnIbdfG0o+//nCfQnQW+mHBt33fYSfTcuP+QI9AfRBTVyUfl2VXjVp0y
n8RcZdZ+POO3bBGPIBYpcPzFZG8K3yAqWaE6FSwbpcocYRXHYpZD8sopmKRDCfntgEu4lXbk36tB
nY9dShEXswLLADer6GF9TKCJ/J+VAiiJHHvcHL47fidzvwhEkODMYaRpy8TECF2oOSRKo2Ef5zp0
qRwxTbpGEs2VHf0Cr52JzTysHZ34iL2fm7hnq6UeAkq0z2xBKOuboPVOxw9mSvOOmD3dO+jNDGVM
zU6VhMaggraX/MtFZBrJCeKWesjn+90fM8D6m2GNkemGNA4PivrCLkFB2iT+B+4Q5DWwlSifbMGu
9TmdYePRBdFu2rhPNXVK7BuK5Q73Ss9ZCypwyTqsoU7BCp/gdhqO0uCnTnwuY8Q5dTbB3RTn0NVj
aKYN4S1/ov2ueHKhVYU9Oqh81FsJ3e45aPSiBzqkmW4LUOhQuXMFibqptY2zzkyqXKRt/37kqENM
ObdJL+BofEFkHC4bWX6HuLCRMVWfORSgTMyzm2Z8JlwUQjmc/wMoCmYPmgWdcXcN9/GrtfO3Y1f4
wNMyvcLal5euhPO6Lk4R6eg7Kjpnpo4ixF1m3zUaprHCwYV1hvwwBIa9JpGS/FNYhZFjMPtMyND+
z+R1PxOPEfP/GuMlv15v/veg39aZZfrwIRdqWp0kc+kxTjduKB8STtQ47z+31tyvy4O0/jMDfE4g
sB65ow6rzlX1k6BP2ngJdLp35jwnJj4kCtj4hMD4lSRTk8Tn70GL2625Od32PVZkLcd67V/UnQ4r
uGwDG/xEYgbYDX6tgWMEJBctqJ5d2bG0zJ3XlBBpkEOMk2qg/Sx0eJm1lSF31UUTAvFJhNiS+3Iw
EMlsok1o5xjf+3AA+bU4Sv7zuvkxVoyz7FMWTO+FcWWcjZuPpdU6MaKDSy1QbGaXBr9UU4IQ9pmz
5xgvQBmMAyujWvw2r0X4HSgUUfiF9A6/KqTethlayfMLSds1PF0ukFDH3XsmEh3ZMuD7vNJp6Dtf
QmdfoadwvhmDPo+TyBFVe1TXbmR5AUoFqWtsB4OdGrEopLYmUZW1feBlIc3nLz+zW1n2HPBHZYZq
StY/q89XlyhJ4CSMxqTqsE1NjZAB/qweWlEwC50O0G51mCY9CXFchl5AiSbFGHt32NnxpxCABC4B
eKyYyCGnOUISnCyZfqbukKVtcxDEQsl/eeMTZSUCmDkYkNfhKhK0dpj5+/+WCxlDZPbLUuVSlxm/
nFufcz7O1nOLZpGEXEB4Yg2XLRp/0uFJbp+YUwRlx2yvpPBlA0fdbVu2AZY3Ctcy4fujgSvQqBFe
6EEpz3Eu6v0LIcxPB9fFqtu5e88QR4PIwDxA8DokxCXOeeB8bIYAi+ktY1aFh1MNuxZPvz2oMj7Q
FHAK6HtXI59kXnxjH0ndK3HsPGGHgYlH8GL7ldvn4hLSUl5i0z46HKexPi2KeQETKxk2Tp6vbotD
7yp/MQURqUnu/JPcHO2z8ghod7OpgdVkqQo7NEJgtKoCg8LVXqO25V5otvsOZjIHUxMk+oAqukdy
Kzwgn++h9VDYypRbTO2T8hlwaXoxdCOmLINV5AonJkfN9NwRqQUka5DnmnZ8ao/645wqKogy+PV5
a07pwyN0HukkV6zmR0qIdLpmQ3gkhDKDe9U7A5R4F3N6if6XPsoc7Hj0xz9XB+eg0FJVZtcy/bUP
cRg3W1hyLsQOGtPuGzGZh1FmFdXhe0lfhDLvrOGVtfUHhwj54eyVMSgMGDA5qLCyhF9UDoZvYBnd
4CGfj9AZnAR/zAxU2tpXHHmd12XEDhJJwsGLHlAW+PTdTtL7NXZOAvoLcMHlUuUa1UFN7NjolV01
+GK15cSAHt7RTvZpZFiMDHlWOK110YFdEx5VtBWbuPfKt0AS1nKgq5g2vkLc0d7WPewCNOnr4bfF
dIICTRPEXI06nrZOJvCtRNbUHsl3SIYw7CaxZVR6IGlc2sBQs/XpCtKmxiGTAhrYIDsu7wCa98BQ
bmk3GDz3XluAyGwH/khlmmS4hDDPX022bfoYXoiWSt97RuonmX7KOeDw9jRKx9H3234LwuQezp3b
XXYJEyOELnEZKXZkCiwFU7jwzv+J+lDdh3P1iQ/boa8+v+Lbe7054y3GJy57cl+bacHkXvT7oIk7
oF8h9Jlsrgo9itVx2KmhtO3zCkOBG/8rL+5KhOrWrtJhKljGwrUfbLLC7h/q3jxJn1k26RumEHdH
X3k4T8Nvi0JiW8yPlUemG2nTHyWL3Ej+dP/EswCKAcLZYoQTvpCUtpIN6Whu4TEJFZBus+cpkJjv
g11cJE8wrdFkPYiaa0jHcF/I4l0A8OTihs9uQEgGo3sbssPz/msbw2ZxBCyKZgvVtpR8opvIuSvn
+Tx8/d0aOKGYfCu0sG/8g2TS3ADYbSvd9W8/bPwDvW6QdVT8egpcT+mazj0ghG7yI7WxycLfO3nr
8Rv2C8XtE2ivvojbcI/FEXOMYS5h06IX9dz6H/A5bpcdcnf7WpoK5nrfD03z+9WG1OwSXe2T5ZcV
/kkylaJYi09pJQuJ4xA7g9YwiPLMgea8vxnx5E9Aoof5FlfAjqL+MafaGh31DrFn6Nj0+mMn2IhM
1u6uYLPG/NCNUtjbEFi40/ZawThvv+PUdE6vU5Km/l02P5o6n0y9G25uw/AujtqE9q2CI4SUgwA9
vzlejz/gAh45a3yR7i9e9YL7ldkarTa2qfbh6TBkSQzeqCg4+lJZgOhpnBMp/TVeHz9hYc5Ae0aY
D5lsXQFGzlhDhQNJ7zf07b2JOWt7ULO8C3E+Sa4hra/hKyScsvCeYOwcBsRFwu9JlycfNATxmZvu
+pwagxMEQHtJyu2qUV/iLLo4pjVGKA9pmKVDBT4OCIRCrrL+1NKjqjpgEKR1uPTPCl9Nz4UL9UiG
VLpqI0He4YbcF5u0xJV5zYYvMmFGzmkplbUtaTrGGJ18uV3af43i0ptaQeTswiAG0Jj7J65OzH/M
zVWhco8QrnazZfQpbnFGBLxuYx1hgcH7qbIKOkDK0uCsGOeyXUyl3kg4YIGuTcRSte0XuZ/KB+BO
S/nnGNgiHiG0GVZtZDTiUGkp/yalDzoQ9w4yNha25QMUwflSV8UP0KZLxeYPb1rrnLRGVburTgyR
kHd3nlibxnhRp8FzrsVpRhqGIxQp05rZW8zBAm0MJt+YuvAXCAIshmuwClTZgGWSxMmXkSLLJYQQ
GKMWKo22n6+gQq/xUYsFf00nG/JcXi9Bn4IGTmaY6aTtMjAfklEe61o4oiUCFctcVuMCXGTUqUx3
EfA4j/4c2RbI8qiOuLMT6apXMv4/fpDnZ5SRUPgtIeFbdoGCUTfyTVmbr++K3Oc2mNc4U9mYxDYv
7TYh8auWWdFHhmUx+AVwe6q32CTxMGtYrQLkLacc92s40t4r0D8GeNCld41zA0tZlaz3KBTdyRQB
pZUUvIFkuLlytF4j9z37kmRBSOyaUCuuS7IYkhC98oqnym/27usJkH/GalBCwXvQ4kfpx0bogOkz
6hO31fxW9HDIVW4biAuKmoCMYi38KOJFatt/fc/mAFHzK3LmIe1LuI0lNgy2Bl2Cy4MMvV2OwH1d
zs2ZFwhanlykv9lo6+5vPoDmtT/mkQkdvdzeWj88WprPb66StcPR4XwU+FWaHQTCyb8CbGoQZfYN
m7DQAJ9S1tpWWOOr4tRzmGOLSI3hFv7IzpCoFwb8dlVaLbKDiZbGPaC3N7qCNV7FCI2V3o7DDia4
pzz77ofyhXqwcUo5EJoKg1YzNNrQ+dBjZkS/FGV/n9sS+3VaZtgzCNB7B6QXqPN+eLr0Ur2ttwFY
zTHDDaMK65d5lLyy1AL2Y+jx6xxnD+3sY10+OWx8aoxUR2U88tIlB5Zs2BWElvo0PDNHZp5d87KQ
CjTQt/tV5MJqNJOTXOgEuywbW5fNNfb4juE1L5VYTCMqgtf/5fk0ABpp65xYARP37I/pKilNZii9
MhRJihqLB6j243b175Vp+wd3IdjwR51DzQ4tBf54AOIJ9338V0KDfjP81c8U2E0dq0of10LIIjMo
T5cWc5CUwWBQnE69OOAo3sx0O1sQ+6qncM3tzJze5uUJo83FNXjpZwIsdm/BQJ9HqlKdwS1yRoyb
SenPoQpc1hmSodTsgp+q3oiOeIxRn3up1wLGKyaFHW7SZpXmJvAjoMqKRHlAxi0yxB3xUjcbs0Xn
YRq8V430Fa5voFjL9NJ+6ZBkCmH9Oi1GDkHSm9vGC2ESXhilnlY5qSc3sjBsU65f+1Dfmxj6aNSq
GwCMzIeGnmP5Lrc50utGO6as2YA3JHXQmYOTJd6Pz0qwe5Qu2bGVP6I/l/3gGEYuKTo7ItB9ns56
Vkj8m+RY6WhXUrzGUhD75hduMWKQJjVXmteeeXZBRVrYN7Txl/F/UmoAggmfMDSfHdI67fzL2a3r
VoEqeiVi10+Yc/uJXVEg97dkF1ii0fkqB9eco9q5r9BZPaWWK1vkWf+GhrYw2hI69fSqjW3Nltr6
n+UWaym5twK8YZCyM5h/CEK7Dpu1g4xtSMOWpdWDFe3qid5UZyfcOFUGUhWQ9KOFsh/6qVzJ7mIm
NcO2FW8kOxjg4KPC2M3Q4GmK/0sLE53UR3lfJUFIn8h5FG79AWm6Q/BUb+7VFzwX2qnMKJQwWpk0
BMrlP7PEMAq0SDs5IQENzTOMWx/BsGUnFYcogEPH8QovRb5Q0/g8wFNRd+uNr2+Ucb3Wq1NnknhD
OkPyU188to9chEtKZtUXQ3h9bwZS/m7XWk/Cuk6yuWtzUW+Dd+IwBYdggn9K3zNKHYHfb4Sy96Ol
PClx0AVJTYD9G67QqyIyokLtlo05ePSH++KjBEwAG+1ZO313/2V2CYXZCiQUzbElTXHZOAV2HrAM
+q1nqm5XoPSzcsPsjQlVwnkMH7zYwe3w8FJKcfpEHerE4b2d89m9dgf2vd2AhYb++mRbUg+rYNv5
qzShZt9EgI34x7+8dMnv9cjZbNT4L3FHb62/q9kquP0JXmCusABnhWnNC8NyBapqkh5YKt98KePr
m5dJ5Uh/fGNS+2k4WNK9qrn8Q14cdvIpTdQT9MfN1P9EmLsxxPoSWAoz2OHhT2NXWi37DsqVasxx
JQfWMHakj+Q4EB8eSk8kqJcUF4jUa9A1SIE99yxSIJqxKClF/SL8rTiltik0q6se+heOlhnPv6Ha
M0kRpwbqEnC88e5pWWGUk/HXG1OdhO0PgorGo7Fwo2FVQkd8dSRbiylFPM2xRFyd1Z9IvmWzMn0T
0gq5QE/ZGJPR2rRZ8k6VVgwM7WDEaejehgHSuHI0xi7t3ba/9oxWYkd0ugyEdWZtaS1ypTODwTox
iwMftYrJAB8NPjU0F2fiL4zKws6S2WN3WiDRXnd+9S/zVJJlvN+efFLvt2SWLk+pc5Rdb6IcJP6Y
GPmdP9J9etKE5oqrYagG6xWkEJ/hYlTH9qo8/gPHmQnfMiqzSfsrHFernTwzRQwgIcJW6mmNg7Lj
U+gAEJOb06T9AXnj5NcP5RCZjY3cV+oJxWySVkTH/YqPSC4X6EOl8Tj5/fhV2v043JpDiHbJyX5X
WuRJ9Ebj8P6wII3lTSDHr9SjoOH9O0SCNR0HVZPfbjqiPZLE8ndA540q45Dn6oj2x+ynWpZgAmhK
+VcM0pFnOAzadmvf8PxKBqEZv+0Q/Y6HyaC/ZonGByc8LF5ZX/N6ZwUM73/b+MKFKZWFFNdZS/3h
OCOpKZaIPQeXGw7SzRehJEATuewsdZawTKALy/9+rRnmrnLn/X2I3kj4v8MrOIjxNiLSf2UcsNof
YTruAYq1mxhx5pcLnKm+2eKof/cB/rd/lEtRvhHlMBvnvOaIoCf3wlX9rC2cKitfvglVvgNid/SU
xgfG1GmLCFiF1c/ZbP765P2GrUOk6HCwgMc0arOB/YgV7wy440KqC+yXBpoC/E/FNag2JzAInc/C
tNLYwQmYzrMkUwLIJfmgyWod1VrhY/w3NWEFQpZ3v8dxma4nxcvfus3UQZNJQsqYuVW/PN6RumxT
6uCBH6gBZ5i0J0EPgW1vQSub1Sz6HiHqb+s17GmkbqP1DIzZ+AOkUEaCvnxtfoqYo42zEUJwI8gY
LgCNrXa72jNmI1cfkhp4aqAB4YxHYfK3fXLL6CWqDKR+nRvISd2EO4udk/zWAdxHoM81LU8NcGas
ia9iVxfgMt3X32l8pcGh8D/2UBna7AW4jjpBK3sePR6Cb3pVQuqvUGHC4lysZhBz+NMPMeCffz8D
5h99bFdVLy1R4QH7sPbrLAZCFYCaK5To8+Ny+mmu6/nSinus+pnl8qk5MZ8vHFqgmB1aYuH5thDc
psdOrGjJUQJUBY3gyttJI5vw3hLtTFTxjczKe5QUjelfaQGxM+Q/sVmQh2PktMhf/NI6gLP4mC47
NLR0RGbFMEsHafwxX5e1xYNKmFGZ3SL9x+zwZPPpfaQDLuvxs29mlyyiflU34X8kkPv61cLldqsE
h9DvSAwchGXy5QgHTJxkmUTutLreFzMU9h7OlwqMl7/Q8b+A4XfILynQt9y0mfMwVRJEmwgV9t+w
pffB6F3D6ZXAexK2EZbencAsY2UO4fI3deGEdcrId8SCeOrIhNBqTZdQ2Zapaa071CrBUTj3QZ+h
d+CtZi2n5Akf0SiqTND0IJMp/vyik3uir809b5D6ekic+BJqZ3P3JDxQCGk52aCtJjqqfECWBR9z
C+56eAZUrQFtyZ+HPX8rNq/VglbBKOneCLb64H+AVuqnlKrr/734Vlo0vbsDlbyRh/4HGRiVvGMv
4Zjb+8+ssfxjvjs6YzuztmQNo+Y1/vFBrULk+RoY8hjpk6PAGLUClK9a2UI3Tzt2Twx8x3wqcPC6
IAbDy1wPCxHCOOzDpPwaDOYlTqZ1a1oh66oJYz0Zvp22AghNiCK34npgm+W/MxCxaH1OX+KZSxsS
j6RBFbvlJZRlh9237b78g36uyviZRyaDJ25FEYf8jLmQfnqXoSSMFcgFR4Gh3c8kff/k8UE8s4SZ
6Zvwc0bB4FZoAMXQxqMppY4sXNY3Gd66PUYMoVxeg1BYfzVyKLrztxw5dwQRbMmh7UNLkg5QHpFh
s6upExnUIDfzs4yqbDQxOnk6bLIOiMKfUAWt8lE1CthAoHyVAKrJRc96mKcjyMkDe8rXgNzdPngo
LdvZJpvfKZWrCNdFznCBGDiqEW6HouZRS6F0rR60VLzuiZ9W1iuwZvB840ciKaEnK82Rd1rYz8hb
EBJLQi3i0fMEmH7GHJ90FecZVqKASOKsLG/857sLHa780T25L3STCQgTU8qKVaqk1rUdXOz2thVI
YOpQV6D6aurJk+91980XnU077y1+xfOhEbg9Aey1/kSN2zf4IOV9BZlAeP5WTdGQtPdUf/DWxoav
6cHspYSymYaxHR1v9tNsq2feJTHdlE+WFikVZA4a46tyvGlxxN2BvJl8COgZ75sT4wt48cGzf4+z
7146herhhTtSIyURqdi8Myxqztc+/b+Na1EmGpfHQZbX1eVkPytzn3/yd2LcM78957JHZXt6XLkA
RooqJslbaTeOchdN6RRNc00VW3G+RxJt2oXJo41F1YKMV3NQklPHKjgaSzgZQd1Jh8/gmIswIhNu
0pczRZsOv45PhYUUHnSyPapOv+vyzBlcVCoX5nIZ4A5Is8umtb85aLRmM+72sFX8gPqBIiq5tSkM
T23xKwTTggIZgcrGRMm2DUs9GQovXzj4ICT8x8pCA/7rjzRSDwxPQLYT+7tXPsjow0fmtJryq9Zh
XZDbXTdtJHtmr6jt+Jez5rR9lTIK/fPpVoc/UHreVl2RWCSerSDdQqPXFVqDVrr9kGWbJqb2IIsv
/vuWqsar2m1aTpDgzl6n6DzibiM9057UVkJjrvcAgvdJqUGWuTAH90QsKOaA66I+qfyDtDDq45Ij
wy5n+/EyDgfBrs0rkQWQpCm38efqdhBmDcKTWOggckn2oOeAQoc3HYWj99GidTaAi5RJ4SLt93TS
m0D/8AmjAx2w5PXM8DLIrA96pvCscD4VP5/IEgjKcIbJVuSVhp6KdE8eEr/GAxEhHkoVsbQyg+20
+P0v1+8ePEUZ5g6OpGRrNHpJP0Tro8xrvHs+KuBJmGz8bq+WAs9CvU2LCcoWq6qkg0AX+bpsupTy
UXpN4lnJ+rVI5s9Iglys4t9DAQqet2OT9G8QAU6CmuTFn4QygNjyncsp1lyb3Lu2Hfs7J+Q5cVA5
BU6odu0jSaEATcSLxkz/6HbNIzSUX12PT94AGj1djIfqKRoLHxk4VIjI/zvIiy1o0Z7PN3L9CGL4
j/GVu0zm36a2hXweCLE78S/G6F1su2isNIR2ioW65dv/FJOZlv7GwC4E+Z1pTJNaFxInX1Px3b5o
uHVCHFcPMBWHckYAsYWL6I4vb09qqtqzjwpLN54j9PgYY3uWLK7Uyf0wVRLAU//oTv3J/BZ255ug
EzqtG/lQe8J2ERlx8yX2F73xYfHbTy6Vbvk0n3aBosPFn4LZVoxMGvJRt0KLy0SNUdygBKTCAO7w
n9nNvojO76aJfeyABeXMn2HsjzgtExb877nprS7+y5A3tQxKWtmgWG1JG76IzSmC+wPIW9eZx6yf
2cMfzQByLPMeB4Yu9+wFWM+iBQSuW8IrbrpUR8nX1IPimmKUXfp+G5Y+MKBqlDfJqA9JDV1DXO2e
OqnV4yFmDvcG2D1KnkwH8zaGw85LKDVvEdaMP7gG/PaOQqDc+nQ23N5hQJJLGv61G/xuf6e1VUnU
8pJUY+FsXvYWDrm8IXSQWZ6jn10eswtNU4YIaIvssfSeJYACfX6ExobMsTJ7PfxavuCUg62RyhUD
QrER0u80qj3GDaEDHCTM4pUJ2vnkMGYKy61MnL+MiZR/TT4U9NncoZI0QFSVCvFl7sLikaZm81zN
BhkfGulXoBERzoLk4F6wt72Z3N8Xejbr+8tZKBfvaqtkLJCq0ixZru3pqfnPtZmi+Q/M814gnrzu
J7K0bukdBo0vV5Rsvrz0NGnDeqfBj72KJxJCL9ZZXkFm1Bexh0Cb7G+Dl2wEeuVxABSp/MGnt3yN
c4sEql+cNRCoH9ZD6lwDhxiVbT69T8UxhG12/ZHRORvcETQlYU3fXiypdayr19asB+bzTK8+eRbu
lSDQ030+p68ePoWC4vKZ9McCEgOMe0whhm1cD3uYO7iREDZCEKD2D+YgnbSW5Vpb9RKEbrbMrTN2
GDR2Jtppv+R54NxW3wUSX1WEpi04Wgq4gssivxga/fhbY+KI2fFc5dUzh/H71nD6zWl49+MtLqfx
d6FMPe2J4beme/4KdW2SxI4xuwWIaoVnUSK2B1qY7SKFjU53H2HAWMGBvdr4ipWf/DCLRDaSIadc
StWakz6aUtu4d8V3LzQGja7gUEZtsftJ2WhgZsZ31/7RwtK+dzKheFsUyUhDkj4SMhtillNec6TM
Q7YHpe6Ro27jffHXLZm1Fm4detTto+opuHfSwZ86Y4+KpRYqrHAFgW0F+gXOBM8dUm9KpQswLM0I
jge6jX/9EVIH/1TMMYK3ElLYxj/v7DtUKKlW/DUt44aFBHOA4+k2pp6a7X5y7R61ZtiYiRaqz7IV
TAZNAHaLZlhZhu9NtK8TjEHLhaPvvfwlcuJi/kh9729hcEoYETl1argoKbXbMgqMFPngJyslEoeU
Y6UioS81uTV2XzG/KKzSUt4+L1OhRUu4dhtIyOZpv2vY1AIhlIJ3UHOWO29rbgCYZpNNMYcUYJYI
79zCi11ugDGBjtCmxoPC5O4W0glE/EIXO6CrFr+kGJcVHbbPT16uue0C0d0FuNsKFIUl6Qq8Pq2G
F1w4y3AYF1f5ixb4JHe4Z7aM9rwefHnynlmthC3o0pcZDK9nAayHIkroIkwQQBfR4PEmMWurARPD
9evI9/0PsIha6qibvNQ3XBwERVUOdpONnW+s0GLlL1RIJOwmMlVD4AAKtj47RYsd+mTrItz4x8kQ
F8UQFELJ5pPoZ+VsXl1mkKphnpvMLsuTcPpVWP8HKWDlmxPDRhaZ3v/Cn92L+Mr05EO3HwsN+IVf
5LRkUE6jTcUDYbMsN2J1tMXsexI/kwhtp35IRFdwK9tgM1HvSj1WGTemA99RHtiIIBN1zjmhErA/
cLjYObKGBHDYJ2GiwzA9Hb3pwhsEg2CYsiaS65zSu/tkSxRclQoUe9tR45dZEGBKzGCz0htKFaPe
Q1v9vxneuDkProUJzqJrSazjl/Zoe+Ha1CqDaN5WT7RG/bHyRDxdo0TGHawxrUlLdrBYrO92fc26
dEsW8uW31xxg9uLAg4JawO6IMhqpQSXj5OHreAb1ZrjT8Fl8F4ZMG2jxqf3Fjho2KOA3CCdIKR4L
CEGYHV3WkhNphquWACfa8Ka4dDxzil2LzG/AWSQ65KGEVUhf3Q3e6AiRuVkPqtT9myz+vKxtwz+/
s6qFnJFQ36qwLjbIbk9ao6HXNnF4A7XDXsgYCeR+93CXp/82Vpi/Ur+jLSD5iOfT2tYLnhEJ39fk
Pc0kzaSPOvGXiCn/shD4WeWYhgNWgYFnSCEUmYWPREKl7/HwQzFH5z4pamm1perUUYRFtLV2qr1r
2aG0wjXm9g2UtGTb/F6tSvTn4JjzzI8ClSRQYPepKygwzI/Yqb4kY3A8KUATdA0ooEFi2P7Ylda6
sRidJmi/WtyaWTnCe40GHA8W9QAJgRh+8dwLHZqc50xDP9kL3w1IyuvWOPuqQBCSuSMnPYkru8rP
RiNZHl6bcmt/iTCosGqNklaHpweminkDNVZCXeqL6HlABjDrHRvbIl5saURIc6AueHHj1elJl2aY
TY2v0k1vRtcL2HAdA0IA5w+2UU0RhCSKETFmHavxT+eZK4WybxSeqIwUB8TY6SrPrwJuLojA7IpJ
w9ua6G7HjylEVHT2Ykby2p9DkQQF2jH5x9n+5AkotfpUXCb7KLxQMeiuVf2uFM5GxxjRggzHoA03
9lDaCjL0wwGbw7cbBeD1eVeFOxNzGKVuFB0Yr8l1Uf/DUB0lzO5BLIhQIy1+oJxpBhSMGAkiD7N0
qjtc1F6yY8nBgW4pTWGbA079kAawbz/hNuFg5W93MQ28+t6ET62ti9vwftmjDVv5YcXU/ajOJQdM
hivBClWKbW99fG1pX9nqWblRnvuT6uFylNT0yKg1NLZTiy5BqLcSP9BNFOAsq8hsq/iaZ7tGCph0
JxImeD5P+7Yra5mjKD+qvQOivHwSydvEbijQkZLpcHt+z/k+rCBlonAW8VjoUoOAmVqtrY2xOqAI
fZb5N947kEBWfNl6e/a384LToklkiUhY4ya94TBNynxM/AUPc6Pe1xPi9qegb3l/blDKZ98C5cTC
/h3yzQpU7tZz3UNOtzJTabRrXRTVwTM7Q+R98aL9Ak7iTJZMJN7Hx+wZtwMk7+B6HvG6v1onJxVo
w5frf/orp/Y6Jv0eQMYE4xCJVjoq6IoHS/NWOFF0dlwXHJjOtNIsfECbVBqwZBIknyYD/eOAOI1y
wAllKolifUpbIDOzOuEKw7Ra4MpOM+nFxnVax5M49J+WPpp6uWle9PyzUbkjM+IFy3Ekdk2APLbt
u3FQP5hzWoeEzsiydms0+qu1foyW1KFDdwwePxSa+lnZsB6IDfFOh/MTfOEs0EkChrsOsVKBYnYl
t3CxHs/4OdxNxYPp09CZcFMW2dkljyfaDiBe40qlk9/6H2ciJCi8P6EQMHauFhGjSrSzAhPmsu6h
eQdlAFN5tTZYIroXm0eoYYZP4IXimcW97DRLr77tsPcEbhwZIMHZq5ATlQEKFxfJspIdT8DITpL2
9SXtPQ6tBkEBGZADBpPBmz+DASMsZYussxbO1HBnF16b5uZlaj/chcEtp+gOwVF11BGzBZi914L9
rFBuDyUXaevvBiipeKcZ/Pl80dCTZ7R2EjjwQkEDh98CYP2A/mPyrdIFABNRcYRJa/BUnBmN3WI4
LanYYGYf97TqH4rzidtiRvkTqDcSd8ZLS08CFGdhl2FN7ooAHEFCZsDlPdcb7JZcT1oi8BlMo9vo
n1zHe1CDp42u9HHJxw2UH0fqoQgBCFjmoxln5Wmr879j94pt0IdZ+lnfb+aLfms/8LhjrN1+v7Ax
Z9uVwCORDxktwcEKtu85y41+jsWnEjkwCFhQ42bBs8W88Sy16LcVjio2zZxydCDxLYFpoJoNXysc
loj9Dpcj6E9IV8lv/dFNhwr7W1F9vgFUjaO84T6ULhbytsJLxQS695ynbuhjBAG+fkm+AAPVFK54
LDd7rTsHjBlSAUfcsELKpX7goToHGWDP0uSrRHITXKZvjoCIDIhMRHunBLb1U9Amw0Z9hU3a6aX7
1ccsigaF76PJUKNCj+kKzE9Eu/uLmSI3jN4/YhUqjGPhSOw8EIh/JEomy74CvBaAlKo30qQLzro1
8ineakiIebk7p0P8REELea2U0YxmbksMtw10pSSaj8UxDXrBCLoUXB6Zi/p6vf3ND4NvQ7nC03It
1p7UbPZAr6w0eM27B+dBfUHLF3ND7v6sB9Fxmx9AnROLNsCNjLcQh88mBMrnJD6EKOwzuXdSKg/S
HL8+plUheDt/yo6JFEGLGWnZbZI/ItNmzXj81xmaVMe0Cs8NrYHOpJOxMKXZznxOvjpMlb3iURvy
R3EzfSXGANQOayUvUV1n8hrxd9Ugfhq6H4vUwuSvU3XFCSNuXQ+rRYG68ZiwSDZuEnA1gfifNGdP
nj/URv1mQ5Z60pcKCs5dYmihox8LVosnYWPvb1ll5eua747sUXKY8nodJCgciKL/M5Gu4CwDgMMa
QO0uzEMiEc9cqQiGwMZTZappRp9QGashJz/mFqPHHkcfnfkh0PF6u6tA39NT9N0jxTDDo+ULVezq
XVLB1uCLAjPbvjH7mYecMofhLbSLpk1dPq1yOzrojUzQRY52kY9IL09hkJ5VUpFHCIlprJ5wca5f
MA9zg8ioHfVEcrvZOAmNUwoJsM2dM9k7g2w0jPZl6PWP1Aexrbi0GHpdog+rjMfA3DKv2X7yaTe1
Hqap+Xxr1xOek3bt76/06xfCFSU12EW8ZEQ4wtH7QqjSZKpR0zjJf2KRQT92JEiuYqrqWexn9o7m
WGnYr6Si7RO5WtJigZpdKVbwqHRxZj18RJu/shywgQTVPceCnxy9/DKLBVOww4o/BSkgZ68kdnWi
ECXWpkW8mRDT8DUu0+C7JjoISNzo4D/G/i2lPDxWS321Y1sDk03hR7uknDavK7afqVvx3djEwO8q
d2bVSCR/tsdh1VAkpPczM0vAMH/tHR67gZPFD/EOR+7lgZS17ai3FyUFaV4ZrK8e26/T22fDVPnT
pZLZ6gwl5fGMaSlrD0jJnWKPXBkWrl7mxvlEiMF8WxA7hvJRPi0fISfvzQz5KYc63/EjGW78FVQI
uxPpmWpnNuwPk7E8X9qVwnSOSvo1BA9pKJv9kAvYe9fzoNrG/m6Od14Yay+fCKkqxGOGS/EJTjb0
PwZnKiZeU3KKgWVlrspxMgIogR/+OgvikKFWzmQ6AB6/gjfV2EDCQJLPmwMWrlzaXgp42jtxAAc3
6mAy9hmZfXdlfpmEfLsqhN0iBti6/ve4PyNxx7LWOiW/Cvrckdt5ZYxWXa3YuYcRFG3/hW1+G6FL
Pn09bumr2fuh2G3x3XH4xRySkjW2u+uEAYMxR04GCLNCscFc0uSP6iU+klc2x99qJCfaoxrcaZOK
mMEQB9seYSxr/U6KErW6cd1xwy0ARG7mXBwAawh27p0H7rvNTpIKdlAe+GxO70BWWbMiGi7QZBPg
01pdXUyxZK8LSRaTqoQ6BLH4f0JhSfUQJn+8PiVbJ6nNUBsEAPREWTkPrdsMmpewhZVYjWffkjFl
2qFEyrPV0nXeaxeVkY3x474Efvyx7vLd8Snwt9ugq+rKyZ3nFCV06uowxqCoeB2Wxf6YkDvlbSRy
jPlIpRD9Y+5+pFusTRTWcCS+30VvZvYODrdg9gxLKW0deT4fP5o5VWmu7Pw+JR+r+3xukg5TNtSb
ms6BykQzQz2zQT7O/71SJXmsXDXnG7CXBuHifqfme/jjgPgyprGG2wg1ZtBQUdd8Qsvwnmib6Quu
IZ4Y6VfttTZFsekzrZ/oV79B6imFCA9n/mQ6N+wIaD6frwQ6hviTsgvjCXJGq/fxhKSJaXaw5609
kOj116mv7fz7kZ0Vq+qrrD01j7MaW+nmQ6yu4NpOfjHy4I0jxJTQ4VS+Fh+RkIlf0PhcDXWlcEfZ
vciRsC2e/UF7JPyA8DJ4IqRAe6jpf+Pd/HxQPYfNm2uPG0vdAT5J7SpUbhzBHm8au+HfqVocxtwU
uhm7bCrRI2180J2eRnFIonYY7cmI2uQ2Y5re9l56PXVAjMGSGuLzCx5TVYlfY9BUH7Cs+7Z6IA+d
GcyE9ml7I/mjl2irHfb4zO2FdDIrUmKucTuIH8wtFWqPhgjEKq6+uMnQsOApf5dJPYjuKHx0MHhB
Rh0GbUF/+e5PYYLQPGyU/tS/TzGAUbluUDK69J03Km8DT8HLiqV4i7W2YZHojLnNPapLZMtCCWHX
s8TejDckGx7qBrOF06Sn2v0dE8O0D6ysqhTO9nM6yb9Jw1qiEZeKbzCm6qgJlhdqoioI63Z8SEtd
WuTqX85aKa52qyNqUtO6p/coD4uO34k7/dV4l29uLE3/BgBBAM0//ci7K9Kx0lJkN5cThTTAdmfs
Lt8TfK9fZ87jeUI1gTZy1f6Eh6tUhhc5/mSgfmDQp1pzupBWH7uy9iW7bVQv/KAkTeSSXDEHFaKj
K930O8nJzRkpeFdOzoPBgygbNVQbtpBitJ0Vb0nf2+vyVsZmt3EA4AKR1YlmdYAZsb2+kHcCT8nz
O4buTuouTpVtHKIuRiCFbBICm/BMwzrGDORkYhBuxNWh3bxbMKBIhigU7c9DwDKV+KalyZOBkQz9
z6LCfXEHmVRVGfhfm01OdNCXmorwpdsJGdiBwYnwJQkGQusrFXconrR7GBlVBpRYxAMJ1lHtRHzT
jNHC+IMio9Vj+Nub87oGSaErEeHxZBV/s8t2gFv7PtGIPGpznGZJip/gfaxe/tGESfJ0A3L2IuR0
o4WfSC1DHfECyhhLgxIxDNj1CDoV86G7l+j9UeFuj3ddw3ChOdTz4S7x6ye6GCS9jSMeqYjyduOg
/Z+1cYDgm6Ceb5kd3aLAXJJLddS2kWBL37s+r/Gj0+n+xYNMXQIQR8BdbbbFqb/CcLLrxpvwywel
XLM0F/rbb0iAmHSub89kHJw0Uvz/b5MmyQibmfXAS31rxYA+rKTatmMOOavY1ByCMTezdERvclKl
/CNJ0H/thlPQD2gk5vdKMne3Mkc3kU9d5cTL9FW8+0kb4f50UILTBjAh/m0bZbcIGXPOrn7wIxcG
jec6UfZ9ADfxfh9oDD/2Lua3MhB0MCU+bMpIbEkW8JpOiPYVDVXEd4b52HIvG6eP7pmXClK4nFTw
vamA2W49lPuV9KrpSd/5/3+busw1MxLSAtMpRh73YecKA4i8pmyBaRViOpMhLCCyn46g2IT6S2rd
72HC14P8ifIL0zjJU4frqcnhAW6JibVbtZbA7cUkSCoLHYX1dIRwMEoUCwo38sYn396Dpd4p5MXT
R7ljTAxWNscPM9TmekDjdx8joDny25QT7V/n3xnQtu0rL0NRuvv7o+plQwiHj4mKrm51C4K4QQvZ
osX7Nr/Obb81t7UCUyjtP+iJ/2gdbl52PgFe8j19etGyVHnCeLss9y0Dhs8QHWzZeEKninIv7Vkt
JTyIrK+S8rg6JfvhAtQHaQGvf8KE4uQ7crqufG4Pr9wFIiRFvNa0Uk5W0nShKBwBod+Aj9Ns+3XG
6XwYTTx6zYCfMOl90HcuApfqHN1iLiwqmOHzH9Vxd5HKaxz94XznofwiSw5LFh+K8L5cX9Z6e5CY
U/R3W0I5i0/RVoDQjfH9OXE4xFcPInYVq9a2ujmXGkiLxEXq4ggRQ48/yxCqLeN4J5ZfD+mOy0xE
1OpE/EyvWn8KapneB+SkMi5jqqEm/b34yTySR5aZmQCTvuy1H2JBwmdECQnc/gE9Q122COqJVzyL
wrhzakKYx38gtK3Q03uZN/XtAaLOW9SRqGXebuSu+N54YPBCAWP1JSGm8YWujsNZFcsG8lP+Hns/
zpWFlaC/GF+aZTn3GO6T3GUCiZY+o1wHZpYQldK1D8o+IEarQB1DWZoYHCNrrN7az7428gTT+2ga
f58ZhZxSupbD0Xsz8ddSP/al4kpSyTDfNA9AUWTZV19QfDWUuj0bLfsYKQOej/tVEwbvQFds1FYR
Pz9VGFZa9GGDO6UbkduzWjvXVIMCUJb8cq6pQ9O+a1o8Wwh8IeLr37S3HvnIFe14OfuHKxtPS/Om
EP0O0MQsodFDpe4+UDQLLpVpPs1QImz2zVc+JgTHPGpiT4GG3TRAus5VIkH781QjgCwh1uGrYxmx
6w+Jbte5yNtQ8a+Wrt6O8ivokO+rtaSxXtIhh+Wlc8LmLPh8pHWoMy9Kp2HlUgz31yo/u682GvPu
n9CLE3wgSVxq+J8cO/J3CBP0jtkuqWZkjqJyjhtPpnNE5gAiKdOxL5cMejgCFbYjKvJlegCc9m/Y
T2t+QApb0b1DA+s1BOpDYUDN0kzaFMKcFYwGqJ4zzkKGTmRZcW4KDU+IRGXIeT6iUIpoVVkemQr+
X5prL5+QALw3/fxlSLXd9NbeNNleiN3izA5hPb1msQ45bNnAtTTU2vFIF+y1Nfz/iY3VQhiL+OuQ
m+4Yq0Yvkx30C0ieMIsE9vqnBG1swusHixZekwHhupp5aku1V0gO8pHRgxNpt5Ix7DZ65cJeyLYo
HSdVOoeP87xlyRWQUUHhm+TdkwPUUXVJK67t8rctKSwpfF8sgPUn+k75eNwZ0TqS7rYB1CPV4Ec7
0wGr8kbZmzGXUNyH2i7LbRJeSxL4xoRoDBk99MPFieZDTcHTeoHZdgjLsNOCUP8eiEbmL3NpTYJi
0FyM6GFL6k3iqyv84YYG9sr+kMsy8RcRKyBSrtd6Nfqd11TWi0HjGFfOP96y1iJI6GPTFtnnanog
VgQRyisY/0vsTjA2I/Dg9UivIqtOv7l7WKBxzbkMkStrsIjgXwz2INjdp+1t+jGksgBoY4TOsH9C
5PoqrmL0KI3gaDBkCbfAzzI4OBQcWd4elfvBIqrV6O2yis6AccoSROE+0BsJAKmMgGFhreCg4wZ7
SOndllu7IoMk1uIds7s9NCj588q988vk60MlRYjbEkVfX4+jztrPgmsqzVOBi2YwYEvQ2BBGqGIC
8cf503Y2ci/s4Z/GnOk4h9PBji9MT5NYKcwUNoT3P3UpVqUrGBMNQ9Ka4TBkPTxQWPIPtC6MNH+J
tMiPAZY/3BNQ8OQboaxfi3ULMBXS0Tc3puLxjAhZu7bsatqtHMLr+9Z+z/N+WmvTtx76LSVd92DQ
k7jL4OngqrNStDnwFXl0KE55j7t/Prx7kzqeIAzT5ibFxRRU+4+5jLsA2P0w1KfA7+ecRRwz1ntV
JHXPGjHGxCTpek/ML5Gr3fRh5gC2Dx4r4zdMQtCzJUp39awJga8xMRvDkFI+9CU//Kr9huh0oLu2
jrCFugVTFpfmbAOP5BBTREMQDBAy8Cl0FoFI8dICs55F4OcV2ZINr1ZmuhfWGUWf9zwF9iVsUSlb
JrCN/DvZ4A5QfvYrwKOrU9xLyb4zUHKnIDxsHj/98nZXNtBoisFIu4ErvBkfOsCpPKCutz9jIBTx
Z4BBFE9pSRiaylYym9c+gfVjwlLPA7OdQPg7g6VekO16j3CyrBW70GIMKLBdg+iORY8FegfoPzN/
gRBskaDp3T7yJSHiUrOlztMJbElh5tqLVKxEuC0LvmvYKe9UkHzOxJQZ08X5dnfkPg1qy+s2o5KB
A+HhsC5XGNfyN7DHY61onRxYgkIXFNSp6Xk4WSvCsczFZyffWdBQyCQjInvWBGq76ARIaQr8fkbF
J4r2XpAcvIoWkItagXui/vQAfLjg+332LffDtkh05/0R+8CdFKQMe9b8fDXubv0iIKEhG2f8dKSj
xCmXfnKqY2NDbLlT19I71pelyp8D/IpeNX3o1yG9VNQmUXh7wyP5EDyNkrhGldS+dCgG8ZFkwlq8
iguSDGnT/M/1QfRg8Zao9Q6/0v4Udloq/0CU4Xk7Z2X8BQfvyrRKEEHuKwgHfMl3VjiMzUzRUZmz
MmY1scahLOciVnOoZ6kL8rTVlsBrG0Lj8PFde3/C8GSbma/Jp0FkHrnZUldDhYNHaqtzaSnRfjTJ
2trnUbsHd67F5915T+6381ZJwdmfrapnHriOz4YPt/O3JUZPh0yxYBey48s+pPlrfbG+I7abnl4G
09t/MS3vesG0AMHAGRms7kIQq+5S+st8KTZKhsTat71eL7EO/K8J8tbQ0Le+kOZMF3lBBXkBcfTn
IEXrvCs2FS1uRgyM7Jfgam0hT9zAbmxFYqNcyEmy7xHJ5r+rjezh6CLR8HtsW8J2Ty5HVmp6UJBG
yN2t10Z5YFqUoNwvpOqu0zEaJuzbuisaFLRZr+kv0XgKn3v7oLEXNdDscpa0Vy8WZy3iTuCpLEiO
t4ckIB9fcjz4BRRVtyA5h3/Vfhh7gG8H4xCpbCb2xrVZ3pgcCdWKyX/ObW3CHpfmlNjEuaKpwdEq
Wal6sTwK5+xPXLZNo9LXGENz4sSFxhlf08GDUjGtjPDvc8hpidyJpkTrnbgFFUtzVeypIKdZj697
y+RYKb8MSu6xn7+40HTlJEs7gw72jmGpaTHcIBTSLz3cYF4+fP2lq8fe9FJFHmkSRqvwwtM3GfpK
qCxr/YDOQuvRo1KpzKgB33pqalP9uz1mM5MenOI5gmxDRpCLq+gxTnELbKhd460U0Qn4E/AXF+8G
CNqrp7kMEDlzd4M0pLZVfPJqFt5jdh1P2TcKFyZmBi/vgx24braAtRdlUFICTedAnQx7nqzHhtMW
6gCglFYVctZ7a3eyEEN89kBTUfHDHl22gTSiWaRi7XvzjtLf0kT2kDXLrZmQYoLsnDMH9eIhw92d
d5yhrsWca0Iatw8HLVFVwxDjFqZKq8VvvqwcPLNUQ9iQ9K/L3l8Q7KUKUQIYVV7EDceRal1jdJwY
gXhH4jSV86bR7UInQxckAAO++7sSpxaDlTHv+IzjmSbFr1rI84RFFKuoxo5Rw2WEu91BkBbz1Fb0
HBEvUHgw5V6TZ2vGa7sQXuuvkbfxvD4A8COK4JG9PHZdoGyoPg55lBK5l3ABiSlXjRU8M3hfSQ0U
AN7RJcvXhC5LOpkRw/sTYg0ecwE0v0Ii9uKpuAatcJD4ydIk4YKQyBuWlYiyRDMPxTb17qoshUpK
uPtl+S3tuPhMF/K4/wrM4bp3Mct1L/4f4+M92pWoj39H0SnEe/QD2Vfp3kVMbIBQikP0Rsfclrdq
c5rHL1j4Ntya99GgMjgN36Vz0upwFCRKvrcpTZYiO8BGNHZ/zSd+TGkNIGnEDkgPX0N31Fg81Udk
RDfEQxWsCKL/0PmxCgpOfEGVXUVwW1JxbPcWO9cfVB9Ltf0clkfSocUOQBzbgpqlHlZpiEqj3rlR
REXqVYIyrTzj/wSY9gnE9o3CfgdyFT9uUs6/sQ5ObdOTsMy6EK33K4gI8Af8LhHgG4AYCwW3NXuR
7Gr2+5jPgnvwOltW4R3dsanHsrj0EwTed6XpukbS+16XsqCMaknAJaFI7OyUkQDryRypsIhfxNlh
0IUFSx0fiR2bVMXiGNgmG9jkFhhE60khkn8QafJzX7WRzFFVmw4aZO/uISIxohf8yZsxnx/gfjs9
lqmAJSCkHntADalp5sx6+2gVFxzttzpSqiGxPD7N6Bw3siJgr7BVYVP+JqYuaE+2Wh7x4MFmlq1P
P3Oh3HL3GAWvIbSO3HCtkWrJCJaM/wwvPu60BoKoEvdedv1zpyc8G9FfCVSzZRrsOrtOXQzZiv99
X0uu+hPJhNTiJAw6VkF/JVhzRC2B8VZiINIlZF7h5UD60KRhEgfba3hp2T1nntfrHrJ44xqG9LIz
vdEwpN9ZXNScT9sFjBR1phI0K/8xzsuD6rpQ2wCVk9nj2ZafkihMQAJK5x3umWhS58iGxE8CSjoK
bTuthWX/h4t1qtJnEy9P7RCvINTMODOxC3hGf4YshlW0EYbmf7UdmeCXShmC+gZq6TIIP94Aa9PG
Selu88f/C7VUdAyESHaU02LfJPWojf5hg5tXToUVrX2KpG5KrxftoX1/Xa8dBqF11lm0EGed8XCo
QJyW/YGQUI4y8JKBJRqZf1X5lfHzlJgPpUKdA6UWqdlpqPAfmsTB9Mq22RakW+l0FuSjChSfurFz
GoCViHt1bGXUXbommmLJVR6kf9fiTf2ptmQ4YQH3J07BTe7/QQy0UChq8Qq7KETkgBqjn5owKGAL
strMni3CTZSU0LlX9hdZPvh7QTyHNcDE4NYbmvGqUFq7yvfQpRsy9jn+9y9XAUw+OzlOrbVRF/A3
XCqnyk9qsxHv7hCqar4YY8rZrFndpfWf4gZ416AdxuDoKDnbEREPAaELN/5KjkwTxVCMLCPQ00Nc
msRBYpKsrfXowhd1VlazYHWMHGUFK8DpLWcy3l7yXn1X+OwBRtLOeaXlEVsOsd96STf2CJTvD5S0
ziCRN92NsCe1kRX/pKXR95fOFGACousE65kG+3OzLoFgUf8ZZ1oLIDma3DFcicXl95RZnuSiub/R
fvD38J6PG1dUgAN5J1pp9XfKvNexSbSCyBSOFLyXJZx9jjfhu5actJO5wzA6Fs9IuwjYt5vrdPt0
GfyvxNYruI+dqrTcetKAlJ+8u/+1zijEBWyZ86hhDqaabJjs7wGWQDoLTnHyjSO1OKQ+LM0GrXjB
why2jX44g+CTYouZe4RHG+LkS/mWbeELhD1hIC214Z+n0MQKFAdZWBZbyziTZPvbjJP/jaYa9g+k
AOvX4FSl2eGIJWph6LJvCPaGL4hzBvfLjsAAaVOfVVcLbTL6N4harQAJVLghWu1hShrJRHacCLBZ
pd686C3jeHG5OgLqXHTcoc4BgLqwA9ycWzO9m8qrcXzVAN4Djzbv1VXIGeTPJ1D1dPWRxpVvR6hb
naVqpPgnuF7/ZhwRh16n5czjbehSdrEG0/0scPj0P347CTa8nOjQLQvS9YI9nmWFJNQWBotBo0WC
GFgFGr9msmDPtjorYeUAyEV/824INNhe8iyuu85SBSxXYeBqjZZ5KZk5vHaQ/KEa0T7LNjIQirfa
MjxzWotRbF+B8OJTCicszHgpQvWW7OfTlYWyS4+VWCCs/OPuFmJGBEJaGUq+FmtApJzCctW3Lgri
HOA4md5ddVWBY/tpaGLmBuCbEwBgKb7z06kRaXWRVRilWSIPRcpxrSki2DdHzA3dmn8ZJqh+jqrN
r5pDPUE8GOkcxf8yNjxyyNuA8I/tbJNwLagDttkJbZYXmoLDVQVRVQud9OJt0bHSkCIUclGX7ijp
N/IOsoJ5l3xSwUWLCgeCpqt2qh+ALgV2lAadEG4gD+/9S/4nASdTn54MAZpYWNyHOee7gdD/JN+9
bl966yCv3YWkA7E0njZMS59jL1K7XJIj8DB1oVfMEX7FrQDfwvkdfa1u0pNHqxP7sJHoH9f4dbTS
Au37r0iGVb9E9JBjBsDmQCHQmZzJCO7rF9hfx6v+JjCzll6I/Fe86fEJczkSqzi+esaBgvSj27jb
qQ7lMPqGxw0KlUDHlycs2XPtPuPlnc8i4hUkO5NzqM+/3+mVun97r+0DtqWdF33iAQYeotIohj0u
b6D+0idOZec1R++oadMhhtPU1ISIfwsYXhNKeOIHWPLSHowjDpw8AHKyr0XbbnFl/jPLayDfPPdw
ogwgUYfubLsagLlTrmvqZvQoFeAxvv9ete0iPpxOpXUr7wQC/v8MC8J0rOISnUJ42AyZR+GkFzKI
uBfCW8jlkHWpaagK70snMCb4yn1CMq7BzqJAKG1Lj3nDCEm6ESCZg2NolrkuiH849WT9HkKEaTdN
szC3/sf5dvt08lgD2XpDTmKAAZ6Mj7kAQn1/gfvspG4H0lCSN+Gl8fyoQlAuMi1d4aspYshiYeNd
mBoUsMDBrE5Uz7O5zNGVy50UC/YiCwW7v6TI2v1bssKYa7dQ8pxtgJGT2IgGWVDI557xeVkEQNGm
sCTXGynCNsZinlV+qTBmSyziLSEAaAEX5AJmczz/bLlFPoIj3NaymNVQy9hInBlmKKzIyujzQcAn
4syRKQmCMCKs+W/9zvTHBvDTCcicWfMD7M2Xddn5XpzmY5zaqQCpSG4q3WIZD9GfDHbB/WEUfNSI
q82QAyETU/CJqzUO6NCwF2cgjaJTNZGQp6D2b6RCQn7zueVwx1DLpzvS2/dBpPhpYRT0uhkTSgTz
8s6r9crftI64pApFNxArr/YDAn3caWmh6Z20dNBIBIap0vjipfFr98woDBb/SfLs9D2DkWB7QRJw
tCBrgHwetu4He3ppg9tTPANq+/wjIMCAKao68EBLDxaqrgV2aaaYU4n0Xj+ZES8qCWWSjPAt2Xd9
FPN1dqDERiibrf2zHVHWOYEt104o+l0bErHBKz59vlJrM91xXdBquEcuT4vBp/+N00k/jCF/98ve
PbqC7qXYyiBlDkFi4VNj77ZwU44DitsDDBAZtNGpepQds5iBv3vR9gpTsVBl457QQFr1e60cx2eH
fu15DVpXhLVSR2bp44XwCaQlNdE6k8fo3loeFGvwK/99Nz1kd0OPKATDAbMSh/c38pbFJ93xXIeC
fsub0QONLl1VPAacMs4R1yVQ2CQRr3jiig7eOX9bVMJchOvz1G6xjy4zzACbhRknE8sigB0RCrwS
RvWniWneLuT2nPM8bqlLamPKm8AAMESaUCj6u0oChLCFGXhEbwYUmQ1DQbVENFJMuOo1Vx7urk3X
7r7wk2+LPM9ORBnKAr07mtEgYN9DqGIMmhSBy06KuAtlAKORtGaLF8yzZA6ERf6GdOkmRf/vAhuL
Mu7K4CCPBIO0LCMP4JcrfHpvkHWfwri4FPSU4gFRiVOzWzVo3qM3VrwYC2/TKqc9F0ScSUXCj8DJ
+caf9DTcuXKpElJFcAVLpxuk9uqK/QM7b3lOQoqS7kPLmxjRc+/fRnE5I2+pX3R1QHxpMDvQMVCf
Gegs7LDBbqWsD+jBcZvi1i+9WIZrFZJfEfdiN951HJAUejvwtEhvvNdvb+Bi5yPPZhVGgaobdWup
XuCAkneVO8MJUIUAUh0+n20XaiNOzFQ0FnBbYl+NgFmyi6V47/jv7tO+jsAwg56cRfk4myMAh1ku
6Ir4JbEcfwpt6mWFoWFE+UYufRKMrM+srXoL3Pkt8ovT40Iki/JccDRBWtvdKLEegaeYc7bYOVc/
x7U+F84WKzPepv13Tvq166ZaisMM564BhMleLjmvHjFzOJkNhrd8p4uqscSHSX8wl52nC0nL6Zxx
uLgvTB6kH3e0gtFEANPJ9nsIsp0BWTI3BIc6FUd6E86jZDgyxXWl5uLYzFJATdKPbLF9IOLSywLy
3aAogdodU9BbC8eEVA0CrxYwqyU80majnslSeKPT48cpRbS1qywvxoeJWrPPkqsOQdXacFj6/68j
cc8puKgvZ4kta+qkLkbOR+8THRez23eDpbZhHQC9nToyYKZwzySFhj6FQ+aKLMli7WyZBJQfJwfy
M9t+ZX3qB9HdX8HZV+fRtvL8Ij/LvRtTR+62aEtO71i08wwuOnNwc2bQ7IQzYRt3VApmIrBNQgeF
UDVsF2c25i1oVdf2/eMBveRxJKzigvCnEsssHXrJft0WmkNU6Cg61IzKR2dqdcej2QA+pf9v6Vjx
90nd9UpVh4l12QRytqhLde+tI6m+EdkTWwluUMxeFMU964KesjfpaokD7pqrR4bu+Y20KEf4niHx
cKngctdZpmAY06VGSJcU3wqD9TTFIi2ixY3aPdC/lvqnd8Q7XxadfpW9Uj1+lhYXFSW66MpcpVDW
2W2pjs5UOLhyWyMlQK3DkhTFzXbhO2X4uHVvfYLC1i3O299Lng/J9YBpWJsRYvGSc9Zmyl1jvF9z
nqY/nYOR5pnwU4RMy74jE5JGpUj94paV0M4XJ70AuMnEDV2kF6OHE7thvEtxFaBmeYX0J9qGDrcW
EncEa7ky3HT4kHk44iQE3KIXz4ZeFs8RsPVArY5omA24xAAPzpLJULxWOEXjfFFXs1vRa7NTnJQ/
Yvgmj8UsBe1MKFHf7sBSvBn4I0dwOmAq1meYtLZbp0cPQNnI2yTf9tcLNgFN6qwmB8P0Qv8N2c7F
flQylvKM5d2siXWpv3gwbhYqxuBaC7X+LbZ96+/5oZ1nkf1lyiJWGPH0vaY+7h9yOBt135XQHODf
vy28PsKEwHDfy/VJl++Vo8u0Rb1h5zIvZ7kMdCSNsgCP6yxrUKiY+EQ734rk77Jr480TclXayxvp
vNXjPszoP/x0UCbtkxhEFQYIV5f/BaIagKLOgo/hXk2foRRTBoC+mEh0xoWzMV0XsJPCIHTeof3O
oK6lJGJXih//pC6ZEDWsT/+E+huq5fFLh0rT8bb46VE6LBUizHqpbiZR1Y2ktFLXkYod6e4OvnrU
uJvTMvgS6pId3hyFCUfEKuRmmdppKrFeX5v1lN5I3/MTo1mJkrj8WQbIn4PqB+x2T6JoBTjM/wlJ
LfHbGYEnowpBQ4ab4K9dO9j9BqA4pGgMKtZpdKTpl3DIKgBHWp8o/KWsWvUT0G0lebd6HlWfH0Dy
rWEDOAfHMeJSq4xPbIrg2EIjyOxN3uWEpxSHJhgJfuxUdYgl+Qq3ZKuYI+ZtabZHgCOMnk4xCgWH
F5ywKT96Nt/0aCbJOo98PRmTvfTGDiEOn2p3e5EHW8tDayIcR0TXQwTFs8XYsbja2KWe6ZWPz+c3
SSHtHL5m8xbfXLY/s8ZQUx4+2EaeXiLtUDrXUvm55qDAURYmXY/ucOepRaH/zdz36d7wNbcT+fEK
ypyHsCYSVCnoTtyTEe3ycSxeZPdfKJEzHqL2rQytk4fBWdPqWEuOESatrzbLqudKdUAjb1/6ZUZz
7Mb2gRt6R7vDzP3SgpKgXAnoJIEBcZD+Yh9pkasMPi+EGOj72yl70ULKatADcztaIDxIXZFV63pL
+zWKzPW9fT8AIRmj3x+5nlf+pM4chsQFWsXsQInxdR912IqtKtEO0TgjbIHEp4xWsCBxGP+R3kEx
xQfRg+dtaaXg/sunMSQBdWXSUFFU95fESqOS+ZAzvmMuWcvCZ/sEJEoYj3K6NTLQmM8Ve1aVnyvI
f+gVFmpWcgWtxixlVJldrn1ULDFsbAmREoZXHBB6M7pljWkTZbmiJQ21ZBqqjgGedJQzFoGIQp+C
4ywBvAn6Ln1DYFDB7l+8xjsK0OpbQD6p4+qUtAAfRFQ37j38pZgKgkjyNt/VC3SeBtMXS5461JHQ
cakPBODrEmeqnCL/Sf2pZdre9ecFIH/Dh7xt5uR4TV/bwt9K9qXC1anny8Jvp/ydJnAWBJ2k7awR
MO/ywOmI2c+MW5q7AitbRbBTIOVUYYsMpTcnncmSGYMk5ubTiIG3gRHWWQZzMVjjztZ3mUBPGlX5
NnP+i9LQ8iR4u6mhIFvQ1OuAqQk+M4QCuAPILSalydIDWR2463hgCWc410bOVR7EUg4yqF5rh0sk
JsaveW2eXs3MVZ8GtffRdrsPwH1dEa170c62M64JDv68hMST9asKvlOLzGdSPMzZZyMCY2Xp3p+i
dJIKe5NzEk/YgxjkD/Y/aM2y/q4JPhGqdxYYwMz42ejGWYuOkXK3LBBz8EpZnRmY50bOnJ9P7OIs
7387wTKAMBWdC6nTNjF/MK7WxI2xFH6AHwoqC3ciXO6rL+v9aluztQDVZf/UVA5LDfIW53VHW4P7
JxULYDPOQS45LQNmr/GYTEg1G6zMm+VE+CB/hvhxwmpXQFmDUPCx9qBzW3sjOEJtp/8+UvaETrMd
5uOhjntFwXQtruPzkBmmCRYvF86gkRIrKMwH32K4mHJeNLUHCrGganHGWOjeaOOzVSshvGoV1eKa
w5JfA7T6cNRvtJ3r9W7tCDeRi2MrIrGv6KYsITUNFUnAdOJilC4kcPyHqyBWOiDMgMulbVn+ze/F
ydkIZlOgG3zayxiAMIiQrb/D5qNFxqhxRLH2HLI/sor0Kz74Sa6rY3I0rfsxa7ofGwZhpd8O1mx/
XSoJz9+epvKbmU0GfF4XVxQZChDmZV2cMuaCJBPSvGy99fUlIYSyApELHeZrIDCnc/VQnq6ufIbC
L+TdUVGIOlA14x7Cm+LCn6o8NLSQl+z0KXgU5xE1eHACBk/8Wu6h5DKjx5xzIY/a9hoU1DFO1Xg8
RKold/bLk6NmTR7IwprxYbw4Ze/HBHaEYHATV9Na1QpYi75H/DmngXcKH2dwtStipUj7KQHP44Xv
eZiOTpvXlsaoioVbKGqmKp0oLg3B0xw3Sebfauk6ArQ+i+X78iRvDhmaD63pyFavmNY8Ic/dpFVk
kV+7NfSWyEtJAA0wTidBqPR+Wak6OhMGQIriU5H+hQqF1RaU634Bh5FaB6SROv94w+MswDlfMu03
WAt4IcmzmyB1WCB/KIAAnkVwUcNzzx1x1ZIy+4W+xMC1skpk0KSM5aYKR9rHQMCWIA7LTT8BOU3I
eG+2QaFCLVYPChaVFS4RV+/II4l+7DHIeqDiQkFn/WGB9P67OfVtOcxpjMJzXIOUk1Cw2LgL4UO2
GCqSu8jXa3qTz0aAzZRn59zRFA1J+ocRzAerVi0Td680xSXqeYk+31vxg3Tr0XrEf9GbyqboTa+b
K7StTyMkMJVR3OSzvSLNmTgGILHWq0DNKwTM1ptuxks6S/5UXeMvVaXR/MmcaNUQwZEH3zIDgEfp
oOsn4qPkiTHyv6tyb6YjWSBuxSuDFNFpUqSATQse3pYk1gdQVngSrEacrXcpRDynHQLAs5qNSXxf
3COQMsoNka1uHMuNajPkXijlI4VD6n1m/NLL4cMmg+hEcaxKcma7O7wQpYQD2JDjXDPHjaN9FHRA
+n845HV3+8iXRP1ZFpvZcYxS9sDJQMUDjHD1/B9duvI+dK7ErLfWH67ZWKmDDU18ZiIT93nApBHd
YOHHQZssSB9lgeW41zOZp4sLHj+XYopIwpU0L9Q9CZZ1tpafrtQfic5MldOTZ1pUIc5d97QuJjaV
imzibpFTWTMnwNEIOWuP0Ii/eoJqDd5iJ4FmcAkGsgfKFT30XHHbpJyzR68kFLU1+Q+q9s/eY2tR
j/AmY7NugPnT71VcjcjwzeAuLhoTJkEf8MVq40k5Y+n7Gdcek+/mU3kxwhR/8Q1Isxj29bjm9mDS
qKw1i/pnsF+aCNG9S3rEK4WoQVVS9muS7m6dNEnSBfb4iZFeUVV60V9B8bp1+TRdmxZXwo4G+yHS
ERyMplP8+umdpT2cevX9jc2CQxe1rmvKTFkuuzXX06N9SKtMZtYjFRHw9MB27UM8ZnWylnH9zsFE
R5CKR5xTOoVeZK3Ou3TfJJ2fx3BPzzWinnnmpAAYy4Q4J/5n8qkb0+jkOJJA27Bz3ml5QxLY5njm
CIjUBPdEmFaXzfWZsSh3fp+4BRssiuFe6yxSpGhBVl6lZX2Ob4ballAgFFMUyuKAiSp7CzIirFhi
ifE7O/RV62IUWwRxDpbA97BL0X+rIAPtW2s9Fs9W4IuhAp96rSi5esbGZFXwOiQ5Aym5eCzAn7uV
6kj2Lt6RwIFRoEp7PMaSbZt7FbfMkReMBp+pmUfNIgejPorXEq1UdnYX0DwaBZg+7d3qoDkPuB2G
bG6zrI9l+fZjmuyd5b03bCcCQyETisrZ2t9GgDeo+cTwav6r/xCPJ5G+mwoa06dM8usfCpkHph3B
jKIPioloSwbFuf4bJl9MrBMACY9SPSuzA9H1mO6Jn5G6x+CxvSlq51SXKAeGy5rOsXgm02sopMCW
rtglJAspTJO+1tkqVR01x7njpFflgllnLWrNobIHTTfDknFSXBrvhH2DfU8okm+e4d2H+xlGxajN
foXguiyaIK8Zbqb6SOLyZ/UO2WH81l6AdirJQzrWP7qW/t1LcfktFJSeLYykq8c3IUgKQLxdCAYK
p03DXdR3WmUfJETbSklTTu3/lyEIWqulLEfYk8YQEgSOyVnWVV5wdeNnNBFdAIsLXsOoCNVWKzDJ
s/UBP2dhwxCz4AHL/xTVW+XSfPjkImEmkLb27Jzk9FSPdrLXjuvowCeQwuoKx3ST0mGzQApSWl6j
GORyAl9i5vyCgyTcIAuFFgXoPEZsmLtKcZeas4O6GVVEl8TOBnNjLnozid41+e003oOKSPxnbcak
Hfy7kmGfVUy3EDLp6xf9KWM6hLgmyXXQhOOqEcfjsElRZZpyBGyHX3YQPtcUMCJfSmKroy1a3TXp
UeIqOwfAwrYQap9y+P0uhYUsbIhPNNjuywWYte66b0iIhwO2tXpxubxyF8F4F+KIoLBI5Kl4ga30
LZpaWY9C4ig3Ex74z8+pMxtoc0ro23aZeLWmTOMXXGUjxU6SDXeXcy2CWthDc+kKOxXAU6sczHwc
3aHGohRjGOpYTURj5bF9jsGfpFFhnWfopBRnupyAVdgIAPir//GhwiaKXwSBhQKMrSgzusYHOdId
/X8Xovf6jyqJIiSQD6fPBseIINFnjWVgyyzf8oTtVzJZky91CYyxp6P21Mx7JbCJqNQjFYESbKH/
f9D5FmWI7p5I82XbpgCGftEUW0BZOvuDdTsyZKaTUFDzjMm54lZoOwNGAXKBQCW3Kx1MASv5GonN
Umju6vWrn4FAV0NF9/oL29m85LuOXCH3pfjLLpmb3tkQX1DwW5GnXxW7llRAwrIKCEmREcQX+seT
iSptRmh5MIutXg+pjcEU02sfZwHttndz/A2fn2zcpIYa4+AFfDt3tE0TKADwISdSUHcrYMORga1i
DHFPrIc8kh8Ud/Bd5jTWOF5WlLQEJ6pQi4hbLY0ECIHfJgird/QOMXEb6vEcrBoQBC69YiNmj1RN
NmKA4vDc6iximOSZsLWnoD1+ZLOoL7pQVXHLJNQlQnkFQzp8ceTh02Bcv4ssEEhHzQxW6G0uG1fV
MQ1XdOat6R8kO1ynnQQtlJaN1ie1haemBa8VIYgExMEv/qhSf0m9vA/kEoMUaGFLSs7wCUjA3Odn
f1u3AGoGobaUAF240Jclrrh3776yAz7XmgWNqfACNMnCJKjIfPs1MAs45v7uUzyfIknIzREfwGgS
cAHC0rZSpDegzs63kvYDDPOk9rf7bmYHRs7jyYUUA7xH1QhsG7UHSkV6/ZW29Gz7imo8lz3gv6cn
wXdbDITE9N5BpxSYPGcVGM4Bgs+a8yeUIHXGQ8kPH7xv33rNMQrWMPvk6kbPPRKuoOBJk+TMwXLK
XzWA0iYcE1zGX7d699/cxM05YN59RSQ2giRWh8Rqoo5HLJhTlH6AmZTrwAfzwwGF9FiRhABFLukv
ENG5Ga8riizkOA3Dm8XFwAKB/NW/bHbb7IOUlgAtMxRc4qWXGQ+S4LwTZ+QJBQJV48ZFSy5tih2O
7BOCsndOAw7TA+WmbPBxvpOcoLCiH4NNNOUb7WSsiwiqyW4FjR+c6QFsSx3vKoX9VVcTI7FIzdlV
SaerBxWuwb8X5tPO1rMHStKyys4EBPQJnWXjEbgB75/VKF1k2erRqPOwyW9irBfQ9dMac9zH7A22
vsZCrtfI/9SmtmJoHzYoW4+MocQeyKCZEt35I2ZxcpR4W9GqjK1VuFWEuZFXCL9MZO+ahmGFxP3v
2QUcMk7YWvg8/zpkDVpEzGw9YYjoE6gGD3yv/Ds6cWsfnl6VDry5FeV8bN6sLG7fx3p/BSqf8DEt
c5vndK7CRTsEtuGeSjXXU4ZQ/eMsGWW14sE5CaUTBdyj3kmg5vNfxOf0g/fNPLXVl9z1+iRRH9ai
H+GpzbHt2bq4cmSgzxDUPA1zrtLHEDf7Xd3GadfQs2++GTQkUzA3+ZNf2hWNd5vZHgUfuG6zoYBM
MASOKQ8kuDQ7P8KMJyaN5TqZyc7ucgeNBEtXBDg0+Sc+Q0ARami29+xmwVPHQOSmkzZKTGwEsVO5
JP+o1s343r2MzDTgCn2NJzX9dXme3r2F0oBQ5Rbg2cTX6HrrY7iGMf9+hDAX9jPQ3fItBBY6RPYY
o5KMFkjPK2f/fAKOr88O7AXoWUTslwNDjfH7k2wMHRYhhHXSSMH4O+BF/eDHUxkQ5GIviLSTvQhm
edux1WNi+SX6lYrprEXDEaJf8QLCe3H6U2UbC3pOTiODYPdR7ViBJZuY5yvRQua8JF4iIUBMQuCx
gy2/jXlmKItJIE6O20sr8HLC/JKWRFQATR8QdPEFUsZtUF58AxbOw9b9fxyp1t3xSAp49BtPsgWH
s0p2CrxenY+irvz0rdU3bHCl6wOqaIa0/ichu1CkrTHwBqg3ALM5aB3zGZLXqef6Bec4uXyxEPXl
e5Gl3YCYAHT6LvImoGDImgMYNUADkU/tPH9AA4d1Q7QdSXXUtHOh59TTI6x4yM3qgstwTJQnwS1q
7vYlPVzcuQpMKCpetVz940C7/ffdYiJ/j1lhYlix0wtnRradoKnPMHLuFP1ggYyIxKPUH3Ko+VRp
hQi3zD9I4/92cVBRp4MyV8iRE3HRNJQhmS8QgjXmABCxm2QCIJTQoq5CEvTmx3IFe7Vhqskqbi4h
lDj96dvk4cZng6b1eHkClOMALs98ZPDZMT/tnoe5GYCZBZQgvWVwFt3CDD03XPDBnH8VF0bUl8Ly
aiH7ahKwasc9TPKCgRTX8Z2gTl+gGzEknMLzrTjS5RNc1lKQTgQNjZ6sn912BVd3syaEyNKieHJU
V5T1z8deEwTJoX6LkB9AchONzTjvGRCtaejJ5nXlDoGBJx5EGMII4T5oO2gU2Xe5k3bmtQZAv3Ca
oTG44JKVxL9giPEfcpDvRmS+H7K1qdfZBk/SIftBPUXAV0hTqS2GAl4/pdgF3Di5/Ug8WPgv/IiR
0U0GzFyPFehgl182ZZpgqIDYp4Vyaf0V+fCrczyJDoDSMR/swmY0p9YOPG9PGpN+e8SElsXEbFNf
e8sSFtll/IyoW3Y0WSJhrER8in7Ck2cLDJ+T6yDN8FcqUPyhn9gHjdaZ24a69ARb8GTEvmxn9oCn
kbgNnnrh5D/SuN1dbGAaL2VN2J+xx2kGv+AeA9hpIX0qpKD2YrO7mGdqA5miMTzO3nfgHm7I49VE
q8wkp0jMJIOVSieQztbJ/1RxH9Cfvfnjuyc2y3IGadZzJSnTq/U/R/NzPxEWwdllIiTNtI2nr9sH
IBbC0uMLmh4p1fG8y0UgtFHLURSHg/OBdv+s+6+DfLhnIeQwH4Zl/JuilmMS+96hM921MggX1ZXl
ZM4wFM5j4yDBNjWCXLqUmO+w5QIXGkr6qix4k0DHfU0E4msXPAPgWMPaHCBx87JlBE6UQCmQCqtx
GTFwV1Q+AISJDdjSdV+/iSEbw5903oBJLavjsB2XBSJM3YIc34z3XGLisaGey0eZTmJjNzggVOTt
hOSU7tNl5fhDPoGZ7CSw8Onun91vXf5VXmW10LGUbGxjWrHxs3hzpfOcebXvm1kC5+j6oajRRCqw
9VLytabQHtUyq5zMWI35xwyZeWyHr655BAPLE8rM4zl5++S9Z52/kIQI6SG+TKtInSvnJOBlMAs8
lYqBgywMpRiBFBhTDz+OLCaHhR7tu91bmFSBkHfLUoM/A8HTB/GxemtJ1wN3LpMMNcnddtxMA5jr
2171RWQ9CFwGbFnXufpHXfHR39i2xD7BtQ8sW0IuwtdvyOJuZvp9Sm3hVAOsUkDUyipcpbrEA7Q8
WQqxFffbXxAinZ4mhn3lItgqqLXLEpKBBJhe92PPxWcXn4XbQDtrhVJwkOvoNb/tyJySSwBmi/i+
OjQLcK5/4B7oHE4g4hi3RlItgnRsO5TtE3I81HH1KqTM6X0GxxBi9ZSv5a6Ufyl3hilZ6+CHO0ML
uanqL6kp8QkRnIesa1U3cmqDyNM7SqxRacgJwXaCqKt/yeSfbznO3+aFp6P9E116rrd3VaFYutq1
72QvgX4fqDrkYzOxYCnAFQwFzy/6AJEJt/UTCjkBod3Cf//w3289CQ87mHvOvON33CJvmBbxGnR+
uOTS4j2G3T2GZt7CD+tEWUskQZLCi31RYwAhGpBpnbdQH732FUf+UJhZosA/wLkAsABnYAUmk2D+
8uKhydXly9c8k1w/jQcyI9MzSc26nR4O3cLrROzQM57Njegou4I/aiCqafzghgVX2B9xtS/fNHkR
yNN0he2/T2ghAnkgbX+ErIusPj1xakh76LItn6+Mp1UhGOoTQmOq6OZyET4koccR1XDWatwLqpir
tLvIJf/rLm2olxQN+cMq8BogiWA7oNIHRhf8fL8YOweO+DdXbff4jVSPkFi2p0vLselLgPaqwItQ
GPfCOVp84NO9v1SzGdbwh7zcSV+vIcnTa9MUv203NgnNUeL2WmOYxTXRr9xIATgh7hyjm5Tzqzjk
Ful+38FgnMTSNt391I4QfETJ9zkw7kmc/0W2y5QDoj54UZ7ZTDm4mYiPXjwe1YmcS59QYnwTgjWa
i94HUrAeOiS/Tg8mrmveQPMWYwVPrnxmcLYbSCdC357SKOTPHc0RJ/AP7Huwn53wQU8Zl6NCCyRD
uwFKlsyoxYRmE9oDJQxvXafrVDkt2ZdXOMZNyL7abz+p8pUz61mz9LTuZ9kwtNhqHsOE0v1/5wup
Z7c/Vrz6d9uUpuMIxvHW8t2gQfwR5j09x9kGUDgYPCxunQ5wnmBojkIAAKwavek79wpwGooRBSzK
UMLAl+JcbDCtP6k/d1gjNrSlIv0Rclt2cMdRnhRB8uCiwU2javyMh8goGiB0g4PVLEnALRyJueyS
oroahaqM5ocgUZpbVQO3LUxUJl0LO0ZFCq3WGt0IwWrDWfIMEdMLEefNtK4XuAb2KVJdJ80cKcZM
racXm1pyQHq0OHiS/BMSbCZiQR7a7pIlGlw+TrDFPcBkuJAtQpPvmiHfJZ5uSbvjcwi2p9w7OV2U
tafyfWusnOeRro5NRbsE/KBbOwUn55EN4ixPboBuK/Ey6poPtHscrD/kUS5QFjGXIqXujAb2Jhj5
kxMM1uA9IX/hSOWg6hsL/awFZkS5wPoAkjhbNyPVUA0otxNfr7ny5QEAZsauFZS6nuQCmGrL5VqZ
TuE0C/jwL5VgyVI18zWbAslgJuyH6qgvkrerA1bEAH9Yj3pkUg/le4OtBOjyKXGGsLTpW66nsz3z
ngI2dv1gG7qCU5DiZLm6P58wNgVlFd5vPN2fMUwlMpNchLY+0nefajvzzA0RyeZO1q9hSfJYUrW5
dIZ5GE2d6/rJbBQqDWruMeAjI+8B7n+M9E9eJ2b9Tbjs1g6xNy/FPiNLb/XkiArNZBJvK3UzqPFt
rFn6PGskWGqB/JfD2W+2D+kpl8wmHtrvvbyRf6l4w3TT+oMaGQpOZeK+2g/12pmOuUGWGqHLBUUf
AwEEol4UWnvtuRAfUh0z3bbBO2fGSDHFGfyVlETBIDPC9R52ZC9Bww9wTzxOvZUCzj/FNANwtvhH
ewG9Bmz3leree5SosmC3LakQiPpEzIQFC/a/ZZHDX7UMmbWh6wjRyvt6WUa7+pi/yzeGS3yFRBIz
+qCbl7b8qp6A+G2ZQVtGqRkdtYhFQbIuSEGadTZMM+LGpOu/4REbnpHc4eJk0bvWFslSa98SDyGh
bkntTeBK4U+qZM5j3g7qPsiT5iw3lcTsRW12tAXLk+xKT0G+cJIoM/Y2abeJNgr917QOpniC1cBo
4dg2qAYDILoas80bRVnHSa3MylEtYzSE3gC2uq5NQMuXVz9YQ6HPS8bjT7Z38c+npC16liY5wEE6
VZXM2jIHGw0hpjiDrmt2Wuu/YHmnd+w3moizxPe/4UeCnufYyRVNBdl5JvWgGSk9nOVfueTyMODY
9gb2TuP8+MJKgEAA6pvLLFgXtjTBcS8GzC/JDCsLF+LAC+piYzI/7n5riBcIt7Ch4QKZhMzGUYrr
bz6RWME8MwLzbdW5g1sO6q0Ku98NGHiqfgi/qQ8BFrbMrqjSpof9fLAK7pXqnTtvVWQCQvz6g/Rh
FkdR4NB3MQZ+vsa2ZuPXyVUA9UBlgBRrhrdfs9JQ0RwR3sq5Z7ufNhQ8Bxn3vUDojneOsrnmbTZV
LFdj2T/MQrqkAaXB8zdYm4EMx6O1BIbTlxGKFN95OpDpka+ddZdg5Bqxxw3rcfBi0UB4jqjiifvI
iwal+EBFo8UOuwzwd5GF4UxrIQQozLa7DMSqT3f+DYuYBLAhue+nEIVu22TgDag3vVHeesNK6PtL
CA9Rb/zt3kcG3zkvJZwA7N+RV5jhQIL5aMsOg0UmXnKy8WvU8uoz9uwvyLU7JoQT+GwuuB69qJGh
4KMIXYI+12ceA3w74Kl9jTgn01jcqJJU1vW8ilBcG5GPmyitTBdTlKyL4Oma0bVvrMu9p7625rDY
T2AQBecbMQYtcw0EIq11EjEYpQF0OVt157wRmX52apbSb2f6KAvG7jxBlE50lkcn5aizjf/+7Nre
QsE4bbuKGYL6OQuypa+QSAwfiPc1ERXI/fU0FPZuYMn9TtTOym8WUkSo3G4SZfNmEbl2Jcby65pi
ddReOZNNmJkS0PZ72/g6jGgmePbvKmWs9vkMo7MdPYwM1+vvtKWuiu0OekVO+7mEetsuriUxVcCF
TUmLt/CnOcj28QYK+2IR/2pXRa1R26rkMsamZQ08kYBA0UrjFMKcvjNbT9nivJ96CDVFZ6rqMqBW
xhg4aezM55Fa52et8hE279ci/QB2NQ6/xGIUMDWrE8E4DkJZoMSqoSkI8ijfm6M5oS3mKMWSNK2O
chBD5h35OwU9mejnm86OvLFjs8qk0up2RDwtvnrdU25bh97GVua/X9vFrRPocUwmv1rxVtIkZ8ol
rp57UXEWz87j/adJihI8o32QQpXQqyZJ5LIgER2p20Q4f+ikrYXlkscW7IOnos07hDGIamHBFTra
MNlhThcWH3+d7xrnSLd83KFqNYn2JxJjKvdf1tlp5+jTTo3IqoqweKlxDF/TMJvFnKdQOYT0lJZT
z3eWz3q/RB3UYkPSEC42Oh+8bvQsid3NDvQ43lArZ6VtJhkbC4BxBEyKFUOQzAPf82PhC9AUHHud
emTo/hZzHfAyAAbVpLXrwRc3Xc2J5Uxb/nsP/ElIZ1rNGHV04HVOpKq0j55dKlSazwBR8p2K/cke
x5bIBWi/Yik8mOIUEt4tp0KJDOUgrtskQtol7G/bhrG0MvanlZ5/HBk/AdTc7TKn5N2m+yu/oYin
VALqPSvMfu7qEvSPt0ToZf6DO4MfDxorajU9tUCPmul6EijJRJ0vIO9SeZj2DZ4FA/baeEgnTCCs
gf6WDewBVkq0POnDhl0teXSz46NYLuLYEW9RcniuRNokHjrdplAyTHfzieOPUIL1KQMsH9jJTY8l
FjpjtiQYp518kBNyyHI9JggC005lGdLYquVbiurOiL1G02iKDjlWHnPCRBOjhOYK40fH7ORDFglR
CEInYkBNJ/albarQ7dn63+j0OUcEDLe6cDFX+OINWK+3jQkqOhx3h5W6cL/rB+P6H3FDsf0FML8K
O/eTtIvdbE7dADJPCvWsAG6ByoOibTeFtUGKIpa8gJlFf0Rv/LOkeX4RLPIXBlHKkNavU73Q/u4k
48jP+anvIudKQoC5k0JSBfdITjw0XsESb/KkprzrBJshQyd2S3azBSQ6SxnEn9BKaXs7UrI3Imjq
vUr6V7fkYIV0BX+FFb8LDeIunoYyptyh3+vsatsF1eK/UqYMMEdDtEHthv6cTyX2qybL4YelLPSI
dMZzPFdwzpzuakxGLKty9+7OL2BwNkeSIYgWI4vXIQ/0eGpUmJjco6eAlKoSeWm9xVp+6qZcmXj3
9gkf8yi1q0REnJ4z7bkK6Il5QV9m+TcUHYNJCHnUDL5aNh6xcHwh978UMCwMnKX1AYkXXfiZpRPC
sXHeMlqNN1TcC2cGX/g2PUhSmxAwS/pOLxg1MCXHNUZwXcYAk9Rssvu9ncO/q4YX9BPbg3I/JyRt
PVuig+h5tqJvQJdSADyuJGWI3X2BUPTpgGyXifWk7/dxbLPgE6ljEMgWCPx7ZYUCFMxxMxQAQzl1
yju2oapji0v+USjlUNXQ+v7ON+Fu2oth3v2w3NLk663zpP0IeN+ATm3Lp7SmYy2lfbRHQo9SA8Tz
b8SRXdJAvvCtD1MkrINd4Y6PqjN6g/6D8Mq8DuNwz6bEA2/QFIFJuBS9y8MUu+s5g8C8AN6s//A+
VTNpcEz/l9o7jAew1GKO+94jmZ3p5BPlgBnnur4n0qwrmmw6JBy4doQPPCamjN1dCd+OKFw3MJLV
7dz9wSl76o4s7ymVGEvdqa011dk239Za429o9q1sgRHaPbfj5gaSsPK8EO9+7A0ewlRN9fT5WwUu
+hJvDHM3eegIczUt9op2/0eNIso3hhWKRtjIgipHPsssm+EsSoHznc6cqqKnDhaRX0iWiEUa6ZzB
Z8lPa74/F/00XuOLqFqQ2TgMkl/J5SEIpzROFfptRVE+OV8M9yJ140dPPIpfE73fzTKv/Kj8o0oo
Vv9Y1VPkD+lf4LB7bBta2IsywIZoV6NdBwR1bTCxnLT2UbIYTAfVNpSjsSEWRDj0eV5qkKIPqLMh
y5hz/Fp5jEtNbNZAJkPDMnyyD0WaS+U9ctZjeFB7HR7kK1t+VUu7CzFChjRHoeE6G1K7yCqxacO3
qM3Hv88gapEzbf93riiSRfSSsCJd4e9AZxEy4uKFKdD6e+62PHtFkW+WD04+1ZCQjogr/iZ9Zi89
5vXneSt4GgmgaTAs7zxUemb6MjzIEkEpTRYrNs5CzIJ+Ld5uodQYIUPxDb3QdHyo6AgH9NwgPu9Y
iZuDuIM9qph8jq/5F+Yx5pXKeo7US2K07unazXJvLksAMdBqdfK1sBUQmZHqjOphsb8OsklZkDYV
/NaxBYYCMiktWHomLt41XZrn7dYw6qfBCvMbbQ2wd5cXuY7rF+wz6jEl7mFzZNxtcZCh6AhM1rd/
8RTo77Zdas/LMRoShYM2HFzpr4UULRGGcepPqHk04bJxbFmB64zguRnoddGDxDHMayIFgcPh9Esc
wuNox61q1XXdYrkMlhAHn4poWz7/nMa3DL8LnjsAn8MB/wrFG5uOILTJ2avnQWXswfFlbN3CHWf7
UOhTd8l+dp5bhirHBB1AhurHpwkCDDHI7rxpIkHDKjx21UOtcKpT+Hy7doqffjaHShs3UyuzMnaj
FAgVslHDGFRY6Fm5JoLmQEmMlPbUAzKcvVGvVmgWZGQ1D7b9yNtIRr4HtdItl8jp/J2iRP1IO/23
X5j12DMXyAvm6r5s55GTggXbUEj5uoP6nvqo6mHA/fJPGXLLkkY0I6WMN0NZrB2tYMRsHeWRv7nC
N4e8969jgZMFaKhe+93iqU7MOlsY9WQSJPoT/hCCGIxp3s8HnAk5b2YpJEu7oDIBLXf83QwHlAir
eQ/HwTEYNUep6RReF65mJhZdSONweNpZbBDy4GRxoQQ2WapC7+Tupwau5tk2aHYQyVlk+13UoLVx
iLqQeGcZ74CbjglFD66BmkCe1s7RHeOdXS1/azgUy7YdRqoAYLsxHUbJJLABoT7z2JT0u3TamQha
TZoUeaxK60uIRE6MvGwejbTc1FJYBnWTpPf083RwhykFq1huz08qnX+nE3yFumZC9+dFrVGa0CrL
7C4Ml/hOnfUHV0P81sIBGWXovLnLaHwTFJxRBz4LL3OvrT0HWcxRx0iuaE+NfbB2Dqa7jHQ9aibp
HVd13PQhFJCnR12JGHNRZGN6ZtY87ZxUmUNp+HHLfo3eEl1NiDbkzxE0XQQKKT8joqjvv2UzFN04
WEyAQdUGLh/gH7Fglh93Qs5weMqffbmfcd+jqpBBLuZRXipzqi38cL4RvFVzRvO0eqGMzpbQrRY4
yPmFf5rxDR7icIDIxITzgxpbEJ4V+F85qKXa0eEEnJq7kkCIDVNqJADZx1oPD2Iu8qS3k1pmWwTt
UuNSCI8OZoRi7EnzM2QfzwtZ8EJmKW+71sez6nGPlfFRSvgt0VzJkPckm8A8TphoUSr3sIQTIgwX
EMqj3VuFDxxOdlfMwcnyFpVNnLhXeOdWQ021lvUKY3338rEN8jFu28GrtxwobbdUhiB6XyF18Gyb
QtX+1qmXLBPAvS7ZBLDilck/zItDRTcTsq+W2WqkZY8YCV9rPfZTBbqlntIKIYw9Yi5B01jesWnq
Sjvu2kaahQTI+PaEgVw7bvE/dVF7GmjcWMkZuL4VDb1BKo7L50dNgfBhlR6nunZWGJwL5HHk0rTn
59gomCnOVdvMxHoZvJ2VJv68g1HznHjOk6p1CRUBSDkyuJdKfYYEwDKv6BV71X9sgJtidVY3iVtx
wN4iQK4sVGkyUIsf4UpbsVKJb6C4Nkbr5tNDD4tUOjb2WHKhcEL7BUeU0oR854YEeSxg4sTXPRyF
8ucxLQlL7dIYxlRmuNb2KQc0wHSZ8egq37B9OVTB0FLixp3/DNhhBvZpv9eDS+77vpQOxvIoizhs
MzyUzwhByBUJRGf4NkZKhZ+RJPbyT+LtfE0tvdxjOpfDrIOX75lDo7ObqXBs4t2SoPHlKCynlg+f
RMqFhWbekoqkUw6h4UC2oTZQQgHcfIoTAkwtsS3dSqfQJyJL1cw/HLEdYoEKML+dvF09e0kpgXEH
4E3ae9Lf21/KYwaB4+F0Wnpizy8C/DDuMkuKpdSYPufjHmoY6EIjV0StZMKjHG1cFOYr9x4aRTW1
XePEL3Z12uDIssItk+XFPXVF8SdiNZBlwvkWAShLPQOKEU9GPxQx9ICj5sZVsCG2kvxvmJC4oX+x
7ithdf16DHDqg4yRcctm+/jghNAVlNdweSOyzduM6XGCIcP3R0jPmNQ9WUW3IqO8Cew8o690nB0x
2Mv48DRG2DPbNNi9/r6/q3vlXWi6dzn4ixAHctGHJtAlCeokTqzufDwa0UY6zIjJZwn0UF7sZuo4
s1/CvQrtSLEdgTGX6GmXWot3WOO6xZSAVQ9HQ6ViaYD6ukxKtGTt0PqNSHsaIigoRWDThjv+13MZ
ol7UUWtiL5QHQEf7ziztGHZi7J0VrVY0bSRLYdculWG4YCShk5NJp5nNGmTLyZQXxmqw03H902ot
Jn3eg0NVvQ6/wN/Ph07v97E/ocMN59CiTohG7vqHro1JrD1oaElRVaARn1GCpva8UVWnJ1tkEdS7
4h1Sy4V7HkLzeVOxfsr2dJ2sukATgpYmN0x/BbxxrTZOpGt6whh6ESQUxCKtto1f3y/YMWZwoBmr
TZfkMv7q3q5S3mw1Wxnc33tqkkbyUQf5diW2UdpytmPO9OtSOmfnenPNbFM8GL0cbMpLnZYyhUDS
jetD4zPCUyk+dVEyNet71GJuckgvnep4v6Ja275BbXcuSCmPAW+3gHrmBnjNtJrKrOvCdFPQ+XLj
kT5XmKyPAAmemn+IRH+Jh2HHN5Sn+nqYIYiUwBdbE+1fdSlf93RdxNvHNzwHz5onEUjZhaiCyZaP
x4igmdoHoiLBDUbf6hgLtYKwngGGu+Uwy+u+Q1LYsNwXi0eob6h9B0dXVQH6B9dlmG6y2NGEjwAw
M7Yu3MZmEJeM3css3/8N1V9rZ3TJKD4cE+yoEhncYT+EHGWyCppg4J+wF96ro7PXPKckPfgH7HGn
i3G3QyV5DeJjvhRTN6XOEAYIYxR4m6H4Zsfr8mmndppuTn2DL7+abXP76EPgbEy8H4KzJUgHZimn
5hx6xsbGhvKY5wX+LJrHygiSQWhV+ycM1ovcyRYeGswTfczsA55k6C9CfdGl41E3HF14/aGfdFNo
bk4UXX0bAuL/xsryT8qCwr68E6bEgKxQaaB+tLGUKSstejsHevmoMM8W0Q7f05w5Z2BqtBhky0Sd
ftIFU1xtG1cCYFVQe1xEcmmRZV0SwU9M+LBZ3sjMr8S1pttFmYLug8A3dJW7kmZmm2todfju1HO0
OayccizW6RMpDkGMUAfi5Mfg9PoxS7HCXtjeONS8XylqzEZtqCjpewLphujjLtvQdgzgtHrvwitd
sZQdEfZoDAdjQysGrD30UYlWx7oI+L4KM1BBc6Eo/bJXrtn46RPkbQPj6E+pX1ol5QUgcO9mAh+Z
fBGIC8T5MWpH8wkwRkiG7lgh9AEJB59sLOkFEj2Hdr8dAlj5Zv1AeAHl4Gk1+VPqu6UZvC6xmAvG
XFRF7ddT2Fl6CVV7zbX05hYjubWN9gUwzeZfBFvMfBasWzixcQakUCs50KqeAi+bDoFzkzZBacLX
VTRocPGikobJxRATl+nU/O6rT7Ps6fuA53jxm9m5sGj6VLO6Eq+1lqEJqnEPApzE86dDstv++noq
SWbWtPV9gXf9cfzuhOD/xjiLdIA662LzxrkQuxnykkCFW9MPnRpMPicaRxXr+wNEku/mPgxEj9Zb
xLK+BghveH82a4fMlRkx1Ft8bLOQHfOnrBL6FHs/hIW9XxDRZyh//Frl+S/g6+irfnWHoii4hsb2
g7A+QCPvPN9mhEztmXgx2Hy4r/JERLjKwKfF4U8JNntYYZJoCUtJ9EyufYfQz9WDzdpVPiwR1YWO
gxCogNeRfWlaj3voSm2TcnNUXs/YMi1u/JuhnhdSdSkTkDuR5mkQBzo+FxATEtmYWVr5M8iFmdPc
FOZX7FTeFaaElv3hugzFjEWeHlI4mbHz6b7UcuykwMjuWp3Ip0eLWj2AkJRSX/iArxZ5CgIaM2yK
YDQQ+bctl5+g8bWIaJXOzlckjttr+hddGsn7yoUT3DzW25Y0HuVRcD40c6y6tAJxZYrF2Up2Q6Rd
F3VEAfIpV/OdBVWQVj8vKSuA5HdVLDKst13zJZIcrr2+N4aIAPilSqtQ0NZkdRzi38d8pWWLbiuc
lpZLO567R2zIVQyv6RGiYBiYDOiOnblzyJO6xE3EPCiHwW7PSzxZJTy8H9Or0ciRFdcujE8Ldkmg
FNyJRZe7MWA443OqOSGl0ntosoUdqDui+886gngXwnBgJeTzzUcu8L49QRKgY/spzHs0gmPfqRq7
9DnLiSqIZtjeEi5Y698KLeke52wlARZ66J46svomeXQ+8bNo8zNzMWwK9O+qHjG9w86je7IHZlKZ
WKqRw8JE4Y1ji6Wlfz9sbPrk4dLE6OYMBmDdA7HbYTxS3JsJEzj2KlAhmN5C/wGTpcg2RcZdUiSH
uuwjJkrdKj3aj9Jy1WU1lMWaYCowmYl1Cnycnn+lrz6Kd4liXCVRV9jzdzq/Pd+L0RdYV6LyWuNw
pITvCqeExhPPLLuipIVyhMecxl4GusdCmAAbDeKdJLOSyQ6WvG/aIQkob/rMMLOqJYoDj4FQ7fKS
VcK9FY3X8AFwBazW3LAdjAnkjhgRcxwezH18juTdmvzyFHxZBMptnD6bUmMe8mVSvk5ydQ21iQS1
Q2pmtwXHBgRUbYA8k+3fRs5cB3cJUB9NvOBbeBEYhSx5i1pmA4kdQX7lMnUDRUped2TCxWKBjTck
WmowcHf16qis/4SdDQiG6MawsmXRaAPWOhBy4Yh9wjrFirqB1NCJ0vLa7jCewyTHdVIXD+cXYoEF
raxkjeNiFshSDv4qWEEnwnp/yRNWW/DIKSbOBm2/U6EVmW6AZuHg5Vw9Ef30XJLIsCSen+zPUndC
jkUW9cGOWJg8+fYHOJq+2AYBNwQ3sC5OejmuBX+ScXedNKk3wd2YrSoh5cgviv8+bYaV/mtdyWNn
iPJEcxqj7mT+7TvUSRZM+UfH1E7z0F6crz3I2D6AWI4ow8iu2v8Z+PjsaoRfG0LFJXGnQAEpPoz2
/1fPVf2FmX+lvUg4kJCIAAT3xLcHW4ffKdFykap4HLdXKHdNry5MH1Ez4ZqqLwz/WlFNJ4NcgfrC
wSsqfZ0SojIiUV2CM39wEPd+/mX0ghpqIYEhokF9bW7c+ghrwT3pynwy0DFzfa2qc0Cbc4H4XS76
LNHxxV9joc3whiXs7K+Jo0zrOJ/pQI5iK2UMh3ZAv9EXarULreMCYdawxiHfXsNw7gcq2BF1Uop1
+TmHdr5acaHEJxMOuU3S2qkinQSIaZUBc4FLvbBBfdHvM1IMkU6PzBXqmqAg03ADSONdUUaF7K9P
s/yc7YGH9jO+94nPOmaTjbc0iLeCaZoNgHW+WzwdwNf90PG7emfl94KOZ6nJ9Idu5wzV8cYdDDdH
pK0tPlLHNVqgoh9x7I6U/R9Z08du662Rzu2ujajymXtYragi+ry9wtAVeRBopczCxDDGRj7RHGnk
a0il8BSvFC7i2qnI/UQprIgirxodXFJdtqpxQuA1SIGbjoX8MBqFR45kNEb01vz1CaV4vSqJV/49
4Cz2p9YfVqqe/pUC8TU1Y96gwIXFmgNsusZKLI+b/PwDKkKFLLt5q53bRcH52C1i5QlZj12/GE1c
rwoqNRpMxHsfjpNPwPBLC8+Ev8CSEk1mfXjvoND6HXAMdU4yB+CX/Joc+wEjNDkL/Z3v3tlJ3m87
oOMxHqnKy9FC8EC4HzJ41pMr9Jc38QLYAyKKV1qQKyBQcndHZ3Xk2MtXwjBkCRHIgIMFjICtkmWd
HM3AKECgZ9BexFELsOW8V8CTwPSZZmGTW+MlUv4rhQmX10uEJkoUzl1aj5xMlxSTNafrnB0CLOWB
drmrezTJS0DjmH2TgczNCl9Hs6xe5ZlIsx5/dPByDS7C0B5FctlK0gteIQghiWfhIkWSV1YTvXBr
4BcOvMA+QoJMIvmyE3tKzg3cMz8ssUNdaNE5FFsXPDbFdCnB6/vfSJ9B66/b9rPd/CLtd7cVg29p
/+qRxcuJHcOqJZNw+3l5klLpNL+ZShKdq3174SXHHhm3++k9S6AkChtcIbr8mV/OYhkPkUh99gat
AVyofwiMbSkpGilWo+fqKx547YeR4qP+JSf8U9y+JEesSpwIpl5uHGlgvvahjv4grUjd8/WQst5L
vZAXxrZMDE7XAz0vzyCQhJCJDopD3TRW1AKRtRw5zvqRKBmnLIAH+oiYXHNyNgWu0oAHGzqCEAPH
ZoBiuJLYWOBAD+eLTTVY2rMGpZQon5ufjEeY3MxrIma4+F9WmyDzNLLv8JKJnyGGllqWGbEUJ2Q/
eYb1EeCbJyI2ioxUngprMpyQ9my3t6CSVMydysRe7D/vfREP7ZrANW64PK6o9V5kbXXFhNhNu49V
UV2HU9TsoX9xk1HWnxzYwZwOEh/OSzU+/0M0dg0w+hewpCSLWcIM2y3NBVdGkDXwhMZNMtzvT0Dz
yLT95Zv6dbms/U+PQaSt2ziyZ7Hq47+WTYkHVhxshep4IrgQyJpQhORUtEXgsifqA6FxxZRUDS8C
QqLM5+WE/xFWQ0JELXjUzimbfHFFynkUekFdDsaqK5yfb0GYtOGlqrXcEdgfy5Akud/tO15zqoAW
VjQr1zh2bWeFQ4vZgXxS6rAZYqjangiUUF1W48D/i+ksPLJsOQ9AXWQr9OoztS/E9qaPCjLpttXy
5cQskJvCHwl5U5Oue/KGNn7DU+TcOsSizCUh+UHWvzOsAi2shSs/9CZdzdl99yEOgAhFec0WsgiX
dWHow4qW0yeZ8DvjJxNWPLdKGMp+XbkkeovTwxyqLnVtpvNWaurtiThgK5ISf/gQ+RpHSzVqaF8D
KyR2Vct+OeeKfR26E98p0Ni4a4u4A/YBgokJL3lMffKeai3QCGQ+NHDd+THeGVLhIRzljhKLjURX
2evd5omUHjnR2P6vECeHkJh7qErWBhibtlyPb2Xr+XJ/StQhvWkA5Ia400exbDw9r4S1PEjbflAa
2HM/g2KJHW4/tuTaXLyMguk7DuxA7oipxZ15TTCQqxvLTSAb05Adyc0uCV2TUiFAUqElO/VrMdAa
CyYYEhrkz8l1snt8MfTHzEsDbONM7dFCJqAdxrhfVB8BV1GQMVpzC3HSA803zGkFoMvHins8qrQX
66oZsH6kkfLjA/c6GS+j6ybVJCjBXd1xj0l/DmxlM+/dDyuwD3Q/umHT9n86t8p4edLTUifrPZmP
Smg/iSSEKsAymSeV27OLtkb5sqeXy2xMGLGrS/zsMV+cG4T2EmxSHcvWStGcIIXrc3yvltbEX/u9
l9BVh1LDLcDsbsQdSZxzy4Mr1ooLVdv+JCwXPtmt71iPgVDA460Sd9slcwo9hWDJs0k3S6mMUjXU
DJN66X0O/xNUx6SD5BDPNJIFFTsEtXB9uwwGRE/mISqWj/HnSikxWpgrBJGdfYwj0Z7jsVqi6fmx
Fzxlwu+lhHGyiBQ8kppM+jS05WmnE8zN/ocKGaZpH+BPkdKL0mkEEhNaLIr9dXS0zULJEaTaQkOh
BNaXgh7Q2cbsEziiQ0xC8uxHiTBg5uwBX91YYK6YvJJHcCvgp2j2r3qlzsDq6LoJgcnG25p1V6rD
PrCt6a3rH2T6ltmChIOhQSFxDLqpiOOYCbOtCet/sPtNwwmWTT+F8iFHdM3Tax9HR26ZYRPq2S4R
tW057rhyMYGyuwlW62EYyCcs/lAngggdB5xEwLTMWu86cyEmOeRSsdOLSEJz36yJrK5fC/RDeoZv
kqRPhGoPbGTYOccMPBoDms/VVSbHFgN4n32iDfc4LgfYBAHEiywiD0dYRdS4e+j4LbCyCVeAOp0o
Dpa6413TxIqZesc0NFJWoH1d0ybfZogUmJX0Yb0Npcnu35tLCsYTgF6oQ+cEfLPysGP0YbLKSMnf
lPxch7rBZ5yQvzfyzTOjFdV9dk+AQKZWXswwtNQ8n/po6pwqTifDO2EEReg6OcWpe7C15bm09BH2
Lp2QyiNN0AH662t05zwgjb+62JQ/tpbB7uO/oN0bPPD8Y8DuczgdzFy4yEkDBsJOg+7KbMmpYAEm
Rekxx1YLkOTUWsQOI4JUEkdyuFtm5VQNCrAPyykWJjUAqxkeom98tnY490vNaD1sA/NCpuRFJWFP
Zf7za2ukSx8NvYe1BnVV/WQOXQF1BCBRJLnwYvrQ9OO+TO66lgWUF5tKEQNBBXHdVJKyFWaVt4+t
jPVOr8lw3YTT2Q47J4/bUup7ZnItJ7/YmZndjqno8agEQGdyrAXj1xlV5DO4TC1jlssPTjwt2JxO
QWgV3RH6RG+c4kZznOFNETR4xWFanarX6zYfzw/AXkYC8TyBj0BLdXSyzu2bJZjQ72UYQzuCVdZR
RAtmTnlj2MeC5FD2AtNazRknqP4hYhSOYsbqjPsr6gMkvqfeGvyT3mIKfD7Zpn8h2e8/v/n/7Nw0
ycGfmiGev6fsNJmsGsLh8F3TbZKGnooEgP1XN449MMiW4WW0iMbBzIroAvfFHEuAfjeMK5j021i1
fRv67zDmnw5eclB9jSKzmLa2db2vI8qwY4xD57WR5WOm4skcYJk26+1l06bmZZovFwDT4gTKaNP4
rPZ2H8fLUhyRvm9UvI9FdjHo+Cjx3A1N4C/xJx6GrdiQBu8x+5keFRGq1tx1I6xDgQ+BP0gk0/q8
qUSMdvu3OwVh3qjNCqSluPqI9okyJa7Gm5ZaLjXRbD6c3ZlNwLhWHVUYa60Pq68FbydE3dJ2sEcx
CYhYzL0Qx4b0L3pZCA11hlI4UQ201ixqCxYR2WSRxUjgvOvFTZiM7FhgaNMB2yuSOXI+EWw0j75O
IceTF2JmEfv/xbW2/EeC+/7wqJL37ZNIpCLNPJcNsC2lrm1NEoDzIrU2fsCR3Z+cWH94rC4dGHN1
HsLfW7KrhoNdmtd0IVJyCxwNQJS10nhrRlafwZf8K+oxnRm8JjuHNJAoQoY7vaec/SRSUbsj4mGl
0WnbyMsbcC8KT5rr/S1vuAJXP9FjwqyufdWRmIRQst0+SDtqQxTvDz/QGxEdF8J/ksZKgs90wNCz
9Y3VBxvfbbiOMv69mWnTte4mkwbO38s/f6MIzYdE/n4WGTfhp2WqBGKF7r3aKpeqJYFI6iGtqnre
mq3w1RC+MWq4+bFv2UL1WqEC1EiPjCaBwe07CAyctmoZA9uI6ieMEk2PC9yYfBojs8bKDEEfL6fZ
EmL9sR/2SN0pV+4O95xgbQlEdHMwLPtrwCIneVJlUd3D2gtHUCIOAbgc9b82bRYSIPViR0ImD7fC
R4Kss1bqRR8YUmJhwe0SpAMtRf4FI8HbVk/zgIQlDMnXbASO8FhcqTKXAgJf/OHc+fJpOm8UybrB
gvK997rSfZp2zWxxUGMo4vQ4oCsR+xbbJ+sRMb5c4FJin4SlhvcxCsTyxzqD/0375JqpJmogvHa3
mBAbTZhhgZpKje8igxyeH5nO4oL3MxeKQz0G9Z+UuiWkzHqAJza7pVFEo9LzL7NHGfmNfgs33LdV
I5xY6R/1tAXS+RGEjbTxQzva82JA1A8Pw8GMbqR3oONTo/1Lvmdoru2GD+TpbTWBdf0vHbnKNaDm
Th6f+Fm/WUBi0xJuE3lZjVYtAng4Vx7sqewrHwQkv5iMt/OvS9KToeOCdceKcSZ7DbVqYhoeXHPZ
70ggR6QNELabeqE95UYLs4UgvJ5d+nx1KQ2F6ssFBH6h98n2ZQ0jvl3hnnYjmn3efKLWbAEwCMyN
o4RehNqSaZbVRDYzBz7ao/HRg2sR5AFrHT4GetX3TGtUjDbR7zV04SDoujWf3tcUm57gAoSp9Y1D
/M6/ZpxNZQLw0Gpsg3SlpKyTADqjpjXU65WoivfmiOu9kLw8+6hqWpNw5jxCVrpM0a6knhSRop3g
k/jYQJTdh4s8zRJ+6NewDiCGodFMETQvIFbMxSRHfFSd6y+w7rNrZgsDHFBVNjgqoQBGGcSjM+uo
JkB712Tk7DCGl2uXU4OSSJwzt9qJspvpiXoEbX2Px+fKRp/XN3TKCVUDUMACtWdj3lAQLno0854y
bKT6zyU8tQVPSLFbW3cpD+SJB5B+kKCMBwazGkWPO+K+gKye6VkaTnNj9s99fKtYdq9TBZuT8V0m
3yFst+omb6XAKnurtJUT1qj0xGCT72a/0jSaz3hc65uQRUrTljBc0ZpDpTdTWJL7siedoTnYboqh
piOh3U/PyrlpK+D6KdQUy4OcAbu88BKNVL47vGdxyiUyliyB72nnHXg3Pot23adnlK9DNpEABF9a
zZ1luB0UqFyn9mE1QHfDA4436y4ggTQ44H0fNGsVqVUFG2QeWeWoWR2VPXBwT7vtnQaVckouN/5J
9FpvNbRoE79S1uL5FoXrg/Xuj2nOVHTez7XEOl4QO8nxqJMYe/CSTB/tuLAq52iCudvbGpdD29HA
6nm7O1DQRutZ9QxH6yqw758+v8REiqdvy/DzEXnGIIdsKjuBaIXSJKVoBATF8h4lCWY1XMp2G3BI
2GIB0G0lbcaZJHzqJeVDlY2jHge71LmBLBJQTTmABOMeEKedsxP6suN3qoPxVEkFwT30+KpMzHT1
fxgijxOJbJp5MSTPWGrO054Sp3XQCSlcEMBhqWoAgFppQHALzJqU4wVF7wVJ3U0DE4b9G8Q+qDCi
wTVICEvydFJC8rno0MNL+7jYZNay8NanRTYfIAwecoaVTf7RIOop6bOBb9UXZ5v5HHeCNi9X3iby
hZM84mElh9Kv6TU/55hEHEPrPRYK8t9xry+udMGZP2Bt1W9zr/KaPlHbvepNojWthT1BpuNXwcol
9s5C8BFpVEfM3yoOfmUXpJkBJBnVMHVYEFyFoQ2T0vT9//WMk7rMhAx1/ZxKSmRYbZ9jxnlxqU8O
0cUDoWLzHMwui0vHzkv0pqFO0Tw4Fm1EhHLscETlvtw19qXVubAzqriG89V/nYvy6xCClKdKoZ4l
BYNNKw1KNUldfVV1wUD8AGzue3PtRcBd1QebwcbfrtK5cmHL3Ne4DcWirVWIMHaP/FDKMQ+k71Pg
7Y/G+rwG1biEpAwT05Dl4jfMJhROba3NOVmMt8ponAzfQcw3pHTLLpOgjRT44uZWs6aAdyvvu5Ou
vNovbYXc/9ZFsX7Qx9ft62IE2GQeh7LtR/Vj8gpCVd4V7qqoZiNMhlN6n4U6ghQbzbDoIb8EJC2f
aTxiMosMQ8ib2smp/tDenvQOOskhW1pE1eo7l+A+7A1irGrdTgovy9B9C8PLAr8ciW8Q8oFZQPHS
nZPtKQqDKw4AdACIl8NfLUFqpO6tNyz7Yuca1u5tQkdwB5YC/t42/4e1mKOdoToeiwGh3iZy+zhe
uF0q3onGwimxKyXGK7Ln7z5bF2Lx7mP8bGxGmapCSGU0auaOQY+2fZs0PjaJbhOWvGofB+95+skW
WOLdz1wDVK5TKXugK7FFxPSvrSn7HxKBaisUbxkV9wnCqLCHYrxTmbO/EUNnC2S9B94ZK0Jchoys
0KY9PUSjAxmDYWTuE92BhtAcHBgVKloiMOyU0y8rMNAiylwzcHAg7t5iLMqoQL+21th+LisvC88e
buCAmVGHlHRbiAaxD03+HNKzyuBpXO473LSHajjy0/1I+6RMpePemAKkht435W5pn5qOUW4ut9Kh
5MeW1O6SRqkwrOY+WQvNTelrlx7KynvexiavP5BDQPKWdXW+sm3wHCAON4TcLFRzKLONu1NxgL/U
sgYQpCJVY6Byh+ic/D6HnPcXPqO9p0Yk0o/9+HeUbigWQWlkKM7JokPx/hMXyUgRChiexVwUkmqq
saU1mt0kqESM0BtLxOdlU44jSFZ31y/Tgdt2VnERjP7Of5+rBT5AM3M45vDo5XDA8WoIX5NRa91G
UIM4j14PyE8yt4NifDa0tj+dlTtMmVvC8OGOXdjq2f53Y/9UncGfARETOqD9QAvNiU7Sptddcdyh
vlgguC86HPyTdkdR4QZW5Wmvxe1jUpQHgwiuJhNh90CptsI8iEUTYDNUUdWL7+OMLrsR2qbZXzyk
lZazTWscT4fifK8fEgsEAgO6P2joTbGrSVVhXOCjyaFfXsXlS/4mswE9k+lST/Ya+TbSXCxpI2GK
Q74yXsi2GZDNzu10z0hm8MCOxyQeBeglvpOvhXHNUJTEPCnpQAqktgQJ4k9XnH286GLR6/0WaMEL
jEyiaaoAqRhsGxvdAjXp9U65FsK98qF96wVzzZ1o5qwErJEUlIPKl9blB2AvVqNxMpUao7B6uW+q
h/maL0OSUUZxd2cpHwK43kQGtQfDP/YjXCRq9L0aGwolj2tNN/xCSuJX0/LC8Qb6W3Q07t5YqNCo
uY00Vkg//JjmUEBmeGDcpNOjKxUClX2Fel19quPkwNTqI2vVwSmtmmK5oLHukS5k3ynlL6+js4t0
sCtmgR+ReNQZdvZH4K65tpwWjxLfrC0b6ymCHAajqCL4El3HxHwodPomNa/ZTtE0WKAk655/SAO5
JTSlLFwq3ltk7iYyi97eRU9T/qQ1CILUfIH7scHPTilP5xLWqxjlChIG4fVyjNMgqUZ01/sVTVY/
MQ1TCQBjmjNb/Jj+J/ETOJMBCfdYkEg3gIHdVocwbgJO+Fo5vY+w7dlcktqLRwQtXzwxuizTIyQ6
9eIMzZfkP26SFhCu9Amk+Cg7QhTLOzjRLTAnyxOC9d/yVBAhbmdawYyDAe9ogV9S1K0tKyi51e/S
vBB4OzN1eiUpXIEIqTwRwk/SlNsteGa/qlVkcxpNsJRBj2WVanrqCZBEnIM1hErAPZ9zC93Gu9sF
btHq1oGtGpTZQoMLwZspSC1CjumFZfNVmow1BrB5xMphvLNnJyL9RZ2canr2oujCfr5fR9K0cLwf
5ZrAoKX5fVkWdyyNVuj3YO97UGdj535EIqEFzHcq7J8Q72SeJuv69yXdkvSy61yRYaIG7ifPXk5A
kGnzspidNRe1nVisZI3s5HBPaNgb7/8x0K5sf7duhLKTMlhmGpOoArirRa5q2iEWhJQ036iDPRx/
bNe+d+SceAzmrb6Za4K29nX1KAX9JT1I97ZFAdSUkofsrhZ2TUOOdUayBigXFnAvACyW/CauqN4x
Kk7SMpNGb3Gd2AhbvZKEdepNbK+H9gldyEBmiSJfItiHb7HwH3RDtDWzxHgAcWgbgRNTwiyLKYoX
X6GOFTDCoH1aKBO7YQxltDTCQFqvRcyoncOdX4HLWKTFhzYJtwLwqUW/3es7CGGZdvQP691ZYAc1
7XdyOpuvzloJlt49nIFOzBaTw9do2++laSlA8nYR+m9MLOi+EvQNFbXGg8wp1vJYtKXJoWNCt064
YB4VahRYy8pSYJkexGemxCIvqS48+lwlqv6+7frxDBIO8dh1wEMQkoUY5c/DRfLlLhhZmp3WqQAJ
wv5M0UvYskjaERO90q7fLck5AZhfjZikUhykbBi5VNe//pMW1MRg78vUIdFQd2tKhh/NhpzHofS0
uicLMJRh7rstbUjWSyk+Vlwk6CIwOEPLaWojGKGDdAWjiC54KqCq0GlGDdnjfqJFSoGJPj8SfS1r
8YLlfV7VZasRELBfSYulnY2Rs2ogd61hgL2tnEIeC/QI6tb0DddQuP2LJIBS4rF3fDAPkfUfTiKx
2FPUWmjnMN1LRUBJ7vUnpSqkk/nq3XuKFNnTL6LLom+lw0XcZA/cTIIn4H084zdcsrQqi6RJYv1H
vXXVr1G25L3jwUCKMAV7zDypTolNofNn0zo0EyebDtJSgLDPRVNLK3ZCXffMH975mGMyLwh9KmT1
6BizlymC5aSuLoUbdKHVy+m6MYu9bbOkCGNjCsT24udqb13J17O+c6RVbzaqOFKxVsGO0vtAaXpr
V1YyXSoZWSIcKkLNp9DJEaG6AJIWWE6F+ljsFUapbko76EnD9YmaaT9vXm1Drjqt0XMol2vY08MB
9lDbUzRlYMTo3RnmWpARPlztY25SABvHUA5uGvf/uRmqiOz1YXv55LNh+RZ9uChKln6scylQVk0V
AIPuIxPvUBJqGJSExWRt8fwdnCfIqKJsbynf5AerZEuBl9fT7MLh5YjVaLv9i4+8r/huTbJ3wzv9
4Z72syTBpzCiRWlSZ2z6QyJtX2ZCAZgLRMQs7S+NPbKSf5V7wx8+ur2W+cG/hZ9tXurNjjjKiTYD
2rS8pTCH3zC1CcjP85Q9tAxhi51r6Ia5PolBkcnpi4ugWouKv208TBy7nM7mbzXGHZE9k7x5yyJK
+XPy7KPcDgnntVX0lhypxdKMUMy2NUiIRaiGbJW5Xcj0j89hjvrTINiX8cxX7NiQVEd5bVNrL1g4
VNlqAS+9nK+JRFemQNP+LLceGN9ycQVoGo4DC5ZDYCa0pQEglranPOJIl7SnhH0WYqRCpWW+tmh8
Aa56jNHI0pWqK+apq6BlcYNu6pCPkGIRPIqjDaZs4hyHve/5+ihXRbk8Yi6H+qGgdPZ8hYogkR+Q
g4K4PPp/zgwFK8yCpizF9eY/5EGhAwVEnEJrjfLl1LoDASrlHHoNFunvy/uiuIK5JGSd0T3IrJFy
z/ksvpqo/Cl2w10ujOnFF2UHemTqRQ2Ti6UeVO1bjZfmcnITdbsERXtPeHvIzZDyW4T40WDeowFU
8WSh8bq/P8K8We6SU7S7hpBVdVPen73smLHRMv2Hv4BMsWjI3QHuO0ZnrPz6AYCkduOivwYR+hSu
GOR/s3OtpUHUKY4PikbTRRjJdrLG1XV9ooWo2tUzEhSeRHq+92qY8ojdRiwalBpZVpfU9rRtnY1+
+7JgxPQ4YMmaNpg+W+AIzdA1LogORLPzje+uUXGnjg1Nby0qt3vPswrSjeP3o3dyYrsvf4RLUYPO
9Mmsr0QL/vUm4fIpDtgt/LWaAm3sAugZv0Pq2A7ILS8o1McESFL5QLV8Cy4BDNUT/g345bVc5d1p
zmRsqAC459XJfrgdFvU7LHo69ev/nXeOVuFcW3JnEfXOfVjdBCiNpywzkP4+P8T0sjYnc5XLVoHA
OV/WBR2UkN5eYl762Ske5qad7UyVfZh5zdka1qnki9GZ2zsyuwWDpqVKnvrxxD0pvbB4diRofxp6
iCGvRpaawK6AhG7aH5s2e4DCjfIi/qChggOIueky57yStTXlrxdzupXTrzyw//KNNVSn8tXfjt2I
xHdji0iSsNopkgKeps5naWFVf3+Zvv1Shb4lXmBufgkD5RH1S4sOPi3/NL2hd0sZewXvH4A1IyU6
vRIHUyoyBatLo/f1UfdHr6BVB/15PrHavaSuZnZ9xqr00NU8uyXwHFSoKUpYgxdLIeuXbYZBv/lg
RwzJw7XSi9nZ3uRksnrDJwxh5CE7FaYjD/4UICLHeeCtOBbLenH0GA2o9bl6tDGc9RsKHJDGutn9
+yBY7t1Lik/xpy89gYo+DhHPCYpLEjgb9TBK+KHSIWVebc1ghJb47GjIhs63cLM40UMAQpxsMipW
2uvIkf3NSfo/XBDZS0skLL+T7HvFa+fH0oGEhLiKNNvDgmvtVjaUzGy63E4ILVaLjaHGapjTA6sR
2oLasscGPWKGcJ8QUW2BtdiAu7a6g2HZL2uOd4fjEgOvziTtd1PxoElahELyNphhWO5JUqUQ21dy
xD41/7FTiPTvE0XwuZYSoeFxuV3rpzx/8pMrQ1oHW4HyUVJa7ja09qWUfuUzmAKxd5YClFN/4PdP
WAFjJY+J1H712v09KPBAB0Jc00rJSI7H0zKwzSKFEFs93vYn5H4i2QRmgghy5Qz/hL8eVw6XjbpZ
/oS+5Sikifc0LK1hjJqUKeErbHN/QqOozMz/vibBh4EzgRr5u9D87/iHldEy+7f3gehC4sl2Bqvr
xYb1ltYQQfBbr3vtjb01HQlSNAR4hgiPBnVeZTc7kcCdGoeCVvvqeIf2y1siT8S0wbqOtU18qblY
cbx2uXDJHTgW3WgEmQjSwLAiXXS/+YRu00G8Ox8qHqTCkCs5zMmynrgvpQ1+Aj+jEKbDkbBYZM4V
8Cba7Sx7cH/dIRcKFt+CdldiJ3SQ5S9NlIQ+/GgNa6zeOuACQmcVnrOxJz0+mLu9G23cCxe6cba4
Wnlmn10iOk6yOC9M7BqNzOGs29wM9NQcGdaI4wk35xjylBibAC9h0YdH4hIe5ATenKUG/6vZl1ZZ
8XZIPOEBiqrOB8ReCmh+zN/qIh7Dia51L7kZqEIaAo92uLDeqzRlCuH0Q9c/KOnXm29Lpv4oOvcK
0fDQQ9D8eyhCoXSd6oBYNiTK2WspFaHYkS4i8/DB9uTYBnzp4JiniMToK+eUmn5j5oG4UsYSx432
gxceEipdPXJ5VD3QpnhGIZJiNLLDPAz0hF7NqmYSDvhaHU8I+Nsr0rW7WTfr/PCcd3rPq9vBg4zH
QYJmNT4fnXOQtO9bSmRU+yjptfNr+9nMXch+glY/RjBIGIHA1NkriibWWoNRf8H7UrqYJr42S/o5
FUNFLtu1WW8EbCRdrTWqImG9Dhry0Td5V3EtoYbW7KvIntkjrwtkpAbnIff0yUHIOWuY+4ih5IpI
3kQIxx3WaerI1UrljTy3b0fxesfcVRUblRxvb0L8PnGo0LMN0xqtbfSHs2B2juz+9ELvwAYQsWNO
oXsrXcGSJm/IdBBCYQJ87003NGaW1Es2NX3tmS8jMExR0NIQ/StO13IbBArhkSBwQRRTrhTC8vBW
1di5IlC7e45MeaqlvMMLyp5TX0aQ9OKtDw4/fKR2EAaxIyc9q6Yf7b1ZOr790ArX9MvfSsMuWQkA
HVABjPi02BpBicue+TP9BQHvRa4TJ3GvHed/UFvY9OgOV+poePn3B84khPveinK70+i0VNiFSElu
CVHhN4EJ9ExLgHIYQy2pg5NY1WdCcLt5K+BYwX2U/Vg5RvBaCi5YBSxZXUYUeexupFgqSpxBZOmb
X985wY4GsAYBLZz76LBmbSZAqwcR3FRoxwi9FWXkSKiK5xj63I1UxPm1eN6xWsEMrwZCPuMW4amb
/FWPLNkl6bm7JBqvtmDezef8XBptFlTq5l3UH3IbezPgYGek0x6EivqX12y/NA1zRewtg58/nVt/
+j2TXrXjCUl4Nzs1fJl+7pz3YFt0Te3ia6wR1NKkUki3msfD242R4wXB7jkiWMieKnDa0uzG2Pqm
+sTw5Rb0UglHqbSQFFehanwcpTqeqHk7aBC1TqwHA1Yvhtbd1YE9Lgof2oOnEP51dPK86Q/FK3pu
Y2G65hSMADa3dEEa2P6Bafz4Bsrf4tf0wQ94xMe7qOCwB9oTbjcgA2RtNcWAMZSDrXoq+G6R4U0M
ETIL8jfvAWrhd7aHcBCQTizEqtE52Nx7XoGr2W79mwSQAXoGafoQl0B28Z6DLME8HHL7jiQLsNLd
Q/X6Y1dfhHlZsGODCSmkbuPxoGsdFcTyjEmBbjghXIUXiSkTq3uTLvy9jYQeB6ADJg2UoNWpUxvG
ma12G6hVaTxUEshQ7GFIBUxDXLHmgILmemhQLb5sMnxxVMp28E+pE1g/fQ4i2O6aGWW8pAOFqNg3
IplB9zHds5daAEIjeDolwYbKn+TkxY/e6OoO6GXDX85AVBultpNhsQymnNni0EKPOtX3EdiUI6za
SfAnI6p2fc0xIqxzIAvycwXl2zk7eqEEjCZncjX6u6Z+ugU+Kh5rB0PKrQ2bNudPpqo5z0HZ/4JR
1h+sn55oMNUP+Tr8XOJPbQTQniMC560dUUuTZDbmIARUiqmsoX/69D/Fwh2siRcEr832eE9uV/fU
txAoBTaJbjv9z8csJbZ+4yZIEewmS0ror3RK0XQKoHnhPhNlRHfcFebOBp6rO0QC/2BnQo37nJJa
nk8l1WTiBN24x6YiLfhHSaYUoK6QWywzm6UGAJbKFd91DwfNO7tsT/wf1MGoi+k0rrIZ5sxbOJpx
AkCT4Qt2F69RLqJ72GXBIueiERp8k6dtOoVRRe/i3XFgNUlDyUZzAOFh90JBDeeENiVqnn5MaeFD
t9AhzYyotOf9KalY/jYUx4CKk0qb3nP2+TQg88xRciTaYXOqdpdC+xOq0UKKScy2TPKaQlrev3Mc
BdGg7Tak3EMv3gGlGThlItnOVobwjwgstVkermtnVpZe+ODYqUV/Fb8EVa2XllHFJx02nCpKQcT/
AhsSxmPdqMmZKmE0iZhfEeOOTOgqPN3QwhorNzX+4DdDFd0Lq4mZTfqaykP/XwFuSuI4SGJqJP2D
gnk0UIxXT8vamuDUlKR8n/3FNxer5FNvRNjzFbmbHcKTKGPGf8cXiSBv7FK4LhFqaWnQeb71zfFC
ICrBo85FXI6Stikk4201j8TYztZs3uD2pduPp13bO1CnbJfE71c9n7vUPe2cdGjHMZCtUSWPtcQT
DyjysIsin6AmhbyNXAOI4gnZC4BKc6idHoEvHKt9tkdN7JF1tobQ8g5T7lCqBy6Mqmesa1+M3rOp
kn6Z4bjE47dE5M0hWrLbJp8agvfviMBXjMd5URK0WmjSRNUNYa1PpX9Hrh203yqbZwktolGArK2Q
ChHBwZaBmvpm7lT2qB0YiwphpbicYq5NwgI6jdU4mi2X2dPgk63o1ZpS7MDP2TihVLlYYojIJuBF
6Sqy82Ny0ZceNTHHb4sZdQ0xKoHS1jilqKa0HBwSmfvUWotX5J6wSUD7pquOC/PX6f0spoJpglrJ
U7jpcYrk2YwBaNL54UBKmj73h4VGByniAFm+bG656ALkMAOJyzX17r8NxY1kHKRaTymy6e8i4WPe
CKrgjx0VJTQfZ040ljZJcecYaSmTCr4hlULkaxjYCjnX4X5OdEKNQrLy+xdB+2vtdhVkf3hvHW2P
wexYLRQGZ+5VMIVOLBaOAXfEDPV5wmkbXS0oK/jQPzz7K4DKMXUMA+ECoaRCYKi/qJP/Wcq0E88N
3ZQoiwp0bWkaOiAOdd2pb/qoIkHkLisqdJybJeEdOv4hbztyjYgQ7mgGO6tCUdGXiun+FrDW4eVI
o/DXkhYqGWRUTEpm/ICi52ZH+lKtITk5Qrz9U52uoDkOylrVllBQQSJ0gbNvKZpAM/y21q0Ls/fs
gf7PGzNBsQ7++tbBCm0dqjqiMQMgxNW5L3olYkBrA8JjHfjTJJ7WcslPhbay01c4XDr/mpay7gHz
aOvghSHZSV+8x8nKwmb/0AEMp/EhkdfoazPQc7SQK9oezWVXJxfmJ3qNRyUdUE879K7prNIALY0B
/eVJDv+CSdeP1XN02enBf6/Nr/y5mygsE2P6R2bYQQqHq5p4LvdObWlL/7471gA9Nj2cKfEHPiXB
DLFliWURkDwAFI+OIe4roUa4It617IDWmewH17Im199RBALwgFbsH0Jn7vxDrNqsmB7gk9g1NRUc
K48uUFQM4CU8RLP1b2ebIRdXihMFPAUhiU+qdw9sQR1RcV0WOlPWrnK234MXz+NH+40OiG5T1Ka5
RdawhHIc1c5HbswpkKD2X61RwqGq+4EHxjUHRPmo2uvZ34neVkghnvYIPc6BNg55rLN2RMeImm7P
CpBcr/BW6n/dsRBnCBB71Ssey22FxJd4hOFOgLkLf4hL3CJn+4nW4pwvgkJDGSXWsPP44chhMvEe
FAxodPYm29B3mf2qHN/TDYQpzaQF0aCS+7JHfjnNU8exJf69MQyOupbj8VdVk3e+yrz2SSD4wSGX
olp7YRHXuw6C+J9vym3nkuIQ9vUirbd9Zx3ugBGdkyRuwNGJNarSHH39VtNXb1ri8mRx8feuFZfM
dluSnn/RdRueOSjhHpMJY++1x1WPYA6rqCB6+fhH++wW2v/a0PzwF89LFyB+j22MvZKIfQUJe58V
ldNyM2xUEqplcWgeex0D3kRC0XZ8NDDdyAAzuyS5eGtfHtrjxWIAeic4FDkSM/pZpXr3gKbuL3Yu
ZsLEDI6+T/cdmZf0vQUNnB/W/S/XleSlb/QS2xOwo/6H0QIsfx2ZUiu2ukN3Ot9lOUf/DW/qhJwk
zFjvWCdwdeQYw3uDSMEdBJ3Cm3txw6cFJZJq7Z+QXsbO9SP9KOVXST5VlbysF3JYsW8xYeD7rBvE
3bZo/XPDYjydT/a5SRXhVFYLBB1Ovl8bRYlkHY7RlL/pDSRBKB0WnrYXWfeJxZ8rlRMJfNTcLh8e
4udZPvw0YpXQ8UfIx0UAFOg6ggqJjttpPvwqeZiNUijMwJdf6DFD0m++AB1+jg/rMdFNS1pVd4XG
6pkBcVvRiSY0CXkBINoOE7rZAw1H7UUkIkIZFwsmgXFwnbvkn5B2gBI6cBewYqYKjWCQmEc765Bs
I8+h5P4dPwQOF84jOH3LIwO8R4Sux1y2Pj5uUSXoVO097W3PfC814prrbAPgIMlcTeuwUdKz8Pk/
YOkHLpEg1rOIqboTBMpo0V7+FHC15Y8S9ZCrdZO8wxbuH4ipDCiWUgN/bt335wNNRm3k4wtZ0ksJ
56HuTgxtow84d39Pp+vgPrjmfdbWymAb3BVRaP7h6cAWtgaQVUE9ox1ibwzFMWEbLUE2EkK7+KR3
O4wX0BS+fke0TVTWqDQ8JK3fe0bPTcyzbMd6bSZyVPG8NngP/fMtaH4/ZxSdjApDmr12ws5K8wEs
LTwVbK3+bEEuOM/PV9MQBxO5xDj+Rjhq7LiS5N0nzfFU0pufVu393JQ7J7AWToC/x8oTio8x+RiC
5i7s0ndrBQoRYspceMPxdWzTZfU10ZdoeC1HuUTkZnOstz9/+A7Le7BXhWFfbJmzt98rokfCCxmX
a1d/bMZTUr63XB/uWtwx2m2SzCnQT6CQcqSUOVt3GRpy2flNhgL+KlFEvPZ3leqzwv6ZqpNwKQs9
1blvrBc4qN/Br+s4eQ3Ix/HhcCYewQLfWiraFQRKe6bT1S7svVfEjBAj7uJA5WeX7a/TcNRydsNq
zXK93k8Mq/W9aVo0edfPKAzPZHZilzOMx9ls9ZC3EZiuDMgFhCYxBXI0dGS7KtuJjzMrBg+eSuiu
eob8+jI/bP3coj3JIPb8ZdFJfYRZ+dkrm38Kz8TPetQcuKzBmKHhP3C0hleCwHr07c0tCdtVb2wi
YHw2QNE/4YJS510gs5qWN/ZBbzs/nrEez/v5G/765MJId04idwq5v4CxQg7XG9gCQ6LLfqVItGl0
85IcHK6ffTURoBqeX2xhm0WuWuZgiOgw+B5JyredWzKCp+9/tZJVHrK1XWaD7FX2UXUn+adrK6/6
Dtd8nYpPyeFlAdYDGr7nBg0isalv0Qu1+85enVI108Q/s9ng0JnkJs8FgkgKQ2NkWSz6k4MF8ILj
+Xry566lYEIaTwN5KAKdjTlMTaqoIakpsxT55vFDTbutItPZR+gq5v38Fax1NSjdNRNexWi9FFzY
MCNzIiNnx0+aEV6vpD6GysgvjdIOWSjon8P3Ngt2BrCzXkboH6JrjKhMJ1B/ayJ82y1wKcKwCwu4
ZOvbJjZD52Buh/BCgSS2O4uQDWEeTDt8QjL3vbbkcGLExeOnzSbzMGRU4WakM38Gnw8rXuObSXtK
xhQtV2eDXBUk33iQTEaNDw8wlRWpEsQF12MH65BqKog1HAOKsas1kqHYRbq1B0TdEAabptcrVcnK
4QIfV3bXrsx4BEanIITo3GorZyTTpQsQc2xoAPg5nCqqJicgWIeEEYxekYG1Ni2g/EiR9/Eg+WfA
1svb0d5Wt2zrnBnQZcU3ZICHkVFnkWHigK6tIfuFfq9vU7TGkHo+XBg9Cf3iMna1jNgPb08ft6K5
id4PJOEEqAScMWRMhweNKer0I70FR9hB9j+D54KjPlcbbtqP69JeJlyjbPoHlmr+Xs+hlMhIumzM
MqRRQCxTBPl7fy+pnEUCt2D1kGZSWacoD0muSjU8rHDCDOHRuTm1DlgggFfeDoFrkpPtAFBLR+Un
d/X9xamXhkJGdmg17HqZ7zEoosYtY8xH+8QBUuKQIx5l5Fjjxr3rFEJVFBONrSfkYDij4QwdJhzQ
EpoBALpdSPjuzoH+3+zT4Pmhdz0fvnNhqYfM1Tvyoyv+ntfTfIdunX5a58omq5KA3MsvumyQltL1
R6cP89ralC19HX6Anw6edd9Q9pFk4Rotetlz8NVPUYMnqnxhQJsa+YjOtDVvOZnTE0N19hTrML+E
Ygwx16EpZ8Iwn4E2JuNkE2aijVBqL+4WxKTFJW3J/d3yjK3jjGMla1W7TcbTHyaAaY3pEDbvn2SK
DU8kxAKG2UZOnlQu/8B2v/M+FqAZ6Eih82wTuu2fwE4lczv9vtVjGHUHsQue1SU3ogrC0mZBK3R1
pnAZw0ZBNQs8XMEggLSNUfztocgsBi+4oGi++eNfNvLE1+895Aae7Dcm3cEPU9a8Jc4N+rC0g1w6
fi4ecOJ4Zp17vwNifFCcsJHJN3Wf7L6SOqJNLgiDGPginDAIJOV1MpYOq9/bf/TqtjQAptZjRZ7K
45FMGSpy68JGMqEdEoxKlfvA8vftQnAnz42HrQuRzuvka+/+KM+XR6WEzT45hK2U7NrmBB9ywMU3
60M60yGdNwAFhO+mTg/TWMwgGvz2cFxU2omR+3nWtqzwafasC9vcw89M1VdhuWCaIEGw05kfahmM
2n4ie27C3YHN5Fbn8O6Qt/kR0EVEhZ2iQ7pwgqb4syL6840G+LHvtVrvhqOoe2tEfSVP9nIegR3s
+UN14Dj0NMwNYbOdnWFBYi5zQNNcwT/14Ebz2HUxu2PBLaZMt7uLF7AbpaBs6ejgSHeICBU5eqVc
pOydpcWdRnpty7/q8WMSpzLM61tvNv6F0jMdL1R7erHhrONb2MGXM72MoJvVHhJ85sbbqFHtFXxF
ZCKy5AeUThmCOvgj5I7crk6Y7mr4qiqCqImut+l7FZ2Lyz4EgqIwhEgNkK6BaIcefSTcBcV9ULP7
i9Hp/oly9aeX0Zpy0UupI80Cg85pFVqH7+twP/4EgTXvDUDHzHyJQc/TuN1dHFkW1khk4no9wE07
8Frrghzqp1bBRrTZV3jzpJ44TX+s07pu/WT5jmZVZRfKKnlrRgOe9gQVedicqYCs2ls5wHwA0sJq
MgdQEk880Jn+hw3oVAmQg+MBF+VKKAfWhzhevr0EAdQ002BoRKlI/Z1AHLEul+4nMII3zzokoPCc
GY9l6MI8msBpCktJExy1+ubFkGbZa93+F+5uyyA+c3DyQ3/kqzyL5BQlEeiwZ7HkH2Vrq1ITwwvw
h5EIFnQdWavQYwrs8pwq2iDuwQigVQmWyoulTP5ShBVlpcMMOlgmgGkkWpOPi9dyzJXzqOAEVRfw
rSjzPbvbKN0Aq6j4Niu0QNzVNV0RuGgQtgUOuBSufsGWg+gixi8jbsPuPxMz+mCcWxzz6Ig8UqZb
2PlXyB14LMu0Xv1sfpRTKUiRhxtY2cLJebzMYjl/bFVlG+g3+SDCloPpkc82WsHClwe6ueOz3GAQ
8+O1xB7yRbJNepk27+Nl04QAaM7h30pgACt6DJ9qbKSTRrAx5WHPuF8b02HEutRcpniDJg3Ubos9
fbLbCtvE1ZEJGQ3Wm6lL0qSyNnOt8Te1KJZmqLFQMnGDYYYuOOTOpjgFAfAQHdznMrMErRqmTlEc
cW53JC2c/znD2X7kRre9jOVP+MelE+9o8WZzQNtu33nIVXe74+8b+YF1TX5Wt6+w2H+fzkVTHmLc
yw+wX0w3HZJiYA1CHtvl8/FNcnT1RkIDLRFKKi5HeC0hC65k7HLGi7pXEmGjWozSG+pfFyKTtn4+
tMc22YoDyaOg4GJZ20IxstT8L3OGT5AgClVCLiaINTIjBvZtOCEU6CqXVp3NYdFRmz+I845xQXoU
Qp95Ju1bGUutTo4Rr8fFCwJ39kMnkG9jKgM3nw4fAKv+NxFqwG53xrRnnx6gWSALkQMFyKtBnaQy
+G1xV/Xm4FtpbHi9rD618KCCk4w7M0PW6vMKdplBg6n5+7psDgi2J7RfUma3hk48Wo9LO++rUHUl
ge/0NTC59OwdtPLUAkIQDFu0hyH3eiUp+uRLm5sZUGN3xs3xRBzOJ/k3Zyb7i0Ibxm08in0n/T9I
RUPmFjHR3VuQrw0uMIiUuY6Mmx/ca7Ib4DmY/DNO/ieD4duuBcn/Pf4YykxvX7MB6IPCsevrf/xn
cdfkAnkUR5fa9NK7MHx/Ljs7O2lLaa8W8C6tyah5laKNbtdq4yX+b14ZHGIg2ZFU8tSugBo3GAkb
WRiaeR285SXR4aoGsV1YRzObJ9kSLfzq+99K96fb+rIiGImWr7t3EGdoG9ilVwDBYTHT5H2afzER
umtvaLvc7bysyY70b/0bRwwSX+BtdAVX2Y5EIC/Ny4u50H3P8cfoMs3bo92hYv/TGhC7jRDQ3WAA
rH2fLVBN8Jn48rpkays0Q7HKFC6JcqL7jCZvL6Hq1ucx9olMim83dkJATDxpp0guF6iAQVNwMDj3
wvtKHK1PfEKaDdxEz+Yp53HeJRu7G9IkjJl46irEpI3ahx1tdOtLJF8h2VTLXi9m05lDjHp0wP5N
31PEwsBGxUubfhJSsKRwLyZaiUW4GtFdERphcPy9gEKJtaUq3EZjI19Ct80Hn8yWzuPbMfwGkqg/
jrYdp6OX2qo0QuXRz7ofDRQTYbHfdMuIu2Se+YaSF8WV0VJzvd5i8FrOCoiyXRSsRI2bZfhvmnuZ
lnZ9AeUKDF2WjtIIeBUX2N8WZDhJCNTQEJ2ds6p4xCSCXfYaayoNwJ+i8/Mody8kKBBC18zq27bO
KgC+aVciHJFAIzCbxyzrDESBcwaosSUJIrLpFNtsvPgdBHupi5arA2htBCHjcmY5iJUkUgU7nSwC
RTSHQRJlhrMaG7modHoeFCUELAD1q7U2Ddqe7JC8kx4xhBX0YUXIY+N6d7vfzP8/P1S6APlfRaoE
VJ3wV5r4pHPYUpH326g/vWA8E8z3I0bMmyGk742zDYZ2BDuGoSvax7Z92vho1p74zZx5Z9BOBK1Y
u5D/ieYTAMILP4M61bVcruz0l3eRn3KJmjl5Ywe4S4MlNJ+ZFmuSjxQymHrm0LVH0O4wwE5ZVMe7
yv+DrIRtaoE58WCwDBHXZN0x6WA0ecm5aVi87XAPwv3+BnDbXKGzEaywKpH6LFAo304KVlTiiG2l
CZQSoPlSMtuOipKTSHuIqq6gDtWCTRgdSPJcKdfgy11i+Q3P/cNTs/7iEL/sp6yQieoE8hqtOInx
QTMDQ4YtOAV6AtKnczqK+tni1MH4K78/vhj7cpdt+wQ48EEt9wJ7feG929E5/WYEaNqQ4HJDTDz/
7E8V+A7vyeXgPXzYEMqWGraVbfc1KngVpFWrM2M7Gz7S7WscG6jK7tdq4B/1breM7bRlB9ShVQBD
uj3E/uWoHVu0o0iX7raVMwZW8WafK8KKDNIN/XAZit7M9J6dnjqdBMJsngTdfNCvhvhjeTlqbvDS
gltaMIeeK7ZWMNvqFpiDSn4fANGlnxaBs2Z9qnLKxsvlDUBxptNA7ZmlBNqJ/B93rKhVa6El6UTC
157Ym7aqOCMpvcY3rIDYcpvZUlPZs9GIcaYPFoQCV0nm4gDGX4PVcky02ZtqdyqrgL93EDkfHo3u
4K72OOFPiS3VrC9ln4WZ2Vy4Oc/uIrWCJA02b6bhT109vlJDsPu9c5F8EMXe6dCzK3reWFsl2eiE
7nM1tiyJKX3/HesteEErfccw7fDnl1MrSAXbMNf9ytv7vCpkqpbJjOvmKZQuZZlHzYIQI8tRR9nu
Mx3F3yh3iEUIbyQXiKNi+xTCNAWAH3QFqdJBZ9WX/FkMT/P7VYlnWxoJ8lsK8HSBIjHq8Hdu8F9A
LzBkBRkKRH4doiz6+7by123XfEHAEk+qlwkQO2woiuj9YQtWvm2jf0PI80UYvRMzyE6VpxtRltVq
uWbOiZAvIrIX7heg4UVu5q24ydiPC9hbJlumIn03/ECab/M5mxT1GCkSFEoXDhuGM6N6j9q026P3
c0zyfnQSTm08tBXbZSs05cT06shWY4XRXH52ERWYNBdaiVvu4ZbAYwM7d+CfXqXkHtdZj41KYarB
tyC0Z6mPiuQ29qfQj6iY+uN487b/x2g4SC+zwu9ROs5T+FIc+Ftw7ncGCz0oc+2NhtiDT/y8MtVD
wengfuP0XroL499cFaufU6Q1tb4waISAh9SR1LkbH4BGZx9FR9LfDi0rTis7kfYdIPH2kd7+JR8R
ip2qZmG2YT7VPv2KvoYdx49yP7NoWO/w/ZbUsfRWIIPL4SbXMjgIang7ZPDEacR9Z3gYwRiEozde
uodV8/rz8+xvgkU2bDAyaqLT8QUoKenKONHsBitGU4O3Z1faWiOF5xOic+XukgbXCZSSugoE2oGM
cJwDr4qSnaFvnKTeS4WWO3bB/63VBSU8pQFb5MFMHaOKyOq/mVtZHi0iVG+A4CiyD+FVSVHaLGzI
u7TeRXM26rqRhr8cYV43YtdmzyuNdH3H88jInkQwWRKiJaERHUizk3ziE2yh63+zLN27CE1kjseo
ix+26D3pIOZApq0Pfd8zwx8+jRfsQoLGJ+bLp5jgUNkHfSggwfQM7eu1V2lzNlVsHKN150AdPbMB
03oa0Us0QAMey3YqwqzYhsp4i8aE2UbisitFjy0jfXwbxczRMdzsJuA/raMZMq+Ps/5Xp5+IoBsF
xMtKmlP5A57Al472sKmRasB5ysCsiwJAEs/vehkx+Np5RL8ymYsaHnClgcnU73I7yUKXua4cBjPe
TeXxq77qmcldRXjGGsaZaKFvebfsFJ7KVgdiRoQCEq8D6goxz8vAIShfiMz2fVc0bsXjuc+OCuKZ
NmY45bnZTRHzeSIieipnc4YrLDbdF1ZFx2zuF0SjtX/Bb47RazD0nCt9ecyctKqSN6jttPcU766K
gBZJ3i/bdsFcLxdSkIf6RpVKvMAj3Er4iFz3kod0QPC5ebL8AykxYkiJVE842afvphMIE1zLOsJN
BJGY6QcJJaVZSXM9eq6FtVHxEtCoGmrx2kNK1iU/Fw0neHP84T6/OCD5gWP9MHh1EMdXwrknybRP
uYddDw2d9vRgrCYfqA/XEyutMd5Zs1VX1dMiffTjAQ5l3ASteYNGUGgiQa/qz1rqP7mT+3flGV0R
48ICC9MdK8oRzhrBpsoeFG+fHTmrb0depGnDbVOaW3pOaT1kz1gtyTfoqP6uMrYlza2lDe3lynB1
7mAR0Erocw6fs6VCTkGiL71L/rMv8klg4uzwNGRBMkTVx7hEwBY8lkxfCBgsdWl4Ob27i0beVhM/
IvIvxf2tTIXB4LG67LnmpYp0OaCrrKf4r9p38yBBsaK+v71GI0lrcsJGi5TqDUeQbdl7s+h28Nt/
267o7jdg9awFk1Iok8BDP+0aJ7To5WgB4N0bNtHahgRCjIOPalzSVZEHVwa9wkGgJEt5kxcZMY8H
vwX8ObrZIwKjAmoveKoF8+p6IIbIf4lUf9VRUXU8WIjyEh9W4Z29GHTxOLcuJP2rK4Lb3LVV6tx1
7Wv1o+Ob3yCnTHCmnHPgnQX0qaV5fWF3nCYnLoBhoDajIqAshX5OS6ungCHIfXNOBJ6uyz14k0PR
fz3jCb8qQji3dYe/qny5Tn2IPxWH4R2X2P+jGeXoRKZEFjyZKeituNvyDJ4t1U4nJBrAzr5x4cVe
fjELTCk3y7Jx3XDye3FD8eYniQSdcM8gZDaYDb7H0/AwslKyFwVDCIHY7mIN/Y7FY6aobmv4m7sv
NAOPjfDhgfvaTIZjlG71uPhTkqjrXkRtsZPI9voerxWKuiuI9mC+n5jOyxW5Lk1lAfyzqNvh0JUj
npxvOc5ubDS0Gt/NT/W5zMTJRoDGQX/HFa+eK0PbG7otQl0QvDCqyE2ul3DYHFJpuUy7w2iD4p1J
MSBG7+LLGUVzs8iAJqrMxvcUgOVt7YDo7s+xvOh8wRiOm5zqjgKlDOGh6eDOdzSnXgNjSYLYqL2l
KCig3OW9dR+aRBA5Ud46fmLNSBxg7u8p2nRCFIBXzgrcjcPwH2lVbhSh3LXAq2BPp0lVXLQ8GWq6
j5KTCVjAueE7vvc2K/AhcJbZaRy86B5l4oR/RE3A83yVYLuLyZakmWrzmPTm1VmIWBbiRv5VjjeV
y8bJ9sP8xOiXbUIQDRUFLFxdA6/GPX+ymyW25Tugzn0s6H4KBuiOjYz8P+etXEZT5Hix+/zaS0qA
Pz3tT150fjd0ZskHEBk0x/CuyM175eVG+yQST9ri475FUkivsUTrOpPCSp43G5LU+sOS94kvdqng
d4oz9iU26OSXmTrQ9cda2NErywg/gT9lJI9GNYL2iJLcm/upuTlmmmiaBPDTZ/kLcIiTf6dklCkP
4tFYo5hKMnfmBQwA2RfgpZ+tcGEHmCb7IkW1d/Tj/nOWjKmnJxl28fdut17+fosZj+IpiNdmR2Fs
2fPXzjDW3Hv260GQO/IqHeXAnjHsxY2y01OxRjyMapgsGVonnep2Ri5a0SBoJy5lx90NObKiHSoe
Yo0T34D4L5cuIleUIuUCWgtsYfOGvtA2YShutreNRp5WBlVXSc4l8oLCQJs+HYERujonSTE4yPTo
RlVcU90NXJ5jUEJfS04EM+0IbwNoOQra4BNX241Wqg4m5avD5cOAKmdO5djLo9HId7WY2OlvNo1q
3TsuczwTjouHJEIPrpS5fivOtH9kslWL1qhAkeTwDJFFqiYyVzPIWYNzZjgc1vHot0JWT/iVtqDD
dyrhUoWkxZ3niR25nRMKIzfNTyYiUFrhqLdZHYwQ+MQ+8NimfVgxmeR3xh3U5G+4VK98D3x6yEQ6
qf+9LvRLCua3DUfktKCkZGJ6AM/LMZ9N/1PgSNK+OJAJ4bRuiGtcYoMTfVCiXzqcGgrSPXDFyXAp
NArVeAxGme5mnfOtNXkRRJn/78eDXGbVkTiIjBj6l9ubH5dAOGtgjsUM03NqMjkvapucxLdAs/W9
UOVtuRJNcH/y0mrvte5T5MvN2KCBnUk3quX587cNbk5KWYs/tHzKajWIn0qSnWFlw+Zvio7NFc1z
acn5yuYK3bnjTWsj5/B639v6d9Ui1IoxWXC96OtjEEofhdylIydTdeBxUlTuf5yQt82iRtVLFmZ7
9WHhMXlNeAcG/jkpNubZgwR1UylP31mVE0JpcgPN2Pydtyp9BpyvdiuAKYDt4qE4da5sY+33Ov+4
blndC8alsmEq6fmOcQ6wRp7Q8dl5s4wn3pdTmgOdZcFcaMfRrKrpbZDKvT4IFV8LOqpia8G+ozmN
Rs/V++If3cIuT5HzEyJixySheu3Wg42md5xXN5SWqXXwYKq9T8PgCi2cjBkQs8jFT1RC32PgQbZd
LD7SiN3b5immMb9BCO3N4lJ79Kr/i86XuDxtD8jnVE1LjoKKzqbz2Xdw1K3kgEdf4D9GMU6RlJYc
CcgBqX7+LkcVAxyr0DA3U2c+Cfc0nMV5GTulmNMnkyHcDqbR+zoIcYtGnPS8ErzaftSvqmL0p9Gk
hzyeGEwyLlQ+jlHQ6/LjLAt2FP7zUr9Iq0ARMBCyQ4waqX0ot8H0Dni3oqubvT9JSQZihpAOTyWz
6Xb1T3wtiy/r+4WwrRUSh78b77MfqgDKkQLX/0G3TyQ68zQbM032PxRMr8Jh0imXfF9BdU0Tylay
TX86+g/Fu3lMmO3NTllB/bKnOqNShAcoylFu5dnndHvtTrLIdFJQOdp+4YhmZ1/M9mY0HZIAicDY
WA0jq2DLKjxTC5uRzBHMdtWXpyDetYMiTlngWBmRXKLMfJ/KnvgmOOP0qr57gAUoaL8YG3tQoeaO
MWdHwB/S2sl5yiRkLKiYbL61+hNeRBJlWETx55I5ESuUxWuXW8FroGXf61mnoJcfKX7GHgdyr3rA
tksXca704jHKeY9YZfN9bl9IKLYJ+rlN2v6rrUspfoyKFb79ZBnoSrmHbe86hE3epu5dEFztL837
B4rwVTMW90H81KdeJ5RixYPh2t+2UZN6ob0qcPZ/Ct6UA8cMlMo2jExFL1pONaTMVHuZfZXAXNTq
xmQAPS7vsip+0erCN6GVS4fpkai6jN/EI5BlaETaz5i2AladkTqIBFgGz0FJhghxRWgCrf7I8zlV
DfXO+BB2Mpv16SXH6FYTjIvjP5ocochR/MC/bng7buZJnyfiLeLlOMR/sCw6RjHESZ4LvIjcQPRt
5eZXqnZajAwQThCq4pKIe7G5uhC62PiqF+Ygl8cpknk5pYRq1N7WG7yo5K3NtAQCCXm0Ec2pHQ3d
adE6n+nap4uz0U9TH7okAsNwNYAIHBxSR4OjsMN6N/vy8UmVIUzANkHNJ/M9wJwfDFhPKLVZAeGs
so+TGQxRf0wSNah7xL1T20Mnqw1qymsRp+JyUDWBq2duYM52rJ57lLR11lOa3eF4ZikIV7ZpwwO+
y6GmSv/r/7pg2pXafVXS7jfAOuonSB1rim5X4BSysvne1wiaGsvpgygbkbdsSAD6W9NMFlofezgy
O5ucPFpR5CRGzCXuxFxCkqn/yfgncYrnR3samc/YYeHD6EjLPpAWGh3zXPLMEnZDkLuxZOep3FcK
Gf8wXkBssGXyxXS30OOFeJ8f26v3aB1+o4Hywadg6zvt8Ki4UV1UDtL4oEolf3FY/iisSB3Gha7S
+0L2EvdAsF8CMyaNaL0e9xPwghLBltfweOlAHbmV39zc+2pdGAfqTRPeLHq3PWhnndtE9N+zjCkU
RkhPdWNZZ4F3ZpY/LKBJYJRcD14FPxuzVp/oRnRtrz699PWHQwHipLRZiKNkQriJUo2cVfI1hxCb
r9Ia3H8X8hWiB6H4vNOE8MqyJ0kCAozlRGzgaWbzWxtWoEwpcEBUhvcGlI2GwuYdAAAn+EK7KELK
KBogmAwRO/PVGr1fCF6BZuTZq1HZV9ygXknnIzhm4tLMDjjF7wuDMwGC8MKKmBOVuIAkzi/TmTcj
L6dnXGHA/nzZ50svWjNBxiUWeLh17a2aMB3dLwzzpqRSPHldOVf9H64QphpnDDaKExBtS5/nmp4q
Jb6R7WSuPrBTBakfLKPmLIwGAVEbhMniuuwVW17/MW5NJxAY7hn/VZWtewHVhkP1JUGwk3mTzgd6
TKphWxK0Inqo3z5WkTWVBpedTFqgS6EziK3XI34zUru3XlgWwokjS/e7UHy+MFpybRSTUb2eS223
CvsEmuK9/fDWm2VaG8htKsTS6e33r8WM7E8paeVzMrMqc1HlTv8L0nQgadB3sexCv2aOfbazl0TY
bAmxxEAAPFVqI6nxufyj8vxmbFD+GbIvkvjonl91WGO5CQ0Pb5kjF+pyv0Oqtd4/sXil4UJva825
iuAtRjv9voc5WMgrn6nsLvN37FRFKVZumYzoyrbVwP6m5YaB8JhBvUtnukpAD84UDQIR4RAFmOp7
Kjyo9fTQX1z4BOr+8AcDT1kZWQRBmPJ1psZcC/p9N1ZGdY7l9l37qFwb2cizzHe/f/DB9YdxciCY
O95c6AObViFlXgex05jBz65xDdKqJiBEiu7Ui7anhX2Dy3PrwJ4LCYzL8zXiFXs4FnDmhZZ8MIb5
/ADrPycEsZ9vgJNOKabvbAdAUOB0fBv2SqWdth81OE8Gw5/QfbtgD9NXlqzHsCBXIyG0orfft8UK
Ze1dPK53RgBC644l8n2Vr48C6DWGXXqKPlmKHXOoAxIckdp362x3ISw3Es+M4+Or38JI1TEokUB4
RQlDLMwBgA6v4w7EpaPvLElCqbyT4Fl7Qp5o1MFy4rY5WyFJ7wMU86vHpz9MyX+sWSkd3xsL5dnU
rEkzi9kV/g9XkK7EM4MsYY9TFsvyrnnUVj5fBLGohZXAMmOi8xonJHbm3YYzjTrbBNB4cWAFkRqS
pyGlmbajj5+iuoznC+bwFBRcks5y/twkEK57frYoJYk6A9NSjIg7bAxC0OxS1mF9Ftg5yuIvbFmk
jZafddboFybdfuxzELyLj9F4AOMdgeCTsjIjsmbcdwmwx5nhb1OQze4NzvuQXyHTa1JrmOZIlNB8
IDagAGBtT+zAlDmy7qvOZdmIWpbgNajKfwv2XusXqyKEfTE2ha45ADdd5x/LNSQcwPehgW/qGDqC
fJYqa0FY4UwfR+V1xfGlopPEXpikr/EtfADEeNT0H7DUkSzLEAvnTbD5KlrHt06FniiCLPfXfXUB
r0zuylVCICkEul4h62163MfUU78VNcDaZf3FqzlpwmAB5VQCb3b7a8Dt9e47O7jZcnsCXmXh6Wuo
yjPwJpA2WW5ONKECCPYkI6J9RQFOJ0GhIUvrbmjYsflxryPwnMaYrAV/47eCZHOe+5AjihEduEgE
ufjWZsL5ouiD+j0XbuhKN+r4p4WNhUUwen6JQU7NAgtI/wPIaEassiPb0ZQAGmWhxPkuy7Q7z3qm
I3IBZjKQ9ig0vT4flE83yxqvW2+t/SXyOJtVjQ9prXTa/Bvq9ZLOCRswMtBCLKmfqsPx3zjWKDn0
h2+E3qW/Tk92qjLLwrV2scka8BIsiAp035lVVYoDEZ/8krVj9anlXuzO3Y7/rm2uBbwdq5+v0DXg
sLZjlJh9ey7FKQfMmgCrPMXsjU+7+hZjjs7sWSVKLyx0+7I2ZIiaxcQqS9YEhAwwCgvsu9DN0njT
vWaw07Wqie5crAkJ0lvxLOBDDE7rav8Zl6in6lnDpTy6kF6dIvMprDhMBS05n/6YfL5wKXDjrsws
6COzLhVrzTz4hU9jQExqXXROmwLiy2wZy+mDFss5atdJ3A5kKOUt5aczrcAWTaqmgwQ53OqrBbXu
ZdSWl2l9DDGitlA8cq1iU8op+yqqFsax/WyPqDC77WO3Qqa5SCv0SkeKnj1g2PwZEuT3EEU0QCts
EneuSFqsVoEZhMCHCqq7mpr/JEvowGecPcBmym6fNo4ZODf28U6/GbxjT74R5/YkJhs73NPrKhqa
2gRnr1/3JMiGIucghFw7GivkQ/CtaQP1BRny9qfE9+Nzr90a2ijreDyqUQv2rV2G9T6/TSbKsOxz
Fij+ZU046UpY1NRPn11gPUV3+7D1/AatIMuf31ZpB7RG6gapcu1xQcIvwryD+yEM1IWUfsm+Rh0V
CyVNySc9doWbQ8xAMV3aTHjfrWDbI+owKFxSrxQSqHGnhqGOoIKBR9qLVoeW1vJ97LcW6K19q7vQ
Lb/tgXV18YbepgIbK7LodEMdBwQBmRza1NBXRCu9dqz1SJeJp2ZUFWxZk4mT7/NO/gsATaLYbf5E
relWJyI4IqiMgRx+xDW2CM1TY7ykX9IvrEevERMNuxjcto8v1brl/h87H05NV3un2aHj58zBYJ83
9rJ383aqZl2DBW8Yc7vWbcu8qBq0fpvS8lDq6zawcsqiKOhEEplD2F9d0nhx+ecBAX3u8VhS4iND
OJk8Xk17q06acRDw7UlIgwbOKQFzP82F8CDteaMahiaCvK/HRN1W4g2dUffZSuxcP9Qk9IOTazm6
NaPs3wsAo8Bvx9dcDdHQlWU+1/iDI454KMs6zQ6VK4cj+VbiLSFq2EuXTvJcyaw/Z2r4cQ0rQgZc
MmpdEcSAYvUwWm105mselPeEOUh6kxDchTxqN2TG1vdXfGgrTOO9JFfQAdIk3eiRXmHbuCq1yoS8
U9mc38+pJDipWBCiwjvHbDCkIpQb7QcCVbZnbpllkM4MwlsXcDJ1sEd+6ZBEsylIy9ZBTOJCEiyL
zW3KWWHqgPJsaP5NL8AcpynxbfsNefaDgHGN3OzRO/YIWS8o0VLxLVM9n/qlTXxxxVaPa6tuAw3N
eKHuf4Qv6NyRMANgunjYZEL8fd9CT9Cw06OXr0UGOfQBta+TjylJPb4z5nhV8Q0vIUCXptyfAROP
ckP3nVK8gB8Tzij0LIJgmu9c3ktvZHBxNJ8dYjwaKj73Jjr59pu9hMWTMPxmRzgI1ZJD++WbYYVP
L9E84oUgNnxVsXaGRlExVSXP8cVAOfllazbZGQal28WNbc1muWrAO8lfDWJL5KSsW37C3p/hAfWv
6ZTcHtXqNN5iJy5fn8DXfi3h/3VyCYwZpZ6jC+/dXZnXcyxLZQkjDmH+8cO8pvPv6zafJL3kVnR9
HjAoTQQwDh9386ylhhf70NQkEuQ28U7idh84gD5qJVEdb37C38r/w+YOv3zM/3XdXHhpK45rhOiW
q620VYKYlOUbVy0ocCdm5Td9NpPu65QHqopVCTBANtINi38jdbTAlFRTHQ7cAwOg/NbbjfTcH8zT
Qej2lzvDaiIsxe6wwR1GjPikOcPM9Dx9Ozh8oodW2Cir71AYmtQR/Uq+FQNdenarDyQ994xTZA4c
9assTkfaoguo3dAyCF4V44CIzpL+aZF6Q03r+MY/a/lFF+gkEQBbro9W/lMMg7m7+Nx8R3ZmKrtX
UZo2aRDhRhJuYSiS4SmrXPqz25B91wTaz9S29CVuTgoPGB09icSNprXhshB1lGK6LgR6KGBzjMrG
WG5fKRSN8sBOjLmrIS6CsiFKe5Z3icpad7j+6PRFSppDKYliQCMVT86BzPqD7P42QThZQNTXbHT7
eWihkDcvz2LPimbxvTxdb+yLfEnqn3T6J+9u3cuiq/0Myt+99+AgLprvHY+9oBT78lVwaCmwNuXQ
JT3a8yCw3vKWVJkaXlmcbmb49u36rIH2f7GCsVa+LKIrVmXGgGhnqLPjJXiygoV4hUcspW0jpIHR
PnI4kQPSiZPFcPYVcW2ILthwiAsap24bZ0+ecQLVJs78fNzK+m/SiGOBhqT/KlvtMO/nHFgHc7sp
dXENDrOgS3o0o/IZtM9ogW/Wls/8tVF4/7lo/GjCwg4UrIKLfYdUCoHF/QFdj936ThHNRx5gmV1a
wx9YSDOjT7yizpAFqn9mkPmoIta8q2iEsh9WRiWF0R3jMAosu6y+fDgk+JXjjtLlZUNNQtjzSSIV
FL7wykdLKO0ocOH2N8nmC4oiRLei+WVQZ+eW+L5QW5BkFCIhUHM9SQiPO26GjmugysKmGdsyK4Bd
R3CCdlbX1xX9EEcDQxPMvQG6roTEHPyVAJScVs44V4nAkNomWkG5DlQieLHAisXUJILe3dP4dmRr
/CGqap/LuWs3dgTUw2scrFCSVmvAdZt4sKZM5WA80IdsALdgwhyolNyuJptQ8XWviukowXkTB9W0
l5ereZ8Z9qF0+pPfSidxUfasnjRK8k+Je3NqF19hDSMUr4HjXSmZCfoiS+gWe8BpaGKLD4CwaPmH
oju+iMfSNmAOuaPuGVFbxlgDmLDTbIC7WGpAtK7KATXA9F8tzLbSKs/CC3j8qbcoXp9/c0rkhkTz
F7P13pl08yxwEtd+DOwpJ/zCvgFCedNFxAPw8Jpr2zthCNoshvSPHpdEYRKJ3+HD6YjttDY2vE/k
q3u/1rQtSki5FbtXrF+lPs2bhnF+4kakB9RWlZWe0xUeTYVAGg6k7fesdZDlE5s6mGkwaGuZWv/R
H6Afq6tvZ+NSo4yeh+kodzn82IDBmZTnyK6ohmZeQuiBSR2lSY9R5DPWocNdmCn7BIfB1eIC31w3
BFcttVs1vBB+U2an8OdqQbR0UFLrVMEeTBiL2Zo1nUD7u+us+wvpSZPRi0Jc67kRiFeYRVeW4R2V
j165ftfMOVpRnoEwjQlzi1nSsSeD7h4hrELCpVNxByamTfZ8zKLGpBSThJ6H9fEpy6P4jDfkas50
eg3T3q8ILL2c6EgR5xefdJDirTXZEkSuB5ewvHqpBgcvR5Y1hO/nt+D1jUNo19Bzqguy5Y5z+xNW
CS/MOw9fDGNCeWztkajMhv7O1GxM+HAlP7A9p+dH0KXj2Znb8hv2ZyMxiJOi03W+NeDmZaC2ukKN
LMOLZVyqGG+pFku0Ij07eUPC4LI72+e6mDObvaJGiN5mWVK3zAaQodRYz4m3+0YGermaFLS2aNn1
WoPXk5lw7y8H2WNkvzVAI7ZIgZefwRgpJLN1MJBWUwtRYQENPtEIyh1N0ky2QoSqu95whakzpajJ
mRLj0pKMstBrDx53TB82a297qCeJXn6olwU+K3CDf0OnIOorFoZc4Sdgp4/GDuomigKX0Y82ty5U
qmCTkqSCAeFPbooXV43+GJi4WfwcFnMEwvLcIJVeNnyId7usjBnJ1nUxIK4tplOo3koizm05DJMl
ktIl/nmrkA04z3VyZAlQNYx5J8K96HuJ6ycDZGF8zc+8fOo2ZBGRDiGTG2e0yal2+ywJk4TDETfR
SQzW86RYi5C+Hmu3PunqOe84hkxHDjP434q3wGBzWvk31jA9fJs2pNarP0aQzZVyjgy2iKXEhIQ1
F+IvTpY2Ji5ZA/0TO5Sfi8g4+nzx7cjpm3u9ngxQhGIdTQV1zQXNkwCW5KKUnQ7wX9R7imLTLGKv
D6rHIpqk9EsXbrVInOtbQ6I7teBsIh9PxAtEH73sDvpQVTTP5u1hTbzCAzgCybB9lD7D+tbTdgSw
tFOHix1WsYZ1+CQDjIvBhFI8fzFiOfvBdMl2s7O6/n0WzeJY/Uz99asKiiTKVuN+APGEgCtT1plT
K+L7oqVjTIV6XPguw0VE1wFqAt8yzfF/HRhnlW8APybklP3xLRngUaMiS2e8oMN4bmYMRHlncqaQ
WLk/YySoPIWyG3SojhN102EIYfiBCpJce5XDOwCptoMKdC4Xy4vI090IbGNiUUST6RcyqWBHOUQV
HneXv1AIBA1qTKcMhxNEZEme5AR89q/YeoOVAyAGZwLXnm8KIZbzlIX9+uauTgHqkxIZP8StXFSN
z3Ku7G+t3IDRJUfM6Nt8PRHHK7VSBz2hXHe2ZBx2tCwjJDja1hqCCVs8HT+xnXkJctHtSzxCjEzC
QBX6uzMgrP2t5Hi5QfE4sJDusNEnm4F5XrvGJHHVDeSKaf4Ys2bIk4u6MICLlPclINUuUVQ9kh1E
SsTt3F96YdCASSPeLesEZ+GQJGUE51xSsY+tXhfMU0h8AeJh3dVrZKO24hepcuZMm/PSc8v3fJlg
yd+8/OIx+ss3b3Q3PrwqblM6Ch+A/WQj1J1UxW/b/v/Y5TF+gD4FwmHf+PZog3vOZTVZAXmoMsHE
Dl9rAYV4r6XzKGL27+y7YGRR89zlwGE38ryItvAh21BCZu/OPPjWq3niWjzRaMfPiv45uuQxVLwi
1fRAC0D6jAFQfzLgEe0M9qPoPiYGmNN0XyvlfcLerno3E4s+GX0k5nIKLYVd5u3K6uJwt1fYG6Vr
4Iuv9V16UV9bZbFdyX1amC7DpQgpVy1+8+uED0LTln/eYryuVKQgI+0hB4drSa/xjc4DfE5g2e9N
g9doxJ+zDbF0jUEASR7EiDJpbiDGQTpA+yCumpjq81102pf9yASpht5JCyM9pH3BQXOl/zHfVrNY
8TOlUJuNDwqtPUgfItjxUFfFEblzYXH6NNjfauVo2p1mfwmQdsdMcuBKFm+Wlzvrz45wZymvrOze
XxVy8/pomtHiIhHBO9UeV0no6V4W7Sm/k98IYfIs8AqR+wJhwRO3DLnBDosPndyVfbEVY48C1ULI
kl2Nh38WMwUGnNk1OziG80hOdwfvTT2fqKGtDRCyh+uVflecH6X+HdT8GlflcyOavbOYU+qXFddX
ln8XjkWFuTVbjgoIV9xbnLOciJnFWCg/w+/q1Gtis7ihSECQULwLQolKkoj+vrRe9oGOQTTvgQAq
7zVSRBVYkUPJBI0mT9zvHAfijz1lzByN+A9sn0ESd2eToz2tMrNabp9I9ei+mutdYkx49/3a4o/z
G+Ojqs08RDx1PW0Ve1+o1iRoSIDUGpeY6tNFJpc+Vz4IKPblhBlUq83w9po1youSLGb2dAmARnLR
93K9dwTcfohVtyuz/5CfPS3IZwGHXer7hOHxXsjw4p6yKd1s4lfVbgvr42mSm8n9ammKquxPEwvb
x1kB2OHatgnlwZ50ymBES38mD+fnJYPb7Qzsg7HPFkAz8LqmXAFnUMWBqTCxjCQTYjMIyQ9HBUZR
1DPZPuhl8QBGiB7623YG3f1qz51i+902zoHYjMOHpe4X8lbmELQ3vANJKis/1UWXK8X+Yc2ORwvH
g3VP0NSoGIngr12TJJXN8QmmO1o60WNrQvk456YFqs8wxwxqsNjsdCviHBPaHH6isKJBVHtHwMiX
Q2B+IYMP819YhDQXtQvSC5Dfhjl27JgThqrnpNTICmpK5KHoL7ICxpnf9o46REFk3iUNbf5ig11u
R2CETUMaDctYpXPbSfMXZUmx84zDGEuTx8MOT1jOyzXS/k/HMpIF89DrLs4xJtpElt/bz65hQDRu
BcY+C8tgs2z3CjAogsrY/GAEE8IN0VZVJViNG2niILmPoNza7gSGVlxzFlBVMUFVllZ/4jT3frta
AiThjl7UOrk6cy871HURJzlQSunaN9H1qXOLsPE+t0ekyISKWA3A8BsHdX/7d/cRupq7Ng+on8ob
U0/JPEWczoZQzbkBqZj1kWZtjLHh+UFbfXXaYGffkzAGYMfWEtPYSiQmPHhtJcEpoCRQ1Q0QDzWV
9TpqTdsH3R8c1T2quEltNRyjchcBJjXa9L2G5SI++hJjPLB3CY6aXLo9Kn2aLjqHJMcrNOrblQuq
7Kxf1Ak0+LQwz7KcKg5PO7wU/ja7+N/i81e66VJ+eG8NuEY7BL3ws8SJtFTF1v8NTJiYNtj1J7xF
RZuVAd4BZJ8+wZBmcWABN1SrepHdkZSX50zhGBnFlaNOqamvnN3pLHc0CVXXMyYU8qGOYqgcMaVZ
XbztFcLbiD040LGAEkpARc0lTlE68UkO8ehcVOTrOL/vw/eE8aCmKMUa5SbclnqL3oNNoKHbo14I
yRBfH0ywjA/5QAzD907gMaLFyeOW1ZpF3FgZnct1+Q34HRH9Apb/AT+ITdqTYixkQQdQ5srwgofr
ltEP3hNWCE/1SditpIdQIs91MA7rzTlmsJL3GiVP6l6gBm72H5f8+6GL1nLoDG1/3n7axOsoNY/4
ydXHhfsgCv8gWXE92DxLMWYwbscrCKz0yBQHp9DVXkuO6EYglXDu3e/wx18rS479pmkuMrlv9TXa
vRraih+rWydQFBJmd9cH4hhV3FcctxK0ZF4h/36kik9dUcWTw2fxxaKoIPD6zLhcjyRoFH5zdOh6
fvxL0xgaZlYB0nkhC98DGBXE+ERKE+GxpwGGSpe1SvVyjpZcosWl9hZdWAFzPHcLNvSJ9GcyKhc1
QQ0L4z6jGPfjLAZiO+QluxhxpWR7+EPRKqYWZo4RAhM+vPH8eAeL/hsAinT/RAaPd40ZVtx6YS8S
D8vrb6wtkrktCPNOm4fGJbebaCKO+n6ZH2jnkZRfEmYAaD2BwSItAvLNklW7zJpRAvaElyYtH/k+
TOA34CdWfeZlWNZ7fLbvRbqnAqsAkeiAnxjsZQ1/qqsSfScqqXLa3rOVsF4YEz2QjSMIxUwzvYCd
5UkxGtC0suXqFSziK8a+rLdOOBxUGXJyTDvPyjvHnt6xvPWNBdzfMhxL/qMCO79GLdG5bXr+ggTO
PLWeiVSNSRhz4xw98L9bzNVYM/xgF7KjN8YN+6WGMpY/FegSrFF96ZkamHqqZKjvdP8IBdmH3zmB
hcV7H/fktayFjZ3G38pQyNsofGSCi8hZs3SIw/azsAOk4kbb+UgLWj0FGm54SulQSlRZaMiMb8dq
NSJkxn/th7vqUv02p5aebcRDx2FN4Nou6YVWiAWb5TdgJ/81/8XTQD+nqhwqyLW6xuoJnOFeGBEl
Og1ZgpvgaE0blXaaGulqgl36+hxL5CIkdV/TSdbbvRQ+dtyEpvS9jhL8S3RplCkyChoOBp7XamsK
K1iz6SM+EM6dQI6X4j0Cm8g0vuzdS7fPX1/9mqwS1gNIb+oEPmhN8RFFMdJIItXQdB3ds2knbcG9
F2gsaA8FAg7n/CNOLoagz4MC62jbavFCT28cKxt71yXMre9bK0cRcVz06gZ/j4IcIgyPa/eFivCo
DT1w+YropXJu4CX5tDhJw3Iwy6s6oyexQVM/x6kg16m5HGC77m18rmCSijSPsl8Wqed2URDpHXSB
FqaO16tIT2aGkW24wTysHWYJcF04HDlKdRxzAPQCCC8CkXcJcBQUltljOhVIxk748lNQQ84WuHyR
Yju6PAEHOm2xJNTCINjHPnVn66yq3ENYxBzQiu3Gz5qpNjNabi+ejOadmxK/GGxVsJAIFwzNTFeD
8D1sc1+lK32h01WS0YGQBCkSnHqJtpk5ZWOtD8Wv8cycOOkBvAHS/wFM9AzzbU1EDoF/e2bSHyh+
bsMKpBB2ZaaKHJjyRQnbPkNgFlt0s0Pe6SHUCETm4PmvRV7YH55Bh9bKCRkHhrnqMzA/N1YBz5N8
w9AV4tP91zakQOSqdbR3mTP5XnMJeaPhKzD0HqKEVAIy10H0v2GOLsIuFG80+bFyCbcAE0Q3ssef
FRGPX8dQWq4SC69ytMsKtvibMc/tkRv+kBCc8AtXQv7O9/uxBQniP1zSmP68L0+Ei/wHZqgILdwg
5cUEAVt0ICZfucih3hrO9FNO7POr7co77CILJgewsKbzEiYVnLKdw0DcRlkpggKj22NuEaKW5V60
1FEigCMdWSyiqeE3HdG43KDv4sJHYWfGMKmrascz8J/NvF9m6Q3F6WJmqPWONtsR/GxNVC52ROK+
+yfaqhjQDn/U7RlG4HwyY5kISvlhsXtxhYAOn1Wg/dOVxmQCu+UpM3of1hVMLnEK40C6STj9wuLP
MMeuMmZ1xc6KaPAEwhfKzv8KiLdU0OWnjpBvqpb7B2yAlyTVdh/Kpfk8MdX+IXXGMXwUM5VBFApH
n7wOKtjeocF0CBSOmzZLg6JqJxXVMtPw/V6rwI835utzRAo3G9MPCuqFfVa/oB3hYWLZW/drKTLF
cg+fiOi3W8qz3UvWeo6kDCkoE4Q9/LS9SJX82x08iFbLu/gupfYlStBNaHxy2dHkNgZjY9/wqrFM
SMmnk3pYZ/xp/NWUB7dmJNyDJdGSI6PBK91oYbx7hqlYTkiaJDmK2ToHu1wOzzzZBF2S5Pz6X3EU
yTkZLEMP6Mxld8C7Nl+EtqMb6YiQgOfd+bTyk0XHevwcYvEDWNS2yYefe5Q6q0RSwjw+AYiRXWno
V0FhVVhQYjsc/q/LzrvHruLFpna5W3c0xpHJDMEFSwHFUkhwN1BzgQFe4CVd43ipVyuSgJZWpxeg
o/OXBUi95EZFxRrbxI63ZjasQa7DfBfSckfdmj4/oDAwPpxATrVsbWiSPxMMdbvzq6sMK05qmDiV
I383I0N9IQV29CfxRm73TlLi9O0FKV9KQE3n+eFF53+E6yn/fAzMjqGHkNk1WIwPFYNcc21JnaLO
qMv1XkVo/+nK99mxqKz9kiIuVHSBdHrxOklEOwbIkjVkV20TtHdbE8/q3UfYky9mwmseOUz+TxUr
RvbMSa+KLXawq0GySw/YPKlciFegNwehvXcIGAyRzh4QOqmIxo0iBpwgMUMz+qv0ofdtnQy/S5UX
pv5ISWSxmgfSYCos+josuS51dAn+mOz+7fD9RoxjiZSwb2X/AIc2IKYMkVXbrU8LNTJGvAMMSWNR
U+jqfn7TkPSJAnYT8UeQ6kg80iy6z2ObekeLeZ98rUBhuEBSOm/s1Z0gBstf3LqqVDteZFmSMsYI
tEm2vh0pWaluPhFYoF1csCWDPhLRG+szgcXFlHYXP/w4zCrraQJZFkkS4flBQUmIMXOieuqKoX7L
Uy7ApNDMvVPMWJ021UMdcuRYC2EVdSSBdeRPpJNAh8LfsMRx9kWV+KY9xl8TCfT4OcQGrf1qGHT0
JrRm9fXte2Cjyw/vOQCkAEHRq4LE7XfyMR7anrdpKLdvh1lpK492mc5giEBMV2+igm8t33cN1o4O
6EJ3FMhSUmuRHHt8zFDrgUqiUOeHYuFowU44B6kjh3iYEii3oHlD7xAvFDPH/nB6Ond/BipPCTSW
ByuEWj8stxYQsqU6jb6Hu2gTUyfjjzqMLzabNwf1gO9vZ+vFmGDuDX8/BvkzZwFBksCph+MBqZaQ
BtAR0AEpmLABztqVyJSL4LsVHVTU/w+cRUXDznoy/6LYiwN1+OVP8yGIWXgWAvoPvTgZXuQ85Wip
+OeP+3SugTdb0t/vUkm6CsblotsUNKagBiSf8AoIIoxUrAV58jA0Y2CrJizUxMIgBa3x6Pf4dKlM
Q43CAdUDZtSwZ9q0/CaMKkLopoHjMXoaKU7sOeYduBklbTazSjIwB3xKK8VmCr0+rykZKyRzOlpm
iNnEmTWkE45Fg6eBqCZkuDeQMFyPeKJBzn88dfq2A967FRNxlKIKkEe/3oxdVkdV2iUHrDxPc4YK
qkHFnbqMDmBFxg4sduoRREV8siN2f/UiXM8M3T8f0lwpxpSHRsH4QK904OxnRpfl1UYum236C2/M
YJz4DfC/ypi5qI/AFagOK+HP4p99P8bosX2p9hplb6xNgxaqQlZ3b1lhim3SncMx+bWvEvduSLQe
f741i2ejRjUlA4Tn8OeWLxyPkqokobM212qFd/SekqmoqBbR3BNHpcRMWCbJawOsPXhFHXu1zUcq
ORvFlVVQcP5tx5fmRgkC2CP0IVahmCsN9YClG3fKYGiDjtVGxictudxVviWO2QEdK4NtdOwFrzdg
BS7Nzr86922ZgzbsHAlyYrb2n4EWHP/vz6wcLKF41gUMxzmK8hYYYCMLEOxYty9W/qLoBQqRFdjI
Yvv0ki2z7TN+B/2Itl84T9naL//107E1T+MvDdL9yJNZpwAVP/yG5IImjJCLqf8r1GbLW5uKa3VP
/ByL0gXLsJJx939FHPSP1ebVWdCrS3fvheAlbVwcCVU1cFKlPbJUQaDvflGDPXxcxZtD4EyiRLBo
66DIr/yjFg3N285gcwbjcZEIjdhwWP1GbefFqP+Qn/3RnFsyzgawMHdhgPWkf7pdpFsWm7IS1dKP
WCJRX88izcQi8p5mVF4zKPXGHpQBmRPsQ/hbvW9m5qIUjktWiya8ocwDl6EhsJOYdPpjtpqk083g
DavdQVKD5yktLA8rYawi/deOBcKTC0f7HU1Nzxn4P4x34gjcq5+XitlxIRS+TM3maLjGnJhlR3RH
q1HF2DsDikaTyQbKze6DXRG1Rs1S+SAVAywTgX0HrPFGB1ytxe+ZbgVwhguy4XM309ffMnK8ZZ+c
LZUtP/Mxf1wkt95sfwBDrSgtlRwpYvVYZK66XHoC9wlMw6C+84IpCBKFJAmm99cJvaxrxxViFqSq
JzRtX8352A7iuTQGOTiLe/z7iu8hS0oPfvVmqc7hYz0Cw7kecSBDaqqvwQ9on34gnpFRiNfLjT0g
0weB4M7/9CoJH7bqbaqYbU5b6NUV7obYlqGqJgmrGgu0my1BY70f9iL9utGDkNXAyt/kjprlRIxH
On+kSvngqX/xwOwfCBnyCYNsBCYTeH++x/F3E87MIIFFVah7+V2JChdP6sh/4rxCemBmx7l986Lr
EkZNcWCXNliJHOba3WTunOYYCppYVfWC26Rvy5fmi2b73h0iIznfBbFu12raPLqQ90IgiH+VDZIc
As7hwHCEJrEVeh0ySuH3DkpwkN7sdt83K3dlYKjhE0B3e/F5wsgW6vNNewYwhNRyScThfjdpOCv4
5jPLMSnlv51G/OvKDJaZSYr9ixb6hbOSvHIHMORAb3+W5JlR/UL3EwJF6s4Gx4KYnvgUDZY2kLZJ
+3O/g/wB4fU1ZwtB4C3A+h4SoqNwGOa8oBFHpjxnyhdOkiMq1hodvGXmEGyXrOQJaCK8AF+41pNv
NObCS38Pb8DDWJzDbrE+4lGpkN6jnqJun+HGtWrYHKkxmPNKJWwRAgn3Xs6nLadQknNFho1c2CUr
o0GYq/t4mE5bDDG8rfCgrRSjsiYc7tWoF9wqB+NFeH0HHTS2r25Pd41cPfAU5luGXP2dOxvtGvSv
MUwS+zHSvWOJ9SYXEdUBNXzpWQb65HV5/PmFQOs49ItpvxjKuI9OAGErNH3pOCHQnTcdeCTssDx/
Y1GcwyHha2dNsMXSdCkNtmC2XR/u+wpJSH1k/pko4KhF0A4DKHyfyusyNoshvE2k9fuZSVunChku
psA1XCHT+IgU06W0uqimrtO4Sghc/ffOHfAvY4iVDp8RhbQ1tytqPkrUxEmRizrWVKuaix3t3w+L
cnsIZ+mNaE6Pbua1C1xM2AXu6Eyf41e4l5YH0fLkohQLJpXjiZyDuN5so8hJ9W27YOIq0krgLRH6
CDW55UAIZ/d9bvjDpWVbFr76u656MpgkVNJIdBG0sPxQ3YciYdsmn++lWnRvO+A1L0rG8DvBQu/b
zIKP6kVUjxgeiMEuSoCq2olaxGKIkLeMWNGZrvk6vQTLaDtUl6D/iL8lsJHA7uHDZnjiSEfEgDJj
2MvTOn54TZy7IIq56LLwhFqQSOcW2rqkqYnivZy7LOP8rBxywwtvUon6GxlNJYJ6fGd50CTaPjs3
tY9nE9p3/D9tTkFay61znqnJceGSbBs/a+5tgsHsNfcjmJP14D4SGL5tOwo4050//xZzcgyDnwz/
86RfgLBctVK8scK5FD+gK4IMXQ7ZZV6Ta2ivTRGuVWtRPZp6yniWZw5rmtFqji5QZOCokd4gWZ3W
srWsfja7fxwHqPOpmAu8XxHGAzKaJ5f2W8riVGYo5eUsA57mX4+Dv7FLoDKpGfBdzOENa1sS3AOG
nYbu4DnNO6a98zjOYIXitZ3s3tThh14BItKbqmk+eLfoIpMmRg4AituWBOYvoR01B4zLC9cjtma6
xbay1FVQFIllALKMrGvib0vpBpgYPT0Z/nFJ+xPhqgHQOSHliJEJ0xyMsD/oDjPFVTFOx7jd3EnY
Xd4tiuPuaUw4fSY2G+lmDaQnsb/iUPSc69uTdqAUwOX863c+FZ0+6ux4xWGrWC0akwwd9ltoT9/V
yGGu7gkaJ2nt/9+i4E2AsPqnjqcG/sLnUD2Ds0IqWc7Ay+ZtQ8CmH6qRj4/vAHzW9tWclaMipHtl
ssAwiClDCjY05hKDBvU0JN2QvEsiDEYV8+tKsUVrpWZLzLet7psUmO7LwlIWnQ9nfdC9noZiYhU+
K6VHImI/wKvMk2orGCK+yKQ9trxoEZKXBeN3PSFZcZESP7IuSP3aZRW1/zKnb+H9DVoiGpAp12gu
7eRndmszlAIbkDf1ZdMb0AeTuOYUWtRZ705kQJEu2Iim3U0/EWlEI3TjdK6CGiZ7u6NTzdGIIFmy
gYOZMhi++oo3Kb8dkjffJMHOMgc7dLOiJd6IDO7Qm9heGET59dhgcdhC2YM/fM+9ndEb/z19MIJG
DOTqFsW2zKBFSMO5niQVPCxEjksGK+E4tqQh7EHiAJ4/39Sl25ssLKoXIUQwuosjnKWYaJ5pzaC7
9bPWrqjwvnq29u4MXH6mBRrL8hEzuT78Ew6JKXARwE3urUw14fa+94mzsq83xLS0liqpQMhiBAcv
BCJc52O40LKOrdEgKl0fCNA9EggMEdsRnd6NB4+Mcz7UkWgMjHG2kcy6D+K1lapsDvraG/FIGNFm
jFrzaKsds/qI/FsjdVBQoNqK9qUypfidKe/59EPAMWaph4n3g9GOwu0Orv3ttASwArBD3i+7j3Nc
h7kultvLaKkMRvE3NBMpNqnqTFz7mf2fXsXq564GalJlyZzLV/KejVs5TwQbJNQGLcxdvgrDCOp/
P+xwnBI+1T5+X6SVdrmAGXuQGki96S2Wa7FZxXcP9g0/TaY3C7/REEQC56ydIFeb/idbO/s3pC/1
RJlYTGDFyegvXqbdnYyx945zLcZKpfYtu4LV7jLzcaWquCH25t+GmI6Xnc5FrtSdYcKA4q+tZlo0
XntF6dkKzHwlsYX5iohZwtfPYG1kxqAjvDF47tF7ASH5GEqJsqzO27uwFMZVFsboKcUmLzmvPXns
vzho5GjV1VewnpThmVUsK/e+sWadXXD4l+sIQZ4j5zCsdU1+OjEp5GN/QS0ntNy9e2kWpSdzW2Sm
mteHLLVoiCBHtvCISKiwjloMC4ckfywl9ROSg8IIYI69H2HyNyYh3J4fObYOQNfzf75yGhKgSDjx
6u4sDhF9egpsS1gdqXK1U+ASqVq6xbuEHnE+68WzZ0Ss6o2BOR3zIRZR0ISAf/ZeXF6pybr6Ueni
H/ko3ZvEawuSL0C0izgsM43PzsbxLDd2+uws9WyvrD7tfmTIro4EFlILdFvrNr2WCf94WNz2Iyft
OoV9q1pNz0kGSp8JVK/KGUpdTHW214AHbVoKXYFMTTyFvRqf6M8D579QoYQE0Z19qDV+nB/a20Ts
mdf6u354rRQgiE289ukHzshQ1kFL0pHaUUuSB7z3Ibp65yQb5atJFtK2J7lTbrCJ0gX/rxzr8rd3
yokXqnjRBedaKs9kQxt7vpvy6QAirJ58MV9+Aym1H/UW/WQjZXQ7zlXBS9LL/7V6E/AJtcxWiKgu
wyPsOt38vOcQH9KEahxRTeb7JwJvm5ghsURog+mRhUFgRzHRVpPUC0xgGq+B+LO38LXSbTREK9qB
0sAg2KI51ScZdrm59jjWbBkVAnSChCv9WXhXiPwCFNr/+WzcCkS2ZC4orkVddB07Tn+CqQgd49uc
wY+XNzf6PnRu8UyRu5gHZLKB1uSpikX3sNLa86hoxPTDahY7aQQ55V97RJsfiOs2X3/UTQQKh2FZ
nv4+IJFo0z4N/rdVxL+ETEKfi82ytNA2r9sXTItFAXSBwONW0P7LPuQQ0mv6muF+OGosa92eKbnD
Y9krJMlah55bVm+n+rWCrAykvDgbCQbBe9laA3d4QB1Zq095Jy8PSFdfA7oLx0uOliH4XXMBXw5o
owhnlKnXGlYr3jJz4Afcvu4JOUe0lu/7mI+Wlvp0+bbP6IgfT+IfttiUSrJVmHmilDQLR0NiT7ky
nVji+w0H4iFoNSszZzf05rwtXlXPJ36M9AJsEaATmsy19sc8YfPeyYjJi6ZJbTDZ5UxrmiyfinH6
SgKEIN3HVfsCrG4/Pl4zPihSDn14KFowkKEHOTqhaizfPnLWb8cG+csaSoDZBzZ+3eiroGrNrLbk
TURx3vymdZHhnRBLKZuzPpm6PMZXisyqa9nQxVzXwjOTkAJps9vqrzeINCZBNO4J1lGIx9PvoYGc
xoOL9NbvF+ek/uFnGZI6dhv1ucYjG/6ojAz1KG58Ix0rc69hw6z480iaDOecjke4Sq43m3gqA73c
SQtU3l3BUaNC19McBjd5VYX+g9hj0P+/9DVRarCMIYLOAM/1BZN1Azt0suX1vRLf5a0HhiXryJd1
98SHQpoC+8v6ETz1+UA+tD8XbrQUtl9/74vAT4ZKFldJBgcB7sk+oc/u4WwdP23LyxPXjp7PeSgQ
Snd952xii6rXv/OGnA2us4taA1AAq87+GMtmOc8l3jw4smigijNVi2E+VO0a7DVCfh7SbrsNtY32
PutJzQc3kL38L24AObqXRuyjQcNfFzNKfiTOZG/IapEhoHPm4ufCQ1Iv7EJTqt/23aU+6KfIiX4N
kOIXesqWeAe0Sg2BSFI7VPtAX1jRE+ZnikZtVibn/yAsGNepKNI7N4DDMgWg9+alS3Rr9hM6CqBN
/46kW8ir1IvTEaRQaWHuIBLG/DiNpHVUtxBG7uy1q+Bhz9Y/5TMuXSEJ0NozvGgCyGGG4z1aTtAI
G7sX2tpdYdKq/jHwfAotioW0WEbJQNVhh3wp9zL7XyJMyv4Z0c5sfMHbnpjxGmTPcgoNwYM9uV49
LxXcx+nwFtXFPqBthEGMnpI5l+tuyJ0LzqwBhoazqgBBEGKVBGPDp+lRqmQCkuIW/eWVeOYcS6g3
NRsivUfwsqI5gjExxANnZuqRBr2MxOimAANNcWk1BnIyiaDjKs2l9XK8n4CCsmykJbBQG+kEKvaU
4oPgrM75YQ4jgZQTi93MmzRg8Buhsx3EHGokf2F4/GFineQdgx0om21xVHvJsZwpLfSLdeMc1PyJ
Xias/V9/uWLuchdaHqTt8LvBEbxBVcjJUTeZRWqMLV7I3SgGHl84xaLtSouIxuCS4un9ZRTeRdK3
ZsrTNEm/DxQLiAL5b2fjufNC1WRcygpK66TkYuwOuJiDvaPtmMM4cqho5nL+OM4YF4R9r8sBTYyE
b0HJN5H2CZdzpDlswscoO+ghJb6lz2oCynq5YWNm9TSgueBcgboRrxlH6WSphoyyc8SAm2YOyqYU
ZJXWNWP7lrswGEpdD+wqNssPI5H20fHyKA03gfr4YvFaafLdlBvt5COmBCGkR4kgeaJDfXyLLWvi
Ts29dtwy4FKaT409pESct/IzWbfZlYPO6GtliQYlPygcVEYhrTCnqopCcooqZBEhmtTq02cYajGn
uMmnZT6ozEjdK6n7+gMViqzBhzcjUC03/COK+4y+noQe7+7x8MTWTr/cw4oDpnRQ3AqHtmyRT7Pb
RnSjp6ZJx+QXRGD1V6o08wn+jTH5gau7xx+AywscmZS7SAK+afv4wbU2lVg+JixP9jOspYwDXKat
L2ex9rrBmC9cGeGCEGTJ2Wo7ESgFtVcH4utPu5LzmZm4RIwEAM85t61+0bEVrbBKVZMhVT2RLDbV
irdSwxaFwSGqgeZgU95pTDrYhbj1oqQaA3CQGodP1sRugJ1KlThj95U5IqRA/L6FK2zGLPGZb3iC
MnVNU5z3x/STb3d4nviUP4Fnlw+hZ5ZCRwwP8QGkbJ/uqUZMtEdg8kG7yl3KT1E6KmXpkp5U+Tgl
wzhwJT1tIfNCmMMmuG1RxoOYxtnzh+HJl/6YDfsBOWzF5JG+gunVDMrxy8+Ezq0eOTx8wS+tAd2Q
hM8/nGMbp+Yl/pYeyA2XQ2i4qRDvGOn080irzSmm3Vcqp1uq4BhUgIdRKT435b+cdeyXvukWeFMq
YVsy9JxOxoZxltSrz/LL33iW2BEplxoOiLsJ1wkB3ArRRnJqoFJF9Qodmp1jyWi0vhdxWlEwmMzz
kNX0OJXXd4gElVE7fsdDmNmc2AKDCVV3JVZ7SgKGQDh8B3xcIHFJAyWDkzHMLr4AtWFK8Qgu+KMo
R5c+Mp5cNowY36VrT3aJfqZW+ZtxFwSMlTs/pVlgSq9luS5MoToDPaccWWF0BrMHQ98c/8MY4Tx+
dLW7t/BQ0aMmgRtJUTt/Bc9DkMelHnW9mz2S8q+HzQrTdg67Mss8H1CXtJ1VMkjbbE+hqA+L3xPq
lyJsBwfM/dREiV9n7/LVRKT3seuXFofrOlNEnMPvwtoAy/WFS093+K4WtugTEMChhGT6UB1k75v8
KMgkjwk13JBZ9xWC/pvD2xZPDAkv2+Z+PAjs9eVCu0IjH8Mg4Vx+zCLpeBpSfwQzfW4N22GgmEBe
e2WdNa2sHEy01/ljgJ4oel7jubMdlpsdAzu5JQUKetZZk69ylZneVA4M6FF68Qpmp5VoPXhRaiBu
cOICERQ3K++Xjk/zscNigJjP8SphEbuRJ9zIt+e63fop1nhqmqIvI7wua+vFSPmffxvIoqGlDdGp
GUQ53AEMiXiRx6//eyl8sys95W5GpFyLT6uyHBip51UaJfz/A5X4VSOatuRaKlNIo9gvCtoV5Pju
kCED8q/MaBWlfGFn4V96kRlot/tZ9qkjyTBWV7/jvunFbukq+d0OoMcGWqltc4SLa6bzp2ieAHAL
AmAF3ZP4XvIe164jEoawSkRU1lAPIF56oRSgRzIHr6BQJu6faw+kBaK6lWTZ2kw55z4IEudqrz2x
gVLLRqNAn/mOYwKhtgR4pDWTEVGc2f3WKyGYAl0Hqxph/AD2FDSJsPLKlpJuViGMd/zgUlPbHfuU
UfPfkbhAnNK3k4OYFs5SATV3f4EzYgo83O4GtKoRbDq17PP+XFuvTrXINiG3Hyzwq52IUitoVrPw
WNpyklew/pFMOy69ES40PcB3DNnp4XYCLiydZKW7UmSgIlR0fDIt9Jcb6sdqdRV6KP2CHO1KKI1t
KPOvrZmDagTYnZ2B3g4++MA3xwuOxGh+DyGTS7QQL5jiP6YMt1m+DS7QDwZ4ZI8pB9VawkVAHKpy
6ScdIZyhnDVQnJyNe6ja88Gja6gfnWExspaH6HD4mlxbRx4URvxSMVERLh0rpXsbTRxrYHuCIOnw
08M/tGYF8xDjvGc+aDrlOQwtoXGzdql83FvhcCbpvqLMPl+NpRJO0PLQn2lnK67OEyHneD+QkWg2
1Vo6x/cBeWJfM9B6gWeQ/iMml5ajRPkel4FJKxbQodEIR+kcRgku5ReANpAzaociwFWYB7WWvMxq
fPVKuh5mLs3e83fFYMBjte7LK5gtfvRvvclaDxM3cI35oJNKIaxd9ez8vlfWwJja1L6n0m9b0xQf
ZNl0A9MC0k5/OFtvGTtqf0f0ux5+VTJ+gqJzUO+k28MKV5I4FcrBLSzhvluw1jvouui9XInHElJL
V6hYlGOyuZvFNgZpq29CJzjGLh4Z7vMwGFY+isZciuODsAiSX7h94CNShTiZg3GYg9IY2R3l0sTE
MDLHclRuSJzOdcqHa86II96sb1L4/McpE5inapHl6NLud96lM3TcW9/CosBuNiTzRkIGxsR8aGhP
Jer4VmAUt/ckDxJDv7L/vVycLinmTiH9uddHkzQiFYRJZqiXCeRs211DAcJVpNaPt9ekkE5WmuRY
bIh9AJOPByZF1zvtU4mra1p7JAB4XSfQXlbPYOqtouqBHBWv2pPQzedQX4Jh9GXVbHwGRuz5oB2s
DBZ6/wY3A5Wpf6itNsIpiavTCBtkU5LhH1ncT1/vwHyZ/rAoQJC9I9AXCPMZUCIFzndX64hI0CaR
iA02Ql/8YEYrEh0e7AJjroiY8qbi7UkYVVq06m7Vl2a0ZfXmqpA26BQTfWiFzkwI/NsoqReGgX+6
bLcFzjwczKugkiEUN27qdamZWfq01csqZAyNuEot25I59RZd+QWRV3NdLs5lxr1nFSCj0T7DOYVn
hAR8P4jtTGOE+BCBFcJm41nDz4Tvbu6TwLtO/4ATUDFCkXmagJtbgpdjkr0Uz3O0hZ9jmVvIy3pG
dBRdDySklF9P/Kw2avUzgDy6wztXpvBB23jSMfNS0slNh8wq9piK3loFO90unDXWN0Y3cpgYBRti
WH44eSXA0hGTbCXAw0F6218Gll8sLWmuGt7mOyjO0mfHy1kGh0HteuU66hjTDeIMtaUlj1HkMsZy
/3q2Kz+pmPyNoWFJVJyPBoWKdsld1V3smPV/yrcwP2mGc9QY6cfZFCXCvdq3XMTG40m0/+1OlyE7
ciVgWWerbXJbaO2XwS3VITirbupKlMgW5pFgSHRHmLVGyjxDflleOj4wwQ30VIeolRAjWvi/pV89
qLVqyRx/0zZGN63cL3EIODKKxjKZAn4aoLcHdPVz82q7/w7ceacsJ8Ij8DQiZQpKBocICXgdlIwe
NXd4j73ssVHE/IaDKDBwY8+T2T8qFDKGSlm5wFee+GA3ROoKeGIi5vQdAZwDy4lfq0tQ2PFDGgG6
Ell8idvJl0PUtkFQT2QLSwbyEfXa8ZrtyLPzWYWqckKNptmQWMFa47MvpYqKX+2RD8L02nUPY/5D
JJLTGEuNCuFWOWG/Cu4Y4Gx6SQ6aSrrS7lM7HeqS0VYJfKR1019CpFfyix/BBkyCFrCYdN6CuOmq
YekJG6uag8nLXX8GVfVGMBZOkl8dgT0zQHipTKHToADdQxfuDiuoZOkgS7VPANtrBk/wp8061XcL
Kx6S4cL3D/0ft4f+kx03k8Xa5bE+sDyUc8hM6XDN7WbPQzECYPjn8Cn0pn4h54uc8hPiNY0hBbJd
hKpuaJAXKymaS/L2vmWBWWl1EIpPGMUDpSx9MhYO56AguMVqYz7DD2qciDKp92kPfQt5LJmGBuC5
8oTFwpEXHW/L+WNKw9J831cNqxxvmU/5QrxqmqxdueIFMjFats5TUKOX8BcxA3kmH3HAAAl0lGtV
POTDsltvgo9KLarildeDPOzD3wRn3Jb8dA3LjYnFRwSt8+9kHsyblQIc7nCT+NJM1LEg6esWGJrB
jCa0VJabk/3MpKcmghFErqAhZtvIZtIKbQnQPUebjBy0zABH5u8InQ5xk8MgT8LSYvsNT3Sb5mVs
zirHH3w9ZH01JuqLdyIsdmKYlYl1hjzYqKfGuna68MuUHa/+gaGkCOW4bAmgNQBtkHqeZoZjEpFo
IyOdHmNtedIIVYmOkTusxN4zAOjejmp0YRUdMgd/XFEtLxO+eNBuV/5mbbR0LTu4YJ7yUVffxFmV
FlSvsowc8tn8lWOj/986qAafM09Rj4nNf7Y/TQwoIU/ENl2xFwFxByyvry4SM6Vz+q4UcY6qQPHL
G+4UuAdaD4qaCaK4h3sMCaMR77Hcq7BQBjciUC8L6/HtecJHMkHRzB4wKFuFh2Ofvjpf9tJPGpgR
vkbrv8iJ1pw5zDl0PUWGsfIWZTio0ou3ngRfnN+CB0ECaZ67vC/opE2Q4oySJHfgOtB91q1yb6K+
gsRuIODWJudxW/GD8DV02bSmQolGTABPgYF/2D7BJLNoajVNze/0eSeC22czICi8K+NCSKSCxtGZ
8XwaF5/z5FXpy6jJI1bNg5CgZMf9esJ2lmBzp0gYNSsow/Qk2THGWH5m5/XAiFzcAJXByjYoseYs
TYBVsuBVN5ZufkbbETp2kFu5jk1b8Nf8XOl/kTNi68LiwNU8l0Scwa2gj/bFTtv/A2YRvbV+brZ6
v0IuJyob48rdA9JVbuIuV9FPw3GfN/+dfP07Oa98n7GIui0LmwQf683EzSzrsQidtWXMWS01wXdU
Dzf9yZ/sDLrYphWuwULmBE8ljeno3m9/xImIiH+1J9nYWpOhyP7i0aFddsZSwQvLlPDTcB/61a0e
tgn9yC010rVAN+qBHLklx/hLdvCO5VDJ+ApAgaXRaNH9WZmrgdNxSNpo/P7S7zBR6Gcw7A7YZsq+
S0pTEMgsCagVAEFIfudyGtaGCgK8wLdGVRUT2Ct5v5T4LTY0J630HwH0/aw6RG287cUpzENKtDwB
TUiqRB8UOiWTGVq0PIwTyYoFgOxX+diwm/Oq9ZXoePja/ZnYa9Ri8Rh+223jeNSyALPFjkL62hiP
l5P6lSWbyjqnuYZ05qqHZon7WnCIQHzm/nsVTuenAIfJO2q2p0AAOksQqk4PKfDsNpwQ3HrX2QBL
SS9C95mpoL8ohlyw0R5N5EWB75GrGJFCZ/4kG98MzBXoK9Fr44Lx8DQmins9ce4vpiazNPJwNZCJ
1QwomBOHkuuxDV9Rs0PgHlskq5EN7CX7CdsS+UoLR2lAaMyCRiaN/yNXBeQWn+82RZnZr++3GnDX
sR6lNJ10FKne7tpvnsIA6xoeE8oflt4/i76iM4fh8Qm8zzIvKSJxkzBo5N9RgvocV/jxuLUDlpJp
wV8ePdKmurf6jIstlNSjHDdarWyZn6Cgf0/bFkynxCZpSlHd/4qb/NLNJeAVw1z48FsPlMo7YV45
oU5QO1xs6ddIRZ6/nuQeOfqMvKWyuaS1O9MwJnyMOQU76i8wfqy/R4GiyzqZBLj7C4KbB75G7feO
jxQRGzL2SUbT2zBDlXbahjcBUcjK0CozNGoU1EIvvre64jsspYig7hfwHoBaX0maPecfTqpBDj+b
UuGPrqdz+n9t0RYROl9xM9ITibReD4ucqWsAuFbK3T4aTqj9HTt8adNPDQ8fJb1bt+g3621wnLC+
6jyINMsPe5XMnW4mzthGHjbwCluxWl2iRhFHl5lV4qNKAXvD/akeMO79kPQl5E5uSexviAe/4vyd
BoGivanaw0P1IHSmLscabW32seTgCl/356J933CIhRP2wYbPQLVOK46l9f/W0LLaNVfMPVVtR99+
NYpWxrayCk5UY0BWUvyvOypdnicAvJKQoOdSyCHIuCQe/hCIGx2nMPFe1/8mrTrx+JuVP8nUjZ1S
Yd8WtgckdLmnjflwdJgVhx4psLIyxZalFUmpc2szF+WKPDIQw5ehJj2FfHLloW3fJzKRRcuabK94
DIrBuQbcmPKbbXaie6P6PYfvPrfynIAZJWZLqpKUQMZAyyPR1I1UKYw6I3FywIOwoq/4eY6eZtNo
Sc5MaYSDy5W/SgTZBv+IgfQrGLFFV/UioHNi0xcOsoAha0+zmi5B6lk06KtPkIIsQUVYy/JaexZB
FiWmEYAMwU0kucI764KvANBqyM8u/0lC9jo+wSWF3hbd9ORCvqQ16KkerZkgArWS/FRmMBH0Vlzf
4kprLsK3ehUfprZdjKeNNEtCP4ss3FlkAxSiQsrwnwhwami/mhL/L3Cxr3YJkAogMF9dhoatOaft
+cUzcB4lAC5od+pr+6odcAYq7qqs/Ig146+qpdG0nJudvwXXwzpaoc9ESXdcXIqkVHKADJfgZyWs
UeyGcuHqtQmB32QtUP/FeH4UCn+4N1b3+/67dSJL4lF0QRMf2ZGcLnrK14a6UntlvvgW6D3xuvVZ
/qQiaff1TCqEAS6aXKoAKVR3YA8Q/WmwCNQ7s1Kznvpfc6tJ+IJ5KECJqqq+AxRCoPqmnZq6yLjL
cKs4tcn0niPHSxVh1O6xIl6ytK702qnbRqtuwXdKQXbStPDz23VCMPzq554Y523ziW/FmIB1TrNG
8ldnynU5lExy9QxxAnOiJT0OigFDfd8C56vqADzo7aspTJOAuU3CiJhvlgiUAbu4bK2efa95dEI8
4HjUV69QdOGgFWxYbndh7CN4P6SQlNvomkLlBIveSS9hm4VquCKMxhgMljG4piafvWgUmdURRTdc
zmuOqT+w43cJrSXNij5MvkVwiu2QRpC1WPOyFwDHLVUteNwWyoM7FokAGLKMN/ixZ0SrpOxXM1vH
/mvxUAhIIJ3XBVq3R4uj2yDKWQONZHn6j7WKp9Yp4Dt0uqNbp6gQmkTXNXrsV6dayFGo0wFpT0WR
4JTXtdKQOaq1G4j59oChOMLoJDA2hByUVbWMTaMGOo8VYNr2sOmTCSdccDJVQUSd+2qyfal9ADOT
RFwdXiPavffkpfwBMkFVEHCWdNRclzxgkeGmav1z7OW9DsqcZAGkcogc1PaEOCV4Ik9IUExXBR98
ph1anpbr03VQAbbNIQ2gW9xurd8mzcNleVklY2HkninACzhzqHdvODREpGQ0hprGqv3rK3sy6VZd
ndAenP4jvEA264NaGdogXaJrSyK1V0Cc/DaUTSucL8S9UytLclId/EO2nwOlulO1NCX3Ru2Ohf0p
WJBS9fqSJfQjz1kUnEpVD5yMebibx7h0wr3sFARyd9EIXVymrYdnEm0Jd9FjAlSXO0bEQeQ6Fhwv
9z5K8xVDKYTUVuJQG/kIy9kcoIYVpKry7CoifK2vq3JZYiKQw27+/rONtISWymnSFlCxqObRRuII
SFC+OBKwf5RWZS8IazacX8LC+CYqRuvAfZWitttCdsbz4WOpb5BambqFtq4dS/6b5SnuPo7xpGps
wb8yebtvnVyXW23CVz07gxYHRum6ieYM23ZH86pzyIExXtUAyD6JNrPewCiHwuoKlwZ5hGu2Y2UL
fdtlPyNYeYotHNHnbNXJ2vHXq141eIsdn926h5XWCh3IP2J4G1W/Ccx9llwfP6txxdSycwKZMIr1
hMQ41ATgTcY4kTDPLQzJHFhvfN98zq6veNX4WUOpVuPF++BH9K4KANvmkCqteyJFJ+A1u/sd6+Ok
gAzUpXIZmxQkNtB8hVENJtnkbwQjbrVd1kCXTexhIzgYJdmsh943ebkGBEXcNRk0iSGYD+DobgDp
IJj7+rX5FHW7QRYqhboWg+KsB+macPy6UFL/lSIrxrwGYNgrLdlwNSlYFYHqSFR8aEgWvuEyeUi6
k7kMwBChSAri4DMrjvy3yBfBWROVZpJ6eHa44y/Ux591CzDbcthIfMsRTMzwPzwjS8REY2mJJhl/
bvQqON8NsJPljSFS12iIwn6z93hsK16heA1qfEo3DkVd4ja/8PhIA5IW7yerkCiPFicKXE8Z6gIF
XjTMMB3WLaojMSIpJYIn1AcyihPFGXquulsRciGNrBpOuo88k2HM2xRs8DHmzX57zwyqOa+NMivv
xA/R/eJV8XA7+F+Drl/37pp96nHI+MG9HijB+txEuUlLQMjaz8G9tnN6HOP02zvNAAHxQQms7c/R
+v4+7DtSX9qei3AgAsU7J/LXk46Co1FMZKjC+kKI9Etx8bWCKMgexqXm5QEbYkb1G2QacZlkubgC
G8eD8/Qc0O4DRBWLUVW0QiZgyjfY2EMi04ULaUyJHtdkywaQOhViL+ddf3xrtBolW+wlQ4SySqP1
ZiuQ9raJiGWya6Na0bcbjQf+yiCbJuK0xou2cD2rU84Bj3H8atq2G6JYzmmgmMyG0Otbz7T5Npye
sa9lEQUqXhBSVo7c1ixXKKva7OPAta3LyKA5KwNHVj0sU8Vk26GYWJRllQ1VBvdMB9uZvW0EIgNg
njaxGKzOHkk6gsUHm4MdWtvHg0pWRDnCm8xZmAL2ruJHLETs6A0jdO9gGQX+H1R+o7G9NooS+VUY
EeBBk/xRjsnYU149PEAOQzMf8rNIM51POxi+qfqVroFuhUpDHdo5i/5tgaoa+QwgYLrhsjzLLBgy
3Bh4B7BZ/xeFcnWELEVt41j8eaV5Wby4SN1JA84QDC+q3sz9aXROcrm2AaTbJtCzw1NP/n2kiNMh
i3lwp4X355qXSbECat7RMg0J9aSmJsAGCEDHnVElmm7IrdBOeoUQdK5Ub0SnoPzooor4NvlXb0Sq
FMWaVbvjwimSl1TX6f7b0dy2ar2g4OH8YgakVBJeq5e/oKe7lKRgwwBrnejEorC0NfwiDcnaJyHG
fE5ttle4PSB+9OhkKuIYpcI+RRmoLl+ZrOhtgPmJa+ufnErDIxUxLUdmjEYxKim40MLbVRWo6Naw
zfy5DKOw5xflGRjh6drUS4T88+7FgChBQItvln7SYv717q9PvfKeCCSNgc071SSKupQ//5m1jJ3E
03TB8YW63jyudDpuUmhe847EvvXvidLPRoeQ2VeB4UtczTAqh5b5gadcln9qFnR+IV5jmPKir04i
BVxjXIcJPhBzWwi9GwrKl/AEqneVpbmBc/SqwLugxRYf/rG/CbkAK7vdz1su+XmoS5vBQabCmJqO
y8WmJeiJ65p3cIFmkL+vawhXdGSHeB4YkLxysBTTJSUEC7DaihwxOrjvXcs6uqtiRCp43AHscpUR
tTto0VLRtXdrYNYzEQYKbvI4I3YN5EZi0shhwPZik0Cz4pKhtvgU0C65DT3vYiCFwagjtGUOoS1f
6CGP9hVawRcDeTuE6vzUmsoJFe6fc3skA1eDpZ16U1+ZDKxFbbtOwQEENlawK83zS6eIimAiXkgK
I+BBSw/xtEldWA4BJujgvsrAqRzaJDvxngUN24PV4f0o96eiE39ZNPQoKeP7Ja9mqeTTAMJaWC8l
+2SWoLFalkmOi59k0L0x/pQGwryOan+9uQRS+8mgt1zBIehchSsRTgri+JGuqekTDSlJ3fe37PCp
6DyXT2vwC52UwftHX1wl9tunYac3TWyP0Slj9aLn0vjV3B9bIsb4xoJG1M+93vRGgm75VUbXmh+d
IKBb1A4NBO8U3a8tFL9+2mu3SUjKZRMccOopO/6cj4vJfGOZhHPbWZm3laotrxYjDtcb/GY2fSFo
OegQEJ+J79CR2X+rYlNrrWPtvXsFqAsY1do5c68YcuAIbZRjjEFZqCQqofryfO4hGhY7HyznLSDy
KJTbOC+IiACu8sxRDNx7p4UMA+USxTsSwfmk5EMs7meTMxfxeWP84uAW4emHOW0PRySrXjuvXf0w
19StnOhAIj7km2n0opVxP86FdYc0t0Gb5lHiStdiNAArRdePbk5MqhbzoApz+2BI4VM+tFoP8T7T
TBmiHlNeVZ/b7ei/CRQB3+4CCMEs/bUGw27xfW1tsv1EgxFJMUUdOzENhQ5lKoYmq9h2jUdYpozw
IEr0nwoNQCQNgc5dJyDKBWYzxyl1qOybNkjEXmd41Ad+C+0mjYrp1rpP9DlomWagQH7POJk5srnj
XHCbqaZw/hqTSQRB0FiFnIUpahaVV8r1e/E7LdEo+CKCe3f0/H2HQRFeJqal3XeHuIrpcvOqc6+s
bzJ+q2xwtv5xDPFfTPilcEiTOU0kWmZ/7ebI6ZD+1TIcFI2p4dLvJx381M4tSZ6+gcV6eaEXZ3Ak
Dp9irTDT9Zw56wnTY6IINRNsqLN5EUWXNkc+eoEjcgpCjQ/aKb6QXqrR9eODHajNSUxYLKERaiob
Qq72sSJPKgzLBxRySJpe4WLaJA3XKSfYJZzrKvXfveYNXRMDQu2adsPxQxRm5InnjLRNIivQFVFr
qqqXPeiSA3xN08KUtBV5M3BeDsn5EZNtYRkDgmxVooXCCLjN4G71mcp0Vi0NRr6GushHcE0R3R3J
BUJjQ7CZT4aOBBZyELcYpLRIeVJv7im87mTQCNch07p2WzmnYxGLQOSwMu+YcfYQfQgOcAqpbNj2
v/mjBnHYsgJgGUy5PbAg8hOYlrT+HCOtoDQSMIRIyN2IO/it/qoHN7gQSRpSIrei4dK4TRMEVmG/
ejVp4XacWt6Q/ykNPsRIdW46nJ+zG0ycLWj8PIEsA6kzMPIFhrb1VnZYxsmf/dz6A1uwE+Jb6MH1
9YXYVTLIEL03F/TrhW/F1t1u0LQpg/FhOZLbhHpdln9YsRGZZgUfY9zNcLoTNXXCKQsLWjgt2h4P
axnPJQYfpPsvGcQrOFYEyYjFHMYlVLcojLdMCNJ83xGO/VZTd36mJGZOefLQrK671u+62RmIMcMF
vZ4MS1+j4JbTEkLhVETx085kk5mSKiMuj7wC9m2F3L+rLOWBIDnYwF4/OzHV9vaIR2lTZoaoJ01U
rVcJXYiSm9YGktCrhdvlKvrduCC40zDILdnoaCzZMfqrBy6B+uJe/QDllqpfZxZu/KG7tQoxB7nw
w/r1r4hEYfCc/8XTLKSpEFhwSrqlkmaBkFYZhIADx/Q7ZVy0MwjTMqZNGMiUXtKvXDvX6BWnq9+x
9906/DCCnSzJB4E7fGoCyL4dJm8T7OwvXlyIluYQMcwmzg9mSohYVrDkDgNQ9GtnFNMuZKD4GSxO
NKiXGavPM5WEncLttLR+3I1KbiDRO8Do5l+oTzJay6Riv9pM5AqvEjLFCYBwOEh4Sm+2oXS9zj07
w5wZVZUV1TsIETIPzA1REckXHwFziAaFAT++NssflojDmaoeuvu5w58/bQg9soHBPdfrY85tF5WU
iLPAeQaKRb35pMxxj+TQpxx6gj3HG6duiajYBzt048q1I8s8+KRqKpA6tpnR6GrzHX+uLAkF/+bY
w/pbqAqHZU5RfAqPTDmkBiA8Fsfdc8j4bq2XxVp4YCLAOdfhHQ5ZhhK7uHTxruhd6ne13qkFy0bp
ddo+2BFIPmKRbG/ov0wqsveuFfyofZ0PdY9ojZ1kNdAkBuVmTdVxEmlePaJn1GKMDnQad2mCWD9W
hm6QDwXwJ+jQS5XZ2qbEL++4CpU0tkaJfWWKYYp4KYB5vrYEPGuo31tftnEeZrl753USAU/+jRMp
j1hsB6XkKF8WdnxdE0LSa/q4ngC2Es3rIFE+cKK+XGnEBMhNXh7UJK27i0YIXQjee4XC4+x4M4GW
EC94fCudzSX9Oe5w4a1tNWim0TK1usWRafU3vH68p0VymlKyEhObdkLcsXknzSYbqJ+MChuKinVz
+1w0VESaQKejYpVzhFtwMTqGsJzYKh7EpgtgkBnePbBJ+wPj6E5gWAdtuEdVWUQmel4K+cskrkhg
YzE/qRQ/oy0UjytY2F8JOA66KQ0JlGvDJK7y1FHy4ZCoCLwnoxIXd4bThfuaxevt2ausVfWtt/AE
ItVbKeOcEtfyi15g35oUfVEgpt1ai/sASCbHyCjjasfS2UL4kWCY2SiVRmaRVux7NvvaCKmbFGxL
eMhR8EXBtKQdXfqkaW2whZR0GMr7RCVYr9Ez3tZc4WT2fWT4it/AA04ASY4ZveyIRww6GkCejKl0
6mqyUGAvBR7JnQuHCXm7PejesfF27xKXdhZqgdx07yT+UhKynzMQJVyOL/YH5JmIjoL/gUz/wp9N
SqrBAHJydUSpQVw8C1xVuZS/3+afslWcFDAqQ7IvfEJ9qm16manBiPBwQutTh5uE/ATrIrR7PUfx
46cnb+D/K5pMB8/pnmOaeO5cHIz21EZWTA0k9SuKnShFdVANVZfe+hhRrnfg+/pOYU4q71xvJdfN
EF2KfDf2DggIJJM+XH0wpoo2KerpXZD1osJtbwDAEXATfb56anbIZNm+RkUKHeh2N1g4ZLwQEhJK
hECKlf347uleGsR9R25VGqzfmiSH9i8wtSLY5rGCYcdveLQS2Qw7FmYn14ol+sQjzajuoldiZRzU
47gDWnTXSMTxyoWBtumwRNmzRR71YJewjy+suRiiqy61tmwa4EiqEPhIBZ+fOv1OuQRUIAFI9D0F
TBVS3I9P8HVcx8dbQw9gK/zbfSVGQ6LO5FF4Dti+YwufaqIU3Cmw3UFtp/HuovxiLB2lIR9c5/64
hQYZX/qtoHFSbNcZp8v113Ik2dM28jqJzst+udO+kC6SvSUV/yEBkOWB5Y+l2yNWepmFkf2ahl22
OnIH0ClheBfvkChqrICnyXCR1XkLqtRzqyVJ2BnkvvTgKQMW9EsreBX8jYWxaXQuVCybe+e68COY
x9F6vrE9sBwv/MhwRzzO6ToYyGTPWRqwlELJVkzqYHvxC0CLWHTQCNg8oem2yTQ82SMZv0N7CxLm
SRrx17uDCvp71XfZllpPpLMcji0rPhplYzhEJ03ly+xMVklJZzBtjGKwUv03R9jQECxv2Z+nF0Ug
fE1kQWlPgJ9CItYgsqq1NwrItefYk/sGKOhexC6nU6puEiK0/NAzBoT6D3xg4DZBdlH5J0tck2xW
85spWRFzxcaXYXGiXpQeFxxLeWFedtMFiCbnaygcxtkF9iJAICddtEB9ZsL7+1xTCUEe1cPPF579
LC5zOLLmLmTndefE7affjTSaxVOyg2IkEyg60WFIntEY5agsoxqxiz+SFWyRZbw4yYj1hyKNoz2l
NIjYB/dBzqzEthRDkc9QCMPtcYvkLJD41fDTnoFGg2zvWRObvE6oRbZm3qtsz/hbR8w849GdioJO
9u/T1hxxs2jy7FTfNqYhho7qIWQFlH41lw0T/CnJkaOZsH6S1uXgTLd944mN4JjzBThy4zmYY+ob
WGtnTwIpJQ31sr2RA7E3Uy8sZkfFwAcPgzUz641svnby755BXT0W1DJFZZHC5yiRAHr2fBfwYInc
Tft77xdZsrL31iNO31jvhU5cNQjAaLC95mLStHCI+VmKTvYK8tYN2UgiMC3VPOaIYPNSMosNuggK
z0WSGgM4AgE+geB7sMHYIuxFIiIHgks0pp2S/3Tf07P0PrjBlWykUII3BPvVjA8jKZVdt97oxARH
OjQtgQ6hXDnuP9ezb937Ke7EHzhIu0X3n81uyg2N1U21PWr+786eSj+2zwdEW2KQ4Q86lZOEGDXO
Z3YkyZypp6/hyCIaJxst8h1N3rSlouWysJuj5eAUrqb71hhrqG9LrIq8xdGNJAncFhDPDjrP24hw
uNHkLbpq5ELqXnD6b7JWa5icE58DbsmDTOn2uouw8NXso1V+tDC8Vxv/8v0djUdWxulyoN8t2pIM
b3XrgJjYR8SyPaqZqX0Y2FJDynvss3bYlRchTdh5pmUJoxRAyRTZay4aUMIy0kSiFe4GkKVhSRVd
Wy3ERQffylLm3FLgfVE3IxyZaVeJ0SVKytuEMBmzcrJBMzkmnvqt0tBHwaKfCVo0r9K6A2odaKoA
0DzGKBZVXTXmX2bkAjWJRpdGibdSvpC03go9IlTw/gL7tQPnANaYteQmyCwel73JQXuGUtu5GvEo
Xs+J4RSXvllTnVrFBj2jLx+0mbMu/kv1dDte7v0AZjq0mEOd1uqfYTtPhT9ObEeKHoElzr0u525z
3f75mOSugilhN8cne6c3Hw9tAyS3Pqi2/OnLdPF0TiuqV+yVSW4emfNmCH2ljwJSYLZgw64e3C+z
6E8Mlyty2iOhzDO+kmSDExOQWtTLi7sHaPTnropy35p0ChmlcZjcCYzQwEcJGE6jmFUe4DMEeKWF
71qLA4Slu8V9s9w7rZCh9h9RMXm4jzZiw3G1mWCgGdRSGXujk/T0fZyt40BSUOy94CPAnioHpQqF
Hn6QeIUY3esh3hebfxUp4KUFpWkdFVsyu7UpytSkwuu8QFIAB4aeXj4l99DSA7khs1LRqtuhZNux
X+Ztkx9EaqaoZni6wlVJqDh9P5eu6gjXscsjcX1VYlciN0C7hGEGlfFVMGKB2KZu3aREKGyUBkub
wjl5FAdPh1u11lFBOpMPjgdfpnuj0HYK756NbE8Dt0r4FVgSrPZrGecYpiskj2zlWHUViNHV7jTe
aHJ6qTqxMYviKZUahu+1bacE9X80lOKHKSAuGNpTc0fDtx6IK1/Uodtq+4GMbt13WcbD4kSyvQM0
YN3TO9T3RIi0yFQOhJ4A30yr+jEKGjTjxgjNvT7lNZ29A5V9Oux6sd/PiuLrjNq9g90DzKeSjGkb
srRB/amBLkju3U9Wjn9W8YL440ZrL0bHALRi8PGWLdxMgfQiG0lJltDdr9+EOrMYelsF4/XnCx77
FVtloSo73B1D1/q3u9ST4WyUahHmLu/yWfgAGbIFPcJWCx/luw17QwmMlqjphm900Njw+TkhhSaX
Z0145hIz+aC/7/x7YXE0YbL2aZ3khbL519t2TGK1qVu0y5u+ehlsWio6Ylo7cR8uEOeI1/lV7rqQ
VQeQykiWqfSDNlcu4Q26CK7oi1I1BEeLHi9HQj4empl56V3mvA3wyON1A+ciKOZI7D7Bg3QDyDx/
TMeo07s32eje7DwTxpNkPPXvC/F/dI4Sdl1ME4KGPNCI02CQ4FTUph82nqjV/o3cfOb0RzQ0IjoB
94DJLuTvQ2G+v0XOWmpnoI/+OzFNOr0FA/x2uVwNNS+OJlx1cpYOP+zl8WUzU9Z1X+jfZP0/zTnJ
iFBpYzgoh78yuQvSm18ljTL08OTKh6O1o3wUgfCzPeiJaZzY1x2er/352f9Y/qW8Jgy2nEcDzmn2
Tonoo84KdyXadHTtqFViu1i6UjHeJ+KLNkQg7puI++opQkS3zF71O5Nra8j7t96Dd+3ueHE59anS
L8GYtheONFM135OzAI8etlS+eTg/rrsNYM7+UnmHSvYMZFoBsJzxcxrYR63vYIpbG5zzsLdn9ToK
sO3/pjV7E0byvdZ7d0IqxGRVq8Ayknkx5Z6k11xbM4y/LRDf0gAwMz0ILZRDs5ii1vvokFEzB27e
2+WxyqoegS5eJEjG2ZxgdvV9GH1/XkxjlTq3niakwcXJ3ka+3V16IVhITik0XConsYBxEiZDcS5+
TsKZ09wWCcBMu9epQbMAkQ+pBDXoeLm7Df1kcwB9Uo/WJT7yMpkXJJqpWrPrLBw2N1Qd2BKHUSVW
NVLABTZE7SPq69k57skzxJC2iqhPhhJ46NTPzq9KIT7QqjOSh0/Goj5wYdmqskcnE5W/I8WxOaqb
rl501CX6a9ccEXqUigUlDNCQeAWz9Ftivvj6hbXSg1IuzcBhVigyFCaaqwe8LgwDMR1dIfFFgZSH
F7DEC5g/er4MF1+wiHPe8nNQgDo8m/1InsASrvM8TT/xlw0tXI63Hyx92TdwZsk/VK715pIhcxwE
PwnQVstZd7S6ADVqxqdn9aDZK5xAzy2SnW+ZHPb8ukzVgugETCKMOvi4VXWkOv1jgUuScbw2Q3Bj
ZRgQN5b7a2iCqMAiw6NOThERgApCIO6B0nfC80L0+TA18jmZyC8UvFFgNRVl3gA0UPRbf7jIDJIO
TUJTdBBWOE1XJg5kOutBdo0FIQz2xua+wH7OrHb2vL310/ZUC/Eiu+17MlMAHVFBcFYyDahjdt4K
39tPYV9lWnIm3swMJ9Lb/nnDsQQViyBu32Uo1S8OfKnWAUg9El6O4uiNpiTJaQWMgb3sCwB9cunH
dnaCZBWK7kP+6vzoUnFEREoO4+pxmHwqeDai5Rgij0JtMo3Q4MMSXX1y771tbLP5r4Eh9vpYFfqk
w49P+/9/c4HiWDVCM2k/OJ6cSpNNjqYGZnFT3v0P4PaFwl2dEXzQGPJXfgQGugl2YUkZn8SAiNeP
e3yJn+tmPkGHTBuZ3n2LZu5pbicm4/odKvV2a265CiGZ6EBUzIzvsq0uVXvIOBHnFAA3aEYDMLzW
2FRHOPNB1DGLJj+/Bz0TMt82vBtwmMzCEUmIB6etO0WEOKzxjpKQ2AMDnz79emVEa7PTASMIKV7X
whXWkY07xKnbIZ85wSSYvS6MWL9rw19OVx9SSZ5uUOs1AkK4ZgcCzMK6aNTYDNY0tiCN53p9UrJR
uH7yDa1xrfaEJnULiADjmoTeC9MaJfOZbFRmKskw9IUruyYXOgs6kH35/t2g+KSPXIb3hnFzvvSH
FSxfpwM9m85CpmXyt9+RFDkH97+b8bFHH/X8K1rTGVDtYXdZLiCxzapEthqLCggygRfbLcyJZRls
VdItJInzeRI59jVBJEQ83Z08EBTAm4q31G7vfDclvOnDC9L9ovIAhsnrzLl/yRvpCxGJ3orkrNRU
HU/Bx2mK3o/4k/U38VOw7U4LDi0Qta0fEdfvyubPgE1kqPRSS6z7d0gVg2vlRXIstHRFHAOaeAEw
t7bOSKGLjzXF2g7tdB5E1VFgCIka07iL8Tsj86EiCPUay9Egyb/aFNeF5XrJTOiosvWJNkmfzcoJ
vrnw347J+5Q59Jbu646a1eDjAnzJD4t6MmOjyyiIBtI88ZnJlUQ0AUhGTkoQWhLDyFmQmdjoUQ/m
kFRHpyHpHzb53DRBpGyVBMNeS9z5YhRWgmXLiYI3zes/VrHI1np61gdwNe87ZrVdd/DtCj0+8mSA
R9PQ5wLjOKNQF01vfVnjGm8z1iw2nzyPsi/qXxhIJBow+lFBNCcK+3IJ+mHGCRNOMpM4FcZtzp9C
FYg+BRhY4oOamkL510XB/ExKP7o21d8bLo1edhqSn2vZTzPEd0YzIg30k3Yw8SpuotyA+T/de/Oh
s5Mj4gFkyL69O13JUntpv4XMVw61TYyVwrt6+9n4Oom6nbuy/AAXw3xj464kOcqFHXNt5qVpE54x
pDD+sRWEZE6+Xt4CtJfYmxkyhICU4cSFFYW35WYe0M38n/Rl6WGn8HoglCcXblS9tTWSxwWiQEUm
fd9Puuo15V9/fsTi4DVD9+O1SSyDQ2L5sl2oNzFulhrPou1pdUEXxKThvnZyfWGyH6V0mWPgUGJN
x7d7BZHDPPpU0NDccAM5kCxaO31m7j4IR+gB0/+8aEQAMcyZ7Yo3S+TeYzdgImWE7afGgl2jTu96
94CKxtTnHZFjRzGnRKUB3vfXfntYhZwCD6E8764ITLYhtTyPFL0YU2jr0/04Da23dVZo3q09whSF
bFzPHWMXUuy3Drz2RXIJXoMgaZgM0xa1rx0QkEKJcFxP7qLhrame7JBsau076bBTSnB7MqA3Npxs
O8iDhsj/YMw8Uj/u+jkIZDZs35OPp4jpQYd+E1OBLOKeO19Z6ffKqxtTCovF0YgIM1qUn4dPkkXP
AsPCKFPxba0909YfBRmHH9ygpBacfBWNWaJhkupvJkcVaIt/TguWS+HbuxEFQ3G42CUTLBradIKw
uFW4pzv6G9hfmEn3lmWcYP3J5xyFyToTlH3MyWy6I0o6S46ZwfQ8W/3QOvxZVMZudOxP9X35TKvw
lzq2ERXmU+X8HwzmhBCUO8BTc8u7LAk9RQ/iH75107QU+GKoXwSXUMu8uIlQreJ9w9RnDZIIsm5O
Yk3tHGX1hL+koheU3qnJ4bsqtTz2C4dMsaoiOIJHY80Yq7HCnZs0LRkwD0I9pqjI2BvhWCpcFVKc
cgB/vrCgEfjX0NZ9gCt2UOkbw2R31nXJsOCZPXlrjEE2cYR8bQ5uKunJBGbyUDFyVqT9OxjTAJUB
hnWL0lVgf9du8yB1i1oWBIII4JPIMfKRrllH9swWXTLorMDw215lIgZDYWBMJAHWjM9AJXJcHCSC
cingpISSfc/2DH8jgWCyHtbZ02JHIBPEJ0flzQAMBxcWV4phODSQ2t5RndlIn8pjoQzABll9mkZu
8a0dS26RQyVOq0nj/IK4OVMDsv4hiffHrQPIQAMs3lvT9Bkf7KwlD3WBb5bcUPfkgmLtBDV+/A/r
KpLkxo6LlCQQCPM7apaMaAeP89iwGqysD5+OC8xSy50FMFFdtFxh0XBD9dDx8fZm7CfmIkuGRVpe
fvqJon+c4VB56a0XVIJ5mxyctTRFzPoePZPQliLlsli58e5suCoE/QtNAb9rVMJ5piABBgAFQtEX
Q6X7eWhxUvkJSoFhgiFRT++vxHf/Fg8ohdrpGFR7DFcx/ugt10hq7oP3SbkG6W7IU10ZdUE=
`protect end_protected

