

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
oYYUZ0MeKqJUJoI7DJiuvSB+q5Ix+Iwj9N3EwG3d9aznfrZuw1+Fc2PVy4cVNiksbh9EhD023m7N
/1rZI7UBsA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BmgMGlUziZwp4Aeom40PM0gFb+Lk4HIg7NJ8Ke6/iR/nzJgqwxvBOYZHlsOO/Hp8XOgAeNb9Zd4o
mPFcvStSgKrLqxBJrTC4jOtTOOUVOGECik9X7RElVDiKeZuCTuuYfKks1rnTANMNKsXOPeJj6Svr
YyXA9D2NRP6YkUNuPRY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
1jtnTjcMZBAylJ3gewlkrSdkM4rrC/SF7w+2Gpl8C9SK/D8Tzq+D0qrZVMnmX2MWMKbqqYu6bkIj
sy7Xox+kttnLUyhBRsrBNs6gr3T0xsxsJ7Gnyco/P3Bde80gstdJ+PNfjg9uJOXa0R4ym9WtfNGf
swawtPDRNO3XB4oPqX/YBORxc12Z2+Xzlc5kJQDf1WM1UoKUm0j7+JBzjmig2WrmokL853BM29jT
4Ht91JL1B2bOy9A+fEpZnVLxL5NzuQ9svrSJluHfL94vaMxePXlPq6InH4B+XQp0TAFlIitjElNz
4mBAF7U6zb9GPz8ite7f9+Ofg2sCbTc7qhRaHA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gQeqr96ZiBT2MmGHCpbhB9Ma/ONapmaS0FJH16GFlg7E/VRDUjqbqiiC9oovpVsOBnNDQZNmXNgv
dI/YoLxA/mPd3NXizDTj33SvvwJdHC+sPFJrC6pT5rNUHqY3WkLW4EktYj3xtwACazlM0R3H+N1W
ZL2jtTv4hCIZZw83DISHIwGMevxP0unAXWFpAlJTyOmzC5wsjnlwvjA6I18++KC1ECVIFCC+grSL
XEAA1xdZCU131f12m2UaGi1yGaQH3scoEe37TXsoGUkWCMAn3jD7PddNt1X5zhoSRxPsOfUDmtSO
kCNVtrnPznMY8kVS/SdMToJlnwH2sKbHJZ6YoQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aYbz66wynlNa4RYsWnE11uoqAUkMOGD1rK3oC0qHnHAmOdMhPdz4cV/CAQENwbN3ryQY7/k4qEBR
2l3bOqYxA0+CBRl+jt8CXXxWU8WE2qwf32lPVes4/pVAbKANmE02/Ysj4IR7MGLvUvtr934XOsBK
cCc/KqvEbWgnnzkEdl16nzyz9Je6iY7Ni836+/z9BA/OYPszoNI5lKgO/06ni9esrcL9aCuvKXjM
Vplsu70i86fjOGURYjM2YFmCk8Xng1M6ROF+0KD+TufNMvK1W5if6MPJr/BsB83OF/hzcDKyULpB
p2+Eliq8StuhC0n7jUXEo6ZGATEY2a8DWEYVhQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
B8e2xR5DNyjb6SEEOPCOnfB9/yUC8O8izWpzVz5s4/hfcHkvr1SHS13gqMQDj1DN3uSpaoGxcSIv
a3uLHDL4nIDztAAEPOvl5rp/eCLKhGUauWJKGzgIaInIPCBXw0hsptiyzlIicQEO3rsxoS+LR4e9
ltN4asLfvR5i5+Aru5E=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o08P3wLx4KXr1Q02DiaLH2vPxf0H1jXIwF3rbwsiMxYgYGWIJGF4/mxUFC7J/WeIjcsQFoTUns3o
ZlNZWWRR36HJ1r2GmZoMunV8HAWjNjCUrk6RBWvB/4dYllizQVzRhb+3YUjmiSEMr4rkGsWsR9/t
W+i6luLQskwMDbMnn7puINFUehSDaOzDytgvFigNs9cj7haJi7XjPeMPUBa/JbbTJGFnxz8xzl03
55+BSHF5m9JHUn2eN7uDkExSgYolpcYI1EQnoCH8U6Zfcweg7A+n5SfklkTKUeWInYHoz9tHbIHA
y9aJwNoT7f6uxEt4GVf7oKjEfFlxUe/yajXHuw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 132672)
`protect data_block
5EA5e+7eoltHbXWw3KRYLbaKaZMS2W8yIyZM3gMKf7QJwRko6++T/04ckZ0owBxWtBoO8rzErcx+
NRzXLhME858Tj9AGBbMAwplsfESGnKSghicDaB2xJ/vNPCpaw4iD2qSvlR1ojfpDdci6W1PkZMd1
70/770RzcpqR0Px+lW85P8e3NyOZUVXOoWjsLYGgY5sXtdkweMeG8UTojm/XV0Y+8vzklr6m/AKk
UaEFyEHaGvUGJrgG+i5uDdwTQSwgmAmPgELe9l9bYrelkYldctywoo2PUSKpyQ3c7LM9nbZ0RCu7
DGjwuex81w6oG83iXIBt5YtOv5xo6GLUGFEwXSDPIskoSaA67/R29wDNsCJWcNNU/AZKWENhm1Um
d0hO46tA4/P/sRf2BiZOGUzqT16orveWjYBmOhzSqR8vkpIdJWN5zoRSbhGs/CYtnxVp04p4jdz+
2waYlPPpGO1EHvqewR//n9MmtqyKWbPDF1Upu8jP9fh9/LwNFxKFBr6OILwSvTkXwjB/Nvb2ckRf
G3xymLtj5dELn+czF0k40Ffx1WHoINoIa7PbjKaOSu7/1Xetb9VRy171ryYfp3bu2gkCqoi1MXdD
tw6x5QjbdDv0ee05Uh3fVf6aNbnoefal5ODVKyQ5iOHbMmRTCNmRod2Ma1M4VE3sNK6jfXxaIZPK
Br7Uu9dppWE6vbMAqKR8IVpeVpbSqWHhmw676KDA4zAuyDyZpsIDhpLogcLftCrlr5HywZ5nZdSj
GhKulmyIYsS6bwrHS7avWexiNeWxc+aA3X8OWrp8fQC7vO3s1Ol94TmxMw+2aRfLQ47U2f/E7vl3
bcr0u2ADTNJt2XEDhCGuaVpqAp8Aa/fRvGUYM4VP29pDXlpwjS6t+ONi9A3vq1Yx/OirXdriIOGa
EzNvz+fHbhvOsRJoJRd4TVz6ejmoH5qurS1elMr3FSGxKww/NbzZZACVRCjV4D2UUdhvGE+C6VFp
WqehjikVqvnClRZ3/kPHMREIDlU/0KTSjU59aJ3n3l+5X5jkTaHeGmm6nrPCWI5R6FS8DGcT5Qzp
Ni7ZsnGfRMq9G3ppq7WHuxo5fxntZM3XWKcD+VAKBDjhGSlPE76C3ZdmU+L7OXOk81Xu29RFDwNG
lTx71EOKwHepgKERcdjufLaAv19tKWVcvZeLz1hOeiYt15oNC/eHEAWT2XLKG0383tnAVLPpA3gT
bXQwv11EGFkXNYfYOHvCyk+oEz4IJCyObBbSifwrIqC+IiHaVlJufFw0+2GujZqH22q/SJPQ1IlA
mJS+FIoC8ljqadp9YZuJXKuC+LRdUidyygPgkLpGrT0Sd0ev+oR2h7Sdngazm+bfSKnUkyX7ixuY
HWiw7eVaInmQZAOOHbZz5Gta9YELNvVUJ0Ubh2Ngg7sDs9ZYKsnbYKVyFymoKPIn5iys0AtRNhqR
1wF+n81otn3eVqLkPmrR3qFrQA/LQvTQYTgowDR2eTLZ3TFa9bwC53dB72hjHzagcDOlfuCO8O3/
DzTG4lnYJKk3xWpanDxUVjs43oJkn8I6GDW6L8rpnRWvSwqiMehqDr2EY6pNyPsigOyNdfvshlWn
NOGHHK0slMyc76nv9LPdcI2xogAqaqEcEWBwnHReI5QlF0J7vNLApPjsFmr4xH7/op2bdPclhe6Y
nGwTcb/2+cbsNhcvQLV8hpfhUjISfjv873YfrCnHpcOLjfVj1irfotFkPK3WZoyY4iivX/EPnSPS
q0wo2EYnPq210NvNeHjnVr6vQmImWl9XDyPpakvhB/mnxh9cobLri18/s4/HKJhoFpQXRCL0cl7q
dPNTiXRYx3Oiu3pbKPuMVkX1/46ObX4Jdyx3THFBJJ0IGYW+gl/DdYY/Hl+Q3Am+cZu68l8ecyPC
DuaMaErV66mLuvLggd3RG01rDBg2l1UfkMWQdhGOC1+P+N5d8Z9/Et9oKfySeckC2iCEFmLm5zhe
gUaWe81YinnGzWoRcPZf+rbOn6xVS5oeMZfrIeVpBUnkkOSr71KhMSQypF2nSsaLa47+PQepvWmv
BKK1wg9O7rM+CoQzc8xnQSl8ePtxxQcDxgDcsVYmepbuBT0tc1ehEXaW/bBOT/iFbbSLexUMeWqq
zKNw6dmgqpRGg+8JPCJI24KhjVcODvgyqfR5AYf7rGEesdt0/wU0ylylwCXwAYq3OjG4dEqk5Im3
5n8w9r/w2DRZPENiwBZkJld4b3AY7/9aLVjLRSLq3z837T963BEp2D0ci75Hq5grSlBUyY+SeqPH
M0icvG5962osc8p9GNTJ4W5pGrQRVzZHIMqWVLwUiz8NaHx02D9ymis/Qsw2dP9mUGIl2EzmJGsF
wvcEkASyTlUTkF/RzwoklpME6sPYGVkClzdo1j8nU6txoEgnUEwU5V3RIN6beclLnWrQOGDVEPpo
YUPfx5V0QOCXbuF/UkKniMQDTMRY6rr6x08G3uFv5pI9DCJWxSACG186u8n27X97HQis9xTu2iGJ
SKYClFOxn6OCGQygOLljwIZ/OWo/DBB0yximil8z+BdZ2Diymm5WOBp7nq1INTD0SWWfjHHhJyc5
SAgtAbjkuNd3uqEnnZah1bHWy0Bmx2dIotTWxH/NrSFK0xBlpd4ZltRw8DnWNgQKhtuMiJ5HWpII
3ZsHs4XJc3cyXVelmIfWKE5RH76ijZ2tKMJ6RlEK6EhWWHcOLiWWEaiRHfUzncWS0u8cKkdLoDdb
GcJKvmyPW3kwBIIpUDWNQ/WId+eI20KLY6/2Nexz7n+jTc/F6NjWDgF/7WRQofK2N0sgQOfDnZvZ
CTqo/8T6dRGVL8lJrTtmrTLyWfSj4AIO68kgvs1XzRFviWYy5Y4uoAqwCqi/NG8j2zDgAPxKEAsZ
8Qn+yAKz0gDpgDVqI5Ldfb0BWL6j7oTg10FMPcUnPU+PZq8p9SF2TF0BTaXGFaFT2UizKeiMIc6o
M+KFENoHguPnwfc26eAZd47gEZJ62/kE9Vkg/vSrUqXuyScQGezS6kIhhWEv5MaYR9FI86z4TTpI
MzCWWq01omXT5pK0m+dto/QcCSRl9rT25GjJyyJ0Q7X/wAlVMu7ayUsgju7UbJVztE8UT8sy02/6
H0SXxWjHOLsiUm0id7CUDj1IxnigGY2/AH3j/8MGTUYwPQWVZSgMdc4ycWkW1CzWdMihSkOkubQ3
v4jREhVs5BaRjezrhPnttd+nabKx/aMcKy/uz41PZyIpG7qBjAhbFL6DHVDlELskgOO6BylQEDxQ
kA7AdJUQlhSByH5Va23Zyk95tXgN41p+qclwzyPNR7T3m0aI1Ik9HiYz+yuUoACkElekko6DXR8O
BjayluIEoCz9WHFgePX410fc6I4yUlleOypMw4xMnHCXSS7t1KPOBM5pwnKBMkVZfPZMVfGJyxFb
ojvQbp6oPHOG6opPMNKEQN/kHmqTLfy6qW3IAnEPiP6+9Kx3l7cLxlIYomMCi52pqSjswBJ25u0u
Vd/b91aIcoyaltbqyZgeKVOEO9r939MHEsTlpsYU3wqDEpVpVzlyWcydLU6ihc/QkKQj5vM5ywJu
wuAnMFSatlqJ0we/KD+f1BSlJW7EFjoeGRfpSni0hLzn/YAzRSRpOlVsYF602pD3vZr79EhM/Ekp
bZV0dC2VaHaDxScstdlitNAXYohgIrKWut2g+CnFn20cDPfuF/7tVHna9zsL06/rYD5cy/MF4aGb
NFREeiCP883SJjIvJh0Cn6155L446g/eBJY9H3x/BfQq+ch8oTbOaamRLohhOWV1kkxGqOQpOOrd
wBbLCcGd1eyJsIXwBNDhatyZVOQAirAl/BJCPs0ez9DEa+HHzU8/+5uj4RrVcmQe6Y52Q/+RdxQL
oeeznkPd08x5YMVcFncbC64RkTPkw7Dg9GWCdIQwbFRjHoHzJDWsdXe9Rf3ppQ0wKOBTlpPN3OX1
r+d3SEATpB/YH9cXLBgVWxotUhToEqG2cTfukpm71zMSp9YP9UsGhbKAOXJFZ7HGa/s6rfTQhy07
ULpXkqCM7GEZTeXve8SdEgLSpuorEr3HrOnCaPPtT99VoRnGLJWqZMuN3Z+SeG12CY+znVzuXO9u
7CtyCQHyzrKKi0u7Jmv2VFiBxqTAOagk5uRjFZvZlwr5z2rOWSFiiR0GmbY+U+z2XHKeMmTa8fbW
ni5NiUfKKy68aS+SCOIVfxZSwYUCQl8/Sv46RwBk8wxyaevU3XQAbmRWK8dTGIqGA8PWbYQM3Bei
BRRJCzx4WpQWmF/lq9yKCj8dCNQ5Q5SIWQt8Hnp2SKeufTy8+v/qv/UC/K9ocKuIYJxC8QGLyM1S
LdAgRGi26UK8NPMHyK/2I9mrPmHnBVF40ZNMHS2XVDJtMR5Yr+bKxQYpGyK3ZsIH6PqrMfe/OOnI
GJj5qBwbi9d5PP+DtVZ2iP/zAG7duYG9VteRPkxUY7nOa6D6iDoxJqBzQ6fCybItM4sttp56Nt7u
l4yDeETdVhnnc3syMbuKJ6EkBxWgEkDraJ05HmPWTGtJCiBsRZflT2myESxKVeRcZNFGcsccYhvz
/L36T9aL4wpLuRFnKNOXHsmUiHKPrGpfsEoQkVdFaKgySQyLRpvb94sf+77GjFyVPcFTK7rmdls3
7o3wyoNgMcXK8Yed1g5fV8WQgWZX/1iBjBDAazq42uUq7r+TlDGVk6wYqrdrqBHCvdypD2PEL4pm
qaXLObUlVhU4RVTAsS8q0NJO5Cx/8f9/sBU3ETLPPp9GJNu+8R06STJCyuUZiZ5cOCB2b74cj9HB
bohGWyHpOeWbk6lmn8Toj0ogVf6jxXj3I93Cj6Dj7llDVVhraG7fByB07zUXqYMZZqmvIi0aB3oE
0bVdfE011L/RKuUECk6HhgUX/5X3ksQqUOcCu08LWm1GsQWqVv8NM4Fvpcfs6m76yEEHZlI96O/v
jJaKqy7xTc685vqN9sBGlKywE+dcCjt9X5V+4p5Y/4fLuCN+iANMGecoYD464lasiKDNEoQgTl9i
2pzC4mnflESv2RNvt607RVwIYpggox2ytErdrBXaLPJOkDLm+Tent49alphYfCqV532RSX6r+BBu
vTmXj+HcipZ327Q5SRtdJpDmERk/VZatlo8kqnGzY+Ij+glxepQzSu4AqhCullR2eVdPeopdGSiP
pLr8ERLjlbGlzPNsmQXAvOAxoP5WCJaUS4YY3rYYp0fyW72nPzSV2p2qfNTh4gwYogieZOD8Le8w
7ypkBVEI2DRSh2FsJV1641JmFa05uuL85+NvsbvBe914N7Z1r3gwdNhxFKrpa9S8uKcwg3Dt2E6o
CD1KmK55FXW8PIdGFBHI6fOYD5bnOdrWnOXuSfs4MKeY/iKoKnDJzJzuFdvx1JpY7UY7847bw8ix
mJN6fcoQHKYYmhBkv7ny+I40ohCJIYfgrq/HZApkd40m1wwYfzRroRb2N4KA1RLujgXikIBnyA+y
jf1MKseOjMxCxKhkzohfHZ8f2+uSdl+Kz8IHwlTbsc0qWBVtnE/ihESqsJoXD4IoLvdsGSB2X4yT
UG6A6Nw8uwPBwvxvWDNeufkMpOXhmUiZFA4aFu8V7gC3rkJUpQXNWMnFOS3etZgRhQlvw5U8lA3z
KF+XWyg5Z+7HEW7Om4gLHj0HAqcRys2McAHUPztrXA4DrHo8WIB/eL428GYaqz0h456wMEB630OF
KlrTvD8zZymk8xSubRM9gFCN3CUQ8isWXYD27gdc0GwA0A7VZ+05BrvWO0hCsjrmbz7PYXsqE2pc
CzIlmvguT1OxWSwP9nBqLb8n3NzSxX/0VSloUv0tzl8NilPeB2MbH+/WjCoREVugFmkeWZaJz8FM
VlDEyEX559VriKJP0XOy1Te74Agv6jfYD4IrY2EzQ5f5wTVgoHm8MnP9rQJQ6x/C8c9ArUUvw4F+
KStf876scG9wR6f0+vp9LT0obt7e3aOspZuo5Y2NSHk7K7BpYWUuG8TemOgeUvQF90gd3fkytDDp
srQ40imWOQevLkVF5dKj6Xafka+B0anL9X9Wo8rySnSwdfPZOocY9xtZTu6wKipOYZnVmGfLB0mk
ICdo7LjknZBnGXH6i87ZaPGXZ4o6iGD73q3wuCFQBg9aA9/R8+dcAhrpCtHVb3ynDDz80XHobtFv
mNvqfkbteUZSQxBFnSNIZiPjCdPcx0iR+jCPcys4xVve2oFXCp8S0B44LHbUEFHJnrShz/HX4A6B
kBhz/rE3bq1OOtTjeCwy9X5gnSqXoMVWu7t8FXRqeni/YJMVaSXKdD0Whlvcf6SKigkF/SEPV4Fz
k4IHbEtVp5WbLnHXE2/zSZUlVPcLr5U7ajeFaco+AwCZoTAD1OhFv0K2B4UzF+Hy6xYmtXSbeZER
a3oA828BExdLPtxuS1cVeLWWfYHYxYJoFTX7rr2oyjROqoyEd9sglCGlKUPOhPqhEiHif6AvPAZm
Adkf8aJO7f9WZ28A8zoxubazbaXDpdCN6FRw/w9pgeawecz6uLuFhSKl3Oi53gY9ND1sIzC6TuqE
YIuMBqxVVp+VpsD/sY07VlDCsMBVZzX6rMj5x03z+ILSL0DXya4lha3nQEp0CQ+NhL7JadOlQ7LS
mMXP0CmzvUZ8awFJkVuV/uKOzOpZqwZKOyNKj1Vrg/FWhhFZOn2NJgrHkRMRHS+Tlcm78K/nLdjp
wa2I3s9QxQeyY4hsQTTc5/+/AxjkgQMo66dx2+gnp2UjfBF3WrDe0WwLr6ed3s+xP5zkFuFav6mB
ylD0nxYGZ1J2apF8AKItlN/kBUBG1Gt1zz3T5ZvmjWpKubGWYINDuolxIFYbycC1dKwr+sHj0MB6
wtLjQxfMIKY7tiVTnNywBC/CLELunMt4/KKtW1ZGG5hJSNZzaLPmeh8TNNxoJHvOBx7ANGmdvBJ7
vNcSfAN8C2u/m8zDc+RB6q0NEQdAoR9+EqqhNwCPENT6yX58DTsTwQ/Wx1qC8mTR5k8q+zhdKJi4
7B5+/0XFHqVtaUMuOB+CyFqUtqm+TqFsAGD3ad3sFqpJgR1YqjJqIzOJ9i9X4OAA+o92kXSCi0xD
N1GIClFWRxLDTJJW/vyC7gLMVC2CJ9F+T6jnr+qFtbfbXmU1cSg8bK+qlow/px/Q5dkQod90s8Cw
qBmTdm9djz9jjg/3xHX6fjADD4XJhj0CShsl9NFN5rKejjeeL73S8w7tjDEHw1ovlKi6byq/A/PF
+RI428vYSwe/eiVbJq6RxX+Jrnt2X1zTYCye4omwHYiz7g4yPMoYTEbOncn0S/YUY0RQLZ+JD+GJ
KQfzP1ibSPRcW0/DcZfnhZoFAdvDEzYQio98sEl4npI51Rb6ziBffGj0nY8ulUXN7m0eYz4vq+5E
qmZJ+SLJvDkJYMFNDBK+HionOqN13a8EgltEFwBaJ82EqjVlvPjh33LPIR/dlhPOYffl5U6u0PDl
Exu0/rBKsvb/LFdjmPbvOLvsjJ723qw/rkoYrT31RxpLhE9I6jgD5+aMlVABo35WItXTbRCYXH2Q
sI2RnB58g0uofRVjDQIdaliySxfhfRogJ4bQJqu8NHzAKxK5RWRrOjRoPMM1mLjdOBuujIaQXl09
34Za2p856t7bCV/UVzUp5qvW6+pFqgEOdN+7UmqSfqS/Q62t8JlnDNceJF+VZTGnHu/CLj+8k3Qc
VkFWd/L8v5brl26DfnAR/u1DR8Q/GvEYl5BKJfSOqPY1dLNY1FgHnNp2Nfs6Zeusmz36CsjSj9fQ
arkDnf4LfvnMrBcFhOt+5K3R843TQ5Os5mGIvErpyttlaTjseBnpnzwVSr0EYrDYVVqmpura7d5q
8Cws+V/F6lCzm/MYu/f59uOLpTOp9+U9rw5gPy5J/ZBaP1GAuYhQesqRCpQC7J87DaXQc3EdIXcZ
khRVsw3yzKPPQq3Up1+xdbBLk38DYRjTntsI63lnkL7na2Kluu9JNt0Dn6VvWtgDz3fBZDR9tn0y
PZZ7BvDEf8P7i8rruZ5XicjaZiiW6cL8z+8/64iw6bt2HPidIOepWeBIv+ysrODTdpwJWG5oRACD
5fikawWnpT5eZ5R4XkM/0B8pd8+D56ibXZuvGPd3PGngr/9dq1tkevTKSkJV+U8k+BxC93fn+5q1
jV7zTyZyDBYxhgDZ+DHbLIFg12UVNl45iJ5tP5sju96NiQaRvuw4wbyyxlTeOS/L3ybOOrl+2uYX
uQRBavPXwZTKBuP0IhDzX843bpij93lpSXDg6v/vt9q1udqpUoONOhUqSjdph1HDxWd9bUzmRDqd
Ri5HPoG5cl3+kKDZAEq34kY+qpQ0YepAvN7bQ0z9XFMQEU0JaO+5f9bzuzg9HjmfPHC0Oc6iY4WN
8KEt2t4yJ3l0m/O5LoMlbPZ3h/eEzW0P3aPf3gW92/Nr5Xml18+hY0pQNnVTEsZBVE8V2jokd1LU
Ey4KRUkOXxzJIBEirO/0kdjbMrC7n3Vx6VwWZWxvDlvYVNA4/poEy/mMDfFF8D41bUeockuEqcPC
H19Io8+wpgNOBhVoup9YcvH3pbrzPsgWD4Q5Ms54sS9v5Ywu9DAMPbNj5bHG4ZhhqM5k2iRP3lko
vXwfcHl7p7q1KLW4WMAVvih500IqAIBeaFO5fFiMi+YTUNkK5tufzCG9u0eNBBliA5K28f//PkpO
y8xarXDZqi8IuVeLfB2UzdjlMuje2W91naIvDu7g/sNye6rbo95X5iR1vvRa317F8g3MXJZt5ft3
I5tR7MbToiLKFG9Vy38Za6JhQk8FbRBZCXjQwYubmpgaTPuezy0frRR8NGWphGbNYmdt0Zf7/jTP
taHY1XyWEgXL7oLLEkU8V2Jtw2DLZ2mVgOTHwT74QBsGoTLoGx9NuIXIj2i7/Bkdlr8eS128zDl4
iVETV2mgPMc7R5x68dwMHgB2hAjIfbNz9oMn3mlR9rxY01HBYpS1sQ5Hal4Axff/CTxh8J2jKOXe
rTNbq/wsNHCcBKtNL5S/EvvlAu/5w51D8Q2IsMxo/DMhe7H8KefE7apuCf4JiE3UVxvGSE9snS0n
5rvMyhmioJmPKJt5BfBbkEkmh8crpFNs9c9lNmMOJBoX5UmHKOcfGKRQzFos5BMasSOw22na8yj0
jpVZqWlNMnrNpm89dLMkn9V8j8nZ4gQ2lsIomnz2jgEMyZ7G1ScsOdcJ3QKwGlRcMze7WFQWBgr7
7AhzneGGIvUx0V2JdLOi8SdehYwJ4fbOCPJ6B9JgRMNRwKBFRkn3BJ/EU431QNrTCuxPwMul54C9
ZrGjQ0bH4ZxjbR3u2cSWS3X4DvnrQcoW8DjPi/7exJH7uAH+5MdAmilCBBITHjKAM5+iz53SQygk
OXZRv3I9REV799JhlLaT13H3RosUMCoGIu57MnNYdc0rjhmqL24OS3gi9Xe2JSZbPUJvJCCCrauz
Z81ToKwcEDa6SAugsU9gO2AAanZdycX9avF4TfX1Ekabq1iohZAkzUlNzej9W0EdZU7/l1EcohDN
4u6b7DxO4Zp9wSPgjv7jDhVEYvCkRdqcw4PuA2koMHoTt7plEPLWLrve7/hxLzXS9Xy4Ti25e89g
GmGhRSCKMH0FGJabdgMuc9RLXhx4WhUa8LLvWwk/4Am3zZTHo869C2J6n5nFZ699M59zs0CtTEfd
b355XLVefGw6ajG8hu5w4ZgmemJal2PWvSUaad11ardcDIQ84+wVyXMQX+vkAfrXlk8VzBSUon2Q
vpscA5/3T58Cpj0TZYcQPMiQ4bAnpBLyeQokl/ecolON0TqzhDYUb2LavTjElFYKX/cOJjUV0Dgh
ucvZwMreSzqV0kZl/Nov11KgNnYBjkhx5Cc4vBsBkYDeNRupC9yDaWCttcVoLc5AdaxCMofp0kV1
iXBYtMHyEI5+5DYA3ktLWC7zi4wQDo4h6/43sJxkjocdvNXtPn955AgyVtycNDMLqrZSok1Yll59
i6+fvr1gsldvmNjytxDxWJlP7UaBQKdlOuioUXfRJJ9JyzTQy606Dd/VpHRrsPhJmKKBZBIfHLGL
eLH3pwSBfH1u+tnuJ8Ih2VbUYNdUmUk3KWoF00Q0NowFr4FVb5aF5toJFuExtJRJ2XQZ7AK7BLur
hVwjzirXJMrKuPg9sE+wO3gQWNQdCR0BxUubQZwfy1a2CC/9BsPLIN55/dp9ppgVqFNYe1tS7NqI
WHspkpzMJiuWRrcfOz+V97xQb0JbebdKYNWbKSP5kmFIj6nrRRk1Fb98a0RAKUP8pwaBoT6pVn4X
7hhm9M53N2vFZhBtJLC6euhV+CJqH6KypnxFiw00Aae6y1uQfgRWTKkztD5U/LccgOGAWX+R0iUt
RSsVAMV8M6RGMKCbDcZxk5mUCA0ZAA2bqhkZq+4H8DiBYe5sy7RTMvWGTRsiMU6Py18WIJCR2J4L
3MFqrYFuyYPMwfpiqHU2p+ybCRTqP4dBbG9Rnnr6mcbEy21HES6wW9IIuqjF/atwChu/VwZTNMzd
IhPbn6nxisAqEt+5bI/Rd71KI+U6Q2kG1Fof4JouGXfucDRgA1o4lgb348bbhlWoKEnmhyBaEixw
8IW8cPQ4i9F4zP5hXCAZJ8EMEXBBlIWF71loXGSOHjmifeGy4/sIyvuBM60dDG+JKwbE9IPDOtwn
cLJYPKKFx/z+4uteTNHOAv6C/qLsjetgbHowXiRCorEub19Xa+inp/pB/qoEuuNm2fu1rQkeIy/3
z4XC1PJIqXVmLgzHC+yFTbqA9JnzSSQpJRR6Dtx/cHp4XICEUn/xfi2m4/l1LSwSF8LwrJ7/EtL1
ofTDgEOB96lGgrnOEtiAFK4e91uqyw37gc+9cJgg/7J5w2ApyGmTTQz2ZqT/f5iw34QrFWGqDkEz
UANLZ30DQhB/kGRX2QKu52wSOtfwwDc4w/YGtnTHe2nZ88XclPIvELOOr3X+T8i4aiqLhapYQ3Lg
5TCu0WJbeKGFZteK5teXfhymYyAkZ7UNQJDZkG2bSlJ+DHomserifT8v78MmrVHfUTHIX59b/wK7
ECUuLMyOoW1mNZ73kFInghVTUGUi9qhZWHu4If8YP0mUSfCn4m5j/CfF3lt6o27gOlsifGEhu4nS
R4D8IPki5+2XoAz44HrYlXPHCBJf3EEemVluFNSI4/Zax8tWB1A27TTGtXjhyfn/X0nRvuVPxR//
mnRU2fM1Ct57Gu/RaH7jVzw4X+eYa0IcADcUoq3kFEH1SVQKBx+8pzKeuFoAsljPIlKAurCLzlaf
7GZjZM3EwidVfMYp6D9JwYBXKY5fdr45iGSOJZrNrM9s3+yxd5O2PzvE8Nf5m6Xb82QVCF1gCUs2
wT7h7MU8WPzv+Whg0eze2qUwAFV8Z5OsJWYH86HskKkU7Ir5AKltmhKKUp3HsjxdYiTG7IkdZb0X
8BihzVaXMYCYQo/4kF2cf8EBau5bTjF2xlQKcjK7wq3KunJPR2d/iaLozBvFIXmT+O2lgoQXTbbR
X9AvUc+WHqAP3PtVHGDKNZVNv9LYNq/jnBATiRqbBhgOVdGKWeNG8eZuzrK0i/Q2qpq2JSKA9gg2
NQyd5VNI9Zi7Ktduxjd6Xj0Zyk0b6BbGLRQPsLB1rwGR16f9vF+WSymZi9yt9djHIsj1u8Wq0ZwX
mgEthVEacykN2kzuDsYWj9HAOm3EmKTOSkfZDm7zsl/i3OrhHVXp2erRPynWlfAK9G83SYmjJAzW
6FND2lek//0BY/rUevykgkl4AKZKsVBtbujdln9fy54ElDgISRWU0+UjmySu6QmDV2z4AQBtwoRj
7CJilPmTB/P4/TlfDTUNLT8bXcrfdBVnypyUbkxMIcgeQL66JMhqu3Er1qh8MzipDM3dQVr30fJ8
b9Q3HMotxbYVmdB63Bm4EEqee7DxuXcWnW3p622Vkrn/wo9HnolzIb91JDaSmLzhkFxRR2pGC6kw
8f/FxgziaM1xrMLELOVayPRTcBNZEQBat+qPCcgq59I3SPW/i/PCu2nSsttvpkNARoTKKjDtpNnM
Q4LFPa0us7sYBw/EOtqsp40thEjR+2sRAJ1keKCQz0db7IV6AlFJ3IlWOH9LJv1a1O5G2nmZqN6U
y+0OAH5YG4R9ofiKw6KUj2g5qxCnVkjGNVgHA4PAXXqgOd1dUh0SSQWxvBtfQt6kkNLqVSSKqJW2
xHFOyaVczqX3MvSVq41W2QhPDcZjHa0E5AiTSvEcfdNTqz44FdNF9/ydctLQAPdDCDV9IfdnULKN
UAG2/HcfDdPw9cNrPlQ+gFMm91s3ESx40hZbb99lFAyaoQ1QmDmosZ6bJDkI4o5g2aYxIo8ulel4
MWnEQ5Lx+Fhd8r0mCt0RnxhUTAaBCwGrB8oIyAOL/8phx2Uy14nCN6zYh1F7cZen2AT4YNR19Mhq
9VwVXlB+ZspFVq1o7UcxxoBNSJeXGsWynLo2hjhy5lYX1atcGquK6OyBQh/5fJ5K7xWCuwOmW618
mz87OwTCS4dKw79rPTRn/7f5k66PDpvBwCGt/YawziWlrEfNe9FHoxbJL3uN4Z9Ry1wKEnXm5A+P
iY3jKLGmNK5Omm6ebsFUj/0qGB7guQIc6AhRQ0037VJ9kjYIX94rRaDOq/JvXuWXsU1xjvEHJPPT
esLnMR9cWZl5NJ8QwhxGVPe+9f/I8HqBGnghs1J4SVssHL3Df7KHmWCJhRrRd705x9zlW1ao3dbj
ALY/jK8DnCHQthkdR/6YTILOenIT2VnJqIHhiY8FRYnyM7WKJs0/YxNRHv9DUMqMZB91rPDFEq6U
v1nj4Jc7ajUyotimXGv2d7RRJWG8c7SCGLnE6NRlHVLdnOBJTeWGZzlEWdB9QhwRJNqLM4RHvy6y
1+V6t+WAR7xhy4JO4ijXtjL8a5nrXPHeTs8hYZsUJXZes37+Nc+6SYfQ9r36K0xInx8T3LmANUIW
JI0R7qNV+5NmWZpaqIFB1Pk6j2ZdBGZOWngKGT+XDHX8f4UIoi3O8KchxhkNXyD8uyKgTpivIbar
Q9dpPzYrNnv6x1UB2rRMvF/Bdg1QqMfX4vi36qkHPv9omDy5rQJl4OQVskIzDVmtleVk7v14m0pb
gfpVwfBbApr8n/dJHMBmgCM6tuzlZ/qQuz0NwWzwJVtn7/Pv5I6o35TGl6buCPGIIvMNqlLzlMoD
JUVqKoNvhZDgGxJsAa+9Qme5xhHOT/mkuK0gm6GXx+USYv7mbQfNX+7pMBGoWyMGIzYI+uhkOUJL
6wK/ZzZR0Jhp43XPCTU7qlGhcKq+Y++RjZUWgNO4PDV5qpZtuNtFhCyUpsh+PtszofWhL5Y3srAY
wfWHbKwDFUndp5tnr0VEjCGYaMmsYNzDuxoz6YbKGRvdRbCEJLurt7gK8QQVX+OrAFDgqznijSHP
UAP/NQrEjs9QdkUsThKP3bBdUqa/insdKNd75N6kFBrdHckLXOTW3GOAAD2Z2wutDXVnsQMAX0jK
CLYylMsyR33Sw1Ty8GLq03PdopvzfP8hxJ4eEB/wnNsifIm0IlUMRqIxakdZV2OWTEKFm626Ornt
TQZoC/5eyCl+x8e8cpvowCalX3usYKuIBVGRz5xxjwYlKz2eEgeKPQ4dRA+5XLRJYgI3JahMiIUm
g9GKNrqjAp24oMSb1kKSNlb0GlB6ZtOtVKKBimIx0FVaS+SUcKhcnNGCZXNLupsTqXymeMSElrgb
IljftUKTgyp0KDRqYszfcY3UK/iNObWiAgHEmJ/ZAC6PgRPSnKNxmU6KBkKUHuHbAop3detpKbKl
nKyg8X8rOR2Df/nGjLh5KtgUFf6SxqTYNkITIJ0gRmt1uxkKbFTa1v4VelBe2gLf9Yu4UJeok94Q
utl+qIakdEpAfCixj5kraDPpt+d0/NNL2RyaO4uB4kqTNCNNEkKkcK7VRjUASGFGM7gGGLyfPUeM
9TQwOLngmNCkafGmZ6H4MqpQLCdSEDxJEYZ1pPrGsRkSUYFbGhAtQAxVhIGjyf1BKnKEZXhvfvxe
Bd0A08iWVdBMwm8s80X6s4BtfrbdUk2/F9YK5BZHeqoxdKzDIriJxsubWg7fcWDw6RE6oTRVIxFX
FE9NYRNbwz4FGGI6Z/1MgUeGH1NbCMS0SCRHHi/vAf41vpAlA2q3FzSDxa88pBmWz9z5ObqpdONf
Z5O2C+lpyPquTWfP5WXiEMtWWn4/26YwptFNuPWZkB86q0BninJRroprFGSzZ2tLOqMwh/Rp9gBO
K4LUAR0Z+kaggebVvBwroaqn/wSYb9iaMaWHsC/n21fbtRgGwfS5UqXrQPepiW8p3375tVxwzM1y
gy1qE7kloPsLyGgBZAkeppKQD2sI+wdA+ZDezEm00Jvcv5Vpy4mswXoeSXkQ/4DEi54Eo5zhqoAe
vjLKyBk9zfxsSKxEPVbrnqmmt4uVJC4zKFhgQlS1kjUnEgfMUEIygabn/RfHp3NnVc69KgovhAKp
W+IFEiWvrJ2Ns6+w0ypazLX9zbl3DRL4yM8G7BXLks0OUwzzJSvfSl4XnoG/3CGG3GXb0OFqcI/A
tPVS4B+BcZO3v+3/a4jEoWCvy17fXyK7WKJwoyTjAH3BZjYKZijAdwkBqgDK4lOEvKe4EjA5meD0
kQA08z5Pl6Fohk39dAyjoe4bMqMSEFkJXGGnS6MXH3a70+FJ9DLbv+r+t/8zonl7UgTkmbtQ1fJd
TUBu8s3dKjcYho4o2Ok/hmI3juXP/1KzGs0NvXSsgBH7q4T5bUWRIrO1uVq30Tw17EdJQcmUPZSH
zfbOpBQrJFPFwW//aulX6xKiEGPo/o9oK+bNwKisU2NqWfhs0wLG/hXYtxq182EwRWYdox0fuc5L
JUTarbi1ChykL6t//xCCO/OIJc51PafqoSJnePSxmd/uGutSzSfYmZ1CORZLFNj5IlWnk82POYSw
GjXvgHnzqf5GF809lj8RrZooU56CPWgqL9doazz23l9nXqbjrxfxJ+7wfOhc3XucWe4QBz2R4Coh
mNjM/XeWRNkGkIKtdi63jDw9VxxV6CTkROcemGqWW052A6J4eSnqaeXMGt537C18n+plz0Gs8fm6
O775MUMFVsCyl15pxbuUDVvGuwBdUlXM7OJaf61bZ2kegaVcqsZb4M0T2P66s4rCaIHeO3AskHYX
3kkFmTfRbj/PnaFmKpfUskobfi4PWmLR0xXpO8g/yJKe+UufW/JqpjNGdAlhoScsICZ7aAX1oyYA
vMRNsCZduwzlgf2wLYGjuat15YxSdyYUXtEv98HulOjbTv4YtXDcCEo12CnLDFMtM03PgfZmzfsU
nEiNGrQjLggbRQXOUi5tlfoDQ6chiDkGljZ7yws2V/h8zmSORifeg+2FGeATA9uf+5Qpd1nI+Cfz
F05mE9fAnV/Scs3djEYZHVhwewU7uXbc3pXCUTSZ6xU72mpOXEAtIcTkNGac4sEsw/5jLxyVbwqP
LJSwulG1vhVv6klgskeZqbtaKmuL2PMchpVno2f+z8eypbX6ste/0/n2n9kOkLFapvN0isg39xWl
M7g8/dFAR/v7bwzTeox9Rf+HiOIBiajho93yjAKFWu4gGfk+yxyxPZuk01A1MC5gWHDqfCwf4Eri
TmxzCnqnvEXoh++7qmya0/vN6QoCce03AVfU03tNd8kL1vHENOjBPMHwjVYYhmDK8ykdPGyuZrRQ
P4VyLMMYqUdQjvNoqVXdVHzHDg0SMG2xfYLbh7HOPPsrxpOTqRaYBrUscmdfx3lIZJ0fSIrFJCAc
CuAtEBLjwqFsfbNVlis4P+M2VmzlDuGNegFi928OnD2goObIqB2MyHF1wB4kwffHfWnOVQTjoQlI
P3q5iCd3xYwLpvz68udXXF8w8liVZ8TI9oDGsWFWoRmy7/qt2py3SfXeUhs4BmmjLxZYqVt6NJGX
OdMAU+LPIiwYCNFNWI1Fl3gXwR7mEWO3nP8iUsh/8RiDVMDcdf2kTK/94pQwZ10kcNHac6N5R7+0
B8hjqY1GPmFidjXB9NTolkFsjVwmOoTY876hygvfi8lXZxt6SrLSCbJBkkXb6H9AHfdoFJEi5ti5
M4j2yGFG2/qUSnayiKQ2U+VYERM2mOzbxlZr0rXltcLQvKgaQ7FD30jlKjz3Fl2Y0q2jco+5oPAw
6QJZhfZ/IqNt0AwiGmqG5xy6ma/qAIjOQIe4mdtfszZTAfKTHAuOupuVceX6jz6WreBlowL9mCIN
QAyRI1eWHC8sFr4WeiQpFmAWgsJPGIZ4s1Pk0bB7sCk+o2ZXgWloUc9wvzJpuupKjKl7LUXn+sAY
coFBRVBr9TgRlpSOpzFOmRk4HeKNTR1tShcKOALvsrwi8lo63pYA3LEO+pISvD17/qFf6Gbdacgn
E9IfS0PyCCVlayraQZOfOdTo8yQgd3A7M2l4VaQC8ZIP2ax7ENT3LDP7ZK2aHz2ZpkyeZz0Zf7Yk
ypPhnE+OesHkHU2YoDFL6xTXq5ackU9+GtDFnXIn746NenH0tvB0GoNuY+qX6VwzClQhm9R4zIew
0KTZ4figjuy5BuKDgFPLDoYPGvIHZmNBpkHNZfReT4sISuH4JrWV86mfwwHtUD/mVt9GKKC45oIk
0xvjWQfxMWy8ddDEpaU+l4qrNskiNGkw4abpdGNd8bYDrxULQkRssLptW1oh0azehnsaYanL2orH
Z899D6rMQRyZdKSBJBzBewrpNnNoYww6RRv41ophj5gH453/1hwh9VHhg/55Sgf9U4dqOQpjtmgw
0++Y9lchsERKuboMvy6njetnXu8RFJ7i8Y2/XOTqWfSkNuWz655hCLzkJBNpvyQoGq/f/AhsrgdM
RZ9zcKKPkUSpMaBH7wNlB2eOVlSRrtFE1iV/KFABp/6lMYdJyRCWXvAZs54R7vQUNDQAy+o2RU3G
io/3yMdj/JJZ0jbZ1Idum/8FJBFZbj5Ej3yrSv9yhMdWj7Vp4keO5I6aRBZ7pTPxUEee+lAWlWCe
d+dlF5C03/BrwpjsFH4jQhoA77ocbS5z2E8E7GDuti9XL3HfO+OO5JSj6oauqcNiLgYKoXmc2q8v
yYffPuJZ7rwrBtVtt4FgArm5cS71+S7G+tSvqRCdXi0FyThfhGCthqJ1MnBB07GlONoshPo5jg/W
8gc6feiqiWWXq8UNDG6EQdor3TD72gmjo8xJkSSXXY5VAM31XWyjTzA129ElxIYwqAF50C2rPE52
SBb8+9TNI+RoFEvdzTXE7adaOo02siNbPdm8BhuXq8swcKIvVph7gP0V7MXSo9bRAC9rzE8UXgOu
+kUTQn4vrMh2J7egdSZihgXieAdyex84uQ0kSDHJx4noRsdM0zh+o3R6t56f+23mofCgg+1q9IHs
ROk1NSIPS7URq6ifEoi9/237Qb9KWy9mTLdx1gMCyBh2XQmLB9gSpcPWX/9aCqFq2G0y3Rgg423k
5SQiB8yxSvYJud8uzzvuf6C5j1VmPE6TUWA/W8sLwdPz8JNmpXLPWLYrIGiB6UzMMdbhO74EtET1
O1np2a1H3o7lPOApDo7bfc1siFAs+6PubzNzMYrwnYzWpzipMXSyquPNDtnnyw2VaT5ZjJNe6BXz
ZjQQnBfZi5YqdTIU2IIKLGlhDp7tWHWv8IFzJ/6go8uPVTTxwadEd6YwjqBLtPRigylX2pHGiyb2
hlDRw5RhQmLaqqCwmG1KNnD39d8VbenQHRrSnk5etnPjS2FPTf1sv3pJ0STfvK0LmOoF1pqWIbbi
n5dwo1sLKdTuS2FDPf6cmOFhgz6bCd0O6hJ0Dg+Hr2rb3jfDHGGt0rgqZv7H8W5Y8Ha4BWWy4uYq
sAPRyOHWW2wz5Ym6ZdC9kWMu5SyplX0Ss9gP6/hmtFylBCf2I2lDHndyYBnOkTRe06PlfKH5EeqT
NdBLmvwsVJte8ROzl2TQS2RzcmHEXrX2F33kYY9Q1wlDUh512EaveIiaUVBDD4HkhwxJ4T/g76o5
uEiBFwRvpMZopPfRtQmtyXj64O67N3REcUrufPppiDSXo7cK6V76aLxgAFPQeowSO9+UvcngBUtJ
xpp+LgCXoy4mKPuVNSv9rq9BpG2nPOyvBnHj/gVhO7JdMIP4i0QxqAlM7ZQ6W45GzakIpbanMXeb
6k21gvJwWrBBblqRsPTP44971/LkIiG/H+aH4sB6GBpiGhI8OCddknBE8n3JW/ou7/vNKIzannC2
+o95qUIGCAGL3EcRURz2EfPkUpslceIyZpOS8UKrC1HmdFyUMiSICt1ehrTnR6gcyyRTfqJoSdDd
rhZMUn6dvXUowuPnVYmNcyvSV48mM+EIz5iSnDT1YUTLaQRlVe/tCKxKk3RFt9r4lvA3Uu8dEJrt
HvWlS8nmx4ZDFThRT2VZCfUWcCgcRiYd0SAA8RowTy8yR+jpVx6XeXrVmQviFPYEv+a9vLdAkVDz
VSVXB7J0r+5OHqGqN4nLxQJhbE9EbkscHgBChloE9Lb33rhBVi1eSB4ii+uOqL/K1UoM2gclXtmC
6EMv9MaE0lTAfscsixg0bm33X+DhGkCTeDucCYr/rf+vNaXej4FGN0p+ugfZsWyDuBjnGDOA+BlX
lsjaZCynqPwnVWLTaVCERwQkxHXTmTduQtUPiWrc/X+26BqQxUa9JPYqnsY3OE63UdG0TOw0Rx3v
rf26WHwCiuMo0wm+oZmcS+EhH0rPa1hu6ztu4J4ETLLiZ796KBUxt+EEGkLbhvd1/t1FYaQnbDHr
ycX32Gl9DQENHR0On7yaCTpYpHSUQCbIW8LB8/esXQvwhb6dXMo5nDVkCYiR1pWbv5y+h+ED7z6O
1Dx7hDWIrG/OHSsQQ0d7SWODAr4CcNiko4MLX0PBNvE2u8lIB+tzWbGeF++LftVQXRGNDUvTBm4L
33JxfKJaqBDs7ztjrQHFdQFT4kFm5fYRZryOEZk/g+HQOPXOWZLFrIMKPyzfjpl7PbWSkxFce3EC
7TPXbIEOJbTJ+NiNkunk8bWrgNnKhKPQAOnvVekLkHmDocXPL+S8DFFZ7xwKB3kkLKQmiXR5wYsC
2lR0cc6zPx7WygjCZ/2UIIa4s7eXtI7awRe03RQu0Q0jk5y0Rb1w2SXxPHn7vkOYVtsrjYB5g4Vk
PPRXli8uq4aWs7GlDRIDm5diN1pnU1v6fzFnDnnGoGUueDduxdg/VxCNrwYz3H62OyEmyM6Ehpzo
6WaywY18iMDFkuEZoKyKSzxtEbT+8xrgG5ManHBrITHGA32eI3MKBnLZ4k2S9H7Gxjp+k5ytfihB
BV3Wvj7gj74tpM71g5F6W0SlcqjsgrkPR+z7q/Q0rC7Xmt3r7vTa0Zq6pUDBTcmSLljLwgNqYCx6
msSljwy/iVVFv4Hehix0Doch1L/0v/ewainANbk9/2hIFHqtVrKFJiNb+B5hA8hCOj59v/WOBjc8
0cOiDmwp+5I0/o3Jdb/Fc89KC2cHgHKBr2bgGuzwcEGWReGJsFtDsR4pZkBVgfmq49dy2rFMqPg/
XqwY4yGughLVzuIPKeuT+clOX00yQi5cO9FLgCjjUfOoHkVTQmyUaXsY/0dBiD2qFahufEoYMCWU
XAnu6sTjLB7P8JQG+9ALsGZbUbxq77kK1Hi1wQWamhmzKwf6mKnmhdv7NwQcKfQYMK3NzvfWAq00
7V6YnOSVVxz/iTvMLSa8BKuiCYIHBAqYftf62HNhzqkHMpnCsIbiGGeV2Vtx0NWw/euxhSttKwNs
lXjOGA89Kkx/PI/S9PqxwjnAxIobGtSQpir7a88wdZEZZu1To9llJfMSAddT86Tz3+44/ejmDQKn
SP0qo4PdXvMKKRuQWGsxoTK1jzBe5DbIl+46LPvJjutDSwoN4NwrQFcIk3ks1PCQtGzDSpKt2Fn7
LHXzZkQ8rQEKz6iJOcDVthyvT6kFLqHvzKBoj/LY71FAR4f8ppKbQkJFXd1la5ffu6sHFZmuvCsC
NZ5MW3/iXFIlVFfJmIUYGqaSYPUTQuQdP6c/VOcl7G8gAsiGfaVawnJg6qMu9AQ0g+kDb7hfsbeP
P9BvWTO5IwW56LeHH8rdZ2WvlEPu09i0+kqz9s0Bo80GiHfwHGZsoHke95jb6DWKzOHmwo6Jlg+Z
7S1eRC9oUVdd9Tv3vDl/4pJ82AcKRaMAzYnqjpGJeWEL5HZI9NBze0Z4JFcSfqBf+FJsec1Ts2W0
FE/Rjnr/pdj1trWUvQEun6DymcYAo7l6Ib/DgjVahefqqr479D7NGAsBx0NmNZix6eaYqvX3RmHU
umoxizxJpdCTqCj46/kK1+SwPjvMheEFeSsNzpZ/nIms0JNY5eZtaYArcaTlpKJfDzTjmKPfX+Jv
w1lC67opLVryeE2vgZY+4vfPftMd6WBzlI5o57SopguhNNz+YT8qlDAvNg5gmXeF4Fp0/CNgIIHU
IY+r/2WOEAX5EvKmPJQQeg3UBTUiwiN0Z1PqL5Anx9Qol/yanPXb23HCzAYGyTMJIXBMUtPq45Hc
9i5MpcSO8YteqY0RdwCY/A6jE6B6zrSKPJRaTIR461yxh2uwhhtbTcdsQbKCblHzvATAdTjnaZHI
ILULIY7cF3yTAPaSWT1d+SOSdsjRQzF00ZwWcGcTY0lriOI+ha6SfKsgbevONOLK1/8n713uhhMC
6fOFvxqIs3rzw5qO7Ct0afSwcUng32pgvuVKx20l+vBpVSmiJNLreXJ6puxE6uDgjhDtYnsZ/9oC
PhSRDE3F69m141ouwoZmPM+k3Bxcvi6VF+WI8QHmqndYEgsidGBN72G0bP+ixrPiBB9ajEiPOy3E
imOg6jlsY3HUyH+jGk8YY9OlrYOTLZ8cV/JXHkVkCVURR5ZV8vxitVwxBrqKAulxomw4bgt8Y9Xv
kMO7qm7zJGXWVGYbAz70+Cx9oHWjroghGLaIMiqgqHm6GusUd5pwUXD3Eq6rjtoaigDogGrwlmbt
Z88XvYv0fSuW5MfSuOMeFz9T9XEiQsRbsT44RVZ00Hb/G6e54KkbIp/IKUGqgWJd0LB2diexmKWs
EXrgKIwDQw33mrxmDCKIMwUOrjQ9uhNTW0c/ptf3ApTknwqQ+tWw9vp/at5BZjeo6giTp4Py/5tB
GzY4dZPxGdjFCy9G5EzQkzxNmVraspqe2b2xcoBLI6J04+AQn3oAUb+08qi7G9dtOfWvu0MGL1Un
uuQz7PbYd0oQL7T0dw9Az2kqg/gkRD9q/rL5jnreHYXAOkCsWmkLnASLhyT5ww+D0u60lSWbIxxb
MPT41RJDYNMK2x+6d8X2q1DBL48tNUsQbY7+wnruOjTGMwT5mKRA6Ge62s9om3T0YZyMwUNuGVrK
VPRDTXC0oiDCZakriGkt4X+t994Ld06UUv2iQFHKRwFbHHc8RCj/GYdi1eQ51PJck4XfRjMQFuby
Z9PtQ8V6PArZwxA7Vrxqz6b3C1+wM2rcirtV+2aRf5+JDiJVex6qlhsMRAmWRU+HctESpfsCYvKw
2To6XBXbwiN6pDU+h9zZGLoHG9vEoVWMUm/ACLhsAsFhIpqIsquojxgAPGjo2sJTCvgw8ktzb58j
+w3Wzv5je9V5WfP73CSxuHQh794hCe8ZYCGFGMPdnw6AW6DbGMRoZhFifKzxGUAF0ZvI1c+l7Kf3
JL0nk/8shEKOm48Y7cbDLuJinnMKx2Q5mwx++DNIAji/oM4U648QzNm5mw8VvQ5NfP4oCxhR26Bc
/3sR0lF1jj308aUkL3V7jUu5M+aepGcG7mHfuSivEKZS/+m6L5h4B3YFnRt/aEyFjLzWIIrcQBWh
1MGKsPCMHuEdy1SyRjR2lF4oXpMW3t/WiCkwUz2NuJIYJVPiAxickP6dRJESktXF0nOSCHVPYWp2
e01feErZnf5ZQPAeWsoc9cJL8w+qysFUiG6dF2XDxnb21NmlcBt5dN6G00auUg2daEnvXsFwwHbx
Ey8wysexaPdy5KAPbs4qKeYJZsVe9j5gMvWLh2rBTZ6foP4FUGEuXh1EfmOeMcQA7T6cfF2G/GSR
uIdfZTRD6wIR9blh10Cj1EOR3cCHYJGshw9xhN8h2GzJiBGXSZJJWjOmwgKwvuPLruY3uUL77WzW
/F62uY+zA800im2+yHxMkZcpHk413/KQajSJcz2KgP3X6k5GuZFFJVp/5bAJgAKpFbcrHwvkmo1X
v7VwnpfqnAqvg0CxUX8vT9XnCeYgBElFjwIhyEoztL4PIt7HUHi4q+HUslEoRTcZCgF6es7Va8hA
eSUmwlfs0q/e4ex0Df7szfl6yl1//SrTJn48K9towgX1/5ggvK41aUbflK11GVk/hd2ftAL4AWkj
Rt3e811wcJOOguwG1du4C0SegNoxpPXL/u6W698YGKRBaqXAKG1Ypwk41tUjIZw4s+KI3ZGu6quf
x9DvqPOW8Hs7rch5ex9sqYV+UQhKYlZSQHEw2Rrpm9jLv6+07X5UZYZQALMjddcAAX5fv38EWOr5
2lCpvlW1rrhp7O0glwGLUaKUp5mq/HSnq3mHRI/2JgMOMif3LQXaO+/8iKxeUbHtr6w3XLkDCrxA
BDtlpZhHJz4NHPL8eow13dSjJ64XVUBNK7sfU9mOzavXkJ7STe8PKsaK6BXg0hCP53SS7AVz360p
lAps1Xr4m+InXAgfI7O+/MYXRTa35Fzam9qZXI+/UhKyiOpZlYFT78bWoYQnn0t5VE/uW4P0zi+j
zEWeQUpGL/v4QvWV8q+l3fZIvXhRtK82hchFrb2dsNTd6l1utH4oadDjWYAHS5hfsqtWKUno1NUn
thTLnCfJYPb5wob87PvIMSMi/jfAoaMgOx5sl19GUqD3ktQQmRiCuihwc9m1ttZ4nF3fWtgQgY5W
MOQxGvN7k2a42ihzXeBZkawvbQKIXtMPFbnbfVmAu84flr8W1mtdvyf/QiaP7uEl+F8KEH0cL4D6
k5TyZbROnMnMW6j8ui7dozdVQ/Sj4hxLPUxT/vQXqmruHOpDKtiVRAWRvv+R4qsbAurlt2Y0mSbh
vgUSE50x/YqGvVu8OWpU/oDJ+KPg8ehdD42kl/MJHkWTfx2teyHFE4b1LybaL59BtWuDaKIMRXCc
Hf4SlFey4+XBCAdfmY6hNAncLVWXBbZkC37BXvBfaN0BCqtct6Ml4pP+fET/lq6A7FeVxxyFo+as
q2vHbHbRCUKBKdQ7zqk4a6zTqQTk0FHDo/y2L4h2imv96FUT6Y/e+6ZUVoolnpmSy6TyOkMffjEN
dzc7K5Dse2AaV4s14rnqDS4pmxHMOWHLGg1G8epdXfXkH+Grd5XE5BOlI01RIMt5tZ+Nfq/JrtRM
rnTEPEZp0VoiGmtD6Y/EdTPqJT/Uqz08k5rMMR/sTdfi3qahrkE6yd74I+iOdQ6z2PdPr68/g/7c
JevT311RlC3RqswLw26GPzdILBHt2EkboR9rD8yUpiuOcR4rnEj0a8yBBMt5h+m0R2Ey88NZPu26
c882ySA1+FwFj/rnprxipX0dVTk8G7s4zJiEQNRbXmT+mAwFHTm38rEyVYd3ppyvzdrnZJM+vd9q
vPrkpmCAXj2ZuJjFMtBTdrpVZZyAN9RDT/MpUtD30CouuK2y+euthsYJCxpRkJi7UqWi3bMTHuoH
GmBhj9OGG8RQ137Ear08hutZ/oWFxYPVqayksIrlMDZ+w6X7afMALjU2NK9CwgfGEyXstgp5yzXU
snDixwU7Pt/D4Ndh3AmNZYMaz60HFkjfIiWmZqTneSv9tckff7OQsXZiBPqXXFzBsLMgt8vFSO50
WeZd4LzipR/9EfQxUKsxrEamgINRMu6K3LGLP22imMKYbbkrA/og3dxKrqFOE88IJ+cZIsS541Lt
q62RqGRfgu887jk/+bHdUEoIGoUnSXqOaM2n223Cfdxr6NAxFEQuL6fLu2qhLBCgFGaA/XTE4unI
xI+/EwnjLBXxwnOKQyXTR7oZLeGf1qhZW0lhqzlRipQnBtMhMwmfqt0Cte/nKM1mXAl1f0Zb2eCy
iPo1XIm7TH0qe07AO7AgJYRItajjxZy+xr2bzNhr42iOskUYi04WwPHGkj5H4wjmSVF7D1mp5hp+
/vbHAKPSMIqaHnN+krGB3d6RUjf61IbUwK1so9zyYJ6xeIGi9eJKiTaouUXJUViDnjAQRGYdHN3v
PIZEh5j2R51AOhjAssdrVI+5rISa/7O60E7GQPoQE1KfTZ2TnCpaLeqNEcLCiYpUVrrAe/HtlwSk
a76fOnaCfsSrIJxXjQ/3lH1OvNSRqHrefk9Slh6HnrUQsW2psnVFtGSnFGYOsMKareDIuJTW6Wm9
jWbkBj1Fs4IsNLCo3thoZnd0V7pdjxoVjR2FbxL4o75BxQC2N2PkYLDG0WaKjr0BNxdDbtCADZN9
85elsxWHjBkBiA23aYAk1hoesMFp7l79Gvh2XYs+sFmuWuodUvbdeL8Yp6ha+VdUc3KO00843Hm+
Lz9RCDlv/dWXEq+aY0/iZPx2K3c9uaDH3nYoYUgl3DhtVuUT5FzKayY62vB17Y/TaHnFeTYO8Nx4
zC9HfYI6txRnc4FZdaSaiPq0S/jkKamKf9DIZUra4r++jG/Oea49bwksJ7+z3g8XD/DQgh9f82iG
akTdn0h0QSm9W+Dn5Q/w5dxsiyGgOBLp32R5PlHL49ai5xhoy9O04ttRzqqo5aDKLA+6DMWqJjgZ
a4zAUqFIIzKPYSFuVE5Zi3CQeUfXSCXioJUnj7SOrz5SY/M+SzafLzU5GMIaBQyVG6lLYnBKlAe7
XEemAtDlnB6UptDN9c2hxUtf2cBK7niLPLxcOqI8hcVgueVKTwPl9Q8QhcZjrN3nU8k9Hlhw1UJC
D/e3kjdR3xmiwkttXPOmCect3i0uaSxjOUP/P58+iDNXOlNSx0sldDYqy4L1wpVQoH/Xq8Xz2K5N
BItGoZhCdHweBRzxgwHLSeOcRJ8+EwvUOvbXOjoH59MLVwo3fDcB2x1P3sqzlD5CaHZ/7B+wVYVQ
2kJASx87Wa6/B+sGOB+d3m8SovJEZHcNDuRVLNJyjt7q6uHuA6+/A14YzdT5I5qL0GLae2E4xSPZ
gzjMCPVkiezpm6GvlrBXmgsoUp5/XjZKMaK7yToqpZKHY0Oej89+n3BnGPynNEDG6qyOFdZo+5uL
0AxkE0BGcwIB2vGgwIsigiURtHWMn6ES4xgfYlVUWRPY5aZ8Zk6U2PDr898DkDe2cPZBBCUGZVq/
TK3UZbvcE5pyEUYQ2W4NrZRcSf+mB/+cbLheypq7ADS8HMXZnszTGquRAr1BaNY1s7Dur8HlhAQp
JDzWGqnfS1F22ckA7R63+588EArVKIMbnwkcTnkBYykbJw8YAumxM82pLMfryhNChIW1qr0azuCn
U+qhJjcL4rB3ueir9T2km2pqrdCMMMqtOFKEWWwsZEBpz7igB0apUHzYpMPQWaL1sMMuTng/NVIZ
QJLs/K2CwMSHN7BzydB0Z3kaafJlInet5nk7HdvnNWQL5/LbbkBEZUEXF0bFPEGiYwBVRwD/jRYe
kNITg3HcUyrl3HDS6xM73/KQh52Y8fvMF+FaDZy2ZlCioYmE1PZNce6Kct90bw9yYX5vrCutaczB
8DT7xbqHUgoo0kvHAaVrjfnrbI3QO7SX7CL3344rYJqmM9P03dCI0i6e3T2h5J7u4SqD3SHWGook
7rn+Rqz6ZyOVjOn4BFVBVLHvOcsw+UIKUT4sPxmkG8nt+d8bIfk+I1psiqdrjvLRqoGjzsAPVlYm
rcwnpubPzgxXS1B1DFYEKrHTdWI5qbSDxRgQlnOLKAOn1mEwxF9xYOkuoQFxauVsHjIZmEUYwxCM
em55MDpH2c8/RNImptllcutmBNhjtoHcJFc1fF35CXqV8DUpH+U0K57oBJezvWsKuRnOfbHbGk89
Kbeg6nu/B83Bba/jwFTXWXta/+anAv8P+OzZwdn0aKvPEqKkC9IiYsyrAHhDXwLMpfDF0YM2q2La
ga4iVzrdx/cZ5h+Tz0ZcQWdNOuGbYu3uvh8c3HyP08BLw/akT2mofRmo9C8MiXr1UhOU2KQpg4RW
3uZwrTe7VXdBb4aX8XZ5v9URTnuQZoronuv91cl522wTsi93AT96l3cMrXG1ucgtyyA1ZhYs/hMh
M5zzQJAgfvDdzBRm1CL2sB9UNsxhPOJFF/8a/kSXXDDDDL3+4ryFvIotvjvxxdr+D5lBv2aaY0AA
MwiqaKdtAl1l/heAYWDE4f4u9pTR2MYZ35uzcd1Vxam4yPrOUIOqNC/55b4CzobM2LLcn3bV63go
wl5EU+/fLnzq9rhVYUJhCX09jb02S94iLMHs/99wLket8vERUUHMhDv/drAWgja7MEh/Fwm+MEL0
ziA0Z87zEa9NA6siKfpCA6VBZNw2f5GV1yGyk9QS7Br7KFcTR0589SlmT20hQy8lTMjIQh7URN1I
Klh5sX10OzcCPXk9VhD0VM4RcDge0904RIr8fzhplKf2D7sp0KWN58pKH2rAnnFUFMsP9/2fQ5fS
qiNaoRA175Z+OyG+Es659pU0zRyGgq2IoCekKQu/xYg9kMYd6LLz1jjzMVV4QorV+iZy8rmPLH26
/cCy7YESACGcwS1niS77ZDoXlNQ1yUO2YQz0eezaqgJ1s4M3yrZhrV6UdShFBc0iNWgYlJtGWzJ7
CVAhWTvhmH7kqomcXgBmkhceAY4QvlEbtatwG0XvA2IPWQOXs6jDaCcXUx7bjwsMNR6JCJmPz7ER
3LALEfUdYqsDp0XpjEkCU22/DxOJHx5UXnviNuHj61m+5bKIyqVJlscBj0a6pPDwluGeuO+A+ark
MEau3jMyxLn7u9qxpy0+yMfBkgWWTi7Fs3tEhiZ3kQ3/W9hBj8xF9PTH0JmvQuyWFHcVZZFQLMJT
9F+EFsRgxyy+cRKWLrmgTJAssLoHhobNdWMPFGgIBp+UrnwKxYH3tNJYICxvwPbifpOX4/bIlOwk
1/SFJZui3STZgqIsy7DrSAvbPLLzXhJ6q6JWWjTIC6BiO7spQp6N2mORqvHo1H4uS2Qvy01kBdO+
/FB/UJhvZE2mpvPPsPUVVy/i+HfIsV/AZEPc3Mr11fRYKjD3ABfu4G3Kkl3vcPRcl0MIXVPdhEkI
hdfqe8EQEVjYGOD57xyHxqx46DVfbUBm14LRMTrzcplDpTfNHHoLrPQXBedY1WK/hHdBIpBQp/0D
Ccl6CoJegjhFthIQ6IySN2C7n+ZxvLUSojq2owdrLXFFxTzX6StbE3wgNqykKvtO1+QacIFAx4YP
H4NpjHELrDLuntwDySQeyHOvkywtoeb5awKWK3G6LMu0Wg+p3ydgdaO8EegDEb/tOcCTLSSNWB8H
TRT2czMPC1JpdQToTKvwwIQbS1Yusi0DRCKU2wlAgIjtdiMcQGMv7GzfvwfNtab9mpiT08Rl/clX
EB7rlDm6xmxwlgdkjagPZQ5vNe/7+DV+RQVyKpwj/IBn+/qonGpH3JcECKkYnGykbAQ00HFcQz7u
Dp842z8T6sGhqgVY9sTz1inQAkklobwrq9uQ0qf7uTsGHmKQCfmtIIfyzkwbfILwnzRPIz1/gsHr
pWUhPMAYMonQ4Zr66k4uZghMcDsxMlPKRwDX2IlJPb58J5TO7ha5qA6jpb6dFZ3esGz7D8mRvu6j
M7hjjP19IxCgW9sisfa4IU47edpNqEZgZyZEIxUPRyd7I3TmxyYioNVcTYLehX8ss+n1AX/+oN3h
IQstH6VF1ms8JdN0OR8BzsvgDJ6Emc7xfZ451Ek8Gl/Ay1VgSkdiYxaH2VSJPZLR5j/GOGpzRnJH
4M4GR77svTxb2SQEEATmMyHT2wtCiEdX37oR/9ME7cvFc8zVZV8l4GeteZ8mL4Hg+iX5FhLIXeAD
hRJpIhk8kXsFdY80pgx/Xi1JY2ttN+XNgQOefm1rrrcacMbw3HIZZUPVd2w6fZ9Y9FiRypmZhsvC
JlnVmsyGvOgAPpb9JeeMwQCKIqyZ6UYnCt1g02z4cQ8j+0SP3QLMxcUZ/olh+59mUix66EBmePyU
Znl/aNdXkne9Qekhl3f49C7Pfdkn5gOlGuCiMLH88/0UX1CdqqmaiMdfUZsQuZ6dGtnevy2F06ac
KHHgkQsVR1itIDh70RXX+s697My6q/6SRK1+JOKvZ+z02QcIch6bWotGsl9GCBEQAjwgqEapVjrr
flUcSTUwicWj8dFlmdtYcN046mfAIe49oFrxBHSAd4OkBjhs2HjNTxRkRPQXIRbmnXbKm85DapSN
bF/TGawYVNrfgFHpSXQdPhyO8ECki4yJM9PUwMgr6mTT7H8vUKMz0BiIGflZjvC3mvsqkFBJt2JP
xCLtnDzuyjgrA5pqGaw6U247CDhkYW6Qd/BrlHHRwz0LhsNwN3zJhB53gbILakWjSCGRhtboR1QX
CiUh4oFpR8+DRpnn56QYKnRugYF9EouegLW9/WqHJiWY4xrwMqVMbufn+5phwZiV2rvSHkgYPrAm
/IuiBx8ZN8Kcne72tUWjsuWeHlW01Zt/wkroNisfgWJx6lGHo1Uolf+arF3HKvHM1sSSBFsdyzTi
TTelUF4ehxZE1Z+KR8YpNV7IGQfvJArwsrFBoJqsA/SC5G42WjBeqqj/HJPR/W4Gv93SeHfd6bfi
NwD1QHONBcJuFfB+ut8kIXb4t0q55/bZgro1tpAZaFXXYEkZyO8nAHGHqQAAJHP+ZN+/aN6Cggs7
DSmyBDp3c2nLT8+nAFiM5ZgZElZ1/xVMTR6ytR0CZkdvbEM7XeXWDGe2y5b3I1Siei0l8TNxeHUW
jLEnNzkjwizzKKz5pGodk1ys2BpqZyFrds2cYt0VYq22Kb/8wdCtQLL8HZ8JodC/EyhdoT6ITh49
ozCnmgI1RRUIXJIrzaT5DiWTZy32VTHdDA05JW9e3BQEIADr2BnYzZSeKzuqeAk9QUYVS1Z6AYSv
H+h1aMOaQU8SlM8DSlma+15p4Y7L3aoXmHY5ze4V1feVqQfgd7Hw1OIzT+2Z118EF6MwwXUmQsfc
xCAcWceJEeIOQwFgaB4D7SUpAFvnEhJb2YvuYahOZGtlYLO69BoKwzysToqtWxJoo9Iownhaf4We
JGntQ0P7IOWhEHzp31foPqnihI85QemGm2gtE+nyS4WabqgFYgvvCQKKxTLR1fmW4S4L3/O8a7Ks
c1J7q7idv9r0lKI2SeYGo4MMOX13bZi5dGKj6tlJLSMrT1cUZAuvllBl7GaaRbP8TE4uUu+L6lUK
ipfMYirc4VVVu3iH461uRBPLmgfcikZ3SPKO+dsUiT7CEmUUfquROuDchBZ7VW9S7yrmlfiMKQtL
MPGh4pLi+aUhk9ZT3FP9FwZDb0v+QDD5G+W/wVmndHED5XNPHtmBnX8/EsZ+krN5+UCUSkaxBp62
x9r8XA8dFz9DgmsvXbSf9PEHgIs7y58mKVs/t0Hcwd3RAKKs/LDxnYVxTNPr/RTkNIOEurPNuGpR
fsLZaV8o4yF0e6sLTJrcgZ5udkN5HOzU/Dh/NsXmaRuPFrYIpJqLP9zLqjQN3IuCQ/34duvo5nV+
rP2/dTp8DcXtT2V3OeMRgfMvwPdmZXeABWFPSWj1/S80BBiALWsU+SyYSmMdl6LgPYsgCw+ZlsRX
Re/sLX6bB0puBXwq+pU68QXU2bsid+igutGrCHLSBuw9osKax1Vz3VWAR7feO+1MKH7A8KavWWpe
DwqIXJjQ/Wy8agq7x2d2kyLjQAt35fnYSDU5PMs/KxUmVbnJWce0kvWuZllzHZnEbJX+M8mCHHeZ
CsaeO8XtzyRowym0YzjxzGkk7W3TexJRPzTpDSs/MexQu1/Hb5jLuXs5F2HFTtffDJ3DWFz/r6PR
3cFiziuGrBwV6TIpW1TrVmyZqe1dmDzVVr8btzI5m9Njcb2eHZPbzGPm+JvJeoKj/RbrIj9Ekc9g
K0F9G3I1R9eZe5I5COGzu1n42yON0yhrnO84zv44IwVKFZL0OxQttfKwl47Evip/5Z3cUtOHjAf0
qMv0Yqk3NZNvWapyuaU562T+mIobL/TPY/i2GTkoOhJ2Yht4iV1kFaDa6UbOJ5bZyv0kmmbmfaPo
kLBML7B/TBP3ReTQ/aYDpn60xdlow1mQEFSxSkO4mb28kiwYBZMyiWnRcoX7bO9d3uZnMtOX/rin
29dgVvTxgq3xaVROcXq302QZQVnHTAg/4fG/mMyXfo4qP8l0v0Eb4bX0d3TAAPuLqE33geiCkPKd
II2GcBIMteBO+nBoHBDry6i7uM+9Pm7xDmfjIEslbsroPuPicJtHu5Qt5nCQMmv0QiYLjLxVuI98
e7BwATC41fLXlV88lNdJYIGrOg8bEklZ2XHuHBgv80LaWprZrn6lY1/WALg1ZBvXv0R03c22U6kQ
V30+BD2xRkON8W+jzZwalCvKSIVbstauxfF0Fqh5PBxY1mwQLoa2IHpuwoAiW3NxE8xQ7NufgKIe
xbCxZeyDP7L0LjNbo02yHDeEgN4FQSUWWaX5nKntSRjcH43i5Wm9Glng5a9bo6zIPasgZOeQ4HvX
pFiCBC/P5qBiW7HDjaUUIcSPBJYn9NM7Y3JRfqKwa0JmcZdEvm90VhQOB9xEA3tz1bLyoFZ2jUfM
DJatSr44KuHHMMYzTiTL8ugGqc8eMj+5Nl1qSExEixJGShmLBgY5FS6aUY9S9meg0SjNRUFbA6/g
jGt8NeiEHrTE3cHcu2089CrW0t5h7GJREa+JmhAfWth2WF6o1U8AXJobt8jGbOybveOjDWaOJD6y
a2zgRbzmn6cxH2WnCCAEPNy82y+r50j1vV6kbVC19disIN6mfX0lN49I5Edf8o0oVOYfLoKZhHW2
iipAu0xYkRQsThR22wdT3qPkRTMcYUaGxYUQ3ghEC0SgTCAWTeHtEY8XbPicrGRZvXvhCAVNUo9i
PDnOyuSvOJaOGehpNAyWZnj7Gwy8ldTD7PpI4XjDJXY36TqskuhVRyEWC4wTb5esCgwfc5Bn2deL
YV/Ehi3dHn0jCp4Y4tWIzutJv6/h/wIu1PCNXH52x77tNjtqueslqOoGWgqyD/9A18TeuTa05hb+
ud+WpDreWYmtHjaFTDwGqUIlVw4mHfArchj4MwtLjYqE9F9g58mDtPnoslb1Mrk4Lev3ZLlJh/Z/
l/JzkdfnfEPilPqwJs9KwF4VKHVL+u/zaWKXMfXNlUJI0+o8ua1hQa8cDLSvCbLh8WJ+vn5dLNAf
DLwn0KZqsqbNj8KMrvO1kx+gj65xiELg3/bhhP15Weoych0a8Khn9ypTCrPEAaJr9Bn0zZVg9N/X
PBzPSbdpxyHylt3dconE4cL52JoOs/nVI7wcd1tlcNFDkhtMkQ6eJNwo61R8Wn6x1oVmfc1cOh4T
egUGggT3srsM9zg5+vCsNnRPWSB0tINZ/8W5uPWyh7S6acne4fKzq9hgpYUTXLd5tpkvRg3wxgOL
IE/Cy5MYbZo5irwYFvtT+GB7yh3kcAoK7IuhkCmDw8O1CJIreXbvOcLZCM/q1dJ0qWPSTDnnismv
Z5hMxza0kweVN0M0EqJgLUFrsqbdZuLvOmAEut2Sw422mgMEs4MxcgiExPubCGVkjo+4zYztn61g
MHz295gGhco7bwyCg/dUaM+oBq/Xhx780dDwQX5Cm3F33RPWGsp3bUN47EQAzmqkmh0Ioq8PMr0N
JhDUzI4qjxKIE0stgJ8UOM+5TDYXCAEUCTDzrEV96lWjCUaKi/gpJXD8R6cEw8WIsTqaFVYqzQxC
DjSQSslFS8UAqpx6kAm/7QPmdKO1NAcbcULjvqpDvoYFx6qys+gyj+koxMhuAYv7CYzZ+1qIkBVN
teHhlGiuWidKt6CkyP45GD9rXPko2zlrABVllU9+eeNXrGgTkAv+TLEyHdyTdL7PQEDLziVJ6A7+
/3pvFMIAZzNB9cL4HtjKTEzEEo24IecHBBBCgEC9l8zjEx90t2w38twSixLQM8FDArUJ6Eq1jedP
OL+nZHrnl3/yrlf27AdiCX1vvz37D7XvormLsYVmDwUc9/V7Id+a896bCTkwc5sy8LBCDKdrCA1v
Zr2KqLfuUzHqTLnXKjvZje3vrje7zX1SRpxKaUbgYUd8cRpSH9qEOlPMWMv+Rut9umxhdmCtvTyg
2SRlR1Ry651YWmLYkoK98c3Ad51dgsIhz1Eeb57Y7PfAy2wh/niovIkAk7ZVyhzzWR9qlRkJJ7pW
4XAzyYXhunCuPKCI75t5kjghQiKlg6S6G+Q9YVunY9tqph3jOxwZ/RD9yQyjLfvxptTy+ZG4eZwv
prKUSE9YuubyqygfvJisDG/E4u7zrrPtPtBKCB1XxW7uPACd8aqze3tpwK9EiT7sB29LUjhQOH6O
vEOb2jLxiAu2P6wKqTDzY+GybVYFa80tLjsCdQy28n/DvDY4r5RNhtxfDi00sLb21tLW2DoCLWS2
jHqnnNgLiCwk1QELrgHebCU6uB0QrhCjWuu3bUqKn1uigpPj+QkhVi53dVZmaFA/OfwVFCNHuLQk
PJgKHEHf/HSLiD3wTBH8Ypd0Jp1MAS5KadjUiZKNqh9hxhPmTaVb66cj3c+2hY3yzKPfym5hrLy9
QtTdjfY6zFQLQuUf6Pujw6UJaafVsoNCQc1g0MCuUxBUl6Zw0wklUo9i/FKtVb2NJsWPy48/OnRD
UIiU8ienO0602PjEgMNDNDaAUGYfj0BeIKMyfmx8jt1l1OhPRIWwbE0ECHm32BWS0l01oG4WsVuj
4NX9uVaz0OjCJYvEQSBhaC+t8IiL/xKETIFyrhqDHpdL/3Di+yLM0d+oHpFeCD2eX9TpSmDGriJl
70JSfmPzqtW4qn2YyymMLs5jZTbakawqigRaVmW7PZXVF9AJZlp5UGoSENU9+Pydhl/9B1GkJkOW
Ck/Vg90lbsGnAlP1dP9s9HVkC4BPNBFCuVQXbSEt/IXXE68QbfsKrQ2DAyWURaGa0xko+/Dt6GLQ
RnDD2ckRLH/mrUxQSrMFHwTQC29nOzr935F5t71GlIfUL+SMeGOqfy2tYw6IkVhCu4xzWmmZoxCa
kdIX9Gzs0LbJJesremdoTrZZ/RJH9SqO48oIdfQXuyIA3JT9Prw6AazLLwrcnEEYOjJ2Nv3BlnNS
Mg60QmdyB4zBu78TsQlLHMbHeMCHl6mczmlN+sN4jrTmIsnavD2jGRBY5rOBwbGSMiSONhZIr/lY
Rgnik+BvK2ZrLLDzAvLyr/sWJxPcbMyD31jBrNg9+dD0dMmjtg0btVbUExwe3kNKAqNdELfJxEHD
KiEdrWkVOYpDae942yl1sY5jR3Somh4i2rhRmYvJ0ArR9UFsLe1HpUI+IHsz+0WmOw3AZhy6kdvg
0b7P/MiugYMGf+acpIuJ0plzqjmRlZAR1/qqtQElJUOzUoPKXedWHUSN5hT8OBNPD4KRXT9fRU7Y
k8ALeIF5KvZB8hHL1kPCROqev/30vlf5/kBa9NUY8WPaWjYvXnWtCdu4AvadVcG5Xyq3PH/5/xjz
/D6v1jN6pgMBuYWNK/w5loH6itUf2VMRV+8x5QRSRlhAe63bV2qcMxgg/Lejxct0rKlzvegkwiC9
uCgyNWQYYac4PGkJdBx7AHIriwi6Xmx5M9dtpn5IbHAeGDRGL2n39nEuN2jOYgigRZneBQVRzqSO
z9EjJNGTdPjbpm2TqkPhZRyhic8ftqcHKLeFYI3a8a0hm/wSGzaeei7w7OH+nVGolZB8mX9Ko1eB
tsafnboBJuYxzNopeArLeEdyedcH8TKnOVE29oxXznOb+V4ql1dIWtHhsczRHPl0Gg9p9ZV/Gf4z
rBrKIoF1JHDfdqEFUU42EI1bJ0yCTKRqv6hhSkNyBqCio6G8boIXrNDQjG9zxrUvPGLijZ8TJlrc
Do59SzgchA1JbvROEbs+dI5XkE16rScdNSXdOmODp1BsFGTd6VH06GOPyAea5jbleVBmobNGve6O
DkeOFd/VVNnF3h52OlkwcXYuCi6LsOKZBKt0KjvGFuLfGVuN2DQXZuazbA7KO6HMVM4AbT17KCB2
/SUax6KlFjho43I8eaIn5PwziGPW+gbIfWPybdjDNZg46tdtrcilvpUCre+Hj7o2SPBW/Ncx1HWp
+Jt4K3mIufUCneAPMeHuJPlPGJoKevSUOVvyWm73OzkgOeicA5h7/LI6Dr1SmzM6ELN24W6IEGUo
pDPnT1emPElwsV15V8luFg66dsQjTm9cZL84XUG/7t3+4nl2ebu2ERUmE6Tx1FeAvF+kUN91EREn
pW5xNkDwiF7KZ2OYg1EmUK/A0htqZQq9pk7ZByMDjXEmngVCVO4jhfFOTojtybiwlM7wklmTbGTU
CmzQxOw7LfknTGl+jWP+LezJ5TG3eAv4oYd1PCp/u1HITLPfgQ0N3GkyQvWpdcniksO7/LpZH0Lh
N4rQDJRhkIwNOwicbRCWLJjFuuO/sTI8M+XNcLLvPZdQT9tA2uPQiAVl+YqUF+sfxhSmIBx5GplX
LruHk7E+Q1nO67hhgKltzm0WGloQwNBjxfIgGUdVv4xUYEIBcKLZpTOTZNoCAnhLtPu+7tFPxzJm
JvkPoHJVUmnytR3mQWUCCWNS++Y8TmD0wecbIAsKbarngLTxmJEkseBHP4pidhluPTVOp2SbpMv/
+glPeGr4GQZ/8hiYEFG3oLp2Ant50aIItVBbs6DZTBW19BMtPzC1Gdztg63leVx4nTCgqf4+mlxl
2sunaIlmzrthRXg3KTdiog+jzYH9S5BTxWeX9w7z3NmHnGZUWft6Mri8gHcoeJR0EU19k3/PU4ND
lXHwiZtLeY7roXp/ls4vyjsmYzNeS2nz9uub5SyXhS+RBBntcGYe9msoy548Nd7+82gygyWRRURA
6ShnzPDCm5rJg55aWjzqy4M1T5/kUSekAJrfevP409yQb8uktPtdY0uUTotDhbYqVHyXaidxJG8R
qjEXVHSz8hki0xtKEyfQHGXYgnMwBgEJZRCJIRv/MAk2WyUfQdkJQtGKoxMv+V+ND90DwVZBY3P0
ISx+UAcS0F3wo2dzreZSAu3AE3EwXhza3Og6ojIisgdepzTXfuJBwJznfyRkKXfPJNIy2vcC8uYj
Ygzyb0B8XxEGVdTSgIyzK+zVvY6cXCGaONzPJi6XqpRqa6HW2R6vcqgw0dXuaHPyVQkBKv7WDxia
Zsb3CIY74lCnHtilLWrytn9RxyJAqGvJaGVUGt+HpP0Z+jxro1L2P3NULb6bpVkw1HmP2TFSn1Di
MKxzGNwB+Ka5CY3aAJU363yc4JTWJORpCqMhk5E8MYoyqKLw4nxU7McAag+Wa47m26S2bOwk8Ajr
ruRBU4IB3hWlAnnS1z0IxL3c3704eMmwru5ij5lZWIdu7XwKIWIo9pKaze86G7DAPJz+FyD5v6BT
4+AnQhV46otbpgPaG8DXIyvETUF+a7Tdj/aA/Hx3cfX3CQcK97uR+qrNPM7D6RNZq3KenlcWZq9w
VqLymUJHYuQrx88D5zuGZCPx7OxHvzl57yWZVRmuWvr1v9bUOvmCrNGLUIi1jfStU0zzLzUA8iR+
Qsx0SBgw6yXZyO13mWrB8PXEI7zGHs7AtqeuavA9UUz62weWdPF8YjNI3OByshr41NsvWjkffi5z
Bnib43aX+mL4PF1vVvxG88wIJig/cIfqak+BSaxyG0iRDex9yp8D6TvQVA9nvxgQDZAjTLsik4RI
/HAyCxkxN+7jkoki6dEYr9PDqlPmSxBs5ElpQs6aWreJQafqqWD6pbdKCaZwrgGVUhr5wSeg2jNG
sUXAUiyVQhPXf3YQAH82RUQUcYqikuX5I11FwCjWn1zY4pnapDBPz2QQ8WwYUktPCaQaWpkrK9di
4Bh5N5axNA+Vx+RQMwiiQMm8mt6enwghlmNxBZBzGySgk8dv3epkdQH6zSaIGkv/5QDHR+fKnP5R
UNHet/AM58lzKnJE42givTTVG3r0Pbj0IAYgyxKhzeAX1D/A+GH9SHQBKtGGktVNobF4BrtcHfI+
eLrD7PkhkSnpraXT63vDT+x2ppMFhBby6QqYPhyKn1RjmPC3V/LxO62tOSax4TUQljh0HRPZuKqT
YRXoQOGsJT2L/VVCcIvJTwIJDdzxtYNDtdn3QE+q1W4XWVZJtbTUjkSz98ERqGLWjyextf7Rp/fT
W+DB+BmX9P3OqnVKx/Fkr7mTfHogR+zMqw4JqJOo1WFv661rEEV3P0WIPi/96pN148ancURICFl+
Jy1YWhLwrVf3RzwpS1xslH18YVVPXVZyh0dAnF/6hhB0uKWDIWskLRxvZVzANcg0iNZTqSPBNQEM
WW4lLRimSqFCFFomkmea5VXlFFb8TOPjftFGF01jzl6lkmkcdoTPpi2kiCv6bg3PlFylmWHGqs5Q
HiVcjopED9vkVhAxeZe5PDdX3HZ6WvHZyR7LThC0LqvVfrT2aRyWgbCPv3eTcVAus/N6A6hbCq0k
JrPPHd93niGq1MnNjuddz/E7fSDMHxBVH6dNYQf5JzYrvJDZsNZ5znvPsEIcOkzO4QhT0wBb5kfK
vHUQ8+p7OONsrCDijzN7VpnAWjGIJFYQweApgXC9v2CbkGLogktyHAh9VWv2CeTD6W3MXEJWQ2To
LyAGYgZSBVR+pSCeVXEeQPoiAT2yaN0TtAoN4/SFcGqnkvQ5fwW0jvJPXxomuVLqrDbxT4GjZh1V
UvtDEvPA6rMIiWhYtfq9XqFUc671x9GxmsaftB+i/sLG7cBowg9lnp4J+OLyi4TDh/AhM4+h/CMQ
VdfyErrksZlkEr231ve/7NnbVINa+9svQI/VOeN2bfM+IaOQhcndlq0MiwJQjS/ClQEaRpdWdfn/
Mx3WB78EYYnIYnxCJ20CLFk0knhjogs0Qn/dZipnsNZRVL98jPP1CjjryAnfVlWmRh2Q0EShfyVj
4dD+cMaMfYFlO/chHFtQ0qKy15+tykS8V++rTw0ojkSKcs0pD4b4FCPuvLIYHSk4zFQDTRU05ya8
kGalUPmNJ8uErrScYH2XOhuvC7CNqVc6uUcHxQGnG+ZHD4OdXh4ERxF+2p48mroDbQyy/DqslpaM
aGxPeIRD2rORTOI4p9RzRfDX2NkKlkv+rThHl6RcF8BaMGSUm42IK+HtOCe+OR8BLtsO61Ws0On3
T4wV4JRuGYbM/2qy546+SpsRDDEtvKIpSe5iAdb1aj4ksHrsB8k+NthN2eU//pas5hXJ+CspuhSY
SiRpl0g4jNUlKatxiFUeMHS+MuL7+TIi7MR2u0Zzv/ef9Ey1PjPlE2NBlt+5XOckhzD1MMhifg47
VSR/SVyp0+h9qqWftSdmP6iKb/b1+rDaUQ8qDFbaTTFsC+/45TgSSDaj16dfQ2U1KfHZSfLsyLx3
j5A57623UKgUrhBGIG75Ms6K2OgLvhXdYIjhhAoqqvbzx8+KrAtyFMlbOc76B2qevbyLzmldotCl
oWv6jMLpSYPQv6AUq7G/Z0bHCCrVUGeD8kecCXBqfoBMXujezsSpoKjWVnQ1W7NG+r5FSAoNRVyB
tWqeaRGBEgtz1yd3rY1xBNGXellAXyrIREA8uvzgP8yFUeOvfwmm5kYEoa3hzx7CZxWQXguTXDdt
zHUK6GP3BfIdiJQlY23dPRCS+YVLsgVXNSjM7rh4KwZ/iCJLeQ87Hy8bbShPgdunc0wI1iIyAoGA
MtOdHii3vXv33ehr86y4P4kAPre5eKDqf+Q/RFrUIWPhAtPqEsQnwnEtLg0346R7uN+jDtJuXtMk
EjFnq4D2bvS7l+XCi10BfPB7sU65+m6uAZGwJoAMnk2K/2INQDx5fgF4vk6ivJFAqW9RacTLZ6M/
sA+ANcjaN8UMIFgxndmJgp29zfx6SFIOoA5ejhOK/YJlMBkH6c6cKXDN5wgbmY0QlnEZQga9CG9x
UibTCbdD87UCQZ0j9XZLnfNT2dOaquSfGoNdXLVnD3KJWlumL63VawDSrjG5a+Di1sQ0yM9DsD4h
v8SQPpVj6Vpkt5uFQDQizuf7s91lHuh9jgJYUYzuGZtj8lx0OaBfG63rnVzdFE9dIX63qKZSwhGK
MHPKlfq0mJKmm0YBr6DZs+DyKAzMZhF55E0yGCyFA833SEn1ttvH9lm0fMbqVMGtENHJGAE+OYOH
Hj+lDmflS+8b4BZITaA9LzY7drwta2Ob/vTJmevK/8O9h9VY0K8Yp6fRDqK+OQOEi/rpGFGD+95F
YH9bvOYSTRIHbdqZmbPz1VBnAf+TpYM6voiht/xb+AncGhzftx88u7KTr2IYJ3vnbuMMjuwfjns2
3ZEdBo+Im4DkGJO672fMQGKEVfZl66LoYnj66XpD6f9S6bYNOisLi28d+FapRZ8Lcbe+SaaNDIRf
TZuyK2GGJ8/1BHpLRQYuWTEqU+UlSHxHJsRWenoIxjiCrQ6vb4909qhlN3ZrTP7vAoyfWre+M0E3
uINC14KqIxFYhxfDW4uhx1tyH9+y7xpuLhbx4PbqngrqqY5X5riPQpBTmeplRNSHEyQLsn79xseB
b2Kf8ZAW8SnXaJ1JkYDCNnMvgPRlqhy5db/hrKld45PTyEaTnf1fRzZ9SRvan4sW1KmrvfJPYpP/
honr4pNmwrWpPhPmiUlEdFJDcuULMVa/j1fp89tHMeetEUoBdZlqEMIIhmUhCVyo4Q7M+gQ+WDD5
t1nTLik2O0OoeBfr/GPVQCyitIog3raGz6xCYniiNHle4fqFAS+I9ffcTKksjFxSk8HYHMliZLxB
BAnRoD0Kytl+QsBsrRHGKd1lQiC9G560J2+knH3Pl1tW1WE8NeDBdllKBNA3LVWZ/Kl4Pxy6fz9C
8snktCFDeAPNsXRcMFWoGq8L/Jh3DMKN/Spgrd04RuZ12kY1AE0AnXzR7m0YR2oFiWVZRIXf80S3
OEpARi6xN9iR2a8jsJeZtMailPcmzAP65+0mp9tyoJeOPmJaDgwp7tYSrx52JoKD110SAgMIu1jB
PxaKdTKrXHfpz6+YCZfB4bjINb6TEOaLHgYhm+AjTKhFq2SVLqodnwr0OSuKA1p/BVLMimqqeoYp
mGCZkdoNvwOXckJySdavYJh89taD8wPMY6wHEdQQp7+tlFFG0+5wBqjkEVPgZ0kHpKLgsio/1IMG
0Wz2xaGGPYa31TF8OWcUNDa+eV4oP4Qm9aRfAAx88p/0XdNpSmeFjBnPdSuTBuh0xKTgx1BbpWGx
lVYnVZlCVDBiaZowlHJ9pAtFxb+vyPrRgcxfJ/Z1RntHGl1ITXdIhmN49V25lp0xTPWobwXYSjnk
JPYnbc2lxNXFEyfUQ8zjFid/Rbm0WHhxdQk25TpSSTPCpBjhiBhIc+ktNhQxdG+XgxVk04isw2LD
Idowv4QsvxqRx0W2r2nvNt4evgZwqajRE3aunmXkRw9C3p6yTRdJMOmpXwM4IjH26l8qcmJYHXrj
qtzO9AOK8SRPO83+vczCPu8mtPNAUpveAhjlNVBEiWxrmz6qlzcaOwDpBdc3oLvqhyotaLvEw+Q8
EVXcfBCQrDrcDqN+qoV7UEHnh7sZTEcwhmkqKlVJ6UVZU5qH3SVS+uE0ZZIhqEv0284f+dvU7djc
oMWSIF3vLBveIG2w20cCx4cFBRqmhvcHkQDatjIpA1biKOFsUlJiNnL6U07QpGVD8MaXn4YnPvjM
r7dQ4qS1ZBJ7lWVTaiQO0/5qtnCwKSut24f+eW8W/d5lJySi14ZszR8prjFAk3sk4OfhBSkKG1Dx
ur0iAyKn92m0zbenUDuFAEnCUUdP3KvqOHpKEpnKQPcZHqsfZvLNf2gvouNvbc+iWQ3NSB0O7aFK
M+DT7Zdh4Z7/HtrgmlAjNWpFacdryCVUSS1FAR3qAE98BM0hm4xy9lvjiNGU8pBWnFpeGv1MqYYQ
ETSQSInOiX6fXbPWD1Tr6zEzFsupV49LyYbkRvG3x9KyJTBxU5iayCruJnH57/GNRtiukj93tWc1
m5VbP6obrJdHBV7UPFZlBrhYkIwmkoeqmN1bwHzrzS4s3EeYsX5gwqHyTF1FsXuLxRiBbngbfbth
+Gp7gFPMCMFQ+8RIshQ8efh22lIlxFdp5XVU6CN5qCi+UKJKH0FtWULci9qn5Qymc5OidRQONkqU
Uw98JwyvtQW9+sIOFbTns1eslVpq7Dbuzp8WaVblLu3IGJp60sIXNRvN2GUUfNT7wrhcX4RzAmjf
CL/QulbzXXQLGKc3w7mFaAIk+t62P9Lm8By+JNkStQL58QBcBQkFFEJ03BAt4ps/9db95hhw7Cmp
krlYsbE6w5RyyainRG9Ggbf7HHDVsuA3AAYAXAArID6jIc4phyTkGRdW650JAOx1lH0Cxlg6g6aK
Oq3rapWMcbLjYJhBv+IHV8/XLghybM6WoWkFrJNBpsXsdpQ4NsMzXjWbku/1J4BHaHrhGOT4OeLx
RNPEhhlEzG1SiJvLL1n1VBjFVMAQZZIN4vISoNzmSXGnrtkTZODVP54QLhsVuYraBqjozJi1MDRE
jpyb07V8OEKP6X2+LsYAhTHY1Lm9wyduag2MJaSVxwnZP50TqjUdllo+ztWKpYmrcVaHx/BPuJCf
RNEjTbks++KswhxIw6Q6ZPgt8uI+nLUHkznF+RHgpC+pPncnno3sfVM/phDDzDP/evMYWghxx8DZ
8B/l29YLkWwK1X/MgOEHr8mfP5g3IaWg+UQdPpxqUZfSyuPYNcPrEWQ28Za6OxYDqowjPQKBsBnv
HVE35POfIhC8KpV8Fuk5AhbsyUgkDJvZM9n2p13IkDUULjueXWP2XioD8+gRk6qlbyyzZObcXDiR
hqbEuRBgpSTuY0sP3k2FXXE61QpbleqUJ1lXiXeazhy2ZmBorHCyeI4QSzRPsYJdzTSGuc5MGu3k
WncM4qcI/deusabI8ML8uJiDCMFmP+WANzHiuIZLUoJPWQmstpBQk1eZQQwfi6XyTIGcWavWbRSN
PbUYsdf7mYQQl7nMwC6+AORRjR+gWXMeAhef2cT94i9RHsHdFdZSmmZYWVRSGq+VZCGyCgl1aC2P
ocVnXEwrrafuadixnazw9hsBZkH1Mh8GkFYxznGneTtjEBgOPZItASp1KT25sjZv8kx0zwazF2yy
i4yYijKqCFYu1vVJCIuk7KmTa5fqcG4NOlCUBqRyHW6G9mPnXSVlErSSayZGvuZGeQbJk6AJyugx
IDz4MavZhyNmcO2sGEfdJnfc2Boe4iUa9zTtdAd+dDW9dtjmjTS/tnnXmtULcE1qO1R2S3L0wyiZ
krLhWPHinPNZObcpA174BDwzfW2wQdm1eu5V/qEtlaeTFXZw5V+YBMdf2Ej8EMEk4TjTULeiI3+J
8b/Ogb6ton28M/90PjBCtPARuk6HTbEmzMQ6a2f52fYM1JywTNPdfBtXb3lEdXzJuO+VX+kV4DGf
znRQ4mHhHkZzxQ2g2JZd4SZd866JriYXhdV76QWgsjBj3EID0UUbnbaR2EeyDw/eheCsEu5SIGS8
2kFJ3y8E65XUFxqz4KsBfcTV90P285j4gPqLuBC1pZrnm114mW0D7NiaimRXNLF2pZNsFVKG4uMc
btHNPWRQMm+EGm5SIqXXmab970AR7OSpwfY3RcCqX4qYF1eYG96ugDQifInKg9T5L/x6nDErD1UX
n7LC5Y9xx9T3bveMapUn1/NLngwVuBKnDFjUTbB4xgnYl09Hdi4eSzyohZ6+pWvNtMctTdutxP2X
MLj+7dL9kASIWaGgVCSn59eHrWOGAp+H2qDipXzEGYomNx/UY9Z6Ep1oFhvnUKillkWDkF9P/Nf+
50HreWOarruISyfHdUMMPRrx/4F+1iu4GpCM+xOIgDaHWfktpoEraFMISq3Y46Tar7t7QiXA0Nzg
UaiiAwp7LGArswqs/eA0rHp5HVMu1wyeH0oYrWlt4l5/VdQCF0+w/vE7+Q/2iis+UxYR0OnIa0dO
zu7OgXZHXlVt7Cjtx5g0czYtK2Uy19KgYV10lxP729H+Sh76tyrTXbIkl6Bll4CyQaKCJkfdnbxf
ylynzd6+fvRkrPhKgygsynNMME3nAZWQ0MSnwVGYMWd68NcKRVEGI0ywHW4Y/HWDIxOcWjLq889B
yH2b4/H8zQKTFFGydz/tiG1fY8Gd9ymEYLQldNhiqy/drreCc6RNgKCHs6gRdT1VZEyUKj+rNXaY
rWvOcZg9BUruaU3R/T7V+q67o1c9aqlg1ToYk8HdhgBbejGnfye+C94FlaePhlc3p2lAWsVFzoo8
ffuMo6gu0T/JR2mV3nT0YDr3dTR3ZlYgsu/DbZi8ujVYAGZ12+H/VWYWs2Nv6dl1m8tadABniS17
YYQWG3jBrwYTV1/O3fHRpyzfa3u1W1tFho6idsLRED8uupVeDFVIDBYtE5i2ozKsJWLhiMQbSMas
YFtORHyCo/0wMj0xMCzlVZLMlfAkUG/DRL6CHqklFwGOGIRYpW4rHjzp8tFPUeGT2NvIhUifQ6UX
fESd1PLc04z3v2G9Svml9pflSzq06BinVKueWN7STL+iCzqbYkl3IfaqbqSyQ80LG8UQS9SkH3Ws
rfXKOiqCa7LO+1fNOuUMx+yAl1W5QHirJFBdp/VnHv1molxnEkEoXGxOUChFpmMLhUmaOG64hYBb
Xt2HddSx1PklCErUrl6a1RaSxpoznakjnFGZWvSHe5SmZP57+FWuJaILPWG0wWqeBxauELzvno2V
iXuTlqAVE/s92ml/7GDgu0ia5M2OpkNMSPF9BfN88ZxPVIAvhu3CmSob9m9QH1+zL/a1H19RsgUz
9ub0JfMkRIKQBRK5/kTMxPRa3q+qruF5DEyiTzvHSk9Y3vWkP1e+i4snlNlJ/ZHa0cvdsK84QQit
jDB++gFUTk80xUyqnIVgTUVjsmDYsjz3jXzFZYF07cP06HwGynNYZMS5NSyCFP6t+F5x5azk6YMm
/BeW5TKQKevqESl3ENBLicdIo4U3gAlGwxH+sP10jUoT+2Jk7lRQ5pAaBtndam3I2DmYYjLlMb/s
M1lcHDrNOudSGg6AE/7Tdml4ZT6q1nCS0bufruuvd7L0nnKpIO59/eDSrOHjy/ZooBVKnHcw/3UN
pslRjaJJREpfzujCCXuGJ+x+AuTvTP9kftmhgrJOVGNy19mqksycG6YcX5rpZ4P3OpxNpcEFC0ps
kxXa5HDtBBx/J6PyB2ROCNWZviv7BMafLvNM0JpBzyWBArYdNkr5Bc113aXs5LyDNyVe9KxLptKc
q/aMjKS9Wf9Xi9arXgB0NEag9/R3yHfW7YdSFmyWzOPN2NWsuY+j1VozGKQpRxFQe8TD1VUywnsB
3JQI6Q8lMGLd464sPbNshAq3nZ2s7HWHtFpVDlx1PfvK1orzjWeqrliZG2HwY0iZvHghHzh3VLgF
Fsg18mDOzZO2VJMuZHUsCkw0CT95Bf45p0xwjLRED7+ROSpTiWkuZEkiru//tz9dmVg0AiUkYyzu
8AGkuVRdoBcOKD8wU7xbsgh7qO5M0nqo92s5UfWfOpfjBAUfG9joJDNJo9n7e/hWV0HkwM5a1hx1
uMvRuhdzWTEly4Zv9TDjMOAHiXdncQPbsBXIUlzCtsTti9WY3Awfv4n6PUObduNT6XYNqY6pwwKl
rz8HyvwbfaKzh9+WGtKbebzEgFQUz2u5OkGF5nusQ2IKu+S0JibQSWAawobn5lSqHgFe4hzs4AbN
n2ksRndS251/zRDHbn7yJjDD4+aqsfGL7eCo5JNOEUA4vTXg6XMl3bsntkD2Ux3sQyP1YTY9Zits
QdTv8jehDZGcJ0ScD8Ra/wl0C1B5HfeSqyiyt075d/M6HfDnG0gdhCoNxyYY+Y9880/xMmftiFCf
wms5tf/Rzq/ncj/cQvG97ta6Xe1Jon54HyENE/Ey1JKRlA1QsBIIPekZ8AYhZwsersLwT4w/fzmA
C7VEdEGZRWzcYkWPsOu3lahYz1Tp0lInOfV1Tnw5MkL4J+55BYnUd3r6swx9Q0oyuTw2h8/M8CEi
1FHSmLClzyDDMEHo13pVSGRKyBvqzBBjQyLrkWHu3O+Vw+TegDXC2q3NxYni/9SY0PzAYETtdcVF
DZJJpfJGFAiltXCaVx4KiGOv+A3m6470waFSu+symOy5qZ/XT8Ep7xJbtUSKYqHxf3SkbGto3g6l
RsAg+zByVa3FHzl0UxRv8PR9PL2mBhuraM6hvzz4Z4gVPppkIjSjf2NdjTZkCYIiwUX4k6MASguu
jcBPT/2UGYCm3W3QOS25Et/AvZCBrMOD5hY2VMykLwbpZlXB912GD2J+8Lf1+DZDBYEP7/8cJ2cu
2dOFKC4jtx9MSv79z9K064kvWsTqMyQOqjrBzUQv3vHQ6PUPAKCmzW381I+O9s5MVpUh5KZ+8Kl3
PCSy5U+a6A6N6zQAmbiK/9N70njfUZcICXOX8g7D/xPdJ3pObLCFu8f2zKhaklyZUxvf0OgOBu9U
LLL74nVeR5FluZfWlhaf+p/8NYS//KJHKFFQtWEm8rQ2f8h9rAWoiIn3tjZKxJoQyVTNYL/yx4P2
FI+n3GhRv795LlRZO5D1/UjeLi7UxXdP//Ay3N0wPXcHCLS3NQAAGhFCvb36dsZwuEGcvKAUkFZE
bnneGB7rd3IlwGX0tsGiV4XudQuvdRBbgFbK/gXXKI2x7PZSiTU6fqTZiqPfqom0uLXWkIg1Q8bl
0zE65ZLrtaSB3rr3bY8L1+/bdm/dKPkWbbiP+vFVubbt/6BSzfCV7NcZTyoPMXUhy9vPu5AC+c+R
k8JGOLblpjvh4jh2GKDxA5Mzgl8Hml91HeQl/4IepO+7pycG4tOnK9KAGxeVBMltJN9i93/HQ4I+
q9eoelm5ZoA9tq3UMVEiOOGdqKDPm5xjtuXPtGMC1ENDokq5NKT7Y4GV9aA/ulqieMxuM568nKmH
1cJWvqDVk3h8WuBeBS2NSiBtaZnJDck5OO7TYeNP0PHOQuTRgbj7Dx8yO7nHdjLm4llG8CWlaFkX
4LIDbX8ElBPN6a+bH0ZezoT0diiY4DEADQ/LlfQOxZqTpObhIrgcomHc2GaVZkZokY6JT3K9CvKQ
9iigFghJpJ3Tb8671M1vPmV+HWzVyKj1qLV/WgYDk0J86XLbc9tonAOfAT7gzOC/aoeYRszA+nJe
JDnKe4mpt7MaioaLBggsyCQTq6BrNITmuRh181Pv+uLr6IyJrGDyNwkknl3bcMWD1DbFcpxgs1Pe
O4BuPkggmPHylt3VBA2qeLVi868xjnVkGConNo/qOiEvdcRHwCaX4VHVyu5zCphcmogGroKhTmbk
UTJgDVtZIjlfOQB6vzKpVlclRVOPnXiv2GMFh4rSU8jdFabJbl4RroUbwc8iBIy+CQa4dQNfkSXG
AdLPJgkdOVNJlmtusF4Ya6GVA1jU9dbrRn3M2QCrVC88zrejlvXA5z/cNWkulMPLwiQic5vfsJoe
OBjQtQVSi2IPkheor/VgzpfAWdBHb5IYi/5teZ6PzEWqqP4V1tCSTetoJ3gSo/bndz2PrJd8BdkN
c9ANwRLPUkM1itsRLnrpnn0wsCs5eEHDNgoAMLWnIN20t1K6Yf36iRPsytY4vKz5Daa34zUsjnBs
PUVFqMA9p+zH6kMEAAC6gZbaNebDphvd45BSrBJtr7x5PEUfN5LxiPZIUKrj7v8EuVrpCuVt00zV
0rbNInQTU6cUF5jSi2qPvt77FRT/wdQsLJa1z4HH9XJfIetTxFLfce2+CJDid5BfpDOf2zH+KBCf
6PHKY4bqjiRyrRtmhZU1Oe/WkQbB8eY6XewABP4PIa4oTt43bzYl0Y5Xbs2jSS3tKrc5aJamlvB6
YsyhoXIeOSWEwriz0NdodkzXSYI537ClHLHwF58rCLwtkeIVmE5ckJkiCV1UMmcAhqfppWFDGGn+
/jP6NUYWRF6n4hjbl/RpaJheYY8TNvBUqezZfdyhwInKaY+mV8grrw90bKU8WJ09I76xDCeJxhte
5PqIWXp09mQILKP06HF14dCAr1cmD9ldv+di7ykPoCrCRX9GNY+orXyzMM8vlAsumRLtma9b8XVJ
msxaD4LyMvBkQurFkx+SiBwh4ACqkZG1Xyx69+GIo/bVKRSC/EJThL/6jRcehzoQK2WkDpKOIBx9
EX2gAiH+cdRxxCFw1SU2mxbJJwxay2dOeWspYRJNb7zDbvarhd2gCp60O2ERvTGgZ4z7Z3PbNfPV
E7SFNWlP+pUYo20o2Kubu/e95OJ9Rv7mYS0nfvZOOBqLBcQ2vIHKQ4C/s+wl9lMNB5ddh6beDqH3
xmi8pu788XMf3XPGsyOz6WFcN/VpyoV3ZuW/UIx/28I2SuROkE8+BDt8IwoYIL2kHapd6PXoBk0p
G2LYk06aRYu7uBAZD4FmDXjEB21W/zAufJFLpjTBnuuA16mj98r9hQSaO61x4XKWhqWOITRuJPZC
GWGEP9thiZN1j3oRSRAvtd+8I7F3xwZ+foiHQf1QeVMtpDysDx94yDjJtKcNVGxlvfvZnliW3vs5
zxp0c8LCxzvkReEDNJkeoPWm7fMfdbz5b4OJcNMHBTGXxiX4v/CUZ7dGBsNJgi548MBB8blV1jCz
Z8+du1vLOqr0/lHVDV+1+e/uUfLjQn7V9YY902t5oC/uYznp8KS+kqWQ9/smRIWBVheTLkiHWMbi
9DGoP5JEAXY8mGORCbTbjYf8Qkm9jso+JamDsY9u32FaCAFN1LBr+kvQDFfGl/XZy1nXK1ejE/NS
rDg/T7M9dd9j8BCamHSCzoiSRtOExZbg4yD3+ca1C7ULw8z98DPUOuLbRhZcBkeZKIWxMHhppY1h
neWPueo8E8yUtMzBbNiFQG68/UnafJRTdAkbOXoJkf7OnuWCnaGD0httSTsu3svHWzI/GiddYPPv
hMF8KkWNDmX4a4uIBFKsB+NXEE+7cyqG+1gk+jFLFwEk2Qb1SnrE8pMEFPTqOMR/q8vmaodgDIWr
YkfAkJs7+dk71x0FD8mhIS6Itu81ZJuaC9j0sfOodDg8c509DJawQ/7T7EeVlEBW8DxyIi4LJENf
QEirzNaWH1bkSCL275b4xOvaHO3ZOXgO9m/UZ0DdLKyxXiSoYRnJyb7co2Oz8UlpJyGa++H3yJ1N
kfa2zdWUHTJAFJUzKmGGqMcZhbq/fKafczz6jrFwf/i2RzVwxCSj3eUOuhXIaXGASYQ+vvIRt1Gm
OnkXNGDAzXc6EK85mAPYDtBlp2pUsfiGMzAF5aEHqJbhThY7a0KN6+hxBuxwxbPyB8YA6mLlqMKL
PXnYFW352/fOCOPsiaJViIl2v/hyJllQ3YO5IpKS90lIYlr7KaKNeW/JPmV7X7qpyX1f6cAAckTL
wKPx8GINIE5qFC6sWgZ5a0f+s48NRFPqd2dx/59gbb+mmwF0PLWMKFLtJT2/4VF7dR2s3lINdNoR
SvFODUd7zJZrrK2HfShJafzyRDu3W8Ptfigoe6X7ZIxYKchJLUgGJf3T4NFQDFQr2/Nyfbti06k3
ivevQxLmUjw+t0b3RicuZmgT5oFGFF/jLQlMdIYKwBjmVTnwaUg6aHXYPX4B/Dl+soIXCU9mSLr1
9r34lVmSaliEqd5b1MOX/A5TZ/tD1Uv2WkREQI3eK/N2EDNyvXBT2O+xrwk4OwV5Jr/lP0TvLpRx
bpMWuqfaxHfoPEF9L1+nKjJaJCiU9BCPRi4ll47KVFLBvcGpzPpf3hSPCXJNkN7MAqPuGtdoKtCJ
HtpVxDfjUjo0odGDxPiofCvSyvL7cVesepla6Xuv1HvS5cR5BjpQ3ptr1mH4AOaUHi7AQRsL/faJ
MbylTcVxoFpYTtoTp5YaKt/WRtPK78KPx9JSEqB+NNzYVND125ePEF0y0mWwtVNsng/n41d/wMZn
DxRS79ZilbA+h3gcUOIDuV8QdgYR+FojHITk7lQQdci/tC7WnoClV2KPLhwgucZqinAwEtZxLJBW
tdXmVX7XBlBdP9uj8OdP5ounciij+b6Qm5BtRNExriYAhJsCZk6O4PtkdpWNM52PtAESPXP9uVRj
yHkMM2h5lMSLDkx0vsxUpqc/x55FuPJ3ev1Uaabij3EMCZCOcpVW+84W0QksidN8ItN1XRo2VnDy
4HZwAqbM8R8UeC86myoQ2bMmRPFGUYuHKKh6O2slgqZLofGRLI+k7GcI5vfkpr2CKoa4JMydIxrx
cDz2C2+hoMmACq2xQZWse52AHKeLb6dTkx7CrFMVmqIpPaSC/nuloc1AETFZaITpkyVR7HeIWe/d
8RnhQyCIQ60HX+K6TT4ExSOp5+2zsW4AusgMzSjgCsqXGH11glV7Yu3aw56cRxz8hsx3JP02aw+Q
SLP4d6H8cBhmrVPJ43NramJyxvXBTRszo9WZUobLCH1E4IDTpX9F4D1bIS9TWwKn0qxuWlUbuuSQ
tRSZel0rceBVaROecfW5lverUf1VXa7hxB7yJLizHG4AUhwgNzpKfibsZ41JEc9VR/E6orKb76am
s5r9ZC1ab7TnSpYNyXQmSCaY5E7k96GWq4voQKYC8Sgygtex7HUfsjoQBlJxdjnKGyYHV+R2ecZJ
Ms5h4YbMPSd8cDiUymUFW4PJt31pIqePeO4DMJb0VosOEgQHrXk1RzJyPKAdIES2FUkgqPIqRk2X
y7rSB/f2kkBmS/XUonpVGwiR/rWPt4DqLWRThD+qITbrALgaPGue+RWQ7D6DdXeC4HEvSwRBg5Ct
AzqoMTzQGaOiDBjrqKpgPgcgRozIIYbEDGHLhq2QAcMv3zlZWQpfRInsOXfPbV2HagyR0C4cn9DA
jg7zVcDbY62q6+p8qm9aqTez1b1EzyPYvPGGahLxttBr9FYO6MzYD2jbSu3IQQpoJe/WH2sPe8+Z
IckBpu8L53hgdpMJVJVGO0BBlS3JGTLA7VFkRd0vgAXQt/VW6NLZX4F5ygpaLSX++1KyYvnXfK3m
GgU5uLimde/DVfgZ6UewWKVEWuhkcpb0U6Ur3L2/J2Kcu+FOytsU8XZMXyLOnOJZOmvD66uC4gtC
qt3wwr6J30H2dJ6oDOJl8jzK9vWLH2uKp1//k8LrzqpNgp93VWd5TPAJ0Fa7pnBVHWhV/K5AMDxc
BufZAivkkKCfBntG4x79ZFv9/c6RIxehtCvI9WYuHt8BvgaJw0wJIgiwO/mDXW/qxXtxQM2T8kQR
Szfm226SysPsi7IiPuo7yg0zgG+mrlA4xxV1BDlBqKOEY490Z6Ianf4R2o/vMrSA/bE92h2GucNJ
v6pAqEdlG4vr93grvsLbgBjOt7zy8o8rtYNdN9CWSy5EGsybJSaEb8BOZolTWrmf4A2h1dk3XmGn
BFDNm9YDxuFWt7a24k7S8I1C5Shwv8W6PcPD2jcpVajPr9KxmOIzCdjBO4MeCv7de20NSb9CRE5I
CvMThnLR/Ci6YcGGQJzAvDh23+6HgkzqkHwfpsX/3awkneBR6RPC1AqoixJMDzlIuOHOatpi73C+
VUeOOQw3IBieG7jXjL4PM5rMXMTwGPH6EipzcnFNvlCWuhCrNtBvOg+TIFzjXx6vFNvYRYbDHuSu
aEVhVskogWbCQ0yMEs7YMp2LjClSNwTDttvy0Qk5N6Z1ucZE3nklL6Ycst+l58VFOb0pOGGOCkbF
HjCt7+TouDweq1gFOQWKX/gYq95VJihw2CdDD4NIx2UetGmkQEqWV7UwT9Eug2odlAmsHspXp3H5
r5nETP95vxustKn8wjB+Lzcf2b4iRCo2akM05+a2getLV1EPhIhEpu96tojowP+YEXAHFlHNOOmB
XSPTftF3HApRc4bWJ91Q/kcz4ox1ziZxPPzj5t0vgyP5vtNLKtAns71eZkUB9jPldcx03JLWt0Y7
rpaQtEgKxx+dJj3qOQ3Xa9TAH7ZQylUuKoc+ryt7q35DLfaijkSqj2fy0UC/0OeM+TbR4Q5oJji7
cTz5CcLXhODky5BDr4BCZ9UgflbGSj5bxCSFW5tet8rX3GVQNL0r01Y2urv/fkEdQik+LJ1z/e7C
lPaIZSpInubHwVF6lxBeYPRSU4s4ukEASEunZ5c2k4AL8PykvxtmAbHXQUYRKCqmem6euWzTigqf
NsezpMXla2QDe+nV5PXawH4STvBisx7XAe/TlGI7p4FtnfQdB3tza/ZUTQJFlv5mLJPP+2uvY062
wJw4SDxw/wr6sXl59FXxUFkUAiacu4SLqo48rUSsrPoHn0KVv8R57VqyfXAJgpmD+5JpNffN+VPM
Obl5NZFYpkfiT5gphXaoqAMUT/qG2t3ufKhIjdAuyw986hlnExKPLPAM4WuNa4rYaQNyyeiixBcS
GYJuX698V2cB0gbnllLZG4q0d6Lfc2hlFvNenfB4Tna78XdFrWDt5DgrXjIADae51BGrJgZ7neng
U7ATEoqRSt8c+gBBWVVvEk+/UAfN+lQ51/d598GYLf6CL/Lk8vpUX8baqXKiVV0ulA02vNi1Mrr2
G0fyUe2gNZNMoial/eEbthS11OvrYZV9tJfuqGH5d6pqN0iR51BqjsZvu89dW/9sMNhfr8NCK7Of
hzwOC6DCo8H0C7f4rKtUXbd6a72iK1iUYlom9CSfPJfRTRQKh/GkHe4ht2CugDGDqVovr0fDYM35
46F1woKjIHeEV6g8neHtQCeCU9rFevqnjQa8a4MNoTefFk+K5ycX8n9o7DTJ28Zn2Vb90+BAE45D
8QdFuSTCakdVV2E+g1/ieJA2a5/EdZvcM7lN5Si5tThlAeHM/ecHaH7y4bDbl2VANJc0rlw7KMCy
wrSfNZ/2mFbDMDTdBVJrWlT7aS0R0meJipWPw8VItMx4rFMxD7pp3QKa9VKYHuv7Qx9BWE9usCIZ
WSDqc34W1D7LTHRwkT3DFU8TqL2ik9bEklyQhVWjlbXZhlgR1Pi2IoW6JVQyS5HuO8VzS5xEToXb
QHXdrcl8bVU0h4rxkwLXL4QAGjkOSETKPU/rXMyriZB1SW283V5u0UU++gE5Yb9XuDtj71rICTtX
11CqpuZIerHtTsRfGmVL5fo1F1zcB+oa1o1DojgflwOhUuHYVQJB4GW2nAnfglg4UYmbm02HQFhn
aM4Vc3AxgIjS1Usxeq8nWR00I6tY4hJ0LX0LIWjb6B3MobgBP0AwHEI1QNksMlFkR+Q9UPzdLcaR
F1SoNKXHMh3ai0aRfJDcYJZ+l0+p59nff8LW3ExFqoZLAbnm05waI5Lhalig4FpPH1JFIkr+h93B
5xQ9QhCROKb9zaZFzHX3opxSLZejeLLXHutAZjJL2/FTCUWAbQeRfb4w4+8JdSVjQ4BoQjsKblbi
0+25avOpSgNCo9drn1jV3y0OVcK2YQwqT2edWUb/LEmT3xwMXTMZacbkLSzTQbkZfmtpQLZTqjjC
nkebfXudz/hJWPB2lUb9EAjzcQYN81nLhZ6YpbV28m2KVkASHPVzqqafZ9gGSZZJ4nYsghDV1aGO
QAN59ZZXEwhGJLCzwzfzexoLsW4vtkppEUc2QS7TNw6W5xnXm899qTSSUDde3kUy8/NP/TCmdzqi
Q7X5r21uUjVUVjzRME/BZs+e0Y4Nl+UqJQbj5QoXdfH1NDoCPEDjvN0S5MPGeXL7JU4AjBNRRXII
3/+jWaK1NJW8sFETbL4wU8pBjb0HsbM/q1eR26wkQkt60ffOytYnyXy2C+Ie/dz1Sgei57bAmfQf
bv+jD9lsdm1ucisGM4zSbcF63hRzoaXK+ne6FAfs8OPjx4gphsxQ6yb7RXWLgdVFRZ6FZ5+m4NDp
6F1KMAnz5ju/4kqEFLKRfHBm02VlKATDUrOr1us8/Ecv3qWFHLY898OVE3KD0W8tf55CqsX8N0LE
Thbmcwr4MowSQMd1UFJNtpnmKdWLZbiePW46GKpTfFKlT01Gg9K7oVItqz15Ta4e1GAFQIcsSHwH
/uA8v6W+mKonMz2I1WhA5bcg1EPx7X+n2fi5MTGc5SSZlpTVd7vWYeYNOjSxMvdMommENqVUu31I
hL4sG/w5AD0McZEzdA6/laJc4DVxWrvJsHWZqewjJIfYYag5PLoKI60gLMPVGIwd1pauUeGYiq3h
tjXV32m/J9Ibj337anA21hlonxesUnzqsaAcURmkjYtkdvEkUtt7hGwy/zXDzXH8/h+7GLPQEToF
KCJF9ASJrzi74n9HA8xJoVbuWuclOxHF2rB+m8wdMNPdgpFCC03WUy928NTaG84ccPSxptn7ZEpz
9uGxDs2EXd6ndVryzihHtPvAs7PHD6xA7ENbDp+hh3pvMS5IM91MeL2onJw8n092Z18YgO8SGfqz
Kzi/Q+k/Yb4zqLqKr4pM/nW85ByyoyhGPz34YGblPMmzPFmaK7xZXcVkSOY7PzZDDe0tJyT9djRp
QAdpXpZZOB5dZ/T3DMJusqAYyUDhA01cje0qBI2+ueN58eET9hA1/U7jCbegywXH5nlxWMNqNB7i
4wyp36jR9+2U0sWi3h/RJmUMYPVRlYw9pvTrhJbDbqbyAiPH4o8GA7hBhaoe8ujxcvnUm93qrtuH
e4M5wpDrsh85UkwmyY6XZbTfqwBDCFMRRnDRBlx8jA8udV1iuynQbodmm+PaEjzuovn7Flb0Zdqh
1KDKSZdjQxMaBNoOAmncN7BDM/Aqlfy7sAwdol1WjjRyA9pYJy8YLUr/adS8GPmNanMSGV+NLyJv
sS1MkcJukk6ZHd4KCVUvXgFYvwfcIGu35VwICVaaSNPx+Z5jGEv4cjauJIACYHewMbGdv0BhHJhZ
ZMxQUXUdNl1zb+CvWa/wA42ODBf4KBvL7Fj6gBvvOujM9ITXNLGvo9znihB8tMcT59smMbt0Nsir
xDVn87CNFRG1+VhyDq2Prxums59O/UM1YF+F7tVHIgNVAICfpIMEJwd8W0dKCChGWmWU3X6jWjvI
bEDeuCDHIxWjHKW11RNelk7rOpyRlp5bw9Wy+zW5Oqx5bT+HhQgj+2NODl9ah0UVXjdQWU7RGUJK
R4ETcjuS7JsFq4+3C8kDT3YPs40CZVHOvf07s4OZEkQEigMKTT2crEeEv/a+RTQN97YOAOsOw9/H
FaHjHBg/oAQpOt7torNZLcrIvebpUzNEg8JhBjsmNZ+vTFajauUmdn/kJlxY8sdzrPrMhQeCDCMm
GOjZc3PGPSENTTCVMd9EkWkkycF2c7pwLpU4OTEH7+5BeN8WZdMahPbvXlvC5Sn3G3P6ZdOLobNk
Bzpebzw9tWPKCZQEb6BTdd8/riJul5Qokbcl8R7SFdaLYOaBKdura4J+014uq30/dfopPNd7qWdI
QA5xJi0HgqsAQRlea7fnbPXT5q5KyZ1gcMsm2R6qVHL9Yk9NFrQJfDUn26etA2YU8dXN+sMm1XqO
uo6tqGXF2FMISQ2nDErtJaEW7DtdK/QqEc/CM/LAXNiOcysaGe/B6Fra6EPn/T7lovk2vFV/IfZN
juHUtytCPsD38KBXFA0NfVGxTbbM4CGsIraXEfs/yw5/H6jykQpPA78Hxei0BE8YcDphaW18YGYK
utpHsa3f026ILUFh/joPQfJZhBoxtPDBzCzjb/gSQs8XunJc4pSIZHnjXajvt5pBQzLx99i9nQ82
pChCvI69dVg0fIQl8duOe7HIhnIraBiOsECh6UfczgHnNSwMzETjsZ/l+iCxJBzOIyruKjMiK7KG
QA1rjVbJRzGQMuLvv8ZvHMura1PR6WLeEXFcVGEfLXfUcQnTko48lZqRxu7uQ+Pql9DjTwJ+Ep3a
rtaoHALoKn0LxfUk8ekkyvb6AEMhusaiIdvRwpLAh7sDnJHMltOwD8mYxzFl94fW8D943I6BUuQQ
zk9VXl9lqClJgp5QQDCwpRWeE/Av3/T5GSbi9656TbgtYQ+DlnEJmj5NbkV3206YpMM1tm4gFwF/
7EHFLjuYt/+uPAFe8TrwvJmwiAmDIcg0iPn3Z/2C8aMDYfCtbb7eD2KMlUnevAIb5jF31S1AA04e
4u5IqIsG7TQmcaFUsD+JndBk8+/V0ywUCoAXyBRPC3je9+nOe5wwppXplqnSTocpF15A/6qFMc8J
n1NcEigU65XdvSC7DuuvfvEY+G+fqqE9EkMPownhZIzO9u2No7NqKfWm27rsGoaa5vdClPSgxUpY
97Xtz8ldcdV4vIS/vpuGXnI+gwUhGbqzwMW26xRc11IaL8rXhDCXUUbSqyQPj+vk30jLi1/5ki/B
NBPWlxcJrfLTXc6ZlJpKt2Cthyv9ORHCLApwqExbN+Srfi8F8xFoIcRq9aIyDT6X5RW2wgYp7cEk
nD/2JWWarqhmFoSSD07nUf389TcN/k1EKPDt1yItmhvy4exmNTgUs7pPCBpu+z3F0lIR4InYbxS/
GOAonQ8aMr5QxXUmJzBHUN/udSpn9Je0YbTqJCT8IXMQX31+mVhWyWrDDq+ryJ9lzakq0lKS+BE6
7h5aG3p6mwMYFKCYA0BSPxKo0il2Z35/G37rJtinkCksC3mIe7m7l4frmVkUinRvThEc7q0pW+kz
UozOXcDXc0jPjmZh+IA2USkSMBR2iJ1xfUeAUdkCijv61ImRTPyOr+Wbq8V9gOmruT/WqsDeuxfM
iO2oEo8auhaeHpT1XMjWk4jDJZPQR1Rn/Lyx7bNuRPDUgbJQbhG0vvV/sSgvqdZwnJOpwrUs8NI/
Q5XZYvYX24YRuJhy0tdvQbqGkFZCYlB89AD3P4CuVQ563rqy+cP9GLUEL/O+dCVxysjaw4Q9EirQ
Bevats+TuknlPKRV3oz2ejKZErQHroKmMS2Me31w2EdvtEjfTjuLAfdcuYvfnA3Qm8eTHgh/zrg/
EM+8HLXRkmhSGvptQZKvdx8n0uWDvVQOVxhvzgt6GxV6jSDPw+UfA0QciQ53jQ8d9ZqzxeU2O7s4
AWkNl89hhhUZ9VWtH8oueA0EaK8AP5c+uFInH2I+y7tsWrjfJPeUQyhPIqWI1mZex5ayWmE/sDb2
c6oW5Fyhz3EdZxi5mA8XYeoBFz/7gAH8ptnScAVAlwiIyqXZtNHGxTLMuJ0K0nsCfsXeTRd749od
BqD/Jus7Dk0O4T5B4hfT+MCNKE/+LeL3J4Z3qmWD7SyZy7eL1EtT6BKSCTejzgZo1Db9SMSvgG59
udw6hiBJF37rqwp9L75VTZGKFvEmRFRYwTTcOS2ld/E24rEfYZbq9Dd9plU1rl6M90oWmlpUlvck
psu7/+HeO2Vj0FGP3Rgis3RH3r2XOuj4X6kg7ueWcIH/okBdhdzKJ3as2UVku0wypdCO+lEG1H8/
kB8q0CQJQ0/w3IOl1kUjUM33OhGCQXu4znUhbNlk0sd73cvbdu/oNDKGb4SW/e84DLmY/z+D1Qe+
B8OfUdFeZYFdJPGq55qPb+ZWiGh2j5vN/h7NXHn7J5OmvkzuyFkgKkOujh9AcsYl7wrQa9P/awRH
dON+ruFg/yxSk66YdzwSMM5F2GlSYtuD5OwWeOuvl7xnEba0Khpf6zWfnzAO4d9nuucxCQpy8d5z
1p8K+LZf6y7t2HL9E4jjm0jYLixeo++VzH984FgbpEcEOt/R2iQ7jQSDcnC+zlsmKTcwmYs44ZUP
6NRjoHvLPcO7YGxWegFtnG30f33hNjQB48vzdlp3t0OUYZjIACebC2m3z/XH3u/45Zn2FhlICGKc
2dXVqyCHQTMxSb7auioGc7wwPbOXuiWes9z/x8k2el2lS3eLeYl3Prw/Bk6XadSTzNyecgGCgWy7
U9XrcL6Ws+GO4v1sGr7tsk1PDers/wZFXi2K6WulaZsGMpuISbTjeUopbofr8EArWRTFBPPg6YMn
OPryZ6g6GdaA67babC5N7tqgDB/mMEugG3Li59rAwHthuDXEwaA0kj+rwO5J9BVYJ+rGog+VgDD5
Ov9jXsrp3SvxhtYf8Q9+buRnETj+k7XQgCnp67bZiGfjy1f5/ciDodY02KNGkjd/6FBYnVhfctbw
JWWJl29HT2Iat545jobUcPGFosTOmqo+FTK3dGlwH/DFptQ8pn1HfIgBvvzccpeTG06bb7VnIc/l
hFRNTBaVcX1zQA43cBJqbbbtzGl8SXsOslbkrQqL7fgzThhI2oy1DH5duiOLc01hF4bBVkTtjs1O
1S6zdyCG/3RFpsWri7qxdB9fEtoNCXc+GRbc9q+40w+0RAEZIouDBm7IY6+sLSHFAnIWKLEQtxpk
oHFFQSltvwAQwl1t8JivxQqNnD1kT6fkY/z9GiuJ/37QZxHZkBDoJ80ppLRAB55H/dNTfDk4Afn3
Peky1S731T+NB2gRcrll1dgSxsBD7QJE6wQyrEZCvsRAO5IzrvQ6MrJ8ZL8y8CvBB5QdW9reA8EJ
a15EX66Z1Ccoc9+xR7GlZEYOFdAlQmYuEBsaBowxC0mCjTqJu12gpJXfpGTkXKkUV0t6n8wqJLVq
qRJWvXhHweWadyF9MYC6k99KWqyVQta/iE++6RDQxppdmgidkGhilOhgDpGpMNhqqAe6wIQ0yzNj
KP7+AzZgfpl9LpS8SXZ642qrF1MgcGn8Xb5Hvx3VwJqxYPBUdAM+pbuySFy7XM/G3ct/Bf6Mu7Iw
DbDGg8yG0CtnhQpoKusnYh03pDte7QulTlwM/lZhnITzSyyyEfsEdaYeihoiKFYR35DJq4Nkhe/x
o2LOwJGtJ3Fx+ZTePujqqes6s4CrXYwGMDyN3UvCW6h69fbPnOHvNqDlapV7EAprOrMOldkd1SUE
BjURT393wfKiBI2kwLEpm0OcDcf6pe7fTG9qXFs6cAqp69olC3jUi5IIN2ggzb9KZ6YWkYA865iW
TPYrP4iiltOmg9Cvj7WAA0BJWIFUMvyY+YJswszirBd/iLA0op5amKT3sQT9lG+8n6atnJLEVYwq
cRDKcD0posHB9kNsyx0eym1RFYjYO9mKeJj5L/rEhLMixPIcfzEY03GDYJxw8BoKP8SndbOkwHhH
WOTW9UK/qHTxXQzoc8YSXyK/GffJ2ksI9Jhrrv5BhVqXFStYtoZdj1lijuzVsdcwP/D+cJjaBLRP
8q7Mnh08UeJkI121Sz9ku7Xi/C7Pyim6mF3CI8bURMcKm5q0o3px5M+wpbpNV1qZt3T85mpeqLmO
jNReADhez7q5gJ5CLZ/7LyntEqfw5dlQ5bXIuplGcLxwpdZ/uHxj8QaKWz4kow67xHkDtmMP5QJl
mtkm1aJ1CUs6rU1JWtyYN9c/AV0upp/CUWkbFMxcGbl9E1erJ9af2V5XmVvNbbHp3sVNRikpXGhh
G9IlBRqa6IFFrDk/h3ySIqbVinLVhz/JE0h/9N1NlkQ9+1eDk4gO03JT6/sbqVJ/WLNV61L77gHQ
F9x0lLHz86oJK85Bax91znfjzZ6AQvZjRFwchZEiMbMx9M6YK40Pc5RHfcHoulxnrDhooaKzvcfG
CWT93JTuJ4F1onQUEseZmjElg0Xlr2KnmebChQi1pweLry3taYwO5+Ebqi7Ejo7arbZHMBKtrrK6
NPwiItSxZ4E2+F+PEx9zdU0cLADBeoODO+SDY7tQixHxr+OTBM37U9lqnA0AVYSXPAQyFa6oSso5
GsYJ8t+V+QEnp3cZLlE77yLE/QBXlJJOCusuF/2Zm+bAwg2m3CpQINcc9WTBiuNuaiuOHh9t96LS
ElDsQgWp6U9blQjV+6N2IR0OQnA+Qhb2YmhQu+Lf3rlxpua+54++D0NmZFy8Ue/hvX75TJUCcIFP
FoIvY3wYTHZM7fDOEfaKZh4iIV4MixyegPB9E3DUqQk1b5R9X/7lpBTVtmav32Bz6/5a0qB97fUe
9LBkNGu5V9sRZCpdc5N4yMaz86LjcG6XKEIpfX6vy1tcEXuP2f0sJ+qldxMRYXQ4zHHb+1XyiHoK
bsTbu8XWeaRfPUp2wnj2rnbIKNWZafjruIEtHM35TAV0TePwm0y+RGM58cLpEVFi9wSb0sMeMCPL
f4sCKN0sCY7kH6ocsfIqawHn58UrEU0lsWnS0GnR45AEx5bdvF/kYe1EVb/N/F4HGDsBH/6XgJiA
gC1pNEHD8NVmatGoRYHyFbiH8RjH4Lhbl17UfFbu89kmCHdMgyal57heMYFNX+bX1Pi0Sy34JKG2
zMkjacgUZzxsBg3UkfnLusJ91Yj/czveF2RveQtCAo3OXIpKO+0DQKtlodi8M8Xabz583H7jMt/D
zuRxDky/dYlJUEYYZYwJzfozIWZhn9YntqqUuBK71axeuWlXenCdjCvOU9duSQKn6NiqMw9zRqDK
tgeDSq3sP19v0Npz1uz9N3jYb1IClXorhzaftl80H1bXo5V77b28VK0a33FwdddXkvrrA6FwKp01
nNGfsZkdLt1kFaomWzRM7ZbrlEelKO7psRrMRhZft66HtedyX1g2Pa1Pn3sXlRW+6rGzDAthPwSt
516Z3xzzbN/noYF5Uz0vq3h4PlJ0fGMrxvxUguyqbgZ4KEd06T1Yn1+pyrJ44rNwDyLbpB6L7UrI
hqODpbGmqh0gp2LTtcBeRDzx8GRq6mWDGFBEKkXmmsOzHWEArrTa3T3HXbPuKjmnGIP/2efDyt6j
J2fJZRkB1vehD2Dz5rbiL6FyU7+3D/G4gPS+pFao+X76Ml/8MrBhJVuQLRm9MlqdTiDBLn5+OEkH
GovcUudDFiKEuvF7KE5ZbgEwvdGJEI8j02xes26am6vCwkTaGhZy1nEn40d60JrPY0Xh9BSEgeES
N+xii12BfJFxXr9/N37dimb3LuolQqtq6EMou5iVqDo0mfM7oJKHjdVwXbBUDCx1nNldsaZCMH2i
/lrAhei7aBcI4bhT2VUpDqe8n/vTUPm6uDHcOnkrMMl3RIXoH2ngIDnyuayHCEr6kEPNAxOQhybm
z6JPvcC0DT8DJA/lQW4u9PESmleOI+wAcCzxQjJfHL4Sg7WpK9cGBdnB0S1oboxbF5WCY2PPjbcz
EdXue64/cWyTar6t2sVjecm8S4nWRb3T6BKq3lu5QFQlaJ6lhUoyDcUjROHmVptMRxqNUrcvqamc
BlSJybN7FWvXasiVxIQhm9QGtaKmf6ux0PFhYYbvD2k/vvdQl2uqYvfSDt6VBWv/wG4OOiRYCeh6
Pm2t1/P/EO8VRyllbTecZ3IErta/iOMuLewfT9LLkOq+6doaaRmGNyBqZqg1xD+lW6MqrrjSXa90
QQSQniNu4MprZpFWHOCgsCWqCln4jPjXDkCjozs5iHbaiXfCqyrPCTVBwfgWH+725cQDNF1lUXs/
d4OT/yDmR9lTEwZizIFRoFT2OLps6qY2tFzCcQ1O2pbvDypN/JrQYn9CL9BKbwTUnSVlVsS5BMum
mgCPMNA2lXhQ3an9bWsyhRw4CiYFoWlSJ8gAAdeIr85z8WLjSvL1mYdP92ZEqGZI2ehbJ8AyXdec
B9QzlbDF9aZiZIAZclYD1fwsOAyvaFdha3d1NZFNpYU+Mc5Gde39OvuR3LaPPa2IrajJszypFeM8
wGVIBKr8/DhYYdlFjSK84X1G7OcoWitzZH4Lb0oiVQn2rGdhAuR8rGNAE61zfQ/B+ltJa8lB4qYP
jAWuSw5a61c5xEfqHjdcofmOKs2lAOF9vUQG0jaORtmd9/QcGG/J6ftIl2iaN4yLSjuvtx508oIa
zUGl5jgR24Iy3SNE9DwcL5+qIkSS589+xndKFjjsAuLPDWkwHRx/+E9K0kqLG1AvAksEdL+W6KTA
J/DIpAA9zCDa4Oso38J0V9iIKfoRgKFCMa6gpJD8IKWD2bc2VaIOPB6pSTGIa6X+jXSFVoto2f/x
n/ML61BNAlmEj28YPcvirm1lcSjAK5CsEjHRqG3cQk2sU3Dt61356HeEAlMtyowol76ZlnB03GmA
pO3ww6yHxC3CTzrPaNvK6xxlYJc9DGuD+WUslUApsfhqyfSr0CiDe86ZFok1xVyoUblpAiq4Bd+E
9qD2pdhcFGV+S9zf9pzvPZOXdjiVC/YNneBUv5CnzOS44a1Ronu0t5deqV2FK/tpQCCXAlbjZ3Cb
76SLjxN7tR+BiwdN4aZo1+NF3dLBC4vuYsf1n8tN1kl8v3Rup55mqxyeQhUIYViKzM7vv1x6WW/E
6+oKjQaA32Ja6BnWKjEnYR6T9cN0v3MaNH9Cbuho9Gga1E4GYhNA2VaQarqn2Bj3k1/JCPDD5zV4
NDarcUpVIkVVIgFOBQIYwD6+21OejrNh8EEBkFXwIYX9NGqEpxwMM5s2AKv6BfBI2xSqwdNpmXsg
ylhoS7g7ilr8V+Hmj8Wr3w0YIIC0apykasTiX65ZX56kGfeiUF6G6bwP+26oah8iaLetjvoFiTqB
lktXPfArdXetUBeB9XZ0fukwbs9gwKhD+aB+MAcGFniiIWrjnyzvkT0i4L9VFIClCx1y/U6H6SZC
frvOgty8j1wWb9NJA5BWxonDN36425C+ZOeFcX5RfF9PMVTYcO3jGVG4RStaCHvHkZkUoSgv8Ulc
Jtv9VV64nanQrBDuMYQ0UjzgpjQZhCKWGDB+SSPKDXPc5MyNhA7b331dpEmHL7FUBzqq42roGJga
GbvMSlDUKwxUK+Gv83mWmwuErHp5oWmIXrSsLpO9LQGWZn+F1+0mwiDWbkZ2mcRGviUWmH0wXDri
ZSK2zEEeWqeJwIg1ItfoWl95+GfK3z7B73lOKBsegcRXDyxki5HKKz7ZgC7LxMOqB+sbSeHtrVcY
mQKtWuD2rX7/V9GSziL1wai/wptHCkKeRMwhuVFVrRFtXufududB8whehytTFVo7JKkU8rCgzCTm
fQCshLzo7DFv4mBll9oQ5uyE1621i8segK+jhE3iooRcYOvZvJI9YwZLh2OULcc9AhMAZ0059FXY
Kh/5DzJi5EHWMPSalchYicwT2NnjTRo3Dc+AU1Ksclboaz5/1CGFV6Z4EvsfEbGGSf7XMrwFe8t6
3c71PHfDKD41SknflfZ28V5Y1tCNUQW20RWgKElqAaaYhJjXGNPDGLnL39Di57RM4866u7cN2x+/
NeDy2pVNEAtv/4Lm0J4SS2v1EYZHpnSi4WRB7rVjuOxuCf9siATiPyau0T+7eCDi05a/Ig7SusxM
Go6kJiS2RyWSteKA8ctiZaib6RMGWhM1U15q8VlyUfgimUgsr98u/t8BPVuebB6g1+C3CxiJmEtf
1wb2Pgug7JJMwZ/AccL+AroAyi45j9I42LbtG1/KwU8s3VbB4HZ64YMHzomEsW26bEF/KVLpS4Cn
LB8eEFUEnXpAVx8kzcxcYUNO07v0CWNqvBT2gUJtoSAd/7Bi6Iog2DGysRpcSZsPstLQhdlnBRom
g1WdDjqHfSR48NeEfTGkpOVTfMKk624+iTwDsp0jWaeMNMA8LM6s2pn9kk+o8sz8ebOptjCmvjuo
X9OKejMzeD/7d34ialSrIetJ0kNhABDcKa6pHEe7f7WSFIYLdfU0iwwJXvjB4FxUOi1y9U/EZlMc
YyuUpVwEsVoKqy8djOSj31QVz02JH+7hMEkn/WXOBqESFm7zdkg4NRFBT1hHFxvYoTuyZVFDz6Wt
1HrUMrD8JVKOwmxkkjPteSByja8c9mc0fVSGwpfSn1rP+OIWHb7Qs6ENEqmUKG5RcHnsmyuHLDMF
oG+haEVZVe2P7W+mklTHBQOAm0DpNwC/XhNi1J4AkWNMNbGGkAopd2blNqoR0wHqZjtBzOMWhEi8
gCrn2vVJh7E7Jg/MLf8pZFR1kt7UHbKecLxECgYDlhl1UX0RLk73KmFb9T/j2EQuvpPc5BRXUg9o
GaGY4RzsSDp9zzesjtEy315G1Y5D0POnXEmZbGJsrkrKNNwtnX4ATZ3kkaQZaORamA2mQBKWeiEm
zBQ38AOSzeZOCKd6ojIqoZ7DmvXeL5H93cETJBQX7v5FGrp0Vd4BSLJ6Mpf62DOxFug/4C3KcbOC
LNhoMgKeUhGXRhKKXI4rdojX5dlCEvEAXHSEmXyx3wLLOMbAdcoo7+zBlSe9CLmsdNcqjDPkDGa/
n13tFD5nOx/wzGjxqq9rddzVhvLN6MqJheN0l3xjCDRBBXyQkzqgGCLgLyDq64tMj5ZXRU5xAGCC
Zl3fsrFuHwRqXDlXKEVtMDvcclwydoohyCIOlWztgWU5R6CI2GRn1c4Vz78Llcc1ykzdCZqI0E/s
uQCtbrhmutQxbckFIHiqxA+VlGRW52BEgtMleSUBIsdFKjwSh5yCP/PndQ1fgA2oO3nzkpgG+MxR
1XDuZh5z4NO8p55wRKKM/niqrS1tcA2u5booKbYFXLO2iFhN2DBOfVqkhFjbOBx3WDGjpkBclisa
8mIGBaA+jW2A5YC5aVsyfuc8klJDJn64Iv45yrlADMt6cjm1SWD+jjZeT0sMsnTeBtEAzWl7Irej
21uocMwEPQxoFB5AW2gyP8YGv0F8a4ZCLPYI2qiXg8yreAJxQKZf3OJ0+KhlOZ77eSmdZXkcCuZl
qf9rPOm3e3PFj8RbvX3qN2spBXhJdgSbS+uyVN57uu2YJw66g5xdvZKiavpUIOJMpRuPihCEPOgy
/PFC69k5XDCA5a+IoaYgffrhYNXFfHU+FMixHJLz/wWMUJwECMcMTSGAdSIDK6COFyCUtwosVfoK
aEIwasIT0nUKIWwIYFGWGn2nU6C3jh3mxaLHUen2uU1UwEExPOGPj0N1xVONz2CS0ILjqX/TW64M
2HOfItiFvypyBNFxozX6oIlvHNFPxPAWkB6fExFOnOrXWTc4jIh4DERxHCeqc6CTSVsZ2xc/xO5x
PeP778JQCdWYnHMQyXLs94iOaqSdfV9AzjKFwPdmExhMTN5EmhlIHuOAKFM1G70lTw+i6Y1laRMc
Id0MuUXOvGOu86yaMyGiVh5HqkEXCUbpw32v37KjFxhxDKCpA4K35olqS5vuvWEM+FYCFBs3Ps/e
JWRfTdCZxxMDvOv7er9KVaIRh23bUbWpQcPJumiex2k5ucGU7BUKfc7cg+rZPlqap2Jmd+xI/z33
IJJJBp2cIqY+7ocbTpTBcjb1UeLQjaBwW80fmO41g785Lo0ZWgcLVbO1TDfHIBdiAwShoApM09Ze
aveju1/yQSNyYD1wPokUGv+ulTPFR9qRIkSkwfQfBMXJK289XE9/AtikEyfOUd0CLhCHNrwNoSLK
6vVPF+lhV8CzBJ0mGCy3R+Fi6Enf8JjVewYbnA5csvbgWriuxmnvtg/QP5tnJEkKrYW6z6wDCYok
0GjnSc062T/pfSLY5VZ1ytEVrZf91RsX0ihB7rsX4zK3G6vrEpvJgh1/gXSX1Uz8rJ+H/SHtzyPj
RJzUdowX8tClPZEMzeQLRRWtpxx2o309Uo1VsAuxtSvT4MvXyPZjDGDnELb1ZdA+1cwTkHFPlDhv
PBWbpPTzTW21hhcmqmUaj87GlkDQWk8uDhcgnUcWF+IVHWpQXWbIcXtFDDoFMwK6dnSUwSKaXq4g
bzIpGy79QuCFUwkiQ+soZU3f7Gn+hyEsfixYMbLs2eyFaD1vGBmCDLcwmuq5orzwVd48F6h8U13k
HgiQLyFIdVYQcM2afUxQDq99pTLfJ57TpwcQorbUAcBA0YY8AMAk+2DlWx9uq5dQc67k6wwV3WYe
bL93LRpD1CzX5hctwRGleYUcwkl/kC4XNNdlu1523R4il4I2bpji7yxLCW37kLfoLYrwOuL7QkIR
5po26l4jbxL0+C+nYpu+PbXnuVfehP7jyr3ke/xdo1LeIY9lMlv/6Z9DhHpdPgS5rwp1icOGCtM2
HzaTf5TjJRZVcrUnLN42v8XTisOwRLL2vyTlt+ltFph562Uzot5WWMHa9tUyyvHgEucHEuaAfGDc
c86kmbs5Kta8xjseqx55Qj49dyN+O4rxIdUVs6oJbJxeVno7NlfR7nncyMrtsqP+TrpEEP/rDqi2
P9FK8Y85fPnou4Klarubf88bKpPmikcimDclHEHxvI5ZO8d4s7dsgaD6wCIRSNFb/Pa5PHfMmPYN
A5NFwTgo0EP1KjOSIVqHN/v6UUpzT8ZNJGVcqH3+NAfmkXLTA1KzEQm1o2stmtopnidiOq2E17Ar
TO47/L8qZY1m98bXYrFyAQgTM9HFUX1Y4hFBT/WG4WZWKlz/mQR3BWwrgPIE1+KiJou9F1Tpufli
1gMHV1gphmBlDdFnRjbhwHGYSgw0/nRbrckH/abGWibKlMtvLXNRO96l4r9P1wNZUo7Q1td6++fw
lxG06TlIdbgx6R9Cwji0CezbWaKv2QsQH74Llw8rm4lcdnyw9pGiG3g7Uhwjk15m/6IEZDmxjmIj
zh/IDzs8GxyFdUYVX+Y0mkobifrXKGYH37ZdkjESEl+sdxGGQtX7z7PSjlYfCb/BoqSTw35Hmv3M
iA0cAJ0dNcRGZoqZiD4byqI0ePcb2fVRAdWmS3Bd6aVvJqG8n19vJ+nbCjk6LNFdGFklQwjcRSFb
inK59YQrm9zb3YmgSsI3PkdhlK9BzCoTWNgRtK1h0CBA+tippqo5hWaKaig1DWM8I7HUJx9Qsv9k
nfaNDgB5yW/TIrjdNcrcO/Ye86yfHNDtLDRcOzy3guAVRSPq34f5UmUeJpHryTZx4eJfc/VkNuvC
C0EykTQN/hAr59qUcJCh3XLkiqAAf5g6d7qbkFUI1Cb5f3jrjoFPkhIuu0lyJrluHe5f2PEAO1we
1gDRQqAe2U0lll+PRx6fAEtaO8q8aTb7lEklcig0yEhK2b4GajABbCiZfVUky+EAqU8N04Ua98du
9PsY6WDGAs9aoa0DO+Z89/MTIq896RCQ8wIi7kav67vqfXrtX4wypVK7hsBkOmpviVLmEYjDTBYp
zVB6C62gq2Zm5MG5qxohS+gxwEpVcLIsWdFJPrNV1QpveoytYxv64aSiOcrWM0qMa3J5iS0EVbCi
m+bJA3BhJ6gp9Efca0OgdN9e1HCIE5mRE00H/5vX0szN3AyBT0KonMxNvmU+QnyBDIA/R7rKuVNE
kUekSeUsHgngyrkBaNVUPWEq7o/hE5o8Yjsl/ViJAqXLJJtEK6pZf7If+7erpi/W3ol/q0+c7rCO
8Jm721MJ79+ncu0nS51Rx4diwxWUqTZ0TLYfDcak6aoSd4Pw4ctsDnQmpM9HmMp+mwT87dYoI8q0
qRUgKoQ9GDpUjCX9FbdylUA50MgtSigFT1dRyW+t/M1SJb3H3neL2O9emAfSDH8ElsBNzCVxA0Om
ybIJf6I0DB53QUIdEhEe1TjT+PH5GMyf3JG14svSuJNioOVr+fuOTjFMfGH5fdTJIpHwFFdmvLON
zv3IQ2j+LtK6WN7PyzNM1BGov5wc0RvtMC2TDJqCO0cvPi+efYNSIQA9tRl/PVc11Uo+1rYsGveU
pZNgSS/S6KQHNiNPDg/1nu5XgyIFoM59X4wjP16vk0TYr5HV2ieZN+YSBPaPHocCkndeBq3MbAnz
ICV+9DXPs2zAYNqf68zuyjnZYuD0q7BWHW1gVlNBtufc0X4OlpDcWqgdBhBz3pBSqIanaXFSg8q6
ek4gglKeDicQpj2wW1srg9+ngibOvMdKw32pIICt8EtF+F67PPZADhZ5AkzSg4jhD7aGR7FWGf8p
7s9wa/0XEygUr6EN4n3XHZcAD2BGnvu7W77sTRzS8ODqcRzEz6wRrtNXMiATSVKFsh1QlJi7xN1q
zvqIXedFBzNTvfD1sGEf7mrgopJX7Q9VeGTl2mojqS43iahBTAdcJSp3+XtFGKfAIubhBVoLDX8e
iSy+hFpJKt2WaBI2+g4pL+a5vvrgKcJMujuqN9Ur/TAxa5+jzkIRHKNuigafvILeHhX6kH+CFcVN
8JOztWncs2lnwuaJjvTJ2MAAa7HTS5IVcV64FXGWU8zbAVQHAUtbil6OFZywz1Pv6mUwM1RI+qN/
VNz6rWxROLhPf0U5ogrh/qvR1o+XcvCoj7iOtAQ9azrrNBKibmjkwRNbMLSLYud6K9HOhNUse+YV
lwVknPsrVtrbBF8DMJl22UlC3sREvwQRNqeoOgh4DEOA+ge78yWVyGKE48N1/hGvGa2KGJqLNHP5
wVz45uBKIRK5A74JDtD0JjM4XBD8oQiaZITYXNlgK8gYl7ZJtbaI0aPuduv2TVVpeD6wbqK09rTk
cun6XLO1I43WSRUrEqrpruTInULf49ya5zXMp8CJRMss3WIxxqEYDupcFkZ4O/CKbo2p0h6rbFLS
bQqIsGwkIUjcgJOGrR2SGgM5NboB0F2Nwi+rS1FDOEzt+U1ycDCllRw4fPGWhyuH0Ie9m1SuQWc1
lmF3p6+Ufs8wtNxW4m7LejSiNtkQ9BG96D//jLxbHXWcaIdKu0EamUJtuzyp3VCUEAYjKjT0VJ7d
+ugnTDLu2a6stmNhhbiMklNLgbzYDvUUpUTp6+jXTYAPAcdSd+Z4LaD3rrYdH0dHi9s5JQXCQMI1
OD6ZWvn06XRaF6nLf2oeYk0e28b5Fj2COR5d6xYhlef6iIO98Zqn7qMhC4BNCyNw2+fnu8DGK0PZ
dGLYITfNwpgCu2/H8u0I6cwosmDExnDfkVbk7cAGjPyBGJrjQ/avmQlDMDGj5y10XMBtBhQ2mYDX
SY+xQNCJwEBRDsMOPOaP6NbXOYGZp4IWBMZUAZrmr6O7/mvI0zmSjUTZgJ7YemTevGpUMY3GlZYW
rHXK6nMmmIE4YL8ZUJzPbj5IIOb7QAUDlVB+Afmmo8qW8JZyk91rWgrDL5jFb1xxlvUljN6U10EF
P9ZzQWIeq9a3GyMQRW/XlUfShLfyvrk+i65Dm7KW2aQRjWf83lso7NxCCIdPy7Jm6SaRkeAPY9fJ
OnLlJncHrW/WJyt9jwypdTFk9TwCnaz67u7cRHDSBgf7n4y1AroZiQDNy98hNWjd9Ft5KxxrZBuG
NDPcg9EaIhvdwd/AoAVpmze91Mx1Vl6AiqEUrny+p2zsGIeMYYRhJQxAPjcl8u0xAtDbPweoEEf4
1y3GU5l7gPs2e7bUk9Zt1u5ETlriMBIhG4NT0lmtQNNcC/QcUpdMn0qWIbH7Gb44tpr1wms7SbFq
m1PjkQMtEWDdtG5jDFC2LHcGmR/6mUZ+pIBrzFToDNqUU1pTF2rSeBfRti1x8ppFDyWj53g1heRL
cbX7qEhLcnxZLTbBlLsUVHVFpIyICX4pJUR2wMkoZFE8ABgG2KjU6MisfCGnG6DWMi8NZmN6yc00
b09ezqkJKG4m1Mg5tbNNid8Cy2wWCAMLbXGs/wyKZFpJNNXHMQP6p0PQijdTE3ka7RXf0zV2hqYO
mdfh4G5zfSierHXvWxMMC2Fr9uOz3Pl2tmOgCIeNz/kuRkHIiy0u2eQeb7ZZYpGIgUc5x2qa0YGk
oVWkCxAMovhduLJuiBZOVdcPv8WdpYoEw0w/hMjw3pEhY817b4Mg/SX6opAM6qqoem3xuqgqMSym
ct/8BbCrXgshofTmw+opV17yw/u4J1mD1GSE1Pu0QMDiV1Wkna/3JeBJIRB/0MVp8WffDHpR/gXJ
b6e/p34nXl/6NZwtYW9UY+g8wgmc4f5hsyUTsVRStV8KUMEYWa76U8LxzjIWw1g7cjI3BQ89uLI5
LncGIg8UM3xZ+S4KD0yMpPcZCFBJc2Lwzyp9/5Ksfstd78/bIJEfwoFu5lYuxaOnEOvZ4jXCImPx
B/CwrkyoIDw7sFkGxo1CAIH4qn52lvQDUqpZ0wQ29A6bCsCtamciSHtKllzu0Ta2RCEIRpU1VOXA
s8bM/LwllOf2a5A1lQ10E5k7HyA2ym5S89H+H6LL/3zuokjDxMN+xxVSNIn0alLwQUUNeMQEB64A
whJ7nSWFwHWpdfHZTXqUZPNMxWnDMGYagbv6JtSLKf6zO0xp/J6U/GLVWDBnNEkzfNFDHWcWzSm0
NVL7V2sPV9qBVO6ga8K6ljiNCJ33IceFnNRzfOvFdsxNjB7QGW5REAOWFRyohg9CohM5i0IVG9bL
wvNJypTM0dR12nDcfZm5bqOvOvskAPSTsBvH2vynRid2hJkmEi2cKtX6U5VMTs/2coVyjTn8wX42
dS8CQPropwWEUsz43/DZGWp23OJVqYzIqpRxtuLFIruuWpMIjtBC61hznO/BUqcby8v/cjF7Llf1
yhOpWBINK7pj4AtSmMv0eza0vn5lbMSs6nkGiA+nvzLL6iPA23sKcPKf6Tyd292JSFkiI9p236G5
H/98yI88FdoMn8ZeuGEPcf4Sim8oYvyTwOfj7o29iSfvaFtn7eGZy3JAtXjBS4lgLe0jBD+aYIMo
c9gbM5/uxJ8ucBSXWydoTDgsoMklVdlIv65sU7696eNXpFJ0L2XDttJtaYg6aqwqUM1GND4TM7v4
eteqUeetfAY8vYixonNTwvP9xJ5Nl4+j2ps13ZoJluVLcax5Wj6bkOIMWMzItO9zgCgSKojcizap
7GD7HAeQ3VBGtAcLRNa1NUzEISbh/a2TGFLM1qiUiWPYNB3U5ArJjMbN7upXThDDxyytAjAgPeEo
1hZqqsGCnVroTYUYOef6PEg+S6H/ipMpeH7mpf1X6GElgW91j09V7YGgh9555Dz2F58tLZ1KycdA
MSSXGYxQ8nsfl0EXjJijgyeQBf/0MtSKjSjtyk1jM+dKxXthopSsJJPgxzPMUgWOLwAkpEt5oC5v
VYxVYw0gt8rXCyaii0XByvWZHEm8zO7YVG3/z5hWc9WRH280DUFjUatoRjVLBOr94L0keZK6moPn
XcopfMfkkKdRcTTuqkYQFkN3E9fuO/2RjJn6huq6UwNcA5o6hhoqMcsfHFgIj96nJRH2lFgzBqjX
YiP2hX1cH8O2pVpuDagWH0SH6PE2IhDpcngXlDOzt5SYjINcjHnQ2yRxWhME25Qe9sNeESJk5WpR
NidRN1EyAhoNpLfuPLJhAPdHNDirdrSs/UcW8tC3usBSe0rcWIlW/OODEnrsNDp0C/7vtJGjCBsk
CeYuU9hXPrqzBaQJyd80dVRvtFk+LD4kBNFrTnydl06CAlBlUa67hEKzUZD4fnwrTjWXdFEmpDVA
hA5eg1+I+39BWJ4DkVYuLe/2QUZEVc/rdlX3KMC71WHOBWBifUNZmurTRtSLig3BujJWWdxVaw4n
j2oZOXZIgFSPPFrd4f6ybGVBji75MW/sYRnGS+pQUq5NeEr5UMzTFz9k5MSqJxC6HDDS5vAEhuYs
y4A/wKv8T6l3RP1C4jG4kj5dFi5DOQxi+yhHUgWzqQ5xrUVZm68HSbEx7wXe1vWGRoXmSzfX5wW6
8HiXKrAemE8610C1RMNRwYXbf8K1vVe+YBsbmBmSkJQK5d9OtLJ2VFEO4D9/hEoWmJ7bp9u4wpEz
neuwaz9KJhnuxZTHid2sgH8MuN9wGQr9bM8+Rk8VO+rGDIc2vV/70SMk3bTSkBRHIcne4qXZZqls
3i7cvZcugZG0fhSeKP5hltXY5AgUh92CVNmWhLH5i7K2E7tdbg7ILujLIkyzz6WYHOoyV6tsz41i
0zlz+rvjPIfKeeym/O6bc6ElO4oR9hLrlr6KK7iH2INPRLR5bdapgRsTh1SZ6raXyxRnldbrxWzn
Jza9zVnf1v+Xk/8wsybGFxnV0dVtcbNlw4qFWztetLj8LT5mkNBI9vx5klF1OkkUa3f6IZnkFxup
i0NxL8LN3Iwwm0j/pYEe8hSdiYndG+MAPhValQHqKLQ4zT4b2pZp1SNCo1lpxQIpsuuZo+4F9sTf
j/YYNSVhiCeG3JLBwbIX1c/qBeoZErq+YMAY4cRvJmU0gh9gTuWb6JsrF1ffW2+e98pXt4fqE54R
LEMpJEYqStFTurgFs1B9+n0W/s1Y6HnqSDn0/BbVVUCS0UZBe38keuL+2FiK1f3/NHWHSzjXFATi
jayA3RL8IdEnAo+QJW9uh0ZDdydvnc+T+bCMlNdiG3ujdA/UUG4ywll0R1sLJiFNnHb9OHQV9pt7
h+SyMXsVCRh2DMijRVrsOign3SkLqGKZm5/H8v+gv9FY8J+ncZeZkshTEYBksGA+wEWjRtSqyhOO
MPHfk7HrLhgRlWcipcoN4dZeeoV6KmSezQ3EnY+BKjsNK25VVtC04+eeStABP6Z7Dy/peV40edmq
07AwCdPXOPYnbbggKgj9T2fYghA9aUdQZqpPNxqPRC16c61z+F/G4rIPi2lbsTPmHofh9XWnmjte
h6Do09E7efj9yP5uAuykl1I0Rd+WaUgdnNI1QaK+CIfcSehV9omF6MJAkYY7l/thoFKOHZTErZ3R
OWuHTKy7TA0q9cVb05XJtrDfoSxglYR6m2Q8+euostij3gIsFdBXOyJPSbBI1seistZsNcU7PRCG
YWjkP10UgFFMhatIqk4R8FakSTHsqUEPzdWSRz9JpOaLMZdnDKbhrpdIgmPp3TG6RD8a68qCZs9u
K1oEi6tbwfcdf3B/zihMsNZ417S0ry873XrHkARbeOMZi0NW1li+KquLcLSCBcBavXYrA5paSfU6
8Bp1MlSnAv97XefoGv1akvb1rcJA7W46Ru9A43HyP9SOcjij0XK4aH6FsXYHWk1DOVCb1NILSSTS
OJOOmeBSMmglPKMvhxlP0MSlRzBPxtaQQpB8em8d2ThBKQiTzAcEDalRVFT8R6YRaOa2JppaRbO7
lXgO4d7TJJo9uDvxrd+WUb+VhcEEqt9C34WNvbYBeQHiXisGSZra994NNYbRIjvU+vmk7yOIOcO4
GAPrGr2XzYc7DNfHfvHWw21Adouy53FmSr47IiVUFRsO31gygJ5mPQX1PPGyzpa6luWUSs+OLdxt
If0kFGw5EzhQnFonVm2KANHw8bNKjd6M1huiW1wksjaZJr5VQfgCx31c0aqnZgjJ2BsWnjavF9W3
figbzGpyypixmimxpwY0odnflBHOUN7Ik/uuHqlAvDZydia2tviRkVO/D6S4IVvDH2AASF3W98ye
KlymcgQESHkV6kcmyFDmIzQL9ZIEW12Q9QgOWWAbkFsyDpoX/XdPXcD3VZJthDPOJI1d2WT7ZI2Y
jkdqfm/3NqdzJ66jJDUqKlrgshpRHPeDGfDFNX/VSKumRqaPTnaMJAIAo1Lno1HLWafhLrtCrHhU
qNUyh00qYICMkYUJkPB2Pewckq+ri3nds/Z/MbVcHs6S9Fxcl0guIlO/9sRZfGgG/4oUh9AY4+aX
A4X04w3IqAH5E75vR7+ze6MhOFWCLOlqE5J/Ngoerlh53LVwkoD88GBAWkXU8S5hR8ongo/Gwmvk
zBmMDZ04Ju1gzZQGVgqrh6UjEBaNXwkO8XPir74odHtpKY6gn3CpYtRzTzs8JF5kh+dPe3zAciiM
/ORa6/swpONZ9FNYoGAhyBPFoEV2ACDNtdFMKxo0ucZqYQ6CExR1Ho8vlwQaVjksfjqWD7EewpUr
7jSgHjeHnOk1Hrd6uAuW3at1i0pLa1XTVQ83GBuqOfPVkbVSOZnfQs0NQFQMu49P84vc0cA4vSgx
7VtVM9uYJgPdNnh8tee+lZ7JyjK1/kkadViPHo+iOxwF1ZwNFDp0d6xQuHojzRZKfpirC4j25wWC
dchDMuRcP3xEePzHtgp0JGPIMehXZuThJGNn89PeBX58DoRe77SP8zdoKGgN+G5GQPZKqZyYOxtE
4NbvJcA7bKueKIcAh8DAEAfR23Bj0m5X8iLOCzhqq/yp4WPPfKwYhUkEd3+U+znHewqExbYAhqxo
1AYYzc7Uof4okOOVaNKHbjpagCIFtka+nlvroDc/Yt5MQz0rgQT85bqdkbTS6eyZ8vWJtJQ6i4r0
AWoT3BSx8MSzB8XkS82edppXthc7TI0hWBvDStQJeUYxvmb5woAefi+8JnUqMFKBLwHeimtE+xaD
3R65Uk5CSOzzlcyXw0QtlsFMpvSyq82c2m/w3zhvP4Ygfnek0wrWLRhpoDRwQWmMVlVR0DaHgKYz
NiMoLwgC3SCmVxDE95s3/VcFohATTjxgzOpTV7u64sknZWGPT4mRR8ffvbI2UWuelWgHgFDZEJIZ
jZztJc8p/ADnA7hU8mpeMb20fUDnNorG2X5kay5ifRLBJbYmsCTkaNtT7d9i4TMyu9NWgrLMILkx
Ww3OKqKWeVi7b8i0KX8UvHppZD2ya6VHOinPTUpSPlMilRzdcgbei3XFdCry+bjidbyScbZGfJ1e
Gr/6B1BbkfHUjZvGt0qfbZh8qCQF2rX3wQ8l6/ZUW6xDAM3QvY9mhhSR/fSw8dkkbx/4YwJLFmir
PBIlTn3vcTH5KmwtHTqlvy3Cirm+PGw4kPgFB4xDsWTVfblX17e2LBe0hyTZxrhdwRzGteglww72
aJnD7TFaGDxLp71RQT+ru1WYVjBiPfLs6nxrJ64IbvVl4b0SPEaxu64QLouUiwt1v8HQLETMjRpG
7RneHMKkuWNy1rCyK6HS3XvyQ5/cts0CT1gZ/YdSuq7MoYsKO1PmKJ4I2b0XniHeBWM/XczqYO0C
xPWXJLWAiMs7dpOPbJEdcNWSG/P9fozZKycPqPl40M3KAPgARNv76eL3YqPWe74wUwf2Yt/g1K++
E/i3tjYj0FvewneEj+9JbcJDqrhD8tB7Krw9qA0H3OJcINb1pGFWc2xqCV6pRjYI3T13bPsWcQRp
t9cisjfpsJ3yoOhKYhb9t7jXl3UEyG4LqRlpMxfsC3n+eC4/kk3zTdHT2aDSLsDjXY9lLvZ9kttV
KbFiU4tId13V8PLBUV9xG/ce/tm/vOLMPdLJWZNeluxDev4bF0JPYOUNbSbdT+pOZj8bWy/kvtY4
0/HP6n5kcwOxGYXH9tmWtECynoSiGyhbWQzMdQZb0OUBF7Y3gxFWzJYS5TC8M1dNY+HEb56UdTqu
1eNqJrlLV4onhH2sAfsU1r6tMmz18/16PuRInQJgGI7lgwxMPxizF0rdEdhbzDA6u+iu/KpHeAem
N0y3HbvnBbaMTUvSecnKA9Dqq7rDXMYmSKGSt33HsI1PuBE2ehNfPnj23ggGkex/wmShbTkAEdnG
vcx7j6TxgTscYV5S6hfRGIJlriG+MNnVC0ym33QTPYsKaXOfrMEuM1NE5VfVjTaa9ptGslBhBoaS
jymEDWb/2V9ZmHhKVBQitrd8c9ntMrwPsT39gdvL/WMTPxxuY+F6WTIxKaI8mre2S4XW4ps69ATL
suKMHL/AqW9ZaXsb2O/spbeDK3OdFGodgMoEUvAIEdCbaNEiItOnw3nLU+04lQXK9f8wIo1ybZ4E
exwVgTwIei1diuPjnNl2p4g4adyNCO9nb02LsFMekEVGwK7E/yi6hQNuz58VXXiStdIbM9nPRcrn
Y4A9HGw+v9FisexWO5ULEWQCbWgId7gQkvvi41zFsbgM6xKBUoCJmAQaGwSBYtZhRflfuMP3yyqT
ZtNMcABAiYZfBRPtqR6H5ujmkXjz9iS5twslU2cOTNTw8jk2PMpX5Ddp+bP6e/JRLIRqPsP1pNEy
1GfEUBzmkYOdfU6mhmSa15togqd+mFqix+2M/+uw1AC8DJYpzlys8lDhENee6x06VFPJr+j6z8AL
wW+JIVqOEC0mylT5AABHnJq622WL6uqw/iR0DP5L/q9t+hhvO1kXsbog3PO3RqHkAanh0ihfZzZd
Zxnd8ilNUouDyZocv001OYxu6N8TV85Qpui9Yf31xOrg6PXdj1V36x6ArrutpO18uOtf8J/XuXP9
+xadlUTvIY3NiuChzmdkKEHityS2FbfBD2dafeWC1XR2cW752YIccmZvS2GZ1FK9cXo2gQ26xlvc
1hTwjeaoxOY/w4Lz0+SffS5uwGf+NWbl59/B2jWju+IHcwn+fpgVuEOOEgxEVdQ/RDJKIk/Bbzgj
rCyI2lYmBiPhjVXxYPiia1ubJXqVz4p2b+aecYx1mhJxakBMNXlgPcmgrfdnOAp2uiOugTUr6ozU
QRUY06ZJ37x+E+dAO6rkumn4bTB42IWILeefwym+ZC3SR4sT0naBoYRuLPBCwsly0mJzDjuK2Mow
AJ3P6n2f7a/KxqEsU0+ysiGNPiEuwnrbtlObVAZlmAce3eqjp9JNHa1d8YTNUZv/w2j0VuBjlP/g
j6d3zsrRvAYiCtYAoZEjAshIpjZP0LSgOU7BR6bJjRGSjrNqWuxb9maVZW2M07cOs3LWQpDyb8TC
lz6NISphvsWVq4xTZsDCXA5zrY31ZWcxzz4FEj1oAz7XVplQGtSpZjJ0Hc+ooMWGSsYnYSRkrZ9m
u4tq+eGtBmBgbG0tOLct0sBK4KYJIvtd5nMh46f0PPwW6x8E+6CK5j09KtwBW9nKCl2MTlmT9CD6
arSkOPNGEsMEKWhKqc0A0h6uHeOXo5Tp23mnffyeW3J7aZoU7EfgXuT690FoqzV/32RvU4WFxoaT
KdjPpobiugD94U9CL2u8xltHd8/9/QcPea6ioD/wfxZvj0H5PBkY+4kGmz1EWq0LbudVPZIgaJvV
5JlLXPbI0OxBLvKdFonx9bUp0w2QDI/MZIDqDNHj63Yghn+/LDgbYSET6S5+U4p2n3MrBnu91gOH
srvvE5EOSCSZPx+gZLjbfyL38LWR0rivtsfUh6BIG84TgAOAOYU2X4uk3qI4pZFs4uN4XSu86yQd
cO9qT3zWnVIow0+ZD20G4qPaCrMGXjJ4/JRIR6awKhnlZJBag6Y6E4jfhJtXYHH9BRKx6I5q1C9n
jBHqS27MAxDAcma2JaHIJd5tWAPDUQlroxBNCiMF4T+ktdSJuOSjj/DLsrraVaHtO0FIClU2kwi5
rnZTlVzCXQvO5v8SbPsimXlw0F8kylNxv/WDYCGSP9N9lbELT9pVj8atQFRHoclKFdHUmL2E+Kat
lk+gSONO3QmQTbOH0zyI2mt+0TqkU7eCpd+aLJG3T/Pj6fNvU5Ns+/2FrQGVqsfd5aMPedocQzYI
OvJ0uB9lLN/qWQnbApIN01IMNSuiQsNiDjbSrhoLVE9tGBZ/U3QS8Bt60BHv+q4pvpJTObKU1H5T
58XFGk4GJW8Jk/Ks3t0QpqbplPQHQRYS6iv5ou5sUmphgRdWLFVftzXrc2YDfdt1UnCzACgKByA9
ZLhVgF8QgoWmv8FALNuks/zWA1Lrv9ZP7szcdmbPGJ2g4ahkZTIIpFsfeoJZ0nR6YezaHE5HPw2C
1lv3Wh8yvKwe/LzVyHqOgiuDkOQPG40StxoCm3E9owf6c96T1V0m/BG5t7j+RcAlYrk5Zj90BUNU
8My9KsLAICbCfRPrnqdydQkIIl27GPO0evH873KlRokviSByuHQTHa1QmKGCKOV68FFdvLrt27CT
VSbzw38f0F5z6KIfymxwQNJE7PvfN70rOSqTo7iWHit8vdaOxXr8SwAfeXJbqrVm5gii1gJgZvRv
DEpp4sKTbZlTeI1FKl9YXjt4xe3IuKif49zR0LsvLpMtm7MJmTgdtUIizSRAH5tZLFzs2QwgmTHO
R/ua0OqYHIJlouFS9QZcwcsGTK+yhMI5z4IXdDRMw6kl/MZTDjA/NIIDqw/PM1WfeFKKOaR/h2ci
VFrNWDpGfzE/z0PjyW/hbCbGf99D/Nc6+JcBVZDKv9GxXXfOqmvF2xPKuIZ3Thz0kqWIkDwbYg7D
7c0bOxGm1SzTZgnSTHh64v1rX53cWRFlE9Z2kHA2HlshRBwxuToVgMi2VcFR+QKWae2f5ZyDraZW
VOn27IBfGEWOUvgyaxHf5tCCGQ9NowUU5hu7eFwvaziFrZDuK3/hepV0gvmoRzebXmgxWh8CpEPR
Zo51YK1guh5hUW6ZUWBURyN+zjVcebsULj80LEZqAdizyj0pC7GcpvrNZGGw06KzJLX0pozVtM/y
0KX6bfs5ccS7saqRNQAAVutyKL708YSDgQlPW8pj/03gK4srIRJ8TB0+pbdEawFQh4Uc5A6HdrjI
y0omeAtp8UCNbeK+Q8CCNVJd5nhsK2tL/PF0Abk7ZAsNLBNYN7qyRsDLu1qhadMe2c+KzTRghILd
X90b+0cBfFlsGQpMLIcm4zKnPw0rQ94rQE1pO8UIYtUI8n7bYYM+E3QR6q9reCJ2/JNQiBFKuhXu
Qnon6TA+xKS4tlMkGfxu5BTY1fxG1YnK7eAShD/K6vg9pTaeXSLtFZBuWCbiVNHjU2Sf7cc991IW
Owfser+tNUV1phABsP9vtcy88c5elzxRka4buDkHoNhtBKlDQ84b8xv2Mg+3XmwujVRtbnaAqxba
u21A4EcYlPvEFA6TCyDGq9nGnsRDyZyUKUWAUx8fDiQSrvoK+G3ZsW0+Yhap0bLyOUtAbL7WIAsn
anOf2qZvLVYzzFWBe60S750Lv3C8d6tGmDYO3rRQJlKqfpr5zJgBA7f8L8A+5IDOq1f9yL3tq+OP
/zUZ10TdHI99Y6hSeOlvB/8FRAL/5tYWvMscY8lbXcadtDVU7pNhB07LC2jH5BWxdTMAUUv52j3h
zfX8Q+df14H/pbo73daZojbZdFqW+vVYqo5MzDvz1MSoSadd9DDVU5Ag1t5AnWEL2fFQ1BNSHUil
CTeZwucuG2wMhhNdxtcaibBFT+yTytmAkQn+tKBVcFu9R41w2Jhhl1pQFXngrLKYX6YrHFB9Zo4d
yFVy4Oxb+cxFYtOFXzVRJGx3/TdZ1c/lSgrEvJq/t0NnzVBHjQsWpgvBWoIKAJJPM1axdslXixjG
Wc7jLiAGJXyh3YdGBq9IV0NzwURwwYAoNtmhlJ+ksnjumIag87itXkscLF+O9O6+VefsgaskSKPx
JeZl7mv6erNyPj18wENqoaUL2BBvu9o2VmP9BKPvTOGn97+SNdLz4c3xjc5Z63Q6S/JtLfDILhQh
ICFDexTs9h7lG1CI5ZV4Vag/aa+DiuGlgYpha7HcDoV02vYx00ksrr1mz31jR7AAxDh7JPjSgvq+
TJ61789XdcM2MIICJwiQL570NW5OOgGHnpRuIYpdN4q650k9/2ltHhfOLjmjIGO4JsS4q0Y4z4yC
m6Zor2e6TTi2Qi93KVIWq3BqBsGEcISywejbE01EDhtGVT4ThdqEtq7DJ0Ju54/++EBwPEqpvIrV
5hbn+gT47SHacvSYTShBuLH8S0ZeaLw+2vgNYRMd1iVPzqKbth3qNwiL6DLXYBRG+vo4DkFRETAd
uefv86D5roZGZZ+e1mYIbesHe4Dql1OnwBJoXlFjK88FKXVs0J4Hjt6r9y+OE38pLZkb/DGrSahw
sHcHpEQVlVgJmIBdc6o3PVjHxQMgyNExA5p/Nidl129K5KnR2CnJLq4PeKGF5xjfGcT0c7369p+l
D3veKcH5tPNcvA7go8xs0XPlurlCc/onuhj32NVYC7+ia70MhmT6Hc0mjzVENjUQZVU+bHgHfYkm
pmrZmmFHhtc9l/HV0KbpfiSsZKi8W2CM6BznxR3A6Vkx9BU0FosjBjNH0f7i70v8+svL1rQ0iz4H
igZV9GWSSZx0Ij5L0Zt0LIBLuJfp1x1xouNx1hi4tp4qm6GKdRkNIXnQ1vw9Tke9KB4ZekzMjbKa
MB/dB/GcfFH3oDnjUcqPLItTQ/8Mfpe3RNd/XzCycidFt4SMgPjRrV2ui/1STGIm6MrBWizc8I/l
907b4L1TYyvCwlVQaTcP/zdegzLz2gEv8qqgXXLwnRSYOBxbxp/QEUlCY0WAOaJVCLBKPWSSmdp9
917zq8XBEHBNYqLLtQAFZNyIXlTExzoAr/zCvHr99ftMTOe5nwmDj9n6Uc7ul5yexq8R6qk3XCHG
nzWX1GeL0NQuYWJh+tLT2FxdT1nM292+zAm5pBCycJPcLGD0XgurrBS7b124Q/sChsNYq2kZiNVX
EsDlYWPytZJi0ZJzieIoICdi7k/iAraLEucfuzSI3GMWSESnDuHapHAV/immyJ5SWLW478JrW1aW
+fPRDf4lvC44++2xwRcEc9CbtIR7H9ZwItvRFdTvuhb2YlI+5Edu6UUNh7BQBVd4xC3aoXpHDAzx
fD443PLqAdUgYH39Z6TQEtXIKOUHj9j0fXDAX9U8Z66KstdKzQFIMelkZ4bX9Sw3ER4sBasTuTMw
YzZh6z5LTFcyatjqntPkVq1DkN4oRczLlsjZfOxVH7af9WhYoWSh283ufVE1NBSxoi8v5RfPpYly
hdmiqGeg9jpSSYXf2XXAXlETF3bmpfZbKjywvdu9lWjv+JZSl/DOj1jvry8VQCNoHZs4xMXBmByd
FXkCyLl7/vt6CXpb14WNVjpnUn6cbMguaw/qwbnt03ezHcJibeMf5pDOdsnEIFLhtKyDsI58H5un
MFec5GwdNJeS5UGUUQ2NHDaaZNPFS2I/vDt1/gn96RwKIZXNxyxWuNYLb7CZ6uwzPpHMD7sHNll3
V2NWBAj+P50BwTHaknGcn/yv3IR4OXm5nSuk+hpMxAoIFs7REj5oRxMJ3MEEh7oaWHdxxrDBEckH
Di5q3P0f1Ug0smhV2y0eF4Rkv/PvfCpxxhRbYOSEwco4GrGdLoYbxcuvwIWOi4IJDB6uvz/TfUak
XPwbPY+lcdIxcx/BEmyToe1/4oXGBWVYKhumqgVlgXQsqWMaOyn53RIcxDWd1OFlFnumlj3YG8BY
20IVb3LfEnDQTCg9hnYDDMWRTOiOibRfkqrsA48vhuZpO6mmNbfa31WShchx8iJNKHAYnq5aPnxj
7na5qVwY3xnnvOtIyWm8sUZqvbkhCCk2GM99B7jnjDWG3WOses30rBfIBC+7g9A7mwCMeaqeuGjp
aF/BOynO19gc6GRFHU/1KGnP7xVnuEdhQEZdUTNDnjPu6YcH2Pp1yVWlak0q1p2Vur/N4W49wUBP
vR+Gel02jqcs5eC6wM/3vohmVLsMqNFIpG8kq8yMEPi9Gw+c6YFv5O5nAG5l+xLvw47fmHhsrMja
XuqEHOaX6/VHWe2mctawuezxLqZdNwoxpj0wq1igsGTQVw0iCPn/PBng6TKY/jMVKW+WJdNnF4cK
dN/T4IhHVyu3kTNfHWyv+jiDqZDanixYDdt0v9bsWHr5jarb4Hmq2FQHEpx0t4A+XuZ+rQwoCdIN
qdhRzAxuZ655Obrl8KRd4oKhnzRb+x4Gz/ca8PVHV24o0T+YYSzDP/Kgk1EcHGk3w7CflNfj4h5h
p0iKbG34BQiQR8x6HF0XZPfYBr86e5vrImaE2Twqrhos3hDRI1iX4i3UZ/3IpP9aaqkGr85hdjH3
ix97avrgumDQgIy9SHrzwDVjmPgvFyx2JtsiBmoMWrmk9fuvmSGaw0Y/5RmzbGc8dWP6aN1+dOim
vMhIdOzwUBr36n41ZR30+2o3oKE/UL7w93zPP9+tuRV5Xg0v5bSPfb+su2dUk0/+dNc6fqY3DHpz
ZNN1yjj5i1x/ep6jvyaMFdhLh+7AVti6YrojWHaouZiHl+ofdDRcRVBvQ+MRbFTBEHZmBTvqIikh
XTL1xedzVCGzZgK9YFSOZV/vtGKVeQj2pgi/6kntosxovPTcxkNK76b25Y5AEYvAlepa85tDyGio
KVPrgeyO+3qQtnOb41OAP03QqTC2pdUzkG3KI6uNL3Cy4OlenLFUWVnp1CEEaJcMr4VIhfQGYWt8
2S5M3w2n15Q3p0jvnS4JTsRaJiydxtpxlTKYfBukWo+8etJ5SmpPj1MI9SHSIZ+TBK6jXEVr/fjd
pB58gDHbQcoZoKFHFgv5o49kG4BAv47GRi916c+uLpcNoId8c1SL9NC1/sRn1ixNbIebcrZ1VUrM
KSP4wPbNvvHGGspeU2Ai2IqwGBzN+FeElR7jlqBCBMlvhyQYZTa2u8eQzgPBWF3lXrHQYc7AOXPm
ae2UdRSpGADH5EOhX2v2PMYS6SVsl/gPp6H0t5sTDvv6E5C8InZHIht6AsDISi2YEVLK5DAuhuAF
voyVgYFDbEFmRfjfz/MmE26HzpnJq0FT7tXdgi1kNwoBTZwkOmBwtVxm1joVs0iFiv0WSXg1WLbH
5049YnJBydZoBC4VskRWM6YQQ4C7aupb1dVLb2rEAgppeIMRR2V6EPgG3RUVeQEnaHHDComTIJJs
hRmsUEGXXS6ZOdSiOO9p8gNZZ7CWigPVe9mQN2KKtfammhyqjvH6TfJAQ2CZP75WGpZtGdqitgVz
7/6a/oA300FDB9KgeH56w+/v+TTbgNMfQ59EGrY8eJw8+/ewlI1k1dVRNITZ5JopfYx0Fqngf/wt
1Xn8lKmUSNsIH2HgDlH/LQuyuka/7/dAWSBreWxwkgfQ57dW1ABcl6R8/uwPAOnTIEPkHUvMw2/4
vnttvp/g3lMo1E/4ma8owHp+NWPUtXYVqPXdCCuZYdJ9YvkjB+/P05QuBj9Rby3AiybYGdd7kAGY
x4RmqQgmPkjyru6p084fDymTlPnZsQH8Zm7tdw4cLOx7jznv/v2Er/GIpnA/xfH1WIL9BckyN1Pm
k9AFAmc4L/Tjcrm5pKq9JXwPZBmWxpqcBHKZ5KNeQDjIAky5ujxDSfHyrmq45I79qepRM8WaRz6a
UEb83HHX9Nx4MYLRBAZWR/8yPG4cZY0kPHGhtGfM2h76cxtNbGJ3aRVHpgezC5B9EcEoudkx9z9f
7kWpC6L3LG52h5iB0x8cJvOzOEhQhBOLJPL891foOzOPwEJP2w3MDNmtU45ua8xt1w2ZGi3SdSp8
7BxqATyIJcQ7BZKsaoPEqzghjbUxVvEUoe/FwyewC3oH0be0jdyCcZIVER2USVZ3GLBPV0f0zh97
mssq0btxhbFvsX/BEc6pyBuhyImD9voR8dWk/TxM2LzOtelNqE4qoOtR8gFEaUipc89gQntmD67s
VGXp84rLqI/8UIDaZZmvIgNzElj3g9Rm7UeTW4qgPaXv1xqqkbEax0osrSpp3K4pwDfvY1reRsxh
mI6OXDy3g6+oCbjwK0x1jXZfebBGFAz6+lzFIaBvVcdKPWzy72kOUTjNXGs+EX2rP0Iti5yz7Ngx
jxH+lf1JYaHUKfU1KwuDz03jH7cQ+22LWh3sfY+q4FmFVaBIqZ40TDY4OMDxHT3QyDOi3pTqpEMj
Q6E30Sv+OKNQON4EzsV3VdozUJUtiXQgGSZXA/ZL/0rmaIUPNS0gmJwW/sDJzAJp9HO5TYxlO4mH
yDGnra0i8dzX+f9XkFkNKp+F+6VQD6uH9+UkQD9VoAUzp8DYrbiAfrHYvP1M0Ty8Qlfw8J+TZvcE
K27AgHFszrKNwwogMuhClX9BFxX7+RG/3lIDTDk0QahB1dP2ZDPYVe7zs9ViRS0SBENLjTDx+uxc
jBipmgrOj+Q7MrSLircS0MR19XbtqobuHDqjAAdLoSgv0hXymq6M1ySC0rOL1DFlbpBQUpUNDzEn
4obM7g11sT/wrDackGYRPGUkRb7Elb3qbgxRLDsEJAuliadf7P4wZIkV+8op3NSF4VBQVsQgAd43
dmimRl28rKcdcau8ZHqoA2E3icc6bWhkZasOuX3lO6lxtg9QnSiVakOE1WaXydessBCUiL98NmT5
QKxVt8vc0g+BdLTcerOn3IsaKWe5whSVp5IqanbKSRdz74hOZPEkW0B9N3jjVNvafbGIPnD6D6os
wuTVuLcjD62x4kEeGog544oTllyJB3G1p0sFHo6izJXwbsM9HSpBq2zKxfsPxTi6fk7I/b31RI0c
jVSRzB47UD0xGa7f/j5PoICgiVdqOzxJN1JM+PXCoVUF4JAZSs7tPOjawmiEJ8VIsVkEfi/122x4
pOYk6LBOI3tUT+cMSfZWGomMvGQuv5Kez9NWG075NSDF4o97D1O0iOxs/IR4I22qD/WJEYBGeUFZ
YzHidijMNDIO8qs7lGsHp3cJYNHI5ZsXnJcSJySKLDiqrqC8h/BGNguIHUd9GDN6ImLiLEPamNEt
3vUlMSNn0UQBiEE5DCRmA3NmZ6YIwnMEdV+g5J901rBlu1OSSkPnmHhI+bikCKPYVIOZoybv0M14
LjTcAwHj9NPFK5SOb49Ig6Wn9rYbi8BXjI4OicIexdu5NUvrkIZOvLqjmBWEVsnigbrVy4+LarfY
2pLuH5Td177UIc8cQp7OaKcH8FQIKTjn54jxo5ptVe7o8pF2RagjLH8FlczHt3LOrhH/ph/Y2pCd
q8JMZusgX+bYbPpnBCsOGNvpm7+uqiRG1nJw5yErwPax35HOVRgYnyvvdFBVmVgxtDIKpXiKeDGd
ybcfxLfHtWiqwbMSBriE341DFWU6m8xFVVqGbPHw07Bxlc16Y0TgeA406cJUxtF40H3KhecJ83vG
wpj0Cs3UpGuz/oFqqep9R+sLe83z1LCS0NqiLocOvsYJdw3fDBMLbbG/KI7dWLJQHCMZZWX/drFK
WRF7Ls8zPqcAD/kr+2iRiG463Wlm9idaerKQvg1DpWsRJbMonZ9y2KW3CO0Do9p2NXx/SONKJfMr
/GbotioK65xbEtoMOJAtrqo7s1M04t/QYtE3PS6Ya8qaEbz5v9m4dVlkedf/9khLyK+T0VDvVoIF
8Jew3Alo6Trc/idkKYN72D5ulmC56mQls6p2tq26or0rr3DdZS1IZ6KbjLTMsHBX5yOCsEAIogFC
fGl0nOcoGy+98ESNoP1Q4RxAq3XhAt/tBG06iQTN7AMRn7CdE7jsy25vtl2PL+jVRd0zJkOR17lK
9k8j/K2FEx8O/Q6SQlGBqLjFmjM8NFwpNrZgU4s8YtVtTpBfvpt9XfsmihqIwxQ3Oebdk9seMk8v
vfZoPrfOdihCBsE5fdcNGv1ewsQ2Qb0djpLNY1nKjdQEg92LVYIQz0Jjhrrln9bO0UcieekNTQoo
wqDWfiRAwzHXomKnZu4yjxkf6spp934RayOJCk0b1Rkx/JDfNGD4EDSMb3ggXJxEv4JEVbQRgoLp
n4YNPFEPrTBjIaBYE2GOVTffJd+BjxgANfgphkP89R+nuriDMOhcLg6nTx995/lCn+CnmGUJqTRi
VWnoHVxa2ruLnDZ8R7jA+VqYVujhCaQk0X3H2CTSR0fPygSVozJ1nN1OJVcekNORj4la+sySRr7a
8F77IDI8G844u3xoWZzbqlb6+rew8gsHGn13GmdwYMfCn6nwC0X/BAFdlIcYAdppx5lnbqyEwiwt
vjzPF3vNAUn2fA39pywjJp4aOMFrTYAt1t7ioKxNBH/Z/a9jGYvX5qsFS1gRsk/yX7zQpHjoJtJQ
Wj3v7Fbl8PncN6seWxYuuz6N03qi9W1YpusaK2dtWyrm9vZrYrh/p9tR28KTS3qTT/9/JVRY2B3q
vBPfB12kpmtBGCEa7E99y+ecL7cCbQpx5y+UKSJgPU8zZxPyynOcsSu51V+1lH3CSdSxuKEWI7uW
JwXb5UH7g1Ra7Me79bP9J0N+/ydZIjNcNARiCBG0TMHVWj8KjUEuMFGPYawwFR+xRwi4xaXW6WAg
UNP3F6sPEE+8uhh1SgwyO/MAQsRBj/L8Ps5OckEW44wxh/PzqBmIBmdqrLTkUVjbVChjwbaX0nqz
7qTAkrRlSsSCGeB9GTbyLmUQlGZ7WEaaBujQ4R+xwi4Q3xfvf46JxxuDRCz8vzt2JztAjYRZmFPo
A+kKmEHk6gyjiqm6f3JUGN+d/fu9SBsJvA2kVoRLsXTgP7HyQWR3/5wkZQGLa1t1RzeASjKNcX60
E4HRRFIEVD0du2IN96ZCF8+CY3Wl0uKkCMhWha0oFDh3JouzQ6I4i1sBROv9khqPxjfoTWuZfVKs
HTLzDlQvc3NfUWOhZISjY6+84X6numTP1C5Ei6MjZO0bq2OyEm8GNP2EoQHGgFuAHvKfUq7v9yfD
OfQcCTbnUc3IncodjUt3Dcx3L1SEbX2WdjJxuAXlEztbfAoLeLjT5EjLqw/MhUBy3CpIVGnskbnU
dYkEYlkmJd/MXGqUZBvfJQiOoNvgp12FgaWlFYndDrDAEpNpv0TvydeQlPYv/T2b4pF3y/kW1bGB
faxO6pvEqL322AZrDieG5mxe0EtQqeLCZwprMr3qboaBt3k7e2/tvQDezj2WWJnwIqy9XFPfH25H
Tg37phLwz0iTpPByNdHD9dkCUh1ZY/bK8pnnMvsCoPqYJzgZSjBXw7u6GGNZBVeAbMM3/chgGAUD
i4tYgQh5yxT+DyVg3nTIqZjrcXInEVZU4RBZhNIp8k3NNKtmKvweVvnhUwTG2ifxEtxp3u9Ar1Lt
P11zCLMf/8SVWSth1B6pg7QY4P4u487Z7Q4fXH6RyIjudkCloXso2k4/ZRgOvfiIFqJte4qJkfKI
BDTsOp+Q3DCqxerhtHSbiyUwSKRqKjN8iuQNEghfFyUYjD1ztmIfSJYMCtX+nBMIie0n+zwJ82Gd
1pCOT9a9y+q0ymqBnHh6+ZTFUK3mU+d2tWO678tDL2V0Zh9UebOaAEz+hBWMQLQsoARoyz54CsRp
jl7uymmBDB16bnnTGD8Njn+uTK4m5x0dmHF3e7V+JQEDLJj6hvw9N3yjogqy2ejYWpL2Salf3VCg
+k8NebT/YXcwYNvq/kkwtEWoV82S0EOleauYsjaYIoOIiPX4npcRM3h8Tek7glVwjFNURjhZgDZ1
L6DBypTLNub3u1//ft+7BtsasXZCOBveNegz5W9t8kIURinXqagdKYWwr6gQRWllCmULeIkrh6zH
qP8GijOoPphVUY7oyqn9T2OTr5+kGmAYambKPnQoG1FWTTZg4EVXNWL9uBkSJEt4m4kUU4bhq51o
4qaA2giPQSNTLsezY1MVAaHJGDoW11S4TSL13ROnLEKDP2FymooSox+2Vk1oecoLHtXD7+x5j09F
AnUeJPfYgIIoAqZiUXYjiWJbnQBs4g+62gAuN4FN/gWxo8Krmxgh8rxfervMX6a70t6xYWI8999m
9orXtvUgyA/QX4PmezKca/oNTxVulSe7Eg7/wrCkrQcIo1/4+1qyK4wcKVRIKZu15erfhRZwLi/2
osl3noxHFVMpeZasMcPcV0Ojv34I/ETl881OGjrGAu6YLBF7z8QIljy2Qdx90q1vDW7UIA6+FDmf
TXlpJCBMLuHIXxR07PTKNtOlKcCuMS0wYbZuw9lbjwRgDFcRCR5wBiDsAM26ThitLSev5TRO2TxD
ypJ1WjnzKM4mTDQkW0srBJw9OZBh7UxnSyZ08x5TbAgF/RnrcNYMmW/0qlhcVBi7QEC/fUW6Jmth
LOhMrKi1lOahwpJvMwGS0AwOwmf5RUE1h1GKTsXqx8aNfqgMCz2y4LjHLznLbvVye0LgC6QRKBM1
CTf4E+/ETJvWlV59Oc98DXM+39xvPwCKrVpGzkJ4LXBdOQlO9xdpxUTZeuBkLnz+gPacYtwqVdDB
jv3PwjsRPAMt0kzTHlEOjWbH9q4PqboYtjHg4VlwGBzdrifCE1jrDs3icb0a/4zwlH5Z8ozCJOGo
R/gMLTbJOcapPpJtTDq2AGhLQlqaq2Tlq7bJmvARzJgAgV7R+zPWDknx38kZMNVIotZEW2LIE0sb
vyZHMH6GOebN0cM0oaKFtz5lZk9iigWNXtEEC6glV130Saj+ndwg7jsTIiP5ziK2GkE7w64KbpMG
Y7nBYqGlpdVAJhzmgC1ORb+38xIqlY8M89iMjpzmNLUdq7gvqH4OTou9ymkoICnToQFD+c4PcqRk
srk17K8H2/6qTYBSMQrDqcbgCWJOw0Grji+wkLdRChOrLNTs6y9OH1+mFc87hbG4TWg7+rBPIDag
/QTt0PIcpsdnaIVuVGqjMEP5vMwFyyJdEzqGrNyL/29vIuxLs8FEDtyyso9hllHexXGOIJCM4T0B
VDTVPy7BI4dWW21YtVQw+EnlV+wuujHpbAAleSjq1uOnFe8XJcwUN/J3LbN2PZcQi1cnkwPwhHBC
/1Kd9dZgsIzybq/HlfsgpEFCBfGDCPvAogHNQTnKFPY+QWaLu0+f2rIDWj0agu7gy7LsF2HspyS/
jI+/G/rcvBdKW6a//uFYv5Uss0RUhPi/UCuI+DZtRTl5hzD7r+hWY+Jnn0NJWF/IyUpeJxUbXJHp
sZAyWccVX9N7/DKOdvVwJi3Xx6my6DPhg2DgCXl5mY3gtPXc+qSjyDtUXlF/CMhZHaBYVE7xLVvx
Q34J/zRDF5XrUoOcOL1H0wOxS2G507+yEIqRPyuIPh0k22+BxiZab9A+8TCiIZh4USJlMN2eT24d
Ba50mngmwSSCox1BwFaCncMwqSWzF2E0Mfnh7161s/XKvAVar7kxF+grUiStZ8M7hw0roKeRJa4/
0XRJaNKP197dNPrp3ooUiW4/LFOU481+RedAQtLtMx5EGJG7jHLxsx1ZGMpnWp6lakFXVSoKyZpm
YgtbMRSMaf8+BOkwMGGpwK+lvtXg0BbNo+q5h9cRIAW2p6mbjIdxVPVQiMPPQ5p+8gZ9TJcL0IzD
GfEUtz7B5KC34fIkZKYsk1r5WxMY8AortH1UIOAO5iECSJs/ToEjJ3o+qYAAfVSfvdEyM5mGlvH7
wP2oXGUi7bsz2hoWdOg41Z5rSXzyY0zBIf9gqPYws/NMDggA47uP/ZVHTVBSYyDbD6aoPnvsEPEA
naJjDOf3wZt1yOPOUXqQ4ARSusd4e9bm7lymbZIZJwoiT0IFeSYiMx3QAhAok9QLeW6d9I0N8Mxt
47OkdNFXjkc+2u3v86bHFk/UslMkW/8jBYEQhs7VwKMZuUy7DJHZcbSkI5CrMdlkd+nrgmst1Hq6
U2jwTS2/jjN6yx0V500ebIVYZP7suSQoSEzf5xAOWhVsLycC44QvZc4Gu2Tfs6wag4uXgeriThuS
KSiO/b09Dk6XSd0x5z/ufaYa6AsU8DqoRLt9MshxnfK6gyygUJlZMOEzuMz2vbw7cTJAm/D7xLoa
M7rCcmTKftISTyue8xGYV49mtSKDRohrbkhBukdLknHywKVB+8ke8M2Qs6PsjMIVAzDyNcNMVWNt
qT2EfSKBrr/TvJwvuyplxIhxMWfEEUCbOv8jpAOTG/Yh+Y6gQpZJtFsHs5TFEnTVDikMYg8uJz3Q
y5PWeMBFH3qQez0+kOz+Gwkx3B4gc1GDEQkdDyfEys63DW3JHjqoGA0g2FYqWVMJJlF+sPigL/37
q8mPw4HHyLMpkUTY/zc78D48Gkfh/aeE66fipNuE/1NhFjMtf/O9T9sLVxw9SrJihOrJ17FeUW5a
h0Qb+7ctnju7H6cKpa5Px6t3iWkua8dTBm94c1kzQ+TZBTe1HwV/MS6e4tuDemLXX0EIO6LP8NzF
s2gOfSWZ/ZyQh5WO9wI8xWiT+W5lPbpUwrtdoP5sQcVcShAIqhesKFbo2V4UImxVF+/EBDLZ/f9q
mMxWl+MSsKqW1TASPjbBt+7Kv/QPOa/CJrNAzGGKOD1aRljIkVa/duP72YwzwoK4yshVKM7fOj6D
WZVD1Y+hZOivHi0jxMb2WfVoO28lJqz/UOcXjmRfaa74iq58VxBuq54exY9UA4rO+eXUdkwE59D+
XDi7hDsqwKMRNw/itDltAd/8wEbJz2BehnIk8bqePfPL7ySS0S/u45hZkue7B+Qqh6BRXdKsJFsg
j03sRaFkQJSrIK9js0i76GKxk3fpGFOsa861mp20U6xaohO8fd91ZbRUHmAGG9UpQr1qtQZ7eQyn
u0U8qlE2xGntp45vnhAez57sMXNKH3JCvbsKME8u/95qmAX+3VL3f4PCCe505Ns3jTyqCATt1ODb
Bs+OncJ5/cLUkcmqe6DmB8zGfbx+NDIJCpQdxS9W8+LTHyTRD1nAXjBxjubvVLpDr51+EYAqa/I8
WpwvI+kielarJdAyLZZnBX+18FhUGmyU/mu/a8ny3/uzqDxlwRsu0sJx+cShnQLV8AgCpuRunHhu
81awvE/Hzr2M8y0vzuTB7pkn4Z0wxE7yzZiEJW1tS/iQLd4xlsl8Ts2pZxeCgPscuHetW41X5F4u
XmD8b66M6YSp8bZY6tIDM2N0MFjNOBlTdYUZVaE4XhyvfTxzOFlriDBKB4+PTdeIPZLontqeVm+Q
cfDM527gdGVopoec+Dzsoz1P0WNpawO3IP63YyPdTmIhicdSfqzzTF3TmyyGaFbWwicRe0NZjUm2
ROAcoai+RAyGxcVvYD5wMWM8VfuWlSgtSB9cQ9sWKY7CQp1Tp4N8tRbPzVC27pneK5WvIfbR29lW
QKqEFl1UwWseHbiPht3jqyCE5mw43qznoM6zJ5gw+tz1+Z7qXyIVif+t+OW8qfMd6xUPZbBW301u
PrM0gaNlmJmF6MynUtacgw1KQ+iCJZ2T3W8C1yk56/BojJPJhclWGWo82p7yo9r54IQA9QsubFMF
hGnPG7GEYCFOE0pT3EyFIZk3h9autiTY9SbO41LOcWLph4ZsMAlXZ/bw1miwZlzbSg3SIbd2ox66
nJIK7Kt/jbOx6h0IaN/ef4yOdGosTzpNmP5gox0b3snz+jKSrDtCr5rPTDY4josb3tbpufjwPHYj
GRgAQ8NwRWY2TSrybPrt9EQYQOOB5PEHeE/OEpNIXHAUuP88ilEHdcfEO6CN+jROxIPjV+83I6Gb
06PvUZaRcl+fFtmlgZWlQ/yn2d+6Efgqw//DoHpmO6HnHPlrj7icpAlT9bPyFBSE35pOrqQKmZhw
vjV5VuLq/X7MMoQzGuuG+fKg9uSYyiLyeUHpUYd4fA1m7e+MHulYyxTeP4s77T5rTy1R5B730Awn
7H6Nzvjcmutrhx3Dr71EwRfEZGdF9M8NCuwI6YGAtwoH+3NjCmFAQPcyy9/6CoweAOvvoqh5Mi33
Ah8nstUt3vrDnw8OjwGmycCnrTFYUpIHpXwUhKMabtAooJ9lKJ/KvfP5A8eaLvUNTW4svTz/u1ww
E+Iaaz3/WKZ+SeWa4rq6XG9/xPWvYJd+1djUlQGnQeRTucBgk/FohLEV22yp9YFrYUnWKYuv9bpt
M2R6GKLCRri5eNsSyMy8HVw5FJ/VmfjO8UxH1ottGl0ao/ymt5KywMMcv5+dxdYJBwFIck7DqzfW
cu5yeU7E9wvEHTqd6qDJ+CMhNJPxQaLgsUbAg/35vaIYZYjde2BJaeKeQbWJfswi7FvgVov4JW5Z
utQmkQvMxvj3nG5o2rSjBPJOgs9Z2JdG0wqyMa2Xilg6S41d3ZJ7cC3B/4sBAhABeG/5lG1uf7E5
yjKKMxCw7GnirN1V/gzUQ6+6FoMmIiYBmMsVW7T9FwHrSCzvdoRmZvmJukgJ/SIdCYpE86VQf28I
8gtFC8h/mHUxsJbmDe7NXNBoVjWnMfkT7UFj0YtAupe7EAQdXnSy9iyIvR8DcoUH+viHOdPZXlfZ
LU1hHW1q3oi/iaPZJdxK1MgxNRd7kamvs68mU60wIKDPmm5uWXNXFhs5DU+Sj7r1l5E1Vma9XmTA
DxWkqR+k+qT02ZfpxmF1ydC2+xnVthYgrbUIzTZ577BRu7syXlOzrzYvPFly6nsOVfsDVR5EAYAO
Rof320d3yTl+9xenBpTlKuK/CugemtNsUzef6/2jXsyG02kcWzV2ON4pc+TWGJztEhaYZ6x7cEhL
NlQ/DAukQyS6GYzJ4OM5HtPAqXJQIe9ObJfOXOciqY2R9brkPfIiz4OWvB2QpJB3ftlvvZgYcNT4
Zyv8DIn8ZZNrnvDC5vuJAeU8D5J6D+yxxmYeiC28Syxnx3j1Hfrs+NSTG5arpKqdZ35wYn9fIPXF
Y6AaVMIqFcxXKWfa+5YgTvDFiHILXCHv+I8YsGcb6fz09ZUzOIHzce7wcbS2RMz75FIUJ161ANyq
pVQ/HO6KxKb43W0zHrgSIz3Jkh1e/Hnt2niHWChKZeExjb6aDu3Krxx5qCuhioLG52uFAlMXqOWr
gHNd80HRzyb3unegKrsoezeMao8NRy8aei2Go5FCh/lemQZZoGLpj3lXQorteDMa3gEEltQMVmZO
Hva5QpJpcsyn8UFYOZQ8cxigfXM0YTlj6fdWk3XlgSuGRoXc2XylYt+dyH72W7rGJIwsNiucE+ff
jMS3bc7p6bE2nOz+ZrU6/rn8kslnh8yQGvxfG5Q6WF+WNQ/46zUkW02F6LTTJJ1V6nzChN6sVudz
Tl6KVQacvrASe4nWisjLV+QdUAZi0UFzLdUTjTmHt5lU+gbmH5Cxgjv0+5ZykGMkVSDgZHAZI1J2
VKmp46DaKif+N6F55+Xx2Sjwb7F5dwgENJCxHZkkdqWKG22/SqGXQlwl2L/5ZUAMP6Ob+hHISkTi
+dHzk1ckh9L1IW6SADkFn3wqsjhn85u/aqeBBwICqkxJzooOkzieUAob8FOD8DJCgdY33eGsfKWQ
J7PJv32Bv7qGDKTRWPU21l8OJFmDM9TsW7A2oF2gH8h6ZbydnUOxYgmIuUcuP8armqN4Z229Ldui
3nH3WbCTJj2iUIp4kmc8/Htgmc/aRlJZpdeGae/IBeit4T9o7WcXGqWOXAWS8hHcbetahRTa2Ff9
31tWjAfkOgo0L02uRPqy9xboQz6i7OVRtPSByow1ugtQHMZX7mfHz4Pe/jdy7LbnTB7FKDP4g8Oy
rFxhndw3yY62nIxeACg3QDY7heWA3+qg9Y2lXRKlA1SodXPHt68i3stARMAcsWgOJU213nRMLPwm
dPkIoZcHsuGOKaN7WlfCcKkp9uvj1o3fzrWxJoxhcYYCr1gTU1ql2mCF/FAe5zyHWaRtyUEDnpNG
L0dmsWrhWu027uWMifhlrLD85aa1ZSJPAlm4cuLCT+kpgA7gjElH2/uvNx7Upik4L5hFsExjbtOO
OrweoiYU1Y90sdV7CJhHJcqHP/J3WLUlHONERVUVsCIelWK/lndSUdwix/XBff8hbOSBYWU5kpQn
wQIYNeNMG3tWiXMaZJIc/4BzA0uLtS2plt0wQfhtasri43lfHHFoIczcbNgRlqGy5tHPD72fCjr7
4HzEIpVaXjIFUOdDI+VZ2v//kajJCfjwAbtRWMYsuaAN9b24Wnl424h976q11QWzXKUnMbQlqXY/
RoA67RofGc4ICYgdAaAIysHz/ua1IuKukol0qZzVYidAWxLRfo5Bm6KzGChi/VcKyf9+OYSy4AZu
G0/+cevNpe3+5u5D3aU9Fxebja7l91n7lmSJXlE75aNkWGR/aqUtNCjeLgJM2pzpXEOGenkTzupN
dhfJZ5hRhcOT5bsytA71MYTgF4g5TdtjPrY7lnYXGoYAY0ypwgV4NVyqJeLeJ33kzGTUeEqgj8XB
9FlqJ10S6lOriBSZ8Ooa7PUORT9N6QHk5r3RuWy1Dornp5CA1xurAX5kvF+sFjGWGLAntsK/PQZp
eR6KDVQLkCiIlM7BTcEER2gzoBV3rd2ekSxMv7vHHzX4DkXgige2+9hRXMeQKABIgbIOVIBoWgBv
0IW9jPwkNndlTlNqaA4ikE6OyAwnfPiLgCdx7xsTkStkVEw1WdroCWpj9hPVxb5s+em6G69cgiwg
ihDR2xz2z+3GPfQKBkrL0CvxR746TBxYDSPVzQWn4qpKZhg/SIaqcmceZ2Uf66nVFGTWf2qY1E+x
pPXmqmdTZr5b/CPQb5aoY7B/nscTWHZ3vrM9PaFSys2hwVUadvPS6kokhDmm/vAjK9o0Q3vPpnw3
1c2ODESOiqauqBxCMSGhyMHT7OV8+e+90pXnELkDO8Txjg83Z2vO+tYqRzxcAbL4ASi0UR74iZA0
6xrqJR/2pKj/ldOvDK68nyYdV8UINmPiFxc2wCZcTto7DWscWQb6RoKwFZZJ7Pl8HFoo3kdByM3c
ur6MqfiHKkw+QIfV+JRnNU9vLYN5l/E/n//q+PQELNDJt1uqy4N+gf7141ZYAHQxeFlq3sarRAVI
WV1XLyK9HN/XuouDF7K35OcUF+VmbUdjIL0Yp4DLVEb+Ur6CiSb3P4B/g/wpig+YwgtiTqEpZfyH
Iz4RRYy2oUKyVypG72T+XG3DmHSsW51x+3vhJiJUH3nieOSdNEUbHYpMP5IYuyOYEbkVU8rBU8Rv
+hqzNxxYNkgY5SQDD73WKq9FXxnJov8PJSrtiGsviQrxP1O1s7buRUfqq0ZoPRJwinFHFzQVk9kt
5OHbsPfbOofqMcAKZY9cwlf3K4+fhjfqDbGxKXWKfCOG35ZUcXqApaj0Dh7DEWEjrVi+p+zOTxbN
Qx3e0urSNc2Pue2N7lO8zXB0xgSVuRuWef1+xUkLetpRnJKoL7uq+v9/6I3W3LdbbYF6LggkSGJL
waSUvtI/WADQAAU5MZke0Hyr3iiVR3zqMYDrqWkKDG6MUclAJsHClg5+RhOzfw8dbLGLZbGvV0Cb
xLbv16LMYFENOB7N2ddU1Dp74rOx625fX59OrM9or9Ezw4BR5hi0MxJ90kTMhJsLptn71NV2Gm8z
lAc/mVkNNs4nuDT0D1OpPn8SJEl/vjG+DV8rdoU1SxTvup40BWpN5+Sk520fypTKGkAzo9KrUPrr
2lXoqLFL12yA0S3FyQ4/chIRgW6wQ9ksqzpDeCzbA99M7DYBY1fGFq19+BD4lPIuLENqY4M82ky6
rM7vg63gyCg2qPcdgt6vEC38NwZjMVUsIF0n87I+1GkbschYq2b+xkf6ZbZcaE5ELQ3YayUAvnVb
Ek7ZJwAycgxY1jnSgniTKUATE5V/ezroziIvYp5+PSHUyq8vX+bMZF4GzJjE3cd7dsB4qnpidQ5b
dFmpK3nFF670jJzMvttIa1M+v4Ogv3sDzt87lpH6f2n+2byfWqlGBews+cJ768UnId+7gkVSC9Ou
xqxaH0Rnqg6m/JI8LPdfHfN3/ii2p5D2nZP0GHqRMfzQMg08QSgOIJQEcytrNiYJCxogBHU/WWW4
NfvceHmqm4QYZbZaSefuoOx2aSFB53WC3qrfR0kNRxo7jw/3lxN4g+MqSlye1Ybzj9+1aiVvoUG0
sy7yB9wHuFv2UmuU3UWU3UBUahiO1xaj3L3EA3PSZDEBMaXWdAfQfCsYUvpGbpkLOEjUtX6RA8EX
Cf/Hddmr8aHRB1bF+JeWhV5pKSy6EIarMrQOaa8ft17hRDk7mY9TClvFF70/yPzqYUmkMB9JnpA3
77XMV8sdDaYobu/b9Y6e33gFamgC40WvuKRe2C8akfX3rwMRFnPBtbpCB1VYZo76ME6XAXxBlytn
Ry55S8wdEruiScB1HgXP34uyd+KabtVsaxRhondujWrr3ez0fDJileVayUYZ2Msp86Hzsck5Gh9T
hfsfoit9JBwVGsH5qGsGK7nVvP8g/HBSlNAFYZFB8tnHewfkRSp9Ai+g3QvxlhdVGwp0SnVs7ePY
UjHtzMD8U991dWF+F4p9GGvgcCzI+pRcgzfVAWkrto/mJAg/sT5iaMpqHY+mOM1RDRH/gGBIWxnw
kJSILOxfI1BUXOSOt6VtmvbZZR/T7msfKKvPZ3wmk89EMmQvGBxqCpPGdjL0X/cpgdPLfK3HwvEU
7LU55/ORPSTBbCzIUATUd43t8tIK5AWKz0NbZWSsihyYcVCo06DJ/wWyUVkedG/VhtxfAvU512zL
AUq1CYiT/1c7gHUyC9pzr8F+vLw/M7Wb7YPH7vWsRopNpLF7g8u7YC/elZF4bGlc9Fm3iDpA5usm
4P1NnAriqEVs9g4Fe3pdFukCKoTtj674wAf1lQvT/21tqvQC4rLcUJfA3JQI/qr6mdOhuskZgaxn
uzj8Mx5jBKVHBLFgpd7WIqql7OyyrJrVT1KBjCG5hT610BbKw34Cp0k/4E7DCiBJGVGGwUsLk08v
KNz7dNwctHGTPvIq0hghK+ViYKEx78uQmuWUDOOi2NlAD1N+zONUtEM2ooy1oePDadSTXK3KAIF7
vqiUClmyoeOpW4ebI+Q/EIQxiMT9rxEMa4lhtNv7FKwkaW9uLc1Op3q7AbWTyeyezFGJmYbbiNBF
2tvdA8hmhSvIKymdm2DBR3GOmaRKqaCijKIoWtKVR126HP9v3IyNa21mZJrcehhTf380uyMkaKHx
TSxrs36AmXl/V/QBNbiZi3JXaK8iwLKQLVN1eraEx3Rw/P5cJUjTbQT03DPjHrxihGqlKkP5ferd
1kEMlp2K94w+a8wD935Xt23rLKzZPL09dFG2wlB+YFpDlJtP+VIfkSvWEcfNKmhAngr3cQRaJE3o
/AFK7QtZiTsW/6zr8KJYGVc3PYXJ5MJHToW/umY8jedznnDlerHIyiD9MvkvrtqzLZDAxCrrC4yY
To+KpWxKdC0ayAsj5SQ2M/hq6omdzyd/Bk01mE9n+ka+z+TjnkAK6pF10MaAwIag1Bjqjue5RabN
gPFLCLJDw4po5ExYvcS+b6UhjBoofwB9fcDkcB3A8maOKtls6i5YYTrSUuYisV3Iy+++ywji87mg
DUiXzevwLBNhqa5L3nQ+vVEn5+W9Vxrbtl1KZmK+1gkzDHdXORhaPh8RCuQY1y21tp/10KVpEa5j
P6QDuRb7+x45vcmZOiCdtoElhS1VbpdaCfXAnsMgsIToQY3+pqOC8ZdrtJsAKhq0fxoW3v8tjzvQ
PiA/b1ST4m9Da8AJjr9Yo29FSJP0vRIt52qYRQxTJnzd6CLwZAbLUHGcPgC6hR/Hdb2m18DYhh50
Q8kWCm/2f/N99IjIBVi1mU2LuFA/5ZL2usPEDXdSAWrAc7oLCaTke7ifM7xq9DhjWgRzfiJtmv3J
YO22liVTre5ol/fEu5jP2K55ZgUwx/9NMqVLWrKdCN/6gqygMRysaziLBo/msaOhhMt9N887YNgq
LjqrMtu/XH3MJ9z3fHIXO6uCTTn1RGELU3aj4nZYFnJecybYdDN18Oz/R+Zx3mJr7OOLPTqXG/xA
WggXx7L4hW1QaEoRMWyLxfI0Gb6x6eEaCE4LNgn29zMnc4VJacaLuhsCDU9kYJghO83sed56jTTA
lU4JLjsBfGUcCd59pCobCQD0WyQHbA+N/Byyr6KGFTPanNFPrtViSZ98dd6r0yqsu4LQGVMIn7Du
UciXKsuy7uaGjlbiiCaJ5EJ+DTzVwVVmepmbaXAIw4DppbfHF5bDoYKRsEK0BLTA28aWpnMIuN99
uurUyaG9TigO6PnrJx+cAzCcgS0X9sjS6TwPWoXjLxUz/U79kU2ByFx6gxmC0EUv0r3spndMWNAN
oJ//p2HMXvTZ53mJybRurcdvjKTc9U2+2RcCdKMVo/V+wjS+xV2rIF4D6PlY2mUppqvaXKDVcoui
w/VltRsh2u5II/5iuf6Ie8qQtJUYN+obK2q5Is+TCKY+f8X5A5+YnqJSj2yCTwwLFOTsCVW3IvTm
q+ehov+LTD2qJK+KkagrMF8gsYjf3GnoGLuwG50lEX8ud0aOv5z0TNNHYvJv+TkduLeN0GCntgBh
dDmywAiyVU9IZNalPrlXzTCMOPunN5XmNZlhJJ+Dz5NWWbX77tbpdB6fqN3tigK0cDBlsqMxF8Hu
Mq/B6QirTyHjNbyjvkNxAuksU6UgjsOb2JcqBy8StxjrJL361KSLOxXnAtRuM6x9HX3W+XdPVlj4
yOUri8uK7DH6nDrcJCcd8yVKBknNW76X6awqHGTRCXu6BMZOntTxpRb0kerq6FcsS/hiCPRmKI+k
J/QmAF6mjAdMGVVCE2pn07h6MeE5uqJx+5LSjeeh1nUHZZl82jQdeJ4o7MHr/88utfV86ityJNGb
6qLzJGXx4xIJQl/HrMIcIidLWXI5HMrGEc6ydPMIyqblPSHLQ49Z1sU/r2vRQTYM6DhnK5WQ0NjO
U21LQ+ASii4Vacwk8xoq76NVWK6cv+2BmtTMyRuo7Pess01KNVaeil2d3IBstYVIWCu9nMmPm/xt
BZ4ZvYSkt+pFqbpgXfHUGBmRBieyjkRrBfko9rEXOHpUR5ruhjd7z7rUPQFL+qQ1RUevtgpULvCk
nC+WArhNGkg9XpPdfj6baFqV46Ag5fMVMulVqgXqhZFPxZg/io9S9mMZhTWPqsOL9kz7cyNQQNoQ
2Tb8EiQaVQjLBpmGhdo8Q1FToG+yY8yeL9ZsU7j7PONy1Ry74dmip8MXBU1X6xpLG1fHVAqmxi6Y
BlABcsAi89M1LcpB0bB3R5vp9m09pKs1sqgBoM3xqUNNU6TRr0k0Bk4YzG0mBNQxkn4FOfqXJior
s/Ef9AzCv6vZ17o0D9jjcDG2exTeHOr1TzZAgK6EIHsPZivcu6t31M0394hK27w35aDidoy8u2td
Ws0pV3FhhELx19s82Ogk0k2GHuxd+4Lcz1RvanCy4iQnoTboso3y+ioZmlgk9OPqz5aS8Shle180
gBlAMXfYFBkG1awKY9i92FurcAfp5bzIwtTtQNW+6IQtCR3rvNmKKeEo+qUqXHZzDdyL2d9ia4qU
4ii05Q5QXnxz3/zkt11WpFulLlUQLp5Pia6vBaKlnK5PWDI/cImeSnIaNk6Wzxxvj+nxElZJytvM
SyWTLlIvb0J7wEOI1o3grUM7qBB3+WwYOnMNr0LpkiURyJD+31c9Ev5uGHAedcqxEnGsxo3NkbZf
rgLve6LrfiOzTVgCROXB2Fut9pW2SN707jk7/VcnGfMMnsE5YNStvxEoc4Tw7c0fWjIK8I+ztFh5
7c+tBIRnsXdvMMv/2WHW4X3Vrhd02g4hNzNaIjdHEYoNmboD9aatanzvjyGwSSZmb41HMpb1TBU+
2szayTTIYUnEQa9YGR1ZnIwJc19Q130m6rbpiKfq1B1D8sBVRWGYwWrNfnrQVQY9XeUl7mbH20th
YUjFKs2xcQhH3fDWy6XgeET1HIdHH+YWrsW7xu7qDCZKocc+mYClrxMnEjDICfG4pNksAGWWmVOy
wLkGkdUrzj9gImFWs+aSX6+ucgdQV9+GRT6349J4gL1Q8zGvEyJZq1pX8Sm3FTVMdFDjnBElap/Q
u7MrypM94FPASYfiBvSYxIy6txYqs+rrQuOe9p87DffJe2uFjmbPKU9GkFzS9FuIPFAW9R4+qHBH
YZft6xpyD+VErqk0LRrWT35U9003hxzeNNOH8M3O7VRiqKBhL6VtR9U/6017L14M5TqKxo6Mzdqj
hNLWP1fn3P+n0xOWpTUF+71VsS3Nyt8W40ULzF3cjA8WrRKipEtYdyYct21/oPVY/tgT/6ZWxyfF
MzN3kxFuetdsU4lAMuW6XaE8A3OwOD71t8GQThcbUCX+SZvxtKv7UbCfIFG5S8SVt7WFzVO8tqyR
HX7i3VcCbyTrwKXUfQUoqZh5TTRRqvfIWbzN9RRres1abMnTKDQKRIHeFiz/aRHPuVWCLl+GvyjC
fCvk5nVnhgRn1AUPmtnS8tNUDV2IUyc1krrq4hlwggSCsAyQbayWrnRiqM5eabVq+rkGTdHfw7c4
R+pTPVCoof7xNMSLCBOil3gYZcIRw+HVCEUwFb42hwMfXhpIwoAPnHBpyv6/OONoVtFNGEGmR5T1
fn2xnF5DqgMgYzyJCvEAhbDhA97Fim9zVft+7fVj0ocRxNtMCO7ytJY05Nsd6kJnU3H6rt1sYv4u
7tRnZWL8HY7YaW83GC196Rtw9Vw51YQRyEAxiWaePSHCw4Sj3hEbXW4NjW458EqU3FjIPXGZMa5N
0JuApRr3VHDnMv2SsqW7eXwnICa8NrhVt57mxHJxCaJzMvK0XbzpQs67xee4atgpGncGQkT0nKrb
NLjXcm1CTtHYm2yW6VaOVa8T0TrIdlLOiFrIZAXW3GYLiXq2bjeRueAA8MpZkFzHQHFQgHLdtBPm
2iopQFql/C8AKQgKWzusxbRVcdoQXgz02rlUwa2GgNulD7+8da7NeV154LZCdHsk/juM+VWD/UYj
sn/HmRfdAePGBZ5z18SaFuWdCKFULWIx/6/Rzl1U89EsVnroNDbXY206rXgjMq0QEmuhPL/a2WTP
VQhXaiVJ5vhu3DUuVLZUTq8Ze4XqHea5GZkHgqJUWOh/h6RAFSA8OHAo5KvIJlOnhvxgpR0wRsaw
NUXmWT/TU2Ev/IyVcXnXd+0hhzvx812QjZEQX6emcd9xrAH3Ia6iKlBVFxxdXoUwsio9wdqdBT5t
w3GIG35huy9FDSDYx/tVkjOkUvUEPIGVPLL+JhJrhDUKDpXTzdRRb8fcPU5WneOs7BFl2bdcu9Cf
qUE68VZ4Dl9M0Marhntgq+QUNfT3BHODEHO/mGG3aYdkQqaqcBL8j8y15B3e4mKdggrkF9lV0Azs
HIUBumGeuTKkMI9ITm8UxmMBQ/K4XMsBbP/3tYWs8Oyg0qcM17yJxppE4zSW87TuiLvUvcGwe95u
AXUqQj5GzkUuHYDefU+C//DJhtsHnyIkZzrNY+y5/ceZ9KR/04tfWbGpf8QzQ/p3jZHI2tsA39Ea
U3W/rHVCxpSGMETDh1knV+QABCh4K896oFg3iPbtwPYc0hYlackIYRItD9u7XnUAcY2wpIZro2R7
GCpzMFLN5H84j8SZn6qG577QkhPXVcvjO19drxB43MyN7ff3wkO110TndOh8/94UTlMMu6WvvXa3
1dqBH8oX7uiCrDZl5oD0faPegJ4gcBk00ul7CDmyKp3NpA2WHpxGS2qsP5bDohvv+T2WA4qgZbY3
gpF1KrVd0rWhVUB/uldUs/uGq9BwxHQiBzpE63yG9IQ5jgiEVVYsDUFnnYppK+RobmH8+0zcFkp2
DCMzTQawQUO3oPuXtntrMqg3dpjeKf39jxLEttFCKV6D/hS1UZZrfvj2e/maZq9lEQXRDknRifCh
+cywv6n8fMES1u1tGqyddmDMTTg3j7saInyWcEtpg7gef+8Wq+8St2QDT7HgWJh6Kwir3BUmYCOP
/ZPrW/c3IV8XQLtcF9/01X6WwRGxFQyPOpowYjfjezEEjYZI5JRUqIPbPpihOdLMyQNxr7Wunb8c
Qcs7R73jIeVDrhTLKi02ZtpbXcgSo/0zGiAtuhQRvWuEO9LUXuOrXEOVdCqaJSAu0xmG29VQU8Ny
avdkxzx4FiP7ggLvLQoiDaA5YA0J5lU7Oa+h6Msz/8We1n7vWO5PvJuwdTHYfh3UZoMMJ6cY5vOE
6Q1/nxbYXESgbu5McxSeBcFvx9UV5Bk6tQaCjcdorKFqPFSzSG5zMFPfE5/CI/wLhEJeqYRiTqSo
E5QFW/JzgpGGjvwZzOawDNjZlxMcGLM5UmCDRBmlZU4ENO6xUn8kWeXuJD3xvYJfVm8BauFbsPy0
RQas/VI42EPqMz1/AarRL7xH92WiuDeKTMsoacXl99hTC6OIDYyJmqOmLWU1/B87GZZXjYNzGQqq
g1R6bR2y0dRu/ki8nKrkxYLvujXT265oLx8Mgj9Ca3D6eUe0LbwE+QllDt6vPqHZR2LFofx+zofl
Z36tbhxvuweLE4hI8iO8Uoe3ocEbjT37IHGrc3VZDmECKKq72iUrFp4iRmskL6e8ffnt6igRLh1r
msrm8KfgLMikofnMTwtTom69JmcaKhcSHrYMSpzjxJEWAbUw09zRQVh+my2eT6RhTsZqWyH5/EcB
Jh8eeCyIA4Ar3iLTPgLRj+FHRzpss0/Be1M4iXq/Mvxoqlp6I2BohJX2iTBm+JT4TqLm9yOPzV4l
Cs46cC0H8E7ZZXWwlxv3Y3wpAwxCjXQlp/viYrnQ0kSaBLIv46wMoKwNWULHuZbWK8zwQfz2dwZ5
lK7swe/8t7ZkLMuGoiKnYrkdSb4boAZ/dpzMWhqiLRUBUhhz5kvzFxII3n31Td/RYz979ltWFrwW
ezIQf6Lfj3VwTgdLYC+3UHPnF2xJHnWr4zAw/OZkNqdGkJpytX4lABKZr8RdQfln10VcvFfBPMkm
WbTw4/m7nmdvZ523WZWxztWCth9XDYNJM4WKruOyizDK3wZ4d3s5TMf2MRRHCczqwe9vaG60OI7K
7raaXVG3rGsgpfwvbJyFK1YbayNVIvHRviA26Y70py6nbrSZBh3hFRvh/hVYkm+IdjnSEzfw/QQm
Ol3oHkWLUQLugMszrVq3ShrB1+BcQQBzH8fozrkJt0x8weEDZCokOHmo/7pptNK+kC4yJefRjHEt
DGFg1Vk3MgXVI52S7V5biSsQIsTLCn89bj5GtN8R3+bk4ckRnDLcGR1+VGvlBeT7k6VJsFqXKa3l
Lxn/ugyz30ENc5FFfx+bEKj1ciMJeRS6IkalmxLAUL5Bxqw1cXMR9PgbJRqPxNWt6ETTc4BvqXYr
aBO5eQqe781XJnmX6+XgBXMczE7w/8RgvVUkfdFN9Z+mAYA4P1EDS7kmbrRoc4ow+eZ4VRNWlQOT
oi8RU7I85aqV9j2QZZ+nZ7BebgtoVh0DH8bLCqlAIeZXGYV3SbATF0g/YqvM03WDfvnepZA8xpNN
YwkcpaT8XwmdtwpxBsfosoL1W8JiL7Uh7A6ODbCAzAzHhXRXsLVQNRBOCsPTHu9ERY7lWcPruy2O
ihZB77wGof2ZayGcZ8HIgshfkiWBwUea3AGuXjUrGXglVJlFgcFJIcqjhoGH0npwpw8AgYFtPRTy
DL5ClfHYXKAzAHtfZSzZ9X84o158nFQFzaC6B2uQ59UJlE4hBNexcG9mdk48Fbg76/uXkMSZwTfy
L1Ev3GmqRyy45h2GE+HHop3HHGKsZ9/8/IfUl8wgcI2QJHBlDahfESHFmHZcT/45fzjzmv/r9X5e
/fszRE4ZsOCtvF7mbcHqbQ6rsk2ITuOzJmpP3jG5U+CWUcpkDy019gyflyd9QJlX3i6BPocWxmtI
J9Jn6nq2QegFOC5c/vT8XNG2HpUeqX45Fl7ZU477+hnFABMgYxRlbDoC7/LJdArp7qgY95uoauzN
0fPxMLVimXYITwf1EnPzaY/U9D9LEs4eCkd93w0zzvkwDWxTYBVztZI12un27V0AP1Ks4NiJIQtF
CHjyUyyiJctLyUAT8Ap3mnw6HvyNUscCSjKUk8DJrocPBw9qxCh/eS7iqm4xpZydhZhFymstvD7I
ZKWI1vEZrrEVQnmCsIfd5yN44bLHU+mft7aUWk4UrAkBqy9ztFXhhwLAON2zni1+49QLugJB2CmA
LsVGbFSEJu0suLoazhREurQ6PrKg14z1q6WeE2tJOenKlc3XHxdKP/xsFOFJQb69RC1QZKS0W9TC
NKxGsA2TSq8njpeHwRDDFPYbiSNrzKL8nD0uICknvIgzwWtT4WAdL0SclB3bH7dDaD31gX0/4aRe
D4JtgHysx2WGBDw3881DfUj8AG/xcKm8ERML9Dt1KF3cLVRhhWpNV53h3NKyg0hA3zB6yIuVo36W
CLiVwk3Fg+UDBfQxgK91PCYikRGSQC46UBuYuEjxm4zOhOxZqsSsnr6P9X+4RUsBZbbpebex98Cz
a5ZWrXXRLjapKZvABgu+hAFHOTlJiyhzXQnJCFbOMKok4kc7Q3mbpRa+MDqiLypF8yfvS7dgQLoV
sGCnsqrpFzXex5oorecvrfZA+Lltiwh84b0+d4mUBvPLO2zdaCcqdRctEJNPvVVhBBMqF3t0Wjpw
Rn5IXPTr/guh7zILdv1MxrV37eJDMZr6Gpg9cJIw/lgnb/CG6EMY6Zkez6OJvBs81wKrFbDsq76w
0HW/7tJLcz1TMkGvcJ/1ei/EdIGXKrRohaTlx3hUplIxFkuKDDcVDhMZjDBTN0TnamAI8jEXCa7Y
wGk0i0fE8hQe1geSfHwq02HyGTTD3ioYTLeG5QkkRR0+RqGJhAyzruiYERlRz/ozPwhH62TnAVjI
qVTyHtxPBfY6y67Miez88jXPOuu5NV8GcYf/+OUqf0dUHhgPhHKzvN2rFqm5zPE66befjgSBr3Xx
Rh3FPN8TP5Zug4AUqzbE9vNw8fq667+yYOOyK1xOb+Z+Su/sK6CacmIO9EE5cuHfcJsMEYesz22U
7K2ORkpRDn69h7qz+Q71zUXoODtf3JaBrKflpnK7z6Hn60m7sRhNtaP63yliXKcHh2Gsp+nXi7Kf
hV7Pc29dD2D5HmqQyYpW7jG188689edcssyYun3jSDXQaszB/oWSusheczMsnfD+m/S4gP4rxL3c
pXWmOkrVBq74f9qyAlJavOBAh9/NH/05ZD05ShGFThAIuZpMhBlVN8NAZrmipX+75C9bZLlX277X
TzDo32Tl1M+6iPiVGQMyPIgRCiOjp+WAR6wFKE1YEalAKVab+Ywi80mlj2vVGznegt8Fwzb4SMpS
I94Wgm0y5JPUMMWTxoyvZI7EaJRAHM2yK9RrRMBA1w3LdAjN9hltmUeq2yWOj5auM0Z78Qek1iqE
dB4Pu3aoeAPkEr7wNfcNaw1qMYCN6t4HSzK+FlxMq1W5S169BRvRLtbp4+ZA/NneSLGJ3x6vozpB
BErHj53X1BlW/ySc9kKLfB0grloPGojIgWxUf6Fw2nLoy2H76YTrrD1VZpWGoOx7GoxRTlKsCjAU
NG4/nIfQXWESwjlrCmFVzaRfQHv4DjjFwWxkO/Ug5v4ZETERpdmOB0J+jZw+zEyTJodlSfQL4loP
GNEBJFepfcwnYA1JOulXed1c+Cl65IeaEYTrDi37OfJQ/b8IE0PsYD9yUQtBzD06sIMcUQKzbLqo
Ou2QGikBIgFBjpQVZ63gG7JBmNUixGHIUdVO2Y8eCbO1EITm/Ln1Myk/cbUGGGKb2tda4T0IBHg/
y0ib0Q4XHxbm2+lmgmgfNdEXCUu2S+O7yWeXesKPmD1K8ibLJdS0dM1rfA2fPtwVhzkUw/fzKqtU
YLU2gQ4GtELV2cvwoag09vq3B/be3gIO8QSoYsm84K3ezkgQFuED/YxrzAlaAviwhn2B5W60oMrK
Eo8fQ6X8BR90zpMxMfl9oi46ZCJtF0cKil14MQ8RWvxOFpYuvVQYjRyo//Bv48uUy/ZqJjFhvVKB
kqKR2ISHAcZX/yey14x8Ug4xbN5E2XsChC9ZoPanCgm0LazMT8KBSuNvEkKuFMtgZtUnpv2ZIgnz
xSzkyvML4hyh1Cpi0l9OBwZpLZjv3MPsgTtxkrqdnYfZH8UA9q/Go/H0nbpYFy4fQ+oRd7cqga+H
G119VOJakNnTPsfJjyQlV+oVxtZfTHrQTwwSV7v6YDAjKbWsRM6E/8oHKg2Z4uSJfYp/WCpioscw
/xF17PgoMaM/RyQLWU6DhxW8ZLsBgtXwc6b8Pr4iGF0L0nmTnxt2O++r6g78x3h9VZoOitfDX3Vq
SsjPEoJkrJirJVnJcngOHPl+rOmO2Rq0ak15VvVjUZeyFhUhq3fSvMCllkKYthTPJcvaC/fP4T+m
q+SY8jx8pzAK0WZUD4p4/Qf42/blFaIyqabie/R3dhqd8OrpS8CpANVXZpEC6PCv8mg7oIepGIX7
iDHXMMLGLRlwWn5bvElh489Jwme78Ck5UOvq1GsMT8osqCWaEKox4bt/5ZQnA8NaGvVmWSs797Dq
wSRuId3dZG//CqHuSbEWOoHcKdoVEaCxRYh40gZq7pQ00OQTCxByqOA2D+9f0+eJbTMqaaK6lkNx
VPC2eTWdOS6+n0FWZH5V0WHOLyIKLzC/6L6y+KEoaO6cvZFmDsmaYpVptXAvHFLkOEF90f8nnUSi
GCzrCS7GCncPTtMnPjmz1uEufrXwh80fzWsqcXmKLBqrGIWv5F6HAuYeWgwp6IGvRuK8SLKr4Lir
Cv1tN+A8F0naIB0a6L1seu+tXZl4QDlCTrA3vevKIBsYTFhF1wGK8PQmNKsddg5M0ayDUHKtXx/I
GcF2X6kWs1ldFZv1fuFm6LkBQPf79VrvcGVseHh+855puKUxFneIarbu4Jw5JKeQkKdq5x28YlTk
K2Bgix9Zfihk2QaH7cDWJt8UiRfkqQ/TDCVlfn/Frac2PwgOSB/cHth9M/QrYjZ8ITWvBMcYYP1/
3gXmhzMivqyOJydIS2+MlwDtUp4ffc5C9k1Cx1JCjbIFHdY4wYJ40Q39iuPuRdhmNE8i937JpOnm
xKjnhM5nWJ1IjX4wp/UoI1n5j/LzSltvAgxIaUuVp06ynrIOr33blTFUfzZDbNpAMoSxHNpl7GHZ
NcgqYRcZSjxacYnV383rECO6gk8qZRho5OK3csPFDmsB6+XolQc+sNOjVhGbLYWe3xTz1CFg/2pD
3A84Nl5jQW64+MD4EhxYMARCZ7xqjsk75r0Q+VWKQey+NfZyKpGAD2lqqqy5ppwaQbxWfXCEksEI
mTepe0a9tRfxICtTApe5OPE2YMnt7vwPF0P2nj60W42IsCAlHtK9ycCSYeZLV9f819Y374KsPAzt
6O1vshZeQaZfTu4bwWPSFYCkPo6jCagiJvZQEkFkEHhQO19nygoIu3km7K5WGqEfWO5Fd/7HAYAi
eIDDz7AT8KQc82pwQsXtr5UIuNxmU8u8gss2AdMagiRP0foMvFOVQlI+fyihTH/cHHSWqsZFnrbm
cONDExNC7KMsnnw5IGoUa+Gq3ON0d7R3XyaHjYZF8HcCo/BzLvpUUNVghXi/i78nBNrfZwnATUOd
Z57lym9YwkJrKTDT7p/N4EevScHdXWJo+0L1FVt5NvR8ZnXb09hjPFr2/rDXly1g6rzfQtA8ONZ+
FPeaIPyHcEfVLeBT9+k+33Yi3/m8cO+hwZcgYjcrR7MljNcLVyk0qAtUOPbSHMY6RqKeUM1lOgXI
ws/4Dq3Ijees9u5BgpDOWn+6HLhv/s5/sj2YZFv6VzzqHf2eZ1QPalYDe5DHeduY9rWFs/lihZ9R
F93oPQO2nh4+48ZiLR0IP54nxUUQpMgGIxhLH+EpsEj2NneIw916m4vp7nUsdD5SxXRhgK+QUcxA
O5oiaHKbmuSv7xyRZSTSbzMT3qVzd0euplwCDribmivGfvyy7uUu2KG8Re4ukFUpBuF4a25HxbRz
4TOaNbJG6wp82UHqUf8q/hcEN/o0f3dcN3nuCC/8UoMdQumsuDLkvAjPVIn20Hb9kQdS3E4dkYlB
oC0xCiOjNAxAoEY+oC4BFFGzpgjYi7YY1kMRC4SfrJziHFiofhL61HMBN45juopSyDB80kpl7JMX
Leo73zsb3tGS72Z4Sg2zohIBci7pp7A/6RpNdoNvo13vyXRIygmabalClwdsvjVLIdHT0RdfmgAh
+UYIRYCdCtYyXEBxOb+iq5tDiHhKXwY2NUZ7Welr8o75Tann854oCdYPBts7AriC3I+jf9TWGl1i
aKeXl2W0/Q/QZ/VirYxDwyrpkIHdQKkiXzpxxQvZGV7xlNzoBVoEtMzcb7C/D7SARU21nak4wkH1
Ix+OGE5vtA1PPp9+NyR7+w7tp9EEr9IyzZ4LoqurhEemlcH+dvLZQmKJb+c0y3VYTjinMcsSBuHe
/i/MfNPJcvf0L2VAQfUSUzOL48rpNxX9pVKmoU4m96Gx8ycSGy/lea10HCxUBl6CUYqNqGCy2STj
cYyAqqtKhsNZRCf801tDfuoKOya4RVOVjIUoXe32++8xP6UKif8IdnQtyyiNxX7AwPuChj3u6kOR
wjs4Phj30tWpsuyOI9OFfZNnjR6eyxrXM8unl1OXGasXQ+J2j7ssfpF+cVZWrCKrmuBrU0d7yxSI
vtUwnOO4+cMC8d0ul+AjUZCCLPux+UhDlsGyRakr/FVgNXHZ0uIvs14abn0NmVP+OYAlPqJ1BEdp
5oge1pjLwc/fICZFqfSn0tKtfmTZWKIBu/OYOg7mfhUGC7eUflf+lDwmPl1QXbwH2W402pcofuvU
n23EjgGsnW4m/+7PtMlTlc/E9sQAMcgf6HWafEF//xJ7Dr/oAOmQf18zqOgXp2f2ImeMiV+giAT+
k/mCUpltVkEEa4+WVCDWWLpNtfkQLewYK/O3QfHtraM1G1P+2JehzfP6VTHsRvp98oA0Ee7xRa6j
AkstKHDGuJTnkKYP0FFudrgxyyNiqeuWRgeEmsEOaL5b/OT9fSi3ALOsts3Ot2Fjexf+n7+Jeg0G
WPMfEYyHpCrYOLCXbQe0rF9PtXUWMbnWMLyNv6/bY3YIVHkl7qaxeiTlnxISEM9uwCW3idOPZb0F
2LFEVh160IrKQpt4SWDzyHc3maalLJ9uSe1Xoze3mw1d7TSEsevx6Qnxfd0AMDfEiv/jPpwDyaas
2hwnbLetyfukMa7kKX2pZtc/sGrBQti5DNI4AtIVMijvf00ztiNTzfgQ/nAyUBebelN874+iCQE1
HDUtvqr+5MVQSirc4+c6vYc4thZld3aKq4jZpQom0OvGK8Y2vJQSUSM6eTA3lovono0JHVZjFjG5
82vO+tmr9IzY06+Q3o1O28GTkFU+S6RxJ06cL9+CBRDP00vGKkhzouMPtGQqAtyFQ1ySrjiuU/OS
OA57hL1xA2zBqKZ/cOx8Iftrz9o+bppCNgxeORkjh8OXhyBWnyXwxUlPHCjGmYeqweQUTM7YePgW
dhXocPT2JxuAL0WQHU0x8CJD9Uiy1UPAQYXzN9NIqs9tSpArWt9tAizvImy4RdHMzmRyDmlCzt1Y
q9MDoF/gU5w1rX+NNbmhodd/RzNE/ZlIx/HZL/C2khZsvg2XJFJJjKlL5/bFk0PGYFmb1504Tc3w
itbkLr5KHCLfq/bs8mlgvcq/NwPEG9g1YLFX75OcHo+AdDqXpKJ8ryO2atfv+dW9Rmn0WXTVdIv7
qPPCMTJObtqJ9NXCUadhGYT6HY07aH8GcTydrOGI1BeABYZ+4K6S4tyy1d9N79y3AwdgEhr9ckBQ
zsh6OwreMn3p79JhSPjd88n0lRwXdVmZMXD+W4uSMnfoP8syJi7NTzTsiR7/NWTXBdQNCOAKfha+
zkCrdeycENgvDadrY8J8QHfl4pq6nrraVWo/EJd6ZP+QhxoeSH24oJlTrEaM0KKZIYqM5ZpOGYBm
Na5Vtu7kmyht2+itYna4rt37CjKkjUmhUuVPoU2CGWS5qHKtdXX6lwG+tmbKap4W+Zu6F0ukFoQp
Nwyo/Lem4gwWhynEb5wTiDIntAvjBeRdZ7ZIm9dkWSoLKrp+1CGAp96PkIwCaBJ6FO7rtMm7K9lG
ds80XLr/zoa92wY2Ha6lSYebRVYErKX/CoEBuXDFuw50zwT6mxp7VhOQOt1ivMuK5wEUj79WTWHU
qeyq9j/4rrvQlgGpoqKYC1+BV4exwlZOavK4DnWqLUIHGGdBV85zljv0iw4g+ve159xjBARPOYp8
/CKLFKJT3VtVoqSObdALhJ/HZtzXZcDHSDqjcaDAM0Wh571WGYlHdkm5cDKZxTC/5JLAELp8Ti4W
jIjavd2uNcWtY6r1cmwHD7ZZUxKs2R7OOtC2JhXbHiGYEIvCBlwgg2LjE8bcgtUULpGLbx4kOF1V
84+qcqhJBHtgauwmKs7rLg8sqgo0ijJPm0Kv+5iQpfabq4DioCC9g0lcyUbTXqWfL2i4gvR1x2z6
5Yzv6q2avFBNNqmRBO9WS5eyd/wazXFAM0CfA03wbxezfLcgf+IiBnfcSAXTEDL3+WdwhfzmtzGn
2RelHQ0FhtdfJBlhZ+ec3hWFN8zgaPQtvFndPoVIbxHI4/KWXhqQkLoeAPJdIl24fMKku/xOFj4S
OxWo2VUU2jJQKCr0TYzOHkZTyOTK0XXIydx8ZZQJrXmGLgZOo+U2E7D/k4aZVve5jlyRXVOD0S4H
bST5Y7YOHWcXQP2rv5EoWlp9ZkhHXeWNQuObZkdXQj0oi3NngzmqsQ+R530/eI32FAHm5K4PXrHl
+H+MbYURkvkzB9IyBCYmMaUtbg27HoXY1jukxWyx8d8JSLzpaK6FSJRCeOIPZO3sdnkw0MpgF+jR
cvm6TzNQdhhipsO/H4vyQI7c68prIQcPFrdiuFVKSklcKv0WLM9UUQgN70PEe8eb+BV+WKDSbVyS
YnbFlgDeNCrzC2enYHlzsOlqkUS2UWlIYJdVJur4zSTz595uRHEY96S1yXXVbnbxifNeLg63tzd1
2q7z0m87lLBNmN8ggb4hPUYM5ICvtAt4unRp5i+Yq9plZ8ARv9kNl+3wTepYtFPc4iSAHHq6xekN
kkO9gA0FGhM3EyWoIbc4isqiDwLfsJe3Odj1e5ZSgPO7li4Z589xNjT6l6q6mTaxakVdJ4qaPVcV
9bxYd/UvHhXBWQ4ueEtUnsjDD8hEGzwuH7jvhW+86T60vIX6pWuZ0Ih6smEDub00qYnp5rfYe0K2
WXaPQrfanDP5odNyHR7HWgvhOK1BBOs4gFfguVZebtDv1vSFEVyLJZZg4hJ37EMs0EHlp8Zeirei
j5l8IrJImO7T8Uilc76YGWYW+ypaTRcehyAnOIFjD50TTi+yD7tTOzuuuvporam+da6+vb+hRNRT
L3aa2F4fE1F7vKp594k+HZAqvZlxXzC+VS7nBBvw79ePF6N1UndU9geKxNGyGgFXhpm2TpV2R0TK
NdZ9M7fNu+ycqC4B63FObNhASd5Hg8yUeQ4mvCHyqz+lixHRpt+nShlzmvMiLkWb4qdRuchw38dp
ofGbRbc6ok/nwF229d2TQeuA0Doowa2FCoLJNljtw74C32h3SmsUgBKHjFyNahPWazhTkMQ8v+J1
QuuiUUESvCU3guInmEElzeksjgBXdCrH6HeA4JGdyN7q62hLkhhk+TXPu0fMkld3D/igay8hX1gJ
D1eVcRX9ad1tesGH2pZXjz4YuZhpc9xjGEyT3A/l3rWMWIp5ITzRtE2Co4F2xLQpE2hf8cF4m0rt
oh4un6oei9cwfZuEFM8cDnVO/wgwMr7kbpanzGjJa7Sv/V/xCWTQHXQZ9GDAcyEivhu81iXHAqE6
CHuroUxX81R3WTcwmZoAfwYFHyoNq0gmhJ4JMXyCx2DyoIUYzdcW2KRAiSAjPOhkamhuu1ohmN22
tmWPNhZAJJY6zKr1/0bVlNxtOcxXm8nRFr5d7h8cZXJ23le1rnsT1bAaNzW5X291/o04ENIh97bI
1CrIZNhmrc9Q5JNFWCeURm3Xcq9eLkvUsXCzPmXgCyj6E3NPDS7tM1QHebPnNIZyasFt2uTYjy7p
Lwik3OQCHH1c0YzRtQIfqwEAmuelhArk/odJoGRJhsNJ+fqSsRqB82/mzpANlafF8BSa7w/C7odL
hjJoW3Qtbz5oa3QtOqbo35GPJShke+m9UkBxG5OVmRUVurkYtd6SwUvknQYi26NINtX6BcM4/QiB
TsZBnDKPgRqDRrya+NszEWZOjckXNLfV5q+6Azd+JC02N98DBKbJ1H5Xn/wopA7ZEQlDNlCsWSHs
1mdL7Thv8LH2dhNhzp1CIuONJMayergQmQ6eUIL1qXvuPJzM1f6KDDQLYqlNM8Jx7F8kAXXbXRdb
zC9pG4LSQ/GnQ1r7Kqk6cKL3zP12IKp9HJSv9rZNVRdSRBOwMVxyM/wRsdLcf3maMF7USUhFJWUQ
TMKNKbO+TSYfN0hzq2QiOy4fOlImnliu0JFQ4PbxDOXJL1+jTkWvtLnDhJZ1onrGJMprsPV7nNJQ
Sb0GM92z03FsKbmjKDvgwXRpgjQ/RvhvEz/zqwyImpuomPjWgiVzbllVhiu2S1mtcW7WXZuccTrY
ZZdjksabAvrLMRqYujGfjJSRoN2mEuEr6I1u5q1dCE9/jAWySM3sivqcqOBQMu3ZL9s0FwjoAlvL
id1HeLqX3zRKtG/yGyRWUD5cFu+u962pwKmvZCJydvJ0vPC7JGq3IlWe/8+pypQEJWJLn3UCBLpK
SgP6e/f8im1QKALNi36OUJUOCiVPVyvH+SHHARPUC85vdiAZUXDDH0vjE/qO7KGX+v0EgFNEILR6
XsfR0h7053766TYfGC5tYyysl0tjFQj80JT8Yskf6iA+N6XWKTu2iLV39ea8I6Q/NCgNwK/3Z6i6
hkbTbdgJKU07u9pF+sze3GddBejSQiSgrpjeL/k7YfRttfQJOcwI1jNANJ/UurYqo9it7joFSTOq
QZWaYiJ8lGrYPxN+K0Cdh9600VQOIOG/d3QRCYIa/uVsAfeiCvPfZLDvtZ2qny7BZv/SBeuXiKCg
w0glq8kdXHzMCzIlCc5yUzy9fYSwUwuDYcNtfziQNfPMEAZIhw+Ltj3DlfL3RyQzuA53i13FVJWZ
TTZngRTo+/WQG86VkVYusua0VoYhMKJacmNRBPd/qbNVZf+F89nnhmtUP4q+eqrsLOhrO+hylxel
9WLRbkplW8hrWICaigr2F+08F/LZcttYyO0MIM/rCJPIJkOVtki6bY9ae6RbwR3eyuoG90cOpRoR
WzQ+lvTGh1s4LYj0XrnYUZPf3n091+5CTktlPO1/bXehp2ugDlwrQLtSwxvdxL0l6VMLUM4xYknZ
Xaz+CXpqbocVT2z2Ye8MT5AKPa1bmmuPYQLUpwy/SwLBizDyJvGFlHqYnfgc+/AVEXc7f+T09F/F
dy0Wqx7D+r5p387WAy0dt8OzCJqnHo0ArIJzsP5aORbGL+b99tYHuE2MOGm7f70NrlrNR3z/ppLr
TDH332BsMzfUgJTUrFK/Fdqmkht5pKs+Us9WESDLQlsGd5um+9smBVV5yI5tOkELbl1Wc2mM8F++
gVDsv+QpzrMnw94Jc9xTjoWUvH2Oh+EaysUNvDaJubS1T4gV5/eGhrPT5kX9fWG04JkdqHKeRg3n
UKBN/Pa3Frq6mYiYJ2xMXtriyyBU+Ff8ehH7ilMTlxLH/EEbcF3dUStrf/sH1y8EtBKWvAL3ADDr
r6AUsNkxkx8ppyDkxmeBuhT5lrRPfwJA6LnT2B9ueg81Bd5BLaiDfHp7ZCum5qomC/kmPwsWd1/P
C3+5AVkykWq2466KFlbLe6bqm7xEU+eu6EAgJShV966w6LsOmcuBO9czqOhxkavJtDsu4mDQ8CZx
lGKOGY5caHmMBTZ673jdi9mbpWr/2lwzoi11+ST91bzT3CRU1ex4jJeL/jFyDIoW5nkVWnAhR/I2
OZtNirsJwoO9zAL6EMkMzwxsH00Sg2O5tiyxNLlG9TneJIMfIz4V3yBQP+onM6B+tXYuY/jz5jU+
D5WN3Cn2AYbw6+xU9dV9D/2002BdFV2OYJZhIvXjN5m4joSjt4DF7v5kNFd9R+/pwSV6RsFh2JqD
A/UQCBxYOND8Tsah41KBQmr3VX/O31F9aAB21fPe5/Vdm2blWYUjr5qHI4y0YhItANN6klDFFrRP
FBTxnaC7LHSQfK05rqEalgJeUttLSLpwvxHxTyQC0C+BZ5el4NgI94Zh6A0iifl5k480Xso3Nuwi
GPT9PLfQrmxB5vLtvcONlfqLAyq0N43V0uJI7ecrVP7hp/RQtQBBXCYUkS0BYaQUdPln5rmR+VsJ
2wEzK297gLd9xM56PPMA7gzsT0ZC8WRIU91LaBUFhKjQy/m8mnKfCc1lV2A7F9j2Z5P6sXJR0Bgh
uGLmwuYWBcty9M2DEAW0gPY3vJ0QbMaYb2Tpbcs56118Zuo9rgso2tDwWqoMu/udPj14oG/p8wn2
RY4DwcArOQtmGsPpuEwd/PbGdXKXI7T0+MriasRGMBsPgORznA0ygfoOSFLDhVnw8eSiR+hukspt
2W3o1mb/bCZ9W+XfuAoNx3Ke9kVTqqcbkeQURTSjbWsOnKuhtsAOAYdD3s7mkG10XFjo1JallrM8
Jtsah10BtbwVAiTneYjZXOCmKTuNtF93ZWwsJnZotlaBOZmoKfmc63nbaOKHdO7Oy7C1KmH5QY1E
sAY/PLsGZ2H2DvV5v77cLZTOTHbrc0vcfzfPEh0GbdoCwQ8UVHB131eACxL87Dj93LdjGoCWXWWQ
FY7h2POzqVamGd4k499WeCg1DgYV8fJXQ7IxiL0JLEKsfFIJK5vrgbj1gW2ExN0WqMZvUobPG841
f8m1PdDbhBMITYQ+gpCfJRwXo0j3sIHO0hEW6iKR2IShZFd4RQnrXeAVmbLj0BZqHthQtJAohmbJ
og31V2K7+kJHXO55qaAQSO/w02M0h26iNya+SHB+mHRsK4j9Mx/DCKjo7EpivBrdhFg24llQsr96
bPI8k3/fccsWvlrBeMQazD/liOyLQ85fMHUiNo8oq4qvArAHjytGA4AZAyUj3tKmUOX80n/PuOeB
IMfUB2jcxPsTu9ceFMLoS6XdZzwV72SY+Z249qf/aweFrjTBk7BjDDzIbyYRy+OQsPSRWF4eoKXI
2/gWFnqSsxsWvHskAjQKQbSXiP3HQTE6CyiU18L0ZD6Tz7GJgxnKPVV3rlN6XMQHEvCxnwUuo8/G
pVyKLh+H1/rGTAO4cX9cD+g5iQ+L5kcOf/pcsFrRAnk1+BHbKk5OCuOr/ycTZIwQNdRrElj6Zoh7
x96hGI18xzSkpg6FQU0GYHO0pdDe6IGvaUE29GMCV0RUkCbf8WjgdOgUR0b4ZGHsLHp4t5pTfpqW
NjObwcLTXcAAxUBJTXGlACwRITwJMt2h0cSDvu2YiO6nT3LYGzWt87sjGFdJT6Etm0kMtbJ9mPEx
qcx7eBZhZBUM0CiAnnG7dOkwSHRVo/Nsj+7ehgdCBIG5YwFx5vi+MogQO6lwnh5Urzf+Z/GgPkXt
C8pjn8tYUhzUoRjkYHg3GFt6Yr0wXa56gK3DXqq2aqln46UmENHjs4zFelqP1SitfTdOruU3ngB8
6A95BH4zW3K3TCZqLKOrDEqu4ZFXzm9vp6y/ooRz9fSbPA++fh7zCkAGHE3SZvgmT1+BUcGK03EJ
2lpavsPCkRoYAjf5kCrquVXgZwm/xIEuGXX77mCNzHAS8juy8pt+intImCtCeMlcHzCadj13E8cr
oiDyDeCbY0Zt4fkEO8ItPiXLtai6N3Mrh2SyIQTkVswmo/cH0u3FsXdevMiPRTNCZ/k2WZnecmiv
6JRkAFhriUhM+bX0SL80Gau075Iid0E76x/R1KpIo0pFd11kSc1kOwxzw4TBSJCVcJOcNvRaA7vc
0H1WnYqPITXnto/uuHklG4IMXhkNLgxuambXNiSN49Y1+14hr2Q3EAL0FIyzAsHxMf32FIBZBFnN
wZfppzM0Zmc1UYyEvr8hoR2rS+dzkZdmUjAVW3W3negu+xjtBlmMUNBkQOzSPLN5mw3CTy+H6OTe
efzRHivwMqiGDvDNJinegP9+1y9/ou4hOgJADdeN/1pCxIVvDUQatLRDYSOMiDDsRBqFwoa34M9I
s+UqqaDfKm+irfZ0TPSFe2IEFegkfZ6/w+uKjAFB6OoSzm6mbIZCbjhybJczK7UgkQRgx4P19Wj2
UZJcLDGvR7Z4ZYdit/RwMdze2dlfiBcNWo0QG0AjXiq31G/PXMMseiwaVIzF+1sGINRmAy9Hg4+S
7QDoRYb078xZhcay6KXhQrOUcRAeRmc4hLT+hH6L0Wr/2OkqdilACPGcLzj6KUdDt4mSrwHq/DvT
QEiimU5BoV0moHyFBX/EOC6Yc6+kF/PsK8Z4zKk1udzoK3ICJnj9HaoZY2CaABXWFY0k4QhD6MFa
9gVq5/ogCX161AxpFLZaynVTjlHPNz/TJT8ljfb9aNvzJjVruV5Kj81wTREmTu1OqeQC4BsANecy
ByiI4xRqDpxDNn7e9cDVtvuXfG6hQztRBgVyskyUjDg4dsxvKN05oWD0vLbaiVJt9G5NBlFHkWNy
mTpMhmoR9eklgAsPczRJe9bYluI1SLnymf+H1Q+499yOwefRXDi+ohxYiGyw/n7TnoFbSSKRLycV
XkyFczq8EB8iX4GBOc/MA8xk/8l06k54cNNZ9ROQt2U82qh/l8/R4dEm3109/tsIgqJuuRN79dRh
UPJ91H5uf2kSHyHuNnX982K/kFATPh/ObJCoMM1b/Lqxtn98GZuVPHS3Pq23yhEBrj9ynkF5bwj5
98J6OVWM+f0hDqZfqbORQfY6hq6tSz8YmyN9yAI5VxdyywMrUEp1re568W6f2Qgsgrrqxubph0pW
+GPxgQhKqNzgqpzrYmjKen5aXO33O0+OtmWiiG2PsRVHgl7YkRhOvmpqeLEt1x3wjc/o6I6XKF4Q
Q5ZudxvdD+iArG9UEzNlxMARYXqbWn/qcbG/+/sD808gu/kKbBjKV4i2TEIfHWTFK1L94C6hskXd
mu73uJeeRmuki0IgzBEIlCgwyVOkJ0mXXr0+adIk9eRvt/DwbWKXEPRExPen06yiFtUur2dRi5T+
MAFt6HiI5l1EEWF2+S7Ty2jMc8U023ECiUYJpGSjKx1LlIidVPfwyHz9ERw3VypMHXoo9KxsyCqq
/3kw/3ojwyEq4fSpBhLaYSeYosDHm+62ePGGrTIatEsVhqN8tDJ4KcsByg4+a5d3Crtgn/zrukqB
7tMMJLipbowo7gckXD1kUJHMtFTQJtNOVU9LtCmZip1kcrBUW9/JTzWvYX5EKmvErVKUfIx2JTqi
6cKKMDqaQhkUeZ3RUkFLdtEQRfu+Tdvso32wLnVupi5JcKhGyVIpRmTJdYI/IAsATDLq2msttLmW
OVO7bGMrjjH2CHpGMCYYjfxO+mYwi3HjeOygeIYuFVF5i8AQV7LAUmjboM4GIJMmtrLTTNsskJ0w
SbL7paXb6TjZJ1E8XjYLl3wpm6wAec5bilEKSgOMX8wkQ+p1lV+j5lOq0b0uu8ml2yqUdi4vF+Bd
CZLlvc7AD3rnXybpTdY0bPyh1Xs9TvP1poStEvxAb6r/1PnLr5/S/NMTvGjECPV5ifxrFEhXVJcK
rAyRr65JB9SnQZFFyTeYq3CsVQD8AYqBL07iCaQ2pW6xPmFPPknMXPDuRtiiyKWaCxi1HA4C1nFi
TbOlYuw4XxiSBvpXMAeLyjJnbJKu02tiXGqNyoYAyC2/NImQvKc79dpLRkFvx5yvModJnFD9jquA
6olGLqSITLWJ5kUoCkN/qXhSnFm0EwMluXbLlTkBGXW64BIvv5vxkVHq3qPJzCV0HcdvM6CqDFTu
XWLq6IZJ3yUm85xl2tmUzVuF68p5Rf152uMx+Ewhy98P5KjwJaH1ZNv5QS4Fk19GWtCSByIgVFDM
EOESq7pXwfkx+MMpeNj0xV9R+HxKWx7LfF+JntnELHw2TrYEQXXUVD7mnhtSKuzweLQv8zD6aC3i
pLxIHpeDeXG8/oig0BoflvgToSa0NlZrYJlivGFVEwXuPLLKu/kTGQQ7DCv/M0ySCMEeEvctCsGI
K5UuqRamMQ6RhzrJBsnYPu2Q/fP0jhKweor869hhpwGPbbCOilGLDl3gQhPcCouVDxhuUCc0Lgs/
DRiDrFjl/WVC6OcJTFQAx8SzQe3jObbssr4t0RrR4ct+PGMPR22CXhViOwuLDi8XOOqLE29UbM5B
M64+DLIEIbav60kVA8eMx3IDXuAzVF5oMGWJb/AldOe5mALYeIjCjHnO51nuGHnOdTdb0Mpqd60W
lpuUL79So3YBk40Z4LECAH1evRevOLos656fuscn5DOVvo4B43UNa1erVSld7bZP8UetKm8oKm0R
8aDbyEn5S42zCIy2OoeR2U+DSn42EkCm8ksBhiMURgIV55HDONatSf8a9OSGgGHRNSHtXkdQ1ji6
zO2Rt7ZXAEGUmrla6nWKGEaS7NZ5rlw2xuVGAT6RzasJqc0JOzecskpXLGXPq2I+wFl9w0+GRZ32
IKMHgACneqQ1mtZUOZC/sJrYTH+sLzbHf7hXepk3JhrEm7d2iKIc8U0wp1rwP+TwF12HLfdcpKsv
vb+fwyMSzpf6PjIcsOYO0G/nkMuuJMkrs47xPU/7ddREUfnYEuicvlHU1aAXt1OavcTXZScLVdoa
//VXymH8OkpDJ8TgYwyJT/5DDRnNYUfGTynazRM6DNFUgWw3tL7r+hkOkL3R6JI4pDsRQ7oaYhzO
Nx/d0g6gkJztUg2sNXpz244AvuAZI6R9eTisbaQTM0iUpmlG5ZHBBXm1U6l2aNk3CWEtE5VnwtDE
0VkA1IehWhmn/dLjjM6ww58ip9k6YJZxEfxkBNxHbmqG2UkSfHBBLYJcgxhRKVOXy9DDsBYu2/Eg
1u1S04FWiZLNh3D5J3leZ/WErGNsJXZvHO9h6Qps7SuZaaGEQM60LaCb5ODDFvEkiFgMsVkmjdih
j3FE+CosvIBFjJ6p7eGeoMMiYas8KkbBfeDN9wFlsGt4fYyNsMIG4VNhJDn9wY9+6dSF4IVwIvg3
w1WaIoQxVPV+WQ+mU6/TDvS07lv61jDCqCm8kKUFvf4OH/kufFXeLkorr34J1Og8dpjGrK+LIY7h
2UxzMGCCk6huyc3hED7nvKT4ZnYXAen5Q6NihPqXSmtRjA6AldyEILwqqia9XpIe9hZHhdTBShPy
AC+k5A4mBWsLl23qFpXX1Q3dtv5x213mqKVeLhVffFUcDLQzQj5R4ohLPZ85QJiCd+o4UV0SgSpo
LaHkmYdY4Sm4m3jXwb+u0ntR3aD8qNrBu1hlB9ZaDJIXnWqr8qYqFwp1riHed9fLV1iiDdpCJIPV
fFUOoyaVeuzeoZ5mBSmJkBXA923vlbWbL73tXJ8Kn0JPpKJO5G8mtQbbocRBPaWxT0+t6Av+7Tg2
uamWhGLBCmy4q4VlN/209bWhG3cGzdGtIdGuj3QL2XnY23dAL2V9VHVbg+HMzUInQy5qXDJiXdpX
Nk1g0Z5tWR3D/qGgCp7StmIFPE8mlV44kRu9g8SKHHEC+QAdvXa66ONzzah/m7Yn2uvVlteG3VRp
zjpKeozHGRs8AhAjkNRWPeR50VouyOZAFKuegj5gy5R/hSP0V9HnQOPHnSe9XIGafhQx9YQXmCNK
oo8dee8zslHn/Wn4EMPAGsya1umf2FE/xV+fW1IXDx7fZCc5fN9t9QMoVJ1O0lXugGpWk7bnuC6d
g/0GCNlDH+9KM9X1jtmHNmbtpe47bVlY2SiH2hfrmKjo+JQVwijdn0UwBuAPSEyycOR7Y+XGMZKZ
9T4VWERLzDHFvv0mjQr/Ys3D5piJ9R4t0RRI/U4tNO8JhxL01T0LCvdFmvlBUQR/HlXtiMB8EMVh
cnjs3k5uSLLESpJPe24I4KQgmPnxjF9Mw/XFlgGyR4XHF1MpKyFEvG2i3BhLMtljSXHW6/rSgY5d
+DS+7jVwUrMfCPrDhu6JW/QVdsU497yDvj33x4otHFdk1ve+519hxY2LufwTU63WsdJ69vhcbtfE
UY3IDtyRODFCC9Z7Ann9+TC7P0STxW1pwn6SiJY0RVnRsfBDIQsVV/AxjaTEwdgfpSu2UfnBSLFj
tCE0tSgggQadu9GAyb5Ezn9nVBKajgiJmqv4uGOtrWYSP6oCOpM5aYuNSDPfYx7jJ5k0S2hHeInp
CzzZLl4Q83Y3SDRn/n+8zwMch84Eo2ePbztVK9iIvFs4DyyDA27SL40U3UJWiNbEyZTRjrBXjmmx
eXYKHZIYtJBV1ayTWD2p5ANOobLL702UivnOeL1420mGEgTbbFqDCWVCdRTcrAVgReYPFPxjnfSA
dkXHP7CxHqxMrHfb0PsJkVoq43speavXgRmUrr2pHr/9rCGEzt4h4tEV+pHptl7Kap8g4WX0x8E8
ga6dRD4cALhj+ppfJ/7+6VOh9bi3seF3S3PAPKhfYyYuoIBIORI8GOxHM0t6BXxLjXbur/BFNYNm
DtcBo7QkiY6hz8uGbqEwb4pmQGQM4v6jRDawAYHzwiznJBi690IWvAZtk0GzyYhxHkSvHTTDDhGT
Y6U1te3+F8K9MbeMeNazWjKJzZIY5jHGJQabPc+RDYgHrzWDXlgiOcIsQlm9LMK46UvXkRDf5x2Q
019kEhAQ/HQbZkOW/r3t2nCDJkMjok5VRjoba5b8XOWYbuUNJ4dPiwiiLvonLeaq0vpdrcv8yyJt
2AcdHEYt5lPhxaISuJPnzucmUf3DtSy1JzNcz5nnXVMB1ola0H+9fFRH80dkLkEChHRsZMLF827x
Klf7ZsXF9LRVZrntP+AZOy6YOY8IBEekSNGAbKIK5sEFXF+lkKuB5NkKglORYA7XjD9kfASPi2He
IqHN5B+rXoQaT65Mt3o4O96PBskf0go3rbp8bcazFuFUf4G3RFPitnuWOuk9GUn4FRGzeySno3iW
DLrcn6TTimexlyiTqDwevlL/Jg624GjSJAsStpnGOSZXGaxkT7e6hLtkKDlgPS3vr7xC22LA/IGq
v8PlD0bF89/a9R5UjJCDwhJoXvRdJneGLtbZzmywumxBBfNtFa6OrTXDOXIDB/E8+k+m+OsKNerx
yinSuaOVWPtjUjH6T2KIKcbofFaHLt8HM+0R6Vt8hx1t/v8Pc/LZF+CiC2uUQlYhHJbzCXVps05d
QBwy78RmlYpEHoH3jM/vDIYNf4Cn7AH/5sWhXeN3+2rm3nXXsQgZ0Ifq8E20zN+MXkOStE8rzUzK
RrISNFMlMmtCU6C4aoEIHIar7JGuBsxjdYkYnWnzK7eBAsqHIhJUb/KTXRA8YXZm6VGsG7YP+ZWd
ohBoPCcFb+AEWiILWeRfidmlYPm98V7u6O3RQJgNLIeVuIo0Y9Daa+3wTTbhN7h9BsrQ35LTPmvW
DDNV9XOo/UNNJCFmbIE2qOUpYXR2TmXt9qszPDa3qsTkvc93mF4diXNajLfoGft0CQIVjo45CDZG
7qV29h5xjMHbVtZQsdgIMUZxxGkfPnDnvpJml4ldOjpEB8/peOiH5tT2/u1hdYAwbb0v17rjNXph
MzgAcdaLW4qmNZoQqZpxKl/+OyF3BZV1F2Xn6ptSevPD2BCojjVLyuYHtmSHXGnpNzntrfJGJEJ9
c+tS4N2mJ31UyjmbYbE+txxbDTa+pqa02oewhew/9FbflRwgYSv8dITO1LGaipfTzO/shVcV844r
H0NqBgnBetHNoZZ5lxvD/6WpioNZrczHAdnmAHFCuQBpf+qgchtS+FpWQlKiHYCJ66PBdzj4JdKk
K7PiVyhBY0zp9Q4riX00sFBlA0a22rLHAxdTMB2GdV5aGTT0O1R+8C22hH/wsZMbxuvKWh34cBig
+UgIyHSfxCJZ/CDiRmL2pLvw9BYQLyoWtjYkv3zl2b+g2WmaJZGO0VhvRnh9nxOLXdIPTBSkb3e7
Wl5Kap4p6VFbsBDI0klY/un6ZY+Zh8hgs5MRBdb04vqm0b5FUe5kNQ/aDSxc4x4zCHHy+rEV9MDo
IAxwlYOEIgXIol131C+SBZvtawBeHY73y+vdmMqaRsya/2CqBkfdLx9TlQzYQhEXuudgO+rvqaqv
xGZiWIRm+TW3h9Ni1w6ONSuTijRu/NoEjY0Hvdx/WgZP42oGQEApH5wb7eh+a/wxvjlc7QoujJ+m
89rqVU2unZbSQ6AkKbAG7rlLixzzauNH99U/tJsnYRmHbW1+7Uv3qmAjtQx7uMilmUr4VPUyTq7o
DEa1kfmSGaNg2u2IJ/G+8xm4hfW/+iLkhYcqQ1JthiychoSSjl7kDtG5dHMhq+k9SAIJsPsUO/n9
1uZKNsZjFNiNa6lZktAQPJ04jDFiQi3IlserM3Q3pu4lWs/P5M9naT5nzG+Ud0wt7H6+vQGOaaON
ogxK/3zsxksA/3zFa67dlNwbGKvMHolKKP1cPugS78VaUXVKtAR5zvIvduVfJtChLsud2qyYPyV+
lCQR7qBYary8ht/T1BQJjj3MAHAZ9YCoB4lnzMyrPykNqwet7eKiGX38tgn0MhFywyF6WRqqkNrc
rSLsBDyxI8EXdI9Pe2H3rddWrtL1iZA7boBXy1pd9i0dmqR03fM9dnNF8pphBZ/1ujB6e5wG4C2M
GFY02rWle0CzJkBvIxP26zUtBTBRpUqm0ViOsXWm3NkdrabBbfFFEvJxFZ9lH5Opwn9lS9R2MghZ
MgyQNwxeYQbCv+9oJXoqG/auTuuSiXu80YyZhUkCu8WjCQvgSUjy78GTV6aci/E25hnUdKNmD57D
pydLF/+AheTmMsa0sdMYjg4RN61C0n0JfcpCxD/B8MvIqFdFT2L/sgas+tIudTJ4RTQTPQCp1ep3
daKw72lk8by+Pmi6CjQ+EOCuNnfWBJDcsgGeGcJIoRubJVrlvNlcVZQrUSE5t1LE9Pmz0WAEXyxE
YW9lU2HbDd/kWeiBKpJICjbKEd6SsJ8OIExt0xGPafujj4C7Nt8fwk7OD9Sp6isBRRIDrk4hMnbc
FzrObX++iBzzq0QUevb8ButdcCaQutr5UbRkD5504rMFXybKGIRHQnepa07NhWMNrFa63eJb9WPw
Y06b40vI048y2zw88PmBQXI/TowZKlA4we0jGPjfHr9qc40aUpATUKsoiXs9Ifgb10dO3q+hectq
PQ0rqQku8Mx1oVUtDLRfNDya5pAqNl6xMJQdH8WN8C1vZP0bv1VHz3sfGljrtqv4qcgJSZKGss8p
BYbjHdGF7QQV0/GDzSQl56Uzo+SVzuhwSFjRcwzLgrmqNXLyaosaW4r6BIspwuPwKJFPdGsvy222
z20akbh5me4EHBmKL1bqc/dhNBQDyTPuZCvjr7osMF8g+pGOXs8/J3g+qcoXsY+N0OB45GzrkyBk
nnox0yjxRJHaToiaztmrADJXSIxnQZe9bICTbD/vZgQ0ZaeDG+lscxqUw4bF8vq14sIMUQ7MiN2E
GFrLQzz99qqqXOv5Rv98LyWfuFEnPQUz1fZb1HP4MR5TXEi8NF6o9wzonmPvPCkiUH1ZOrShpvZ+
HRuKpHEbvJehFNcF/qMVzf1kqqf8nl7O1pOUs6PZFtXO6Or48kvFSlP/zFJpKTOsTU1PfPNOIfHs
o5ybDqnwYSK4GbI2rkLFIbdlLhnycUe19z2CcA05z3zKrXYOckdsR7mMdiJVWGJMZMjMa1rBVf+j
VB+pdjSc6odDj97UQhZFU1KqwxCpyY8kT2L+nT9uTK/+YCTdOgcKGrDupMvgaSgRz2w8mVH5LxSW
xFJpWrTH5dLIYHIVBz3sLvL6VhPcYXqi4C86DlsseBZyZOU47ESosDgSGRPJACUAv82NDBjlrNlx
Tw4t7qpXIblTaKo6x2A6AhR9NZF5NplxnpVpaXaH7IvuYCzvQ3O9UQbTLffVGla4R0t7STTLW1j2
mppBYl0davmmJ+737lBKQDHIvjo0bpz+6YvibmDthceUhCZEH4U6Kqmllg6fZ/6SDObmrEXG1N7n
t11ZKSzf1XzTbQGk1rEk8OPwERwVrPUFYHVboosZbKC1cwt5Iui0/X1uyAXlI0sTHCZnEblYjD/F
hAEdowLp6u4gJ8nnb4pmt5sQfPbXzu2b82SXBCxAWHJszAPp0/YygHfND6mDVrhFdt5X1sXi7aKl
LF5+3OarLgp9VvPCchuYcvNzR6v7lmfafGswW3tEm+uQLqPpBUy9brsERLgvFPsySVxTD5zL8Xx/
ZigkahyAXQxE2gUBnEMAkZ8sXjwk10J/s2h4/Mji3zQ91brtSaEBFECo4G1mRfscphfRzyLsD50+
7e+Hf8sehLBdky8q2AwZlLM+XRJ7As2knWVrkotXiNA6ra0nWl2uYZvO/lhxnpq8HWWS3fG67oIl
GcAWeeYKJZYkzo++3FqNWgyeeSqyJSMuWgZEQqisy2itLw4NoZ16g5iONYgWEviFSkDYw1V7CWK+
V/wPdx9hwCuArns656qRD8Wocc/BExC8mG87RI2PBXxAQilmhOlbnCAk2VW1K2oRu32JU2VLWvsi
Plr3+3N+n71uUXRX9zGRaBM9ZdoOI7A40yr7iA+lhezf0t+H4boVRwivIymtr6Wh92RplEWuppR8
w3jXq1BbJHzMhVksLwlaRcvmtcoMiQuRfHK2qsXVJFV1d5GoD/9vrumsVBUK0jNnO8No298Cr5FB
lHUfL9YujgMRlbZujG6SHNoFV6DKLQPZfrF72125o89VQeox0O1kuKnDb3nWCS6dsXTOjx8LeSlj
dOPUj2wWe9o3STUUzc2oeVcZPfVEumDg78jZlMe6j/dQtVQWHg3NX8g9PTKCugBEEmoBoV0QQ36s
E/hkz5AEsCTDTZP4yFReJm/N548dxJut4AHebXbiZ8HFkyHsh9K/oUyPkcZS72tpiNjwY8I6qD6I
Cr10uTNfdMH5GID3Rxv+Fn92ZEpJp+uhTG/8m4n7YGSTQRnwUXwTlKCVZs3N2AQCuMYJ+oOAHZMX
7+xEitmLBtO/urcRRv4MPdpQ5YqDvhI2h7FRrRJ5aP3V02XAEUrd1GmFqOR7N79zvbrRPjItXTaR
uJG6vsKh7RZm3zkysnB014Xikos5iKx8SlA6nzBUcnedCxriggofe3kLGE4INJyc7j3ix9BHBabh
sB7j3KXitssaqK2b/X1HEBvqQ7PU59ytGmRMAyKdmKcDnphmix+4sOTmsGta90HPpMCtM8zojVOW
f+YpBuoxHQ2m1PsPywOjQ+RkTYrV9Ef63tSZo9wIDOKJo8MG6+1YbLo2/wiVLcNf3VyL1uTKnMqC
6RdDKEJtY9EBzPpmDj1We3YS2+YRHdCzrEqnHsqjHoyLVKoGxQUia7C56GP4LpGkud+IxAy1Op5g
ubzHoaHFFmfKBHmZP+3x5TKeqPkS6BFA+urtLbwtcxOulclsSI7KaTfgo1s2eHO+LqinRgzJtSxI
aqOg3StHpJx0OgFz8DDVgFqFSn6sHGCYQE2owUAU5UeKjvl7wy/qhbBm8r02JAPaH6RsHc/LABTA
v9uFlc8KZ03YfKc/nbwPsuKBK4EwHTVD8IKaqdTq24ceNJIsfWLabwOmnEI2uRk7lG6Pk0LtjAZQ
ZqIEF6oeLbardQrmQ++nP+KUyYstqkc1v2LwXXu9YU1VkvW/NyCWMxYX691ARh3cYFTDZIL0O42G
F7qr4wm2KxWiolnpX+UsT1rcaGW8TzIyf1+B4KbZhAluH3rFHuOCXL52SmllJvt8ew2RjfEHi84K
J/PDG7SBAg1SIl5q2WALRuJbv3S51Hj5OUxBncIUuTCg64BjAYFK8GOc4gelzYqkrmaoKKlR4/5L
4sNLlje1zxZLBbjyUAHnHERsGYe6doKR+4vKx064gSs2f3z1iXVTKNY0NKOLdQLpmNY/dPVe7cBE
Rg7K9cSXdiYWf8xW96hphAFmZNbzazVvcmkDvR8Gn5uEeOI56aIQZcfqibM8WDI6cdXuP2MR8ynf
IoWm/P1cBBbyFDlTaJloY3ANqtASPhSzTPTTvfTo/fI3yZTOPQNy7zMVb/lVpZq19088x4dUHks9
inGQyz2oyKdIEn1mI22YKpwsEmVcQkaau8T1yJodVwLZF7IM+ZZDhPiP2Kn9Do0wmKFPLHxgsfkM
eEktHmOGByk8dNawaMLKPojSpmn8pGwZ6Fp/3Pk5kdk0QdoS/rfH3valNjsG12W+6qbl+l59/Ela
p3K9GJ1AZvPfzzNlLAUR+5fTONb0Ee1BzjwgQZL+LiGQ9RDdamj+YlRJErPTO/Bh5ciaUSxee9Ga
v+gpaw6SXB1e1UY+UHQpPu61pBAf97gs7J5UCpsnHIsvgp9UeBromYHYi7blXrWYwPekXo03aJL7
YKQ++aUNHQfOFa9HmjkD41FrSWU185oDwVmr/7hPWNE+xjrPrpr/ppU8qG5GeIo8W+ma76P8mMDl
c/PTdoGPp1I4EJZBB3/JQrMD4+ZkGizu6sxjS3Vu3JH7dVV5UHAKrn2tgEJqQqHwAjCr0ku/u0WQ
kun40nmaq9Og+VjFEYcMROwjqEP9B3DRtxABA250dVQ6MK/2mkM3uXkXsb/FVXziuDcCSOlF6oiF
6xTu2/8izvt1tuUKEDff47cSgxhaZ7of6CfsnCA4hPnXkTufSj/oivuXT+jQgYRHUz5apeI6YWhy
/gfGgoosVSaRgBg0mO+m2d8edHIipGf3DJ13KHq19rrfBa6z0s+InuesddXrZ//wpemln9ZBdeSW
fXAtjHlPdmnaCszZvxZy/O3f5TecMhifTR/YTdBhUImw3myHggbTc+Q17XiEiefWMDgWZCxkBjQH
CIYYVVnqfTOVwEp+OlvL+zyTd3UFN8H9bDPXmYCwEVymO1Mro61n4Lf9QBFPyF7D0uk2rYQlSkVr
6pY6jYBLJv641KYyi4cryf3NgrCRkxS8foWfX9VVEr50PA+P/mSrP3GdFG6BVBhz0+swTHoaUziG
Pt+HGnslbm89FrHLeZKMA7VniLvDj9T3PtTKScJx3cY+AKa0Zz2NUSPnV3KQuUnlRJxR3y/V1Pzr
z63GU5oi+nKa0NkXlsFBJiOu4nO6HToqV6lB8s0X8++ccnI7BPkibCy3okmqqsNMAFmpuEQEGglP
sj1cvzO/TdCRNuVcJvaQTNXLJmFKT/cDFwlpbv86so21y7/FlMxTY91+NGfNuL9LT9vLKbWSXnAd
JDMkPRlJtO00t4b95USoiVL6ukhoqSenso5+lxNYo21de/Ws5ZRyMCXpqz76oyavo+4ai4zuYcQw
U7dZQp31X/EkY/tA1aijMHwyEIRMT38uBwqHr6ZEwAs6TAUN3lcmGS4/E+iF6YiQ1EikIWRW5xRE
pCIVJJxRzIy5F7azSuF/UcRuvag42yhg70Lwm9nRnOZ9M5yGF02jAV6jabsbyEJtH+r10paReruR
5Ph5eEOzZoBmHMYFR9Hp9aIc0Qwiaiv2xL4Q8TuWResaEIqW+yyCRBfBdcvzX/xW0cXIuQMMG7sW
UrA+g9fzVHK173d6jmLqldqUdnTnZG/UxxKCbPj5x2VUJUcXG1X4LO2l9Jmp7nTzGfk0Ir1/5SqJ
4LLNFN6XcF3p5k/7jiViWhYysy1WLgG91aaS13S5hVqOJKEk3DYDnj5czAkrCbY5qhcKixvWnH9m
QTDKUfnb0vTYBq2tsxyC8E8dgJlOW2vBYXKQ1n7H1WpSfaBAoNeNDZn/rCR9yvkgu6fvjYr3vJmv
a2Dm77kf9DM7WtVbdbYlUcYRLkEDpzY9zRZVwzwDrUm1R2/W8yOWBJp1kY/tl8UNjvbp4kik4w0U
0CTmuiNDJes1QZ+AipKMgNos8mmzj7EceQNO1dMNuaKXtV73F8JuTKGAnwg16GltWmLKodxOAKWS
aU94M9vuztrsQttlGYj9x88O6W+Jk8W+J3tY9vzHlz2WNFc4I1uHyuSfTMoudpT7A9Xy8TdwMG6c
hy+WuwxLU8IrIkyW3cY9kNx76yW4WBPpPt3MRxRE7EWl+Q9lLssJAP6k0N7NiIBhQNuX8UO0Uxis
HH8d6K3r996YIjczVcKYizJcj9Vjf2OFvYOyS3lHxlVAGgKCdJCHL9gyspIezNaQBEQEaPHEA+cW
3CgEBPUoZlg2hEMG+q/XwglzoW/nWOg6kGW7x2XclsaDKTaP89+b/FIfSD7KM0bd7pCyY7ksHcOn
oeawHY4l5l6SArsgJX0gGhagJjkYvMrWt4/YBG7getMi0AxUckk8pBdAyArbMwBk1tJ3o7YakvU7
KMk6xWr2R55+/PdWQIWVrnPXaidfBJ46Kirr7m8Atkh3Y1ujJcWxj+9tBLnlSoklausKqvA/iV90
OlsBY4S6m0ijFxMOi/Lbnf/AVmW6i9KZiQDZ2JLCW0j6O0Ah1h3yfxD+ptoE9b6F2zxEWMZ/5Xr0
X/ACrYg40KJupDmwtWo4abx/CRr6/zITuoR4eVoVy+fICO7uiJEuMsLZKUN1rRoWHsjg3MpVNBho
V3w6/07Hb/W9+seyCt5I7tfP4CpTbcUCrP8C7188wjW6tK5eo7HrnclVucrAHptOpc744UWfsSNd
UpwxHfXL+bH1IJa+IoK7Qn27oTWlRM3QxjnM/+HPb6oep8wkopk7+bozBqUIC5p4Tx91LPVpqqnN
gTCWH9d23v9TzRV0tx1qS7Vl26iSWqGl7OtCJ0V0cYFffZamYjE3vD9LJVphflXDuFI3s5GO9vAw
/2yl7t6JQwXzkD+CiNcSaJ9ZCHN8/IeN5xLwVTBAoow80OkKfnSyp6H0m2WXRTxdK+5U7MA4Wil9
1PoftftVSyJx4rqqb12z/P2E52FbYV3GFHMO6C42y1uwG0lb8Kis+3UfZPPzlauSPFVRPDTTV4yr
m2TQSajgdxufhdec2+6xBNF5HHy9ybwcvP7qlpeVY8P/fygJOeU1m2f4MXDHeoSUCcHkrUSSSolP
+hzdyaC11qgXglb2FNzZbPQCauZRxBXE1oRGjmyB8GJH+UxgBZVRap/FrN4OqMGRofamiuISCXL4
M8cS8RchXNyZLr9piBj/R6r+vCiFCA9ktisOKiD4sW/FYVBVIoWbBCSegr75sjao0TvD2vJ2pjbj
iM754Xs3FO57lmcIL1LhiD/edb7WIgkXSFWqy/rIIFbX760y4qGl5CIeX2Jd5SBmBX10ae/pVc5C
+JtPgnWYWjkWKKg3yDZN4rRpzQTRS2g2XOu0YsjoCsobBsTzUEmEkdjhsgtA/ng40FHMdgC1VYzd
z0BFgJVGxtvP4g1OdScLliY/znl/EyJvQQMHuKsO4NkhmZJWx7YaflRS0mHnd6PFyfWeIXjwGRCb
YwxKiVEENSOEEfsB3i/O/foa5K6Gi6EBMvasWHxndBBWugbhJ+2tmP84J2zwIUldJ2CyOuQHO7kZ
fpSp4LVbZuNdflEcxK/ZdEockUuBr8G+BXOwdLpS4t3pP/PVXXeyDwaZ4nYUXni4kJeSCasVWDIZ
iV4KTFXtN7KyyFuByzyoonipI1CRK8Rz64NERVJqybTV38SB72ilHh8i2G7nHUENXFXai5QwJ1UW
RUxbMisz9VdayJ2/b/bDPeUpVwSmrwUAbImUzgbTieyvGrIHUeFKDzn6rPVKNKhwxJ3SA3BhTt83
z+M5UTTRdzfqx9xymlLrlInS7CUZnZ4eApdCgGawG8WVp1zhfU/Ghgb6IRpozwFqSsiCJO+3ib5o
bI69qimlc5vIfBsJrfWTExmIpDnQcQpGjSjI0JA79w3DxH3L4ywBP2SaB3Oiuq91rTl0gyDRv2wi
cFyreKQxxqbyH1pQ+BYgtPddMhVvbOhFDugiY85k61auoNqPbRyCjwjUvXaV9oYB2G2OQ6EwKt3d
K2TDBzRCmSZ+6p+TLo1ImpL77ntRBEyzyPuyRft4/gkiupZoCYsCNZh383cf0PdyWK8QspkVPDzd
+GjWKd/nFmKXezY5sxi0SAzqLn07NgAHWM2VeYVcQVJ37Yf9c8MF93yVvRhqxpJg8QqSkhEPCN8a
0KWsuBzgcX1nGzWBkLSpqBc2iNAQz5A98rU9fm0odW0KOOvrS7pPEBGKKXRV+wLJARGV76AJJRga
7iufseIvwkcaUM6qCkmobfSp06K3TWFu0z27ahpWm9CU19kjfP3MsovRq5cvoNVkEcFksXKsynMI
iDrTclqAB4sejLaxr04+5hGC+q/jvtbw3UWtKH49PK2Rlwuab77LacN2y35giysEhbERk61iyN4o
tV5Cy9/55rI6eyMcs75uu0RQ9Ajr6Y3D6Mg1TC88az/qq43HWD2goP8nwGiU9H2B3hpP5Jj359+y
6nXvB77DMGd/mdchRNbSdKWYIFRgOSLRc+ABf73a3t+ASCUpvYixIH4Kg8eFwBVJYf2SC906n0Oa
UH+UcgA0DXV/nMSb9HpCU8wEfB5l+ju/XVyJdEyb25bR1eNn4bqebTm0DqCBAVz9zObltZWkMxFG
Hq1+1uhbhMo5LUwXoDp2ul4u+VOP3x6LBitf5Bc2YyQXOKSdjv7mUlco1TCrqoSdyQgBZ/coZs8c
LdxIOgEq4/kNnwU67fls1wPx9TStsQQETKBOhJ4S6Vc+zZgJ2o1FoFYbVGvhUoDpuGg5TIKptbFY
VDvjOkebNsxTwL1jW+J6xp20DzH6kPJvSK3RS51VTYvuG2j15zSLEnAoaZMRX1fb94IyrFI58zHy
h++YR/D7oDvUVOez1SKAEHEn4XxOjFOic/oqtXjF5YuNgqopTalqJFc1W7pBrQgPmJ6fYQ3zESud
C4YcB/vvDAt+NsjOci/4vzrnWYuWwFwzGpBFRTj9aZhnGJZXy/BK6FbDC1AJ+A4YFxmGh9lvluyo
QPcYQ+DXye/kxYeauoa6wEmn/5ont3+aGGETbv7UXEZC9Kt+CHs4vOR7EcosgZoQ8MajrzOk1iFY
NlCHJTDGddbNslRx9+IjzUM1KVMhPfg1TLBY61Q9ijcdVh5ns5i8XQWdNMmXL4jKVsxaSyJdVIrx
4QrjyfMs7m0viHIOs1xbHAljFQQmwwSnUzPlO0z32TLGicVTZmC9uCSQ7jNQXHjNIAkZasgr77n7
gwd1B0RmOEp+rCTTE80tq879V+j2lWIcQYsPewU/hy7X3XlRc0vrTaj7IxeR7gvOERwmN5odMotS
xKV+D3YSN2NCAmC0Kg7dASVQkzvB4/kvSowHdsEHdAMKVXv3Hd4jsU6ouvJi+HHIfCAv2VorCcUK
Gu+H1zYwiM/zQmf+eQmEFoswUU7gpUbMQsTrAUNNPbgYsitixemY+EFCQpUPrGcoql3Z+37wSyp9
2Sv12jeQ1+vt/P29BKXIvjdyGinlj6m+bFlEinWFvy1ILIofAiiuGbaPX5x6/Q96dcKo7KFIKcd/
fLzdFxk/tac1rawD86DiSdBLS6QMojhItOu8Agjco0+kPBUVzGo9DT8MiNxJqgkM4RsSQH+BY64r
Uwp2W8Hau2CsAz/Jyic1qS7cBlLlG07nXuI3DCRADSUdkVYR72mrwoKLc2JumAf7LZUJn0QwMPsd
853qebWu1H04cZhuBt59UsyN9EEhLGW4LPbPlNU0etU82Drmc0bFV85mprI6+/novQnRzPkbNuJJ
IeMQRZw5hZpp9l/NpeXwUZI+mmxFS18Vxklg3u8gxbYJOgGQEj08zlGuH2Z7pLqGu3aAhPIub27R
6LkZm9r8328tYYzOMNOKwcfq8kb7+fOCj3SS+aFeRsrpr53brwUj2ADREUnMm4dFkN41Fbx1PxU8
J9rc14JleYCpqKaO14gpwt77c5fLK5QwpLNHKQwVMarg3nR/B5RYvDZbqVGT4fyWk/iNKXCGlrhP
smTzstS0CoWPpr3b9vt35WtqMKZ31ueRYDqw1JYR4XkrWrF+K2FU1sPVm/wa6BNfii5WhP9a2Rua
bf91aBc4QdXcdPmUv14jhmjCIVDOJCYnZeXV/mzfEaR1PDZHzT28dH0nXlcPrj6YXSld88xdAhaj
83Pwg3iP5J6x9ZoTEGUhpmExHvecvBSgvSLGJKVqXVuSQjb7sDk8UcSP4aEFwtIzVGUzSkr8X6hn
+XVqh9uBwZTgfmCb/hTpzjCzVc9F4gLAU0TjG3J9hYdBXgyAS55DUn9OXw1+aG7ry5jXcPJWiEdB
yf7SkZ5W+w1ifCHrkC4TIxtwg//pFhJgs9gbvVX9Pbu+2m4BXz2GzOTycVQpJQHFfs8bSm18wyC3
5NRpo+hpFB5HPTa2xVz/C2av8X/bvX5CnvivtgvPNQYwR8/HEQCRTl8KvH9EYfMQe9Ye8cMNc7+5
YPU7Sqg55tSad2IWxG4/vuNzVc9v8T5qHY0uAKFhkkefh/blt0nJEhAigbzavObaCoACXmmUIvEn
WBqjLcoHqkEMgUlNNjGnlulqA0RQgXaooXsw565mdZOYLg4QjFauR6tpyJVXsbWC3ne85rmxAw/p
TmD68pDTwG++Mcn+GpocyHO6p20SQ66/qoghR1iNnCh61ZWwKqVeR1IHQB4/nyLX1Bsf8HFnarhi
ob1QtQuCjUyMQVMbiRLV6D090AgcHGXweEJOYuh2frvTBRmZXwbIY3HjCwlwCTVzHsuNZQAIOBau
A+yEY2L98LV9xonIoFXYfqGpRS3lGSKIW5II2YosAMAoeMccJa/NCI1e7e77lOiz1dvXaLPdXM3n
+7zJ/J0cJQytEA/TyUghoLtxOEMNvRwFRCghyViBPUhd9guT/bttsIaUyioDof9CrN6IRA+QUYnU
lzjAd85NoR+tRnJzpb3W20ngsqFE/6vK+RU8ILddQJEUU95odWaImdu41rT4lLm1AiXIj8Tjtfrs
VuwuoFhfyvFyml8RdDUAeGQUS2kWx4blj9tM3C4wt/73JArGr/2BAGTW4brraFdNfnbps5GGeb1q
CBR3fXCXHG4Uz22b908CsjbCDYgRpQi5V1jmC+EVQ19bWv+db6zuwC98E6EGbkCxMZ4ObAab9nqM
qwsDq8vWTPbHTcWD3ndGyLr3uOuwN2PGOBf04y75QdXxfWtcZbiQLyxeh7isyCpWuqirqZ70XvVl
dvVV8V8HkrIgx0W6x99SPah3wL605vEa0Yqe4EkGAtx99qV7ZCL3vm4nSe8dDYsXsgDHS3bND4Jq
SImwz4cmhrgCQD1IG7WfMfahfE9Aw/SemqgUZCNro6EyHICx6MpEaWqE9CsELqEVstILgphKwiFq
jq8C26mcvjOgCZUFZsLCADKTMQuWoQRJVaYTK3UU3XpHdN7JiX6N6I3zJvkdeIYX1skYEgaz3Q3t
ZDA9NwQxH+Vw/6RS1zbQgdVvAWw+qqTdQ2+9a7Ka6+iGOYNQ8v8eoR11JLaa9Cd7RH3SYLC3LMsH
q8KNAEbcenJId0UeVyH3pD/4U4cDbCPjBQ/MKbgzKd4/CSsPGJm5K7yKb5EmfIyYYKwbIp5wZF0e
lEdA3y0PTZGX4W0CCafr/psR9L/h4HpYpnhyqzSQPNuYh6lKa8Oh4zHsfTagq758VApZFg/qaXGD
SxFFA3XBzqtooUb8QYqr2IFjiaudANQMXIl0rtj1jXkl2nlwOmrJqt+iK92I26KQn4oaOZOXAH4t
VwGn+8vAikYiIS26OUXgw24JEKwFK00jQtkL5kLQs86iWPK6M9FoSPA+4pbE5P71dSwX1/d3CnPX
1FGiHBpL8m06GpemAqqTGJH++PnZph5GgG4fkgJUO2HoOpLPBWWeJ1xRJHab2PT+M18dNBfm0eew
KZz66o80jMlwXhoBz9s1kmk30pnsk5fwYMM6Snt8s6Ji76VgkLVV/ziAvU9uat/MgGJkiEV7m1iz
h6A6E2//x660FENIjVC4xb1eL4TszEjF72bhUSlLpu44/Rf2dl4S54geG9zOS+B5OeSBfYQSE2B6
bnPr3fZ4AS3dELpDnNEvqFdc16h/fU258v6LEc9py9xlOoNgMlqOEu8Wn7TMnskHNYLUMnAzTjtM
J5MBwIMK8epLuSIfUYdWCuzhs3buADu56kudqzmJvD03+ZXzhNOIWXv/awaRXsXn7OKJzowhq+ns
bJagCly0RPvvvigCgtZGoyujvdJuFqMu4lSVKgEs2Q4ccE5TbLiLOEeifo1f0DySx1H69MUb1qXp
ds3pSd32ik0xlXwFUQo6DvOnkXKAEMSomZQzf0kgQ7kyj0xciHNz7Umrmbx72v1PEfRKdJ0OCm41
sqCpxoLp2cGehzBVRlvh0TTx2Ho3OCUfCzkIzC9UZ13r/4RxmehNpsKO/7aYZ/d2RWm+NjQ8/nex
5eUBA9zRMTO1q0CEh31Zev3ktdNLfjeMWBaJDQ8mFtrQ0k2VLIDccsP3HH6w4LWzFo8187StOu2v
6FuDkiqK83g5sz2rx1wtvzQyrAugCiWgG2DRtLihs1VwrB9DRCf+dHlvqSHPjo1cCVTXx9UXQVQk
eSUyRXlUvFjyKW0nCrf+o7nj9FqCKQtQ8bCRGVAHYXOyL8mLzt9v/NXH3T4lnmVnkvG8PuvI8AE3
5dMPvQM9qXMvDNSR9Be0fxd0pCFRPe2CEeYToDa52KyBIFM1iKiUd9T9o2f1moQ3KZJgO/5DG+mh
UyiGF7kDPwKUpnEH7Z4MOTh5+nvzKvpyGzQdJ9U76rGqln1LsBmsbZIyLq0uVSJ56JkpyHgeHNIy
VldYbwHgzO+PU8YiPmLKzAKrFu0xo1Oh00SoCGl4s/ATw5PGzp5GxZe38IWTAIwPdXA23U5xco/o
hzgkteQGAvxnMd/GDYlHBKZT0L+jmAySvLXa9IE9voP05/qRzILn3sEkhiscY6AMcpxjzYSnEJ3z
MI2SyVpRXVe/uYAjOPDFOs6dFhAAWDGSdnB/R6+UiPYOYlN1j2Nt6Tldn0SAXmUM8d1pbSQxEp1S
EtYLceczxTuKEYp921J84qb2eSev04MFUw9FnOZ2rdz/WQu6GlXI+M0ODFxjdoApsfNkaGpSG5k1
r9IkeDFAc0UgwUU961i8VpOkD/M5wZMYLnqGFYvoNYm9EJkZ3wSvdb2ZTzsu86GDSxffYHUcHILx
TlLclYiFV2mWC01x4devcVpqHyluPETmZ2eEVb/BvF0WK/qf5uCuJTBW4BGr7thEgY149l1Gk56C
GB9r07YjqsEkKanvi7t9j8AQe8bFAFjJ8n/OpChdD7gbH4XskE4dyn1TJWPfR7CUQlfCJ5Ut3now
b0KczYYJ4Dq5Sr1DQPJ6jYncr0esJPurrSbOurrXdZRfKO6ukSmtTVrD3nRaZPQFIqJPwXmWqfNb
vmfPr1FeXijYwbo6onlZQdcGutpAECyNhYN2YnGdEnc62kql9efeDHTK1SMGLnn7Ucv65Tpu64sy
BJatHmtb8kdyPYxYeukem1mEQNSpRT4xqr8n8bAlf+Uv+F+nSrBLMxn0z3TPAk0vblmdOeBNwndX
C3tIezCJBTW5iVE3GXlzM3+EATyCGpeLK6U4F6SxUa+9feqn2L8WVZrELf3wYkDcfzSRqtYt5klz
g8vicg4gG/ILayRhKeyCz9CAcpmhSSPhvUDTJ1Wio6J4Wzh7NwQ+YSpC0C+dJKyjsqysmkRpVCet
4Vr4vtTeixMD89LPVcnpJTSOmPkUoRGvUWKX4KPuHtFrJr1MgvRSDLA0lLOcsdq4vT2FSgf3dKTf
4nv/iFko1aW5gR38IUsxLAsqAUGrhwx2GSZWpH481tlHnlL8y33mPjSOptUhKTnd5PwLPWMdGuas
BWFjhuSYIgOvFJTbjPSeGxkM8KXE07C1O/7E/zMcEaK4cC4GH+FRrKmBt/a9tPibAJVzfH+9FoVS
kqxkVbqvMvdufF0hq3vsxBTPV0eMfIyFotx6WNadflzFaHuYR/y6Jum/1j3BP0W84AjsEc0zLgZ6
VZxahHja3kaSIUrB5lnv+qJbC/f6K6u0IEud8eGOXwgYgdKUpDpd5Tblr1fdSWWHn4KZA8Gegk3w
Iwy1tKT6DmXwGVYTU6koZMUPHcwIcoa/OZUV1u9DDdKgv1uD2N6+YFg7z1007jcGH/dNtjuiLsEt
2zgZvYd7lnRhJB/V88ZagvaVm8fYSL/5qI9Fa2uQNzW8VOOzYsA6LhH6vW2PwvPHOvr48AIvBk16
RrxQn2l6xWOD4JkXC0utVtWC8Wekddy4Q/VFbfCYPL9dwnpqU9tpegQvV+KT3vKYrPFtin2uC7Ba
w+gDmX8yZYu7WPqNWdGd6MzCS4ZTjoSnkZbMgmkFZql2eGVGr4Pm8giIWJzFKRsky7CAyvE/kb1T
Vx4UOj5aIpxD59flNpqqfWLcDLMwiBhMEhENoNNlyWrGNeSBrED9K1TicG1WT2bP3FcKgvU3QP8A
Q8w0Qqv8sY4KqUKmIcyBIYGSvvXPVQlNOmZVqwzB+UZYTWSKMlq6Pp4j5YUU9dHrHp9jOZptAp/C
CdsJZ4nzybOiyBVPR43zLSzdPZlojwZgwsm6fX474GS2UUhZY3tWEHh4e/yFs5fmlBKQHgr2q6Re
aA9QSnEIP3krrQsvHqyv8zobXrZUeoF5A9I6Bx0NyOZXUZ5gtBox3cR7fwsT9T3IcQvWEALARkuC
iwczQxKdWARleWNlt+taD4k8bbJFwHAqlkyIaeif+jktn45mizRhT0Si0uUM11ZBHNHM1n3mGgo1
MgXaZslXzzrkhgiz5glgccQZZmsjqjA9AlbhzPG3IoBLiVTkqFSeBKnC2X3Wpzc2p3WcPBvG+coh
w7IVmmSRbU7r2Mo/ZchQ3of3hcqE7qWNwCDZtRgIDsZXU9XsSQ52RQs3zIGfHUdJZFbEiNulbi+6
q0/Tf9d51wdj9lpVXaq0eAO5JiZxL9Oo3gWaQFmHs9ZKn73GWXkH48qcQNI/Ew6Iupe6xhUVw1I1
jnSb/mDl2vrpTfhy0GGyT43mwAKkgWICUahE1pUg2zYK/piPAeVlz4hvkm9+zSFJbs/sdUlaXj9q
640xnhBqtN+FuKoqBntu0Woc2NsG8646p5LqDPZeB5E+QmId2pxmyX0OMuuuh9Xw7cvgEzTa3iMU
4jE8zgjYBt8pDEIyyVUM/wzx7zmyf17OYpVE7v7gz6qfAOh/VEFCcO0h3+A1+pcJyVx+Z5M1h+qo
5IPt6ZXQLgowDz4483lqSA0gDZ0nZNVCeEyePHoq0PUTJASuF9mM6LrAPNaPKrP7byxOuQQOFotw
IpxfZ40A/e6/AUwy7EmFyAZxwn5EDYih7L4tuIYExdUQ+FIrgku8lETKvedrv4KI24mTMPe03yNI
EuzW2l7mw863q1M82zcl7v0uIQGNpVes2UQz+NSc6e7SCfz5C/CHbLiuSA4/KmMWi+KQ3a1oBzCV
yHxS+M//5bSDuag0uuMCQbml2c7gwJWYDbkoqDu77Nd1dRDUgNIiH8UX5CD449I8GSIMrsEpZX5t
7P4x+gdVg1pPcYBBuQtrHfxODMUrQ27KXOKi8sg+IldZBdkgz21A2fzWbXeXn8oq+sySZoWjEgFT
O1RnVdAIFhfoNy/T5dBfmkAUS10BV+fHOBzkdB/vcSNlfewv+HIxweHDM+G4Y0JZ1DGceGFvqFcx
+myqEWubmo0ImZRlpqxjylTsm1CV7bHzlk+c5M5QKpM88JEl9Qp1ER90rR439okjSh4qiA3MwopG
IdWRdWaBpLihwA1BqcZ7i8DsbvFG0J/dHsHce2GRlS134twf/ElBjbQYZ24zazkyjJWY6+0LbOR7
HvfLQqRIKoxyloR36XrgCQX+Fvt1sRxTsTVD/gPXNBNUANkBzKKjoaeXjp1POiTYP946ZiKIWrrp
64/zgmlUJeeT6FKJVdqiiExIv89A1hfIQRqIru2MRwYfeXEJOJMG9YQ64XOrYZlbyQjwYKjZecIZ
+WP9RXga/zY4TjosNWezuVHMmd5q/AkYXjA4Nbac2pW/9Gp4SEUgwXYbB4oTYAKnE4kkLMLGRvz+
QgB8YjJchfbctKUlUngI3GUAKEXQYTzCosl/5JPlmWOgTMcGMMNAaOb8JhZU0AHz36xh5Nqu6GJq
+CRxVoHnKxHRZUCE3x1wZD7AF0u1X25Y7cQnNOsHyTzmK19XHCz13rn9FxfhvnfQFQCKcwMQlFQ4
ktLRT4V+8I0Lxi6Fwpj+kj3GlJVhOKcK9Nn3C9KcrkYprGHiY8pGgS8yY6MotRH1Nnkk9MOf97MM
C99p6J0r0Fv2f6aN4BFsvcladLis5Ru8r24YqTI0n1x1sAWBH4/kVGT4VCv9d+6lqsQ5WEjsWqzj
7EJQprVZA+1CU5R6BWYsxzd+rk2ZYyE/oOKgv0P9oUb6tbW4qAMZN8hbn2MKRgFApFda1Re/qnjo
WScUIC9zJ23I6+s7f114xpL2dmMPlAyetZrEm6Zx0DMZMw7HBC3Zkq9w7rSUehKoMnNeARcKKJ+y
SoN1CT2p51sVB2aRT3byMolJT2A6GO1jUJBmedMQxiIFv/2Th8IemkVgN6Mxr04Zn9WY/crjMu/k
z8tGaeoHGgR62TTFNwFLGmaVTrKwmUdTLt79hZHpOtbcrLW2qF30tbIi5zhUD7jZFEGI7IuCzRC2
9DE4pha/7UYtSQ8U51HC7D/a74s9glbb3tZWPrqu9PQ57ZWcTqHnuqwrlgmR1fXL/f6pFm334tMk
0Kyh5aJYs9hrJdG0iNbu/xNJbcomAFgmNCftBdK91KJSLeBAgdDXOQbOcq2ZuAdVeo2bnkyKZm9S
kwvX35SjwBorhAmTrci0layz10Vtf+R8zXPMvtbKoUGZoa3/fmHvEKbhYbLKH8lYLE993srd3GVM
3md420r4kUt9vNSyeBIQu9HY0g3OB5a9vO80bltL9FF2mx8htLuDy6mvIt7JUxsVVHeaCIgw8ou1
a2BM5G+hAPnmBm4y1ehbsexfE3yFmpYuEHoprBbNLKVU8YeCP56TJgsR1K4oTYaNq2tSAhvmXjaJ
d/gWNb8bhV5nEDb1Fl7LPsNvhEXSv5DUuKElpPpEEyHjbKSF5rnXYe0FrN7veW9DcH+gZYAK1Bjy
J2XQ0986yEzFveQRSXOT2FsLiqv5fopNU6I3tUjka6cgi++1y7hLJyK1YSWhzFKTFjYdXpR9SlTn
fhh3ExMLhSMn04HEsItAHYm6mSWtQeDQEMSZfaEd2955wbPnk+/H6XlHVshsVxngs8VZrqvfHrZ6
lH9cgT2C0NjdP1GFvaHMck12NwtoDzb8aP/evlmd8GGYCdoQTHglqlxMCseHYv8QFvwAU63FkzKh
2drUiKJD1uYisFnEcvR1YYPj+iBXpbquMKebdqNTNqMayZ4XyxECyKMRr5WKnJSlMm8Q5ewC5me7
PPRFVM3EMD62DDqS8uOo7XPa4Ae/hQhTEriNXitQu1TqBxWfChXX+F7idcZD8yjmnwnxxnkCRrYY
oxLWKJQXbDX6p9Qtzjbfv41UXdpDJH7dXITsPWQQ1nlg9kK2MKdUjwdK97bBbB5j/6GwlJyooiyF
IESJX9wOlSg7Sr/YqqslvVsQP35v9VAR7wxpeij2IZ2f+bMqnBNUrM/ag0ynQJHeiM9V5CoXUziF
hwUbx5xcbGkviVytd3uPmYYyM7w9MgmFwEgRn2ALdPA2ZxpcLMrsKazVDQrVSavca5Q82i/xf7FQ
S+XPWT9rkcvmxOCcfwP1iW72dMYgQsEKU/9rSrFbluMAi1zfxd/ygUxlTxNbyI0KxvgAVfxu0kqF
qpMaYCcdjWBtcaEqQld7iPJizXCUkQb+VQI8ri1Q99d/XoJnDEWagbebH6SWcDhq2AEDqPKv2idO
JsXLbcK1XyG9QGh/n06fgUgv5Cd/YUsGo6widRLvxYTvIMd+3a8CMtw7ZoujHGNPedqHH68r2+Gm
ft+2SO9064efNMqB286m6YPm1gmxWDeV/3Ux02LYkuRqIh79ksIOX2npeX9yq7BE6TDF8KMmN60P
uKxVg98441NamNDRU6yNo3zRjbvrFlx+CArOcCRNlx4Qwku2cvQ4Ty4YpPCGtRtn6l5E/STtmGnw
JBOloyRTs0j1Dyr/THEkdyoT76LfNFR/VnlTr+ySMOfPgYcnscv86gQekiJ39Jw5MywgYxVGXmx4
GwNB51N5tYLnHrAo+Sv/suKtmW7ijDe08hMMm2ik9W0cfFx6yfvC8hJpWEePgAI9OPmLhYi0bP0h
ffTFyBetSJoHjl/5kysYxBRhTDdv8gZlNcXFIrM8Ub+OfypgPg3qsKBozpZ6A9DFEbF1a9jgYaaK
H2y/YhFq6NMxVBh3bkZHAXmifvFKtfozGcNuMIms0Qa26M+Kgodm2x+HN9KWTfV8Jaz6b53Cq1K2
zP5CDBH01sRioHGfm+IP95rf7dpF/dIz/V5E/3Q91IE5x71aP6zE/R95I3nSASFzvvv/b5dWWKXg
cXtPd8dnV5QVizctN6T4e41p/PuaG4LFzlg5O34657Q+SUkXRTD0eQmV/jM45ZgY+18AEM1Zo6Yz
Ya6Yw45iBPzJlw2UUXToijEPB8YUa7SHDGIR7gCFIt4Gvz6ZjtvXowZBjM1ji//yhC8VPioIbn54
+rptR1KnysYhHvtr1Kxcm6Zrscgu+dZdR3wLO+w9r6fBNz5ufcnnpXgF1p6nMg+STJcEuUC4nIGj
HdfBmbqWwg8nh3GiIcCMclMjN6m39kOsgj+IJ0xvhZgHYoqMZHpVB543Dwh4/dGOknfwyt+FutQz
knnxLXxI5SnTpAvzXtKRddwYh8uJExQwySOJwktaE1lJx53bpGvzceWiuNtmj1H9rOcKzlMlRhCX
REbTCLnTS43xx6/JTQv81S4D7c64LakXM3uwmaKT2ty6X5/7y2F2gxayZEqBAtXAU71Bh3Cio/jr
SiURnf+xexyySRCAgPNlA53jhdYD6Rss0lJH3lbzKjy+HGWNWAQ7EQk+YIyO9iqUZ4tBjBmhmZ/T
eqEqncn3bD7Stkp7Ivum9Kaq5YCw1sceYpEfkaOcIAMP2yflyPL9/zJnXjHGD2USusWK0KWxLUVx
wHi9LzEzMJOsuRCNZBWgjjrNjufwYT8mi2Bk8DEo25HQUNGdcBPClZxrvWcXVBAXlMFSYcZ6snOd
yBsqOPz+CAcUidCedw75/YUC+E0Z9fhpbnnr/ItLGP3MmegrgAqO6/8E5hg590aiinbrXMq4IiYG
U2d2opO/KYemte2UOvUaygYoU/eC7JvD5hkyUQnAvCBkr+aDFKXiz7rOtUV3CBxt/0IODxKfsqC6
WTlwFYg0MCzkn+Wl91n9Fm4tQx4IJS3bT0sbggRJ5WNfv6cSgU+2v3IfHm+BqJ7SdychrGAtbFyt
+92EvVzGQprHzI4Mbe6erzait3dgRNyd8YIdMIEXf2BTzczGwHwknF1l7mEOv8Fwhm8xEX0L7BHl
Btb3mRv3ekeq7U/lmfXttj5wl2vYMuuiOCVjOF3aq1doTUsiOXS2gcDmRkTGy1ZFESnYQv1KAI43
xBDdOpOLw0EUuHC79ssxodgQpNsz2AfsApN2lrKZdBFU/Fx5d6fxMWmmliHEt01NciUAcFbVJT9Q
QBCp+hZwwicKCiX87wbvXt+y6TJz7a69Qi9OAnU1YwzVOJuX5WUyYOIhb719+OY4ypr20f3Gy4K1
qype80BuR0DeEuHpyWL1Sk2FIuceYbTDs/OTLIg8/TidzxM9Z8tzP4VTjQ24pIBAp7pKIupdA+RW
sSg1asBJMZe7Bpbb767gTrRC+CLSgvRUhZ3IstwXZdUrE1WU4GI9nk4oVDP8bbZuRnFNhVd+Gcbw
a6mmdJ1iBj4+pA5Zwh5VyUWCrxaGpP0U/SlMFEMyOQKeFy+L58/gKjBWJdzlgNEihqCwLC+kT9ii
p/ciBitePpWxI4R+92OeFLSOO01Jv5BXcCQ7udo3Ow22p1dtuT0ykS3NrCd/nLY5MXqvPMDbcsnF
0HIv2sOEfBzCTh6xraxSglb2Qg0vGXo5XeQt9+bIImVemBeDVgS9jUIbM95nZAulzDCEt0ttF0B9
eQwbzIPdLRLwE4+4+sYrFmpgPpMnEdHHAjCwJ52ON6ZWTneqheh+krsUcn9F+nFh/Vvf0UlT7Eua
y/b7yvb/SJHxeezEGzqc/YIhgIcL077sWB2tBpa2tWJD0Yz7qfrAE3B99gLQj46xxWegB3CkzLqk
AnGl3LMLVz2LEby8/bJa2XX1hmGH03G6ui7EIlIH4JDYUrOW5IxvXXeLnQuY4P/tLaOoXIz9bI11
fzRAe4oboQyLWieqHl4IBk/pT0p3QZ7J8RHuEiLgEztuZr4dDI5CboAHlxZ9uOoTIARGod7uALQC
M/Y13BNhgrlIBTb86mnj9W8miN7ySi8jiTDgzYc7vrhyWeACX5fPXct49GSZLn4gcZQlE97tehEN
Tcra18CfKS/PKRyRZ8J1/lrZzVZ/MpI+VFdadJu/hYtyiRxxV1GQYsM8ZOgP7vz8J6fVrTrD+Y9G
mHu0TeAyJxnkB3pHKYc+k7CFpBQ8EvqN+gcITsAaHoCjNsLdECZzs/b4u8p5HsEHVyTsj9LAuBVr
ObdilbxmlYKEWDtJTY3WAmGjtII0yABdP/ob4OIa/Z5kAEq3ND3GDhKX9fpaQlpmOPAkiu9tuEVb
ICtOJGByBbbFUdVc/xuLHdZw2UeBniotGxDiIdMkif1rLMJ/T8U3RHwlzKAFUKn/BgSFZiLGVAoT
PijRdEhoiT5A6SGjKzadokbwJL9WCTlur+9WO1xbqne2YLy3NSDRYvIzVBLjQVU01+a5/nrLDPbv
Gkf0QxezUpyzAG9/U7D3v+kO688jYMpW22q3auEyaNctcF5+W4Pt3nvejoXSJiwza2qt6wk51YxI
2vIV5xMr/3PGRXpnV59NynLKR6dEs/OkGrZ33KPYskYMYPDq9wOJCxuSCWb1fD2Q8BfeE/ilRnpc
iW3pA3W9Aj1SJibVufbzBeFz0Sk4Bxl9Ro0Zz1+r6SWHDYmyznOc5+jdw95vO+Z393KCpkDT/qfU
jRMjVUNheyTj1iYUc2/NWMt1l9mdznfOK6z3t6Emy4Dp6z5zzCVtNWT7yp3tLxGxyjqf93FZ1dS2
l2W5f5sS9jDkfYpXHu35srRPLaeM0bkQSnOnEKZaifjwnf8Sgd3RUapA7yxa/5nieKyIIJgTtkdY
3yQzWe+TllEAgQSjnv7MyIQquHvu2oZn0o4yUH3vPd0wB4U/O3N8f3CRqDHQ29vZnHpTPLE07BMN
8XJU2TQehs9+h4jqLck1acdn3aQ+3EMy2bdRvcT2xKnj1k5QYtYe3LkEnSCy227jQfLZfWG2n7k+
07n2UXLhqboQyn+k6oDojVVpu/PO6iY09ErZaT0MG2unxCP6aHmQyuvpFmjrKKXFIXREBNzxacVB
u80GfHn4qN1GJIvs/xSsXlByxfSyncv5e21Gv2P9NcMCOeiruoc8wE9GK3Rf4tFq9yRzFAaXZ7TP
9b1ZNQh+Q5QPniMRL4ylFlqrE1DuO1uNIGgIA2qBd8+Mo5K1nPSzjPGmMgX5fukkuJatvtRcYoEP
6yU7DdPzHade4q/EZa2uf3mtj+DSBRaa8/Chu8DUGT9RZizFXRwZvMGuLbLDQukWa9DXeUR/AQGN
+ME1kr//SwXfHYpH7Y9G/vt4eP20gIgvVlVL73NrG3+EXNaJ4ZFKMc/jfIB9K/zORU14EZGjQSov
1oj1kjEHtrXn7T5bB5cXM5MyGOL55roxy8m5gubCwT6M6kQ0h9nsBrDMjrD+2JCPBM42Bxn+6k/T
Eu9uoidXMeXEBrgzTHiWrcWGAQ97O03JelD3g9aMPf5s8plaYX4bunAz1P1sb0hFkB9YGB/kMS1f
9wIndKQiF2XX64I8sFA3k1sllW7lZ+BVwgB5QcbyDvxeqWaVSdMb6s8D7Io668Wbrdkpb1gq5Ugf
ER6RuGF7E/GSXGZ0x95RyRn2vh48vZTfcMb3iwcXIX4nNTPsQaK5TOu5MqXCZ+2Sen/oZ5hcprHL
7MUCpQWrVhGnLYwiqhJ2XJ2RLucPfBfdiurS8JHU2TMDn2tF9mRBq8fy3WKNu9vRd7RbSoDbGUYf
7SpQhrIIDoqsKaAXVkE05mApaTKUac9cVaHKtsXxekS47bwajsR7wRZ4JpwMtA9QlTxevdpZYPQZ
XSlAQw+r29kGFq+wuTbZ/5ZcY33hIVrpWB6d0R1gZ2d45xpVwE1ugr+RmLdNZ7HP4dhmrr8evrww
vXbv0t2DHJu0VcmdlmTJutCWuUqorVHfjTLDJmRyJrPmsMP6zGmHaoPWAT2XN/1ugi5Q85jF9R3d
/OYgVOHphm4LWbnrdpY0b0RjxS+g8yDbZUwUEg82mEAvxxUSwNlBNNYqE0X66WRKHbofo2+gdOpP
Tg28la6go9bfIhksIQTHfq/hoxPxk1e/SFbrMBZaSsTAwl+997b4MiGsciJ6YN9sn1zWI6aL26ip
RiegZxJCgBO4c8JIKdyUNWD1GcANHaluEcR/mb3jCQCI3B0zlOVRYJw0lfyWKvq8K+YaeDgzctJs
MJEW08c3mHUwH7+wdmbQOFBeSetBcWFeTJlMaZqUMuer9boVs8qnkzbm0fNDwgHY3JSJgaWGbuMu
OTaMwDO/+kEKbgjXsW0E1oL2t7di01lxHjDT5rv/y/BM3JVL4Z4AMrF8lMKAkZXWaomToGnspAKs
pkvAEo2z1suKutTc35meJY0mJNw/qd6lVnYixhfuDV4uWvodKXHpX2F2ZB2ezLlsuvx4znSSyl3C
YT2cR/Yxg41+H+h2m6GB2lz/gt3PjhgPaLv1lHCCNWnVV7Jb88uLV5f+YXNdOB05OerwLyp2XOqr
VX4eFbSOJVNtfZHvI2w2hqJKK4XZ5TtI3DMnTfDBtelAY3edoi17rCfrq7UsI5kRvNrJLn5e6+HN
ExZCT7qNQ2EXRybFwOdRzI7+cezSV7u+q3hc2M8zH72RMXDyOHrOSJboWm2veZiK3fMGLr0HXG3B
IhvhonVAL6auUPIzbKje0tFmg7QPwea0K0WrM2XKuM7e4ggaEjHzdTrkdpDvQarV6crK+3seqJET
kHI5PbcMKq7lwu7Bm7L4AWHmxj67QKzVc8I8a2UcddeRl6oLYRtvbAqKo5NGCgZ3nCC54fUy4V1M
fE3025YUiT284n/iLAFGdd0h2IN5QX3uk3kUZ5iehw9p6N5P48DfOr7Mz6mtTBIA0hRiWm98OpcD
yKDu5IeNOSQK0F+IdnPvZ63x1F543/CCPmesjLEbVOOJp4BIrIsqRrd8ncLsXu9cyzQ+n5tQ2RQY
Zy95GnfqqkPofb6dpzAE1JkolQNcmGsp5NAC1yK4kb8ru1P2kOU7YJQcxCcshZ0FyIykBC4fuzNJ
S5Ja3fcS7PJMMgvmsyWPEnipe5MpskrrPC9NjpjXIsdtUozbgTN8pasM+5u06AAruUadK5B5irYP
tgDWOxKmUnY15S23b5CkD089wBezjSAdirRpQOSe2ey4ZhEF4x9pjkJ87QmM7EVS8iQl5zWC7pkg
ffLH0ycJQRM+23u4n29vcsj+mnAwjcCCWw3Aj058JauW39DlIsq3cXpQZj9aHagv58RPOocHtu15
Yqgx8PAi8tSBRuf7Zt98Ysa2PCyrSkKZ34ovImMJxrkazpgQgEgH9n+4rj1GRN5p9q98EuHqcNt9
wg98/eOiC9j6eFgt/4Q7u0UJAHfs3/ruIyF1gNRHgjnEqJEMzPXAac6gU1tpCar0CfMWLIADwwRv
cxHjp1qFMBrs3+p5fvtNiIO/00bWJ0pR3U3ypdbJ/KcV0hYDbQCqBTVJUyMxzc6ZVwOTVmhmOGB2
P7SG2kDPuPLoD5TIc7DNJ85vj14LPW7WJk93maQ2j/cZ1z2rKqzAi0t5ohghEKsQDdgEcl2F10Uw
puoD3vlgjeMfvWuDk0s+L9d24QNelVJrKsEv8bofC1I+HmCNc/rDVYWdUAXs4E7rnyM1vis/Y6K1
ezfgOpPRJtxh7rFFUrLAdtSsWtg+/AeaHkMVWjKGUG15lII+7zL/eJ3L02u12hUQsTprjP+YU/C0
rNCF1U0YKkVRfyCIjGjevqTaPcGqb/bblZwMX68EwriOoIDPix+v5IakSi6bezRyzWADcEI6RqiA
qprI8tKfnOJE3Rr93RzvCaKgeYRpUrHCX4XQ2KEvgybU9IqlbEDpdjraO++LKt7mLQxisNR7FnYi
brB+dS2kMaSgGG8nyRZNQlSetUcTapkNtvHBNSefwSrXwLUnqK++T7zR1O6XI3vv+dF8Yy0r3gxt
EsLfitrPPhcamP+k19UjXSTUNWUYk8vK0Rgwa5PeAmv0JlMB1k74I/Mmnab1KqATubmmTqB3g3vg
iAa173dJl2nZZBqKzMWG+sq44qIuiiIIm1j9fCKIP57r5CmjdZSgHNWguJjt8fwzQjvjQyjtV5O0
o5uhJATUiQiLOzFjD1cGYT+d1uN6MzRxqPjcIebtU+E+qRa9Dak8hKsTG2tQrrYMwGjIojoCsoE1
iY0vfiBzZeL3KFRcghcIniziNOdLZmRBRYduitkTMmWJq0gr0ErnATmSQM8kZaLylaApRkThjZ5p
sZxO7YVIWTcAeXa0KC+hC9ZRN02qW65cctAKbuTdVqvYEA3veclXxwpHgq2xVSjUluEBlYvhyyxe
lQjRnWVTVFx6Wgp2e7LlBJucW/aiUMFKcLcWDqQlrSt94ik40XMHh5jL77PXTaTmseoXgaD+fHEi
XGqrUg022J/C/cF/YW3VQKnGRtR3NeNPclrYBgYUijywrknNPn+61UyYzepkKbkPSD15zvVPVSOZ
ZfohviPX879WqdRuV+Ui9HkuunUBlMWf3y+TWAs45pFcngm7a/u/FrDgTzLaBUvtV3zgYcmeFuh4
W3Ls0uQA7fZ59XqmwPowGJXwvjQlLQOHNh1Q+9jduiyZsIvTzD5Edf9IrHMtIu8NMF/1MVTH5Z6+
RoAtD6zvQ6CFlSEOZd3H3ziJFShPC8ixIbWLJF2/8ye9d5VDoXJy4B1FMuOQQD6Y1MuZTLP5JBvZ
5jYg3GIdRl7buhsHVz7YwpkGoUYSpqckpoSGzYE0DyPlK75sbFY5pv/OuP2V6dmZoe4Az4TpKydG
9cFJYyOcWAG+4cMnYoLvIJHGQVaeyjxcED2R6P4Ti65XT/bQ7D6oA8wDNamzYNfIh/K5iVyAHThq
S6SbWfY1kYaw1TpOwDaeB9PHqmkU41yGREuRWDIvQbFUNSnyriHYFA60SqGGY53HE7BD1F4wUgzc
yEWhsG2mLGgZEqX7MzSS7VGyIPPhs+yCVxNYLxZnPYQ8lprCGmTpswrAScife2J/+oEJvAvhceVk
Aep0GiVNt7dv0Slp/Q8FUadjMfn616T8iiJppnQIpIaG6ed0RRxyvMdKrw99z3ueAhpJlF1lPbqA
/V96HDlg/Rz+Nxe7dLuShjIJUWc+nJyl9D6wdHXrZoF3c0ZgUp0Kyn1Js95MgVdzOM4uAetGrPI7
CxNRlmrAUE1TGMftNs/V/Z/ooDzxsLINtKp3MRvF84JNjUz275ZKgkBEqyP474pbTjP3L/dxLwQo
Ia6yuRL8Bc0xMbqqDHJKconeqS5VSrxPlqnUBNjdQmSxGFwntdrFq3AWGLk5805XEQedsFlstpI6
G40OQ0GVDKT1Wi42WfWZ+An65yQivYbegVvmf/+hy7Cpz2v9+ow73gbO0nvGHv6fkY2/lyh3TpGm
WSe5c03xUm3noH5CvvHz0nU9vwyJVvQezz34mkmqMXvRZqCBJoiFaFOdEx8CtFS6l0KjpL1I/50J
C+cYNIzG98WviVIFz9jD0Ocy2er2kHjMUJNu8T4Fa7ETfL+ij/DRmfD/IJ3cHW6kB39RH1B6SxIy
iyIT8ZTeTW5btKr/TkhK33qmCp86ORbntKYLA8cHm/dj4JZxk1KrElDEqMv/ao4C+VW+sVnqerKa
N4Humjy2+p9zadBsy0ILQe+SU96gsIm5dAheJQNrO8YChj0UbBf6HRznXG1atmSIBN44lSwNHBOX
AThJmA7Gum09vzNaRqrstRxgsTip+EZmILxlZScpOnQbsFpZlnFanyVh0IxAyWb5HTt4ZsCR6y+4
uglYAZJmHNqa7y/uDBtEapZRiFMEBVSvNtm8XZoZDwe/jdyjMh4rgZw2N80BtaV7jEtd5JQuLAVb
0V0jzxO096UkZQC63R5nvdlIMfIAvRO/3q4T9yM8UF8fzw7aMKPUtxtu4/wgRX3wHCqF68aB+6NS
aIBmDf4TbtRqhi55YsxvCNybxqQl78IlJIqD5WAQWLJqqZnPOqrQi+UevaYsa0cCZlbGHBjzr60p
hR2DCyVSiyckELZR+obyh/i3VtKCbFeq4MdCSSNZfv+xaqlWu4M8JEZEjwLCbXs7q4+zYAdfu1Zw
Zi1STktuC3r7nA5qcViLO7J6dZYNx5j0aKLDcb/kdkus5aszUGSe8wTbxqOTNroLT4g2tHr0GuKk
yixj9mHLTWTundlSorqIv81YD9nT2ebL7EJms0vNbyEOfk3NYHT2mwK11QrM1T9wd84Yuemd9YI7
w6sZuLPOaJYZkCLxpuy04UCl1SWnP9nmPjrp9TWqZ4WANJWBu7LPhAIzks/Dl9MXEJIQDmsmMXkr
Xrxayz3AqLJmwzQ/1/wwckOuUjeQZap/gy4+NhH5QbBMfab2hw/STSt+V2SawiW5xCdPON5N72GS
8ZxUyWJ03OXdMZaMn5/Z8Zyu1rusN6MSuQMPB2WyFfGowGI5zU0D4cL1Tbp8ppmjY6TLnH4lthej
WCDZag4ZE2fhGj50kSSKid0pd9y7t0XAmQfYc+lA5ZncKPr8snf8i8TTLeQNbhG/osk1JFYHujLa
0UZpG51XzSKP0hoNZi48j5snaIKA8VACb/Y2u0J1BL2jloc3LJdkYyShMWAcM+dDdfTOGMjl5mLI
LMohrkOTqOBgAzokYqR99T4K05L+29DnO99jzYMWU0H3MhH6Z20ksLKcuttFn1bf0IV/VE3jSJoF
qCqwWF4BEPTFhejImZFbd3PYUR1cteAsawhSdwKO2k5NXPskFkUSSeSfJpXiU9njH7rRtu0w3Bb2
g+V81TuJ8kNczh6pYFukeX6q0Zu0iY6+XADS87zCwEHvbitOvzeGc3OOcpqX3qsJ9Dob60UxNtC1
svc9yJV9Qm8WXkFW+CaRo+Sbqq39Y5yp4CQZtyIV/sg4UtTINA0O2QXYyLKrOI1PT+DkqKOaJZH1
xn/KxmS5Tb9fneuAVAn4JU/gnfw4y4bDLD6YPvsQNqU+MFO3Yqfi+1JDeLZB2uhbdYLsPBGamRuQ
N98CV+dqzaFVWaOwPOP5pOu60dJnBH1x0MLjnLeCdaMqtlvrXnK4imHji8Vw6iu6XZv3/cz9lkMG
MLyfvIbAxiIBonPj4J/a2vSe4+13qok4IymEt1aLyyVfB4pYhAVpxvs6LDPWkmhRb2Mf/h2XxVeQ
WmvAEipJytq+reR73Gz55lV58FUc85PntxgxVSzCbNMXsNZ9AC1bcursWOndhhcoIdyLiH0ON9TD
LgDmvK3+VOxMhlc8Ls88wwy9ZhzdKHfNa10RiDFk3AM2tHzXZImKcPfgBMV375F4Xf+2panqnFp5
AyT1RrAGMe0wa6RrzdB1gfBPfdctS5A5lIahiG/v8h4gG70+U7xxV7xPchOPzMlI/UBMc5BRAAfb
FslCgl6AKNNgmjQ4woX2WAEHhXkbXZt01OVd4i1xobPceWDuw+dS7hvrjO3Ik1foxbx8NZLyrhRQ
jR8JckWZ6my32nv112SW4MfjqnzguwPWKfqrD5Vy4cHcwaJtimH3C774z31KjjPDhBjfVo2e4iF3
+PyJntWaIz4YSx3HK9JuVKCGoLabWteJaNM2VZ46Pn1dkCPSfj7x7e7dG2lWgoJMaxNTq/h6BZnp
ctJyo3QBTdwAXX2736pk9Ryene9NS+VxPlA0dIncwr+cxbi+XBP5aFxemSv3c90edegDocJpd3Q8
xfC/MX+2/DOJgGifIpQ2qnHtVCOlmOYUSoAqmw++Mce1zB7xisDndcV3+DeI9hA0zCnlAZvi5bzw
j4g75LWaQIuc6WsrvbM2QEDlaXtb7dvrEk1l5E8M1vRYQgtAzP9kXa0gVJpYexSANveYTczbD9E6
RLDKJm5scZd6vyoN0m4J7WJyG/pgvuRBMIVDcw31lcpwQWQs7iaDQ8uCz/SGs1f5XjZAIo7Tr/qK
8EHc7mcr8Krjx5aMQx5Njbo/K//kEWpMJpLve9H2KFg/taTC//W6ZJpteQ2LazIcHPDJCVW9wpFQ
0+Xd4z5hrfoA8SnfCakJI80B6xQsWCjIyyQDlAj8WieZhps+gzlYyMypRg+dbO+RYDGdy0WxGVNW
I3oDlmtYr+UIpIrnqybdXQhCn2hIs8lxh4nn3CJJXVib5UiReJ7DxBXQhjOrVlb4PijI1c8s/qEF
hQ1KrtTvZcs1FTrbJZnTYTG/q6MNgqIocQ0ZRvz898Ut+t5gl/8NLPZnUYs+ajcbRb3jZvSgfczp
0v3inyNdWApMJKPu4XHeqS6Kgh1tzMP+5VGB9clu6MfrblWoViD9BDY7d2GaSOQNhWP6b8CMlDZz
oSX39SvsTqE2yqnXyoeb8xag2/SSQve9ghilJFZ89OobJuDrTn6BXbx5U5TsOuyxQe66a/g5VRhB
NpaPCgaka1fH57pPWvHLN6dtQdUrEoUPP99V8vqE03erSnIW3ycJ36pN0ZXvDyx0vfZSYxge9qIy
VXQIEbNVPVwKIfXwlsy1GrpUKf7vZAfB5T6MqM+X+kOdXsbNnbKzQpyBGARoAcfW2F0YD/p+WhdT
vtmFIq4DzHSzKB9vH+lrI2BWfOfOUwXLECuq28Z2eVXBIUQYF2efQ3VtxAAeeCp2lKtlALHo2tUQ
YUGLFvSrG6OlGHGdopoBhH+S39BsQ+ExNP+dN/ITLhpHadrnepjFfV4gcrc3+gUh8Z2fpc0E7A/5
D22KP+rJMMyn97nzaBOAl5kDe8+v0YWhIp2RDrDNQpOHEC31U61gqLHRvcVBB9Wws5JEB/dsPGl1
qx7U+xBO78hRigeEqEBLWSTZJ2NtE7KNx8U9N7oF5GtUjprz7cDeY8HBFnOmhLp+bBffsK9lfWjT
q0V1i1GBG38/pX2JDB6ARwrCamcBamK0doPHGOSft8TSz1pE2oPR8nzckndOwzOul2DnuUM3atOL
mSczozozBgz5ZkqL1i0LpyTLR+s068gxoqCNTu5dKlG+qhAVR5gjH8Llv30diNkmAiLd+WZSxQe2
H8XgRkr60egv/PoEAfoNI/ryh0aphPNUYv8BYkIaL8MS2lAO4LZv1RxPLZ7mEcwsPYLRimFRES/J
Cl+sGVx3A2GQRqnxT0v5OQnC/TWKiBuyhH4cBywUwJcwIezBDkqtL6SD/3DTDQyOoZWuySiBkDWN
sJlBqjDB2tWIokiEd6AiWaluMjzwCPZ14b7JWzcxgoDXIDbKFTdF3w+eeZ3jEbytMOjOC+X+ivuQ
dBTA9NADvU43CpZt+baP3g8wzoatbQaIK/QhnKHG2jtgJ3pWPoRfbUyHlPcJc24pwHRure8G0UyK
nIcAFjntRfpV8jEcTSRhfvDqu5nUxmJTHJ5D6TQhAR8RBohDLhjgymDbze2vFBscN9fqp/KVYfne
HAnO5Yl+LIYcSLQUZvZphkhMKnmG6lYp5bVLjd3PCrffoJt+fvkN6QgjBiK7yZl/QJgv1k3yPB4r
clYoBKW/eRCmQ4PsADIiyBQBBFEU+ZPv9JpaPnDwc0HbYSqTyRouNyh91ZwueN5TzbdvGpd//Qpd
cSQ+QWJ5jEIfn/EnNB3/kJc04wO9Ulvs0m0mZnUe/qfMdk1cqsmE2i3fHrAXezaR9rj4hgy18ejC
5QIjEaU0+fWZgHfWltA4w9Uf+atZjT3bnbDunUjk9SOElZ7xOsaT3txZbbq8CpRbacXgawT/CJcg
BBAxnEawemEbLy7UFc7sBGXRH/Cww8gUry0MfdNTQIwaTy7H6DeeTrzzISpHVDU2ENnKMSlCeWX/
ug+2y7JnillcTMw3QCorADlbgtLnoto4A/l0pV1etNcFPYg8U1IIeoxEepgzHOG4xqdFh+diSLdm
Tz04ZHo5Vc5MXmpfkqxUzwBWxcp/fl2bNCoMy7nC1hxxFSWrAZjFko7ms1+Sdt2lw3BhPP62grz6
KL+Xv95XzMWaVJjG/tA7wo8VKM24jllY0CsoYZ+ekog1El0HKWbnnLiORhHzeDbXyTugzqNOZOo0
mbZlyKEvUvdLrBgQldF9nGbPAq4JuwbPVP9sqgUpq5oYpttD3wacY/p+HVPGKlnsHrqT1d3xTSJR
TcjF6n/YNZ0dORyVRM8z06o0QgcodiVuoOI7J4Rr/v8eRMj8iNoTrb54BKceXJ6l/TnfpqlwzL2/
ff3lNp/XZ/TrDR2tpnP7mjqUJ9n1NLKEAhy6ijPgmB9miDnnEW5ncEsvvxuPIVloOk0Czq6dpY+Z
eo2/L4MYwYaAb/CBZNYIGog+0cuFLasGOC//+e76fqMWdrZmrP8qBh2r3Q0DV88PMC6EYUUEGKyK
q9S2y4gUUpgg05H/Sjm201ju3PLbINi/r3mGF0LD2TqAJLu/FPGlIYs5AWfRdG9dsXppm4duOATz
vDDpJdsGwDQPDoWHY6SGbS0veZAH7+yk/CrXhapM5g4zkWL6VA9IXA5IoSkc8C1r9Q+bPJa5Em+N
1QN1sHixuUtoa7cVeXl4VzN8TKNlOo9UQPlRZUjZWSPwyAg0bA56ZYFeOfRgMFw1iZgTCbKusM8L
i6ZzbPm1bCXGO322za+CkigUxNuK62YGuqgd8iIc/2aaCW6fyx6vCWXFdGo09M+kaaTq1g1CixTE
OimQDjYZpkFdiIOr+tewsnt0wkxPM/hwTr/Uzg+OLLKbeAT2EABSk/gUYjE2mvvFDYZepLpgI7qd
/9Ae6qHytro+Wi0QnK0dQ7T3ldnrgPvYI6Vmg/6S5YB7kD+Jynbc5MDNTVZcyL3WMsRyJSXplr51
MBeo4xl416D3Qvx5Ezl8HP0ezxUN0fe4FBBXzbIPXjPHST7RsG+limy7jifg1PuEEtc+dqk5jJaT
5nNSF+CoKiAtEpnJjZXOAcSKGNzy8rLCYhmtWAU11KxW2i3ySHQtF0okLbjuOw31hfIFpCfQxjTx
G/BvQd8tqDWyw5/B4tB9BGjesTE1PqqpBARrOP21XpT9RRAqjGXGt85TUGhCl2RgwmOSic6B5F37
V4Kl0+AD0sMtZutDFMxaFIR2yWc+n9DW2cAnPY9FkfUjljaABxt5UaC71YwX3jt7TOJrFK+Y2CK7
LjFaD1nAullY65OYWAtLHVh/Sgz6hkTcLrgkABk91ZmMyxK+EbQGyUeQYyhiEu+zw5POEVSVYytZ
KggGERIK98CMCJgObfRY1m74mva0c7dZwlj6YWewJoI3OmDeRtLncis+LlMHHsCcBuHBANjpydKz
rQXSRQP3N064rwy580z0oWAkV/2xqLIYcmybi1LyPU6P2bzEJCzpK+8TNRMWk3Sre+XF3U0l5Y9a
f1QoOY1kPOEDhkfxuxEaBx/6cAXMD17Sy6WYbVVyMn0bOaxJk9T+sJwVB6Z8lRWmFql48UjEL3qv
Bqofmx5/SJXpv/ua6/KOU9UWqLGpS9BwHIsvWrXC3IrC5NP1RbUuwplBkcO0jrDM2dfEhjyod93r
DFtHryrFf2XjZhm0DCFhsdxB6DkAtcMRBW6mtU0GqtMvq0LxL7HZF/mJFxJ+kh3iHEZvExBdTN9Y
1XndIgMj/k2AqpqqMjycbl0V1XqGTFfi1+cflkv/vF0y8hs5UtZAuaz+NfjUaWPT/lggPNE6EX5D
UWTvRAYy1aCW9pCSNR8FR61aDcjpfRb/aMUs2Az/ODXUjb3+rdYEUC4+XtX21x9+kj+dh3gnXI6k
NbDAlT4bHvy/Tlb7mssm/gl54qS1d8oXHOEDZfRrjVf9bSGAQUH5MHeFVINQ0/2jKz/Xwi374aoq
KtM07l2xuHS9t14pplRBwT8341bWBmuneGOkgBH14RAOMS1JA6fea6ib/vGURKpPkXvjb5SeN3Mz
XJjWmz6EFjn6z9VXRveM1DxOI8dmDwnFfmVzeV6Uqnl4dGkG7y8G3+vpzypcrqo6TsfB6RSJXRWm
+I8ONVYIKV2bpi9uhaoXah4Rx7SjicMPq762YVuEKJJAhQt6zQyfxiNTVb4BQkyXLmoqTH2RaLGk
O1rOq+gAblEcI+BvPfqiAP1uj0leRN7G+uSvDIjIBMfYQSF2s444/D3MWEav4jChaIyMx/AWXZrZ
Wzop+xrRUQV0w2HPm8uqGiI2A/2Kw1l7S9L0i7I/1KTiI4QA4ftsoKk40TNwVUUdIKKjkHvagnb+
2E5juJ/rS1Bk5Nk9dg3xmA7U6Z2MUyBELyaijv7qRW3pnBWq6p2qeHHLP1Zme0/qyQc7ksRvBfQS
T7NISCE1XGttYoMr9zo+zCRSK/vaJ0sLBzKQDemiFCsAfD2152cCfKRKeSkCDWjfCO+rHK8pWcNi
hfUEwWrd6BmIVTN1U0x9lkUZJEExdiyZpqHZWz8XlStMEkZjOEr1UUZRR3SgmkGovTGOFMm5/OsX
qC+Eju6HnlAEL1pAsezWZsdn7TbQow95vZc+yz/uFqeNp8SQ96OJTtRwm/fShPUFxNaHntKWtuaz
x+dcAuwRTQfdFUX4h8zWa6LdTCtcPz0cOpOVrJQCisk4p7nLImkDxw2Mk40r0Si/T46Y7Vu3Rm2Z
mjoDDaF2ku7YNpPE4r3EB5LBEYx5hfEUXWxXlI2xZlbimwIRD34Rq0Ut6MLH5a27ViG9+ItIrGF0
dzpGooaY3Tp1irmE1neV4dYlMzKEC/oWFelN4HCecGXSA4WHgYQEbwtx/vn5bjBT41Tla/pfVnH2
yRGTfazs5Z2Eqd7pmhRuCJvVALc+0sd51Jq1YZieVgg2GKtrW92XNc6JfBVYGpPZpujwwgYoRrBT
dAcrX7GA4jL0qbXy0ruiIE1tJVI/ihpMm/9wK57wmTUWn5BXaEvEDyXpaxeNXQuqsd5WupmKgAmK
BmGgEpY0pBr14+FrypSWaZmBkvEp7OVVZip3ioUuhh8iESPxihxkDwFJZWYHAKo2bSCZIvkJlnS5
JxWfHf0T2LvKjCjWJrkwi6YMqxYIECl0T/9obGJiL/T5oSXqHADd/w0l0uw51rq2T5n2vidcM3fp
CI+PRag5pX4gdEu2Jz5OHJwhXUvXY4Pnuj97dfDw61IplFbt3ykfQEy9IXrLiSnWftGDYfnPUO9M
uhSoVPPywmFAvyeHjNwsdIkU2qx5Mwf3rH2jnBymvaCD/nfAzMYn6pHgzCTJDcfMMkSUt4TQ6RQc
BmuCoZL5ADHgosSHvF1U/8ywCyAETOpThcs8Q1f7GMGA0S53nEefSKcpWnmXsjhnzYfLG9bxImPp
zqstOAYJDZRvBeZ/j6Zf1hCXUfc2VNQ6FXB2rAwC24eL51hLEwLHpc6jrfUdATd8up4+uEKCCsYP
uT5E3z7i9SZsFpR1Oe5beEuHFD5Oq+FDhtSlYTruyaeEdLBNR/nPjKgJxa1ov8iCvpsgumQ1ixVH
7lUeyKW31Usiw8btJ5sAUFqZcTU8Jfk3CgbaaiuyhSgRvi8seQF7cAJVozkwzP7Ue6GtW22dqtzD
d/CJ17GtcW+vV5Xyd0eYNejW2FrLN/k9Zz4aYRH0pJhtzlbYEl3LbdL6Gm9/DM+iT8QMSyIjCpp4
C9faogKGOk0w9oSZFwerl3WQZ1V3GR6Z8FTgxS8kFHXb2quq1PoSNLT5c7KSGuaHiDLJfBAIKyQu
PabmLx2eCF99pq/hqAwG0CqS+AkQGx1mYpTlNxej51qw2/VmCbit7NqWy8uKzDCs82O6v5htGXdD
TlijvvU7XXVO7vtyGZStsOr17UcprXSCtNpQl1uAWnr1YGRve6dYkp3MJe0gNBbxgjNwedUmYCoq
gqc38kzu9wblTUGK/D8yNyXzJYwm1gS8fk302AzsE5FGUPbUce5KuVJAMOWsWtrQEJB7Anxsdq0z
a5IClTl1lfWXupsCpQWlA8bx0eMdUG6G2GB49BIcX2ESYJcTXapPXP977OcG89lwnh0wM2hXNtrG
ACeRJyOLc23izvCzi1+LIOo7esIkVh2cHO8qxibgduYhxzQrT0lGn/L921bC1nTXPIIAIbYzR/D5
p8WgG5mn9K95QDtj99QN/2cx6YEJw6JEXOm0D8lcCSF2PkdhHifHLnrXexUa/4OStf6ydw++jlMa
zz/X3lQ8PUv+PDSGiVhBdigByqDX2ZA5uURSeIV6g1m6pteIag9AgW435lkjdn0u2t+VSdBqbqS9
asXk6lIH6L1p9WCuIPS3WGgER0koVmKhEBYU2LfK+4jt9OVTMJP1dvZ6CJZEsmpNVCaloP7A/9ta
3HE8VbHUWikwGctGK4X4zEdMvFVtTm5tgHZCiqn/+0jreg3OiIapzVscxhf4N5ziSO12xOigQ0Pv
PdB53HjDIyDbFx++UopppgiLCaBke89FMPqzIheUm9M2toNCX2ZDfhIfiPcz2Vb1fbEQSuLFK/PA
in9hdB3REaSUqq0DlQtOo1Dkiw4CHg2Fxg23xpAwJzdsHMCSXAH8nEbdt3UrtKo2+v2NuwcDoUyS
T7BB3kz5XOLsOx0vWZJwblTpvs18aRFPs1gPAdULhYiNsgwAeEkLhAWtAb2h9JL2PQ0XJlWRqQXE
4dkPEXWDx26g4aut8IcBzM2RQANRe8n1mOW1fsiPqIYGp+/Mm9DaFLO1RPcjWJNiN+uT0bJ5Vbj/
UW/9Etd168Ap7W/WRRZadklxrMWQyvZKvtzA1BvvnThStcTuACrWP21qXHUfVvjVyE9TfzYWo/YZ
xOrVuTmdi0JR4G2IYcdoZm02tr26/1tLSkUKYrT2WYxVzI1Kd/j9CzgV/47Axh0v1ljcS3/RAiBH
vbB1FfxvzUYXEkib1Lnmczn4ZtQsCOtXsy5OnnsfMJO5kzJgmQoBuhXizR2gdW6nUr74FJppw2ZC
2H0B3lfZRX+ZGMcij83N+DWGTTOQhOaqwGJCF3U9PUidStSc9RxozkWK/avN6QydAlor48dSv352
rS6jp3e8l5wwjsgOVq8crTWiNcUoG5EfqjbkXdtFJUcuOwwHJOvR+Nwiphwohe9CMpw6a1JeXurH
l1mraPluVCOFBqxJecBX5fR83cZI1wmqnobQrfo+9OEKXxSEK8t040oP5vv3w0gDEtxm2hHtY/+x
z9AOKID65dKrBiPAvT4jvwSylO3fbNpYlDxrbaSL6PDUOA1xwCumdt+0VMDhU91HL2B841VTGcGZ
JOIu6kgMOx3VlsP8uTWCilgJaDzePy2uZRaHY3rY3rhDyexcCAci6OtEhtMbjkp39Rvq5PkftZK9
tAwWxYHBqtIrbMD7Ir5Kk1hhviAmpHZqWWJ8BnsMb8hbXsw/69PSxexg2qxwD0qi9y73NpAwtD0K
nPTBSZM/IQlO7MPL4nO1dYTWHINFpf+z3/nftE5xvKhSPgbe07fn/rN1948srmLYj+1u0ljw9BmV
fPg/Kg43VfHzPnv9ksP9P0UjidD856D48s1qNnEyLoxYlGQb8GuH0anZN36ZaSBTBL3ZRcXp99Um
akE2PdeaUkfdnuRtJgjdq1Fg1pbnwuGh6MtQhUuB8/UkvlzXDJbcBuWjtVQLWlbzpTnFU7z+xrKp
v9f927EDNQH66s+2cTi4TuUcfukIRB7HJJkYhQgLgja3SzeZbEzEcf0osrhi52brhyJzUDDStzPi
a5OVXnRAtV8j/eq6wt60W3D/ih7r2sXiOHJRY675rOHqEMYrRKy4BFfuUOMxK2oozCf67wZgytRd
o8gN/xSpTupyv8W1C0J+4yqiSL/1X3zwsv28m3u+O/c15XkmkG1cB9yPWa9pV+MwqVmHG2UCn1in
EIk0kZjfgDQj+U1knS8Lmx/HqgJFOHQwBgWhOZ+1F1EvUHQfZZmLp4q76gWsWgR/NweiAWdQVbFC
Mn4ibgPyKr/Yl8KOlOSALF98r+1WohI0rNrlu3zrZbi7Ns2H1pczWGFhRRVCZpU1Ena1ieZRpdI7
V6jwSrTjvpdYG1FtrSK067s9S1FSDa0n6BNxEwrVk1uUNiMZucw6/+0IDu8xPZluRGzbyY+SaVQH
UVdUp2Af8Rf8u9e4/Qx/aRxdmI4WGuxlZ7Jsnu/+JIXKTdc2O9j1EZLGDVJV9Dt5vT3YXdRf/+sD
9RcELU4eW32gk/y9K3TGU2y+nKZRfjuYFEvd3Sd5osi4yeqkq4CF0JMKFviX0SX4Qz7Wt3yyLkGu
i02WynHIJcDJ90/LtUKqgcZTTdjPqAuErpbdsjqAnu951hznzoug4loLMaSWO7BFr/mloKbHVbGG
HRxOgYL7Ec7MkQ2C+n3Rt8B9dqhbOHbkdCdy9hpzXemZ6HERqnWGvlF2YvyZK/YKko2mFuls6yjW
ZlaLQJ5WKDavCd/xg5Q4I4SKfBV/djJwrar2G2lP+ykGBx9t4QpZp7DaBqpBhlmXSLnAufNQRhkO
GX40kbKOlJuE6WcmtQ6gOCEhgI8qYYh7qpgeb46creUZktSNPEqNUqgenekOYtPWJxn15bRrKd5E
mkAZtDKCw2xmAtNVDJwPV+FZrKKDXP0m4IzLzvGmaF3Wu0vlcw2FMSRP5sMXPUNY8YmgfMcCce3V
xf1e1o6deFYZfu0/wIwhNHzkDRAc3m+q3zAKpLhkQMShWyn9sxGhdJA6X+UIMEbGNTEw0ZrktmI8
YXNtTCzqUiEmI1vdNdHmdH4n9BhXWiMzC+CUnD1flB41qbJrpcbaEpyPhL5DlNz1h7Uir6rhpRKh
h9OCoi9l71rlf6A6yyH4VoHJzlb3nGQVhQzpVimfvElsu/ItNXrUXRI2SzAR9J/psQDancN8LX4Y
24EQdLa7vK48MwVvHiU/OQEDGp3QrhmaXoC3bsMzkvIRucPurGbc8LNwTaAkyCJ+0img3UJveKrO
o+n+HaSj0hJW5X24hE0Lp60gv+R7fTOvq6dyDx5FaE9D5wvDolOVYASLFgRf3sWY+tIcFldnDHWZ
Vvimpwy5kRk7MBdjHT3LMg7GOqsJrnXzjDPRFafGvQyyaND1cEjj94gv4nre1ilerRchZN0fB+Ap
9/GoZFBlmHuEA93gx4O4DhlvGXYxnEe+S+T8reBZm8qVAw2caLg2oJBpGZ9/ca5vctvFDd0awTMZ
iFoWnXABs0Rs+5xCqaIEsOUj0npvIuDqcHeZ+tbvUGtI9mBvC2alzPmOFI8XX73R5RTNdeV/nrOx
FSY5vhYTj8y6LGk2Hyw7o9tcUi9LMQt6Ae6JmGYJmHkGJ3TX/NRbjqmqQ38zUZSQp7bOpgzPE1QQ
X+f7+ut9ZIomyhNkpfeD5+fjFY0uJmf+nVdnr4s97VXksWexFra7Z38SUIY+9ITCzLmFFeLQ4HD7
jpEyfZregn2yaieHPQ7pJ9CXxWrXzourjBZCWyEXsokL7iBzCEc9XFRR8O/+9xFsDZ94GYXmVEQ7
pVhGjX6WoeEdaOBqbIysRbcaYBIXhzn3DWcG0iN9m2uhb5Y9Qvj06geFnCZhrUxhM1AaI95qmIDs
0/g6dGWszqumG9fAx2pXli3jUg3N0TLSTdkIzQJJIdPYfxzHpj9t492bX53DWc3h8FXaRZGG5gpl
MYnUtG+4xmq6iN3iubIHpZA4ehopiPYj05uVVFYNiAz/v6uYKemvvjPLdE3gS+XsBCcs1t59/cm+
tmeo14XAmP1ebJbkXnLIwgXDhHheR69dp0LNyu9ku1Z7wiaAKM7qOwxxT+WT/wc5kcJ+Xd2GcfJ0
1/qKAoSxikG92ZLZu4UUSF3MI0NvyEPptCa9W0Wlh6R0a6QReT/ILpBtX1vc5N9Hq8iyd8Dv3S14
NcHnNg6OlIs+crNqAaFfmJr7uX23TO4Pl3AZOCvaNqlBPpl3YhEuJ/8/Pf5nqjOuvuVvUgUFICxE
Q9R/SDreF/3GQY6xUPODPDBIL/SxArKQeS0L4/LatAuhRUhHkw50TiEE7peYXxDUwsKQydZ9i2bn
A9cCPzLkkqmHNKwZ+8+bfVCLDV6nPWuyYL1IUkARCWJSQ0XduofdvBB9EJ0K5RCcFp9VK1/ll8ja
LA/UubZOp7s4bjucPkuTXKklMh2yU7dtJpn+3ouCWq3BVSbwIT75X8Mjs7uV1zGMwTXQoqr20muF
feuSSPPaLbU6ew3+I2dTum2kJRrG5DR7ROAAWxG9s1e935WwFHylxqBgj5BpOee6139L9rbsLz6+
dSGMG460KvN44bylaXCrcQ8d4buPz45iOLZd7Z8qIF8oPB+tith4MsX1mQCDBZjYLscBCNW18PKp
k0wQUIFjducBejhV1cXkPMdQtbAilAMkz77WDuvq2UnTncPD6r5CiMFFyaJnENpP4rbATeX3evLO
70BnceagxFJK4z8x8q2MWfGiN3syWBF8jLVFejK/Xc7/sNb34NqGzxeKHmC2fjsaMQVylKD6ysTU
DP9qKCxNR5wLmmEPRvz+CBwENULZBV/klp6I13P3yJNc6btc0UmgA5CgCMo2qVQwDi/zJ/Xsgg8L
qo4UoLcWKkv78mi/K+t46mfFUE4m0MFBYM7J1WCdMIs2pRC2dZIRkNt08dIvaFWxm/wLKALwhsIz
bHyX8+keHTAymIbm+lfJCVYScNIev+wEfpalKuM63szPDgZSyJj3Kw3hU0YDQw7BDCqh796wZdWr
+tfKlYbfl3OX6Vhy1IkKys2JVhXr3oFB9ecnM8d81ucXCChaycqZdV0m1/56HWWCRzZdTRYHOnIV
QnrIltqjv1cQ1eGp3eUfG/QqZQCsCB0/BQ/c70p/6X9rNWu4/bYa+d01yTOd1RGBbGcXkJYoVkk8
PX/+7Fp3kuWTdbPttAbme3Ssxzu0kB9lFnqDOxe5BmWArxamZ1JetMFSacbttick0j0Y2Ef38jPq
9+u47pSdRNndvkplEWfrDe5cNXWuF4TIAcxVKOExFU7aU++LBwyLooz0p+KG5VRrFY+m4y/7ZQ+b
bLKya5GzjFXO+TqGJn/ZckrQBv7qos5hsOBFib5nOKAqlJxlgjVGJ5wHi9Xg//v81TEnsIoXHhu0
us8YCLAeoQBDty3OaIJVxro/GbvFYhDdmgvZFTI3XwHY//EyzklWb0gEscyUZyICx7RdaeoH0diU
FLkjYZj3BmGG0tPKxmm068/mMnuMswP5qHiaJds8cyysZs8nC97PCfPLYcAv8lvYupfUOKmI412m
dLsQCD+CXz3Aqbg1KWWnTQ2m0Yflco24VYpr5t88J7Vyr7AGVv8HqAA0EThCw9dLsKc0UlIdD+cb
e+vKkQLVlDq2EMuuhY1fpwE8LETBgVzjhyuISPwayUFv9l73H120iF75mgm03XrOwXtIc54JuiYG
M3/wp2zt2JzfgopsEOEckMl0ICCiU9hyoZTRcMfQqhWCX5UUYM/pA3C2xd5yks/HM3ucGDWr+QAF
ROY75bn4XLKIwbSyHo4juJ8idWyp5M0DAB80Zhv/8k+PA1yNhUTvAvtDhI/sCwtN9mz+JRf7Qab6
sTS3kpZBf5kPsUj0ee5uYNA80a9dFzcT2u7GQYhtSc5Zo7aQTQji7n9BeX3R24pajhzLfd3b+wov
46BZ45UOUIf11XGHrGNl0snK7K9z9fFdY5U9izoIc8akaSTUUCGLhLcPbRZf90IfV6jp/6b60RoB
4TsVpus/tSoM13rG/9pgO6BAitHzEo6JedWWvhzQWzjwPy/MO5f87nkGxg5q8n+x+Ajjf2UBzo9s
lwUGF9eY4KHmPKzcVzpNay8UxZVa90j8BxUUsblOfY+B9Ty73ruyfXrjUdlHK0kFcAzLo7fMQ6EV
/FxgWlHrSB/vNOtaIBE0+5o703OfeBDDqXGzbninM86M3BnssYoOnlqpfxIVNMN8g5NhQaM9AoZ4
vjEYgY2lyoKrbT9SVw+30/5cr0SBdwsy4j2agCjrgZAOEwws9mP4lyLibdowFH4dKWGzlu1vrQdo
0RUx2LXGCEw4R8ZeGzmkqO5Hzr+F+mpbgqgnq1hsC8HmX/EW+rcZqs4ReEJAxjWpLkzIdN+yOuwu
o3nDnGW9PA9pIGV3/0HN9QnxvtocEx++y2YHzt50A4968avKFWC6iuq1ZD9Nd8RpLsLjkLyPlXej
Gb7Ve7IAhgR8gDTIAzTBVhU5DPMTsTQUjic2WXX9/6GsTE4QfuLUtRvg3zysqDjdee88bDxwBFpD
AMdlTz1nG0V0Kw+UzTUlXCtQFQ2l/48K38k2W8llikQt+i0AmnSo9Eu/DyR3mdqkOZlxqQpnLevx
enVvmvqj3IN8BPI3IJJ4JUzyEE4chlboE1chbY2TB8MahLc3RccNIQVStB/q6dnQ2Fit2+j9wciG
boEi2R9SVrmf8OE52lyWvEvjpuCnykZg8ICnOIFAfkSAKP+ZF7IfI6/xJ2NCOowR6cv/WqP0BLkg
lX5heBsZ7MSvLsSSqRXiYvR1vakEM/U2GyiSFrvL12FL5VQr0YZfgyFHhWJyowZTzpKNcuTR0nEX
7N4yLQju3uvHWFdE5ANLzz+IxP/j0rRdGnYq2saEDdn/nJzLZmuYpR86gYK5a7S+R3UqoPmv5mK6
nOyE1woYk+a95pauBYr8BSVljpQSPPWl+UaUk47GbNSnkKcYL6ea6mcNbpHFPzLQMTA73PQujp8a
qN9XACph1zWhDIq9sjMsH4VSt2sm0V5JqseqkPoTLXb2r6LIpLEewn5lYS9jTS94rYv+J/sOIxZ6
8mZjjRaNb1DoSqENIHV0iPXCQ4kfahkfOozI+1rHRoLU7VY+pjjTyZvbrKJ/6WYHiCAgILF7yECL
Z+pt09qNbwuh1expM7skPM9o3YEA5BXc5G5va/CWobWEAbpbSjFDfTkGJ6/rB+n5oYytPL4BhYvV
umBFDQUT5zpypYkVr5dI7XItgQJNRFVOgqLEud75KhBrbvX6Mdh/+DKjCP3S0cp/TFc/DepzTUhf
F/VECghYr6kQBmopYAxVTrP/FMuCYqqVrrTBD+PZrSoTl6fQ9OfWnvhap3a2kCV4yC9b9IxKJIwg
WuVtjupm5VLWTZ9NhLqVx1K+eITyyeF8YixGtANG2/AvXz3VAUembF9qoArAqlEmRGvXK6ctlCq5
UQdVUo84OLyCrD4Qc+JzO+KO6tWXVq0oaUTueOXo6uEx4FA1oDkZUShTwd+UbX56Rct3XFJ99+Xn
qGxRErXYYrNxddeKCMDp4rlq0Xe4Fzg+/Hk0HbKyZXCFUne1ZHg2IbW7wa4LDn7cjbJc+F2chcWH
w4KYRgbZiDGj4UaZOZ/hyveat969sqj2gA8tXrafXsFLyNRBNpmcQzGxwpYduKeu+G4Kz7S3jWvf
7WIb3k1bQGSWv90xJMeyN02oGjed0S7KcIbFW3FJnIY3vkYRg9JKdgdTJk3CdK8LqEKw1o29yMo/
OBrUHTh85LFZo8CcuNZn0RdczYKyjIUYPThH4bZRf4ALjnZbZfCaz5SYrZTdu07856Cl59O0qTih
7dlIQIdaBMObzATNay64KAioFUqxLgkOnfWHEAWLB8qNZ4zp+cW69A6zBrPtUwEy97FETnWOS0nJ
CHbrE4rAlKUrp2aAtFmWCiQ4EF270ziRqv0eRb5flzHJAp4eBoiImkeMezOVzpoquE0deaYGm6U9
UO0MiipbdtAKjc4zl9m2JbgDQsNRUHsT4p25iGHxvmUnhb0WLBKVE/ugdQaeJqNLQO/uPJMBQ4DX
mDveiEeJl9uUVQPSl+Qd9ZLBZELdPbw65Xx5oztGyPWJKWupSoZsgsOmkoW4X2lhnctxF13BIu4m
51Rczd6VG+vAO8uJARs8IKcn6ixYsJyIxlpXBR5l23my/dFdNbtWebd1rwRvlja8MW6EsBYw2I17
cbF3QDOO1FLimg+p7xECpigl8Q/178sz7vXrSUn6mkzXO4bDUb8MyZ7E4NsnOaAd2/bAqJqEgZ9t
RFhDBmvLSaCnCrP7va77EKJ5g7LY71DbCSTjQi/bSFYL9SZfMR8XiAKdo459ZlndnxEoMnfgaAVA
sao0BJB/j6RmqvtjUZZPFHu9a40+dsgSXQnq96vBDi4HDJ+EDEyJM1A+DhjegzgN0bHgqejpW4cu
np0zTmeVj+5/9pq30BPekLFhh+ZaRr1gkQ8bg6hUGFLzkhxcK6KWgBmgOvFmAP1wDQAyYQC1ZS28
X7o4/n43V2WMrxhMlzOQQ6kLjQ+YYCaL9Gk3X2z+ko/FER3dkaN2YiUCCDFiO52THMmV5//p4HPw
WwqGQ20mZ/s/+ZcCg1RWgJd/Wan8ofEWfOLn5gsv4rDR8gKN9sS792V/j/oEc6kgQaXH2CsaA6gA
cjAQlIGzzi3ffmHWfzWtYaaWTEaWf5+Awi6756LRIhw5A7bXANffHnj3pfCfrTyIc3voGKcPdbIx
gke3V/OFnb25QAs0sSoFwU/971s1sCgWaQuDcNiUVFimnFwJQM4/YuG24Qtaj/yi/05ovy+Y+V+C
nHYgF6Be4g3mXWtoOqM/D5+AtwHvmzHh2ILd6opSsYNe89mQq0YyouYeYOMWeWAHK41iH0DEqADu
RVC9uplZ9ML7GUwe2Ir08uEPfomZlF00itk3D0bEhluOEoREeXZaGfAvQkq7o/h+AMi3D8JxIKEz
pCzYsCNIIL8Af1LGDQYFV2zDE8hDaIf/GZ5UG8sd82azJUxbai7V2wZCT8cwHzaNDrlzLh8E+u5c
LelWELxZ2IEmD+68dTU04mOcJtTl37qksx+j8TqbZTO9jzZ2kUN/u84+r3624lNb08ZDF89UV7/o
D1/lo0VAH/9Ft79JITiNBzyLSazYb/J2xsN/gQRFu5VNkfny6KN5DsXjt2hllcODAbAU1DGnz3R3
3QXAfrToN60o46jqhkOU38bVnqKIGvRzZZ1FOJ7M5GgRLMEBsMXOBVHiuU2HIuePnXYLrwXS1w7+
P7y4v74Gm1U84ZPJ/vtTrouIlTHfFJcS5mXiT9YRwGp9qcQaRv74/72Cidtzll47GGxDb0JgwPGF
MyalIH3ReDt3rG+gst6duLPNCldsC+MUACiwTim6I2pUqEn1IgxXEHqR1vPYKcU8hoAdLJp5Yam5
k15I1np2If0xAF5r4eNvbfLPVFobwUOoswi8kNACPbKDVJh+8eQ6NtAFUK/9vW8d8tdM7mcf71k9
94x0I/IkgN2LHiVEG7OMJxdp0vpiI64ssiuhToVbNMkXc/IM8HeNPIB07hzmDL/9GFUwiq5tyltO
6tAHgWbefbdNeSYf5VAnckyDTV8/EA+Q/wYuMn/sOpmk8tINtGpYWDhQ9XL5Ja3In98mbyXWOiHg
0sQ8H4bNraOsHMGjB/cRufM2/SkBfBL06Y/0YEfvjADZTgiE6cMipO4zr7VL74YSoGbyIxgvwGVI
Q42tOVkx4Bsd885IYZ7f7fmWKsbSFbkSDj4j78++IAdUy09l/0DM0oHA3SwflzmeaEnL9hh/tgs4
pkyMs1RrH/NOMjOsBepMEFwqstRjFdjcX1n3g3hr6PF1wDwMalCjZpqFdY+2I0IwfY2OtgYhIn1u
Wnx8tFglEfmLjp3XO4mOf4zY3BtOF4WMAB1JBS/GN6MVQ4NEq+L9Ht2VNh4wVpp/ILuucqTCPUZZ
ZdIDhlYyv9eCgTknW9ztgZmX2XEVsIAlD5stWMo8e90L7nJ2n/flOap2PhMNfcAuef6msl82gA3i
WtlG7Kr0HiMITI2TXMHZZZhRWkEqd1B0HMdLLuWOzxio7N8iDZE8u83kJ1c/ndynHt5X7N6AFqtF
6ZbTIU6GqMTHl4BhPTYD6k8uR9CZYOm2cnkaCtdea+q+6LyOyurNU18Iy6H72tGR87195HdXA+yv
pRZEaZ9XZBA5NXHxefBARsWz7P0StPZbI1u9acynMx5x2MyTABfFut18UdI/vTbtU++qxaqmGHUU
CmXPMVJCpjgAwYk6Zq2QOa/WZNT4htueCgk5jB9ulWMYcUbDx3wsy60/R64NIgSci2UILghdWQy1
c0+KboxzExy4RjppnedRONnC78+BmOa2dgQAc501L291UMUPdpiuUnuG22QKJYsYDVaRHBihD1A8
nGvzQeElexGn/kqTxfx5ADbsj93JePylcMPb4B/XcvS6VpZAPs0zHcvD4oN9Qta8QueDc6MZ+BUK
rnUplCEbjEqBszIr7fAUw1ICKHMEX7tJ56CUsT+LzGL4Pq8nbP9PPYSciIO6wdKCUD4ufHKWaUGF
nAxO2fKV+SFqayjzFPSmrUERxJwF1UjpoFMHI4uy/R2XMzv2DbyHPAQRw6SR11IFumAozw+rrO9I
E9QXNo5segdiIMf+zaDO1x0suqaE2U4jawjueD5nHhRmQ2D77fKfY6/8rA4zZzoBxUq10LRM9rJI
zRX1GCAZVEBGZMqutob1TmOtJn4wjdnDZ/oCnupW267kvpreiS7AN2l/4aU9HlASZOywFmancxef
/D+AL32QHSx1YEsVZS3yBrLz3k3aWlHhhcIJmjYbXpFgqo//LYAJet/5dAkRhgpvqYXPSzciR0rh
mL/u2NRGCRt8P1KCbf5Iovzmqn2TRHZF6VjF+1or3XVUqS2NMsod5z2AXJ/139ceGxkr7vlcdiHO
3L/8TJBL1k9P4T48U+rne3hvfXkkKanfHhviqDCiikaouEMdHtG/g0xFyE85+qgZgI9enrW7TGXN
9BOqmC6a3sRUVpCmVUKgu8lKK0C7Df7nMpxA66HJlYJRp9TNQhoI9/HZeqmqizEgbOL6XGq7YlTt
ytz5frAZUVY8ezXM5Wb3rKzWpJPPq5zaEi2D6TqF2e5PUEDmlmduIUosRWqjG2UomGSwNHoEhxlP
Z2pV9ZU5Ktnb2819v+3BNaCSSvmQUacv7z5h1KGM1gPGF6eRBdfl1NtcxFe2zTf09bSVgZ3FRtre
hnTB2u77tXaOW+P6LZAxY0l9CdrzFDcU8iXJk6aDPTfxhXey7W7DnTYQPqAPF0qtb5lsN/HFW9SK
7wV2POnoVYlMJRCWIjzm37RQGSfFLVEWZXtHwRaOJ6S7lblWxK7N8ePs4q7gljFU1eQBi3kSD/ez
Dy0F6hWojPYZJSwhTodcrj0Z2ooT4nBus8dwMcWfXjrX4D+Z1K1bhaHjBGGypzltfo8ZT9cnKcU6
Q/gsY1eIQaJElZLO/hMCEkrNqaLAwnngIycILxm29oMrT/EXgOeolbkk423HyDN+2pZwi2BnLuUg
K2tiBZx3DcOD/TUebVnaiX+ghSlxF03P5PqlQQDqLRGOy4/UDzjxKF2QWQUM9MS0Cp3iOPcMunRy
VqWR/gaPJVnJgguYoSnXXChe92IncYARQGyivEs/x20NjISc7BhwgIvFcFq+ZQSxasCElNtB4eCW
F/Ph15pRHXEkv7FAaa3l74lVyrrBKjE8/+3zYNqY9VLpe7n6Dgvyv9b7XczJ9R8wrb8yfeOfas7G
6yhMzxphWYTsOqcDhho7o9hKvVOsyDnpyX9VFQtiicmXHTLg+oJOEfLZyKDPPJ7aXHRuKQ51xqqc
YeAWS4kVr0TNJCclpumLeStfDrH8RABjFf9oX5Vvli0skzBLbDppu/UsO9lDzSjtNtAhGZkWxfoQ
VKufSBYQhOT/ZCUVcwLDiQaL95vvTdKaMvL4JRDBBdQbDo+m3TuIKDVwX9Sai1Qj+pIIcJW/+6vi
2ep9dyl2k2IaPvvH8qywHCQC0ldDTyKXTi+j8GumpQRbJpd3UGVVkItK6pKZfRhvA3s0wJHkkbqa
i613Yic4kNyD3k+hPRUr+Tkgu+2STzceBodItMp6Rg2wFTOKUpWv2y3Sh86MnXEp912Y8cmPnK6V
Hn+W5B8W2CU1Ft1MreCw7dX+Gi6QUHQ+mqC1b6jbi3yTAWF5uOLFpui6c5Bks8uHK4Xe8a0vSO/S
1/XGX6xeRz3UIu4gLGE/zjIs9GuU5t36jvNII1tjAKjZwAie34BIkPfi3tmh0SA4ReVTFwY6Ddgf
nos9ngV5r8qdLQcbw5U5vBYuJ8vIVAKsSqeUfcjE1bimhPdstzx4mCivQxs1Hd+sYPy8UhKYxHQF
UnpCF2HzIxndVgT8HHD5R/yZIhtrCp3Zwo8a9MrmomcgbFEruaafHsb7VMP/frqJzbGSwd99ZHKW
lslitC6Bl69Gx3ixVpqVAo/hZP092BiCjaSuDTQj1AsmnJcF+fj552PPnBuU9wqO88Vmsz+3fKPt
T5f5Rr/2EYOi8254dQuyj0qI2jiZOAjIblZWc5csFvye22L23yUxfSBpL48MsAIYzsobNupltjSQ
VyK9TgUlvH1cbcH7BEe36Ja8Ia3KFMU61hKaDk67I0ruqt5HYL0wEHtfCteXUA1+TYlG2MLdhmhl
TKUY067pHOCk63BSYtRXaCDqXJldx9nyOk5AHrTM5nter/eiEQb11OnMx2XA7O4eMZ3sd5ulIYNm
SaepKK0l4/qEPuQsxD++7ghOOSwHYtxOwCM+/AvgVxI5HVGtBfz8z+SvVfarnMl1kDj3c6in6WJo
7eK57HStpa5r+EKUnTPibRYjyk2m7H9CUim+ExcEMRhYAQH7DZG4GWhrjEguXv0cOVetIC0qcagq
8qNaioL8iFRHCQCqjRDZmWqJo38RkkXpxOe3g8O8LbTDZRgYNIj/hPhIOFzuPLMrkt0am/Qq+f1Q
/s2PTqFh3FgA4gqA7dHtjmTW6caRrfeM0XcsXsf2xCoRo/patJlTXaQzyFVSWubgcqzWjpXCpwHR
Ruv1X1UxxpUYHUMCXRY9oe62sO2+WZjfjf0mbBUucRIs/8YwsuAPlM7kcCQWvkCEGQdU+SWL6BfW
QfhVzjN8CXjJGUm8w+hZaH+tS4ePsSKOz1Gljc65QiqRDoLoR+0d6Tp5DxUoPs8Yr8xAmwq68MnR
9/sESzIOWBB01avbNtCCKmgcSbqcbxdppRL/ym/VfXpr6dkySmAHsGMOXfgn58S9IWGYYvUd0XRt
UvS39qVXI3OzFgy9UUQGiYVewHI3qZmFynVX1gIOrMUfxwAd+b373IkPG+x1QvdIsuIM/dnIoP5X
CYHBrr1vmKUDeDVsrd/1OZBatEX0iw5cQKmqPjouiypKvyuRNzbEJ6QR8rgPDiuiQHJDoiVNDSfc
/wCRgz1QR9dCI/MsAvqgRDy3IJxqXuj+oOU0idDEvSmPLKzZ18KF+bnTa0QcwQ7mpUJyuE84PQig
EMty+DQ1PynN7SbqHtt5xz3g7a/VjGTRIjFB1KovPcMPDFURIsABPqpT3CrVc4xg2bbAl7O5+61P
uElfQdr4bd2OhmKTL+qOUAX3Z95E8P9A8iy88Tl59xiF0N4Lc1n4+n/NQl5/LnDzjMG4FXMVC7zm
b9bmWE9YAXZEuOQpCqrXkNpfJd0kLgAchbtkFw9pcYrwZyzhDeETvWL+JefhpOvgwK4++o8y+7zO
E/W+4lhW/rDuRcIf1CGXyJC/X3/G0Z/16ajgOgURIzEKAZlCgT/zYL3Br349saKWwPfacugt049Y
Km48f4HLqaIvInfZCTMbtUX6Hx06U3ap/qhfh1Ez8c8fIIV/2N7EP5jEQaLyEkLUjBJOIH+6R4+0
ViCg97doVK7HC1HcDF6orm/6/hVv4G1sGC64Qwm3idhId4kShgTIZpXZ4J7iyJrenVUfv9PVjVTT
mNCKOQk44DB3PGwJNLwynQ4Tf/DRSASlEveo8zCRLoYWjemqRjI87SSNuZrSAz3l2G6eIEtSKVX8
ABOxqS5/LHfTgPf9lKcRPiqpXB0kvI5M19tmoaglNcMos7KOMY/wxvEGP24BXlhmIPsEWowrmo3s
9M8rcX51QFnujN4Almj2Cyp56djGLgG0jiConpC0Z4XZZbz3dwNR11SEnPlZYNMJxuGmJJ0yt8f/
zbzanm/FhQAr9bvRe8TvezW3ettqkSVjfxsto1Rm4XW2bRNFBThJa0x5/wfLzJSueql2retYnzzC
0/PQpotyJwtJIn7k889aWdRVIUgrHOyiU7OOXi4bTQzldeXetmMwhX6koytTRloOGPt1sMPviWFP
0wTEqmuBtR+QRPyEPexiJ7+/GQyyQyr1At28LyUqYKXgbjE2SdJdlVEhrd9TXOaIvvfEKkkEW1VJ
HSTYqyplN/GAAUrPSv86lMGnEwP9WA1w+Yz1WWYpb3DGup4gRSpULFmCfhIp2Ut0pSG03yKUA9A2
gCHV0UEjZlfF/lz5fHGOMZa+tXZU6+DdkEEpnL13Ua0etYdv2HuZ1njH44GiwdNsZUJ4y5A49YZz
ETkuTqB80wLXiHhGRm6pTqLkaZ3WWps4IkjJP5WPCM8MhHcQuo8ztq8rtB5PLfDHliMNg14RR3mj
GGHV4QJTcrTJxIlU78pgecyxUtOq6lZA6YDz3PP44+0zc9coYyJzQacVKoRVZjtAUHVjkK9jOYyt
BfjCK6wl6CovocbqF/TKGNRbvMHC38EmQJpLyyz6vztKKmzXZKd+6V1wh8s61/A7zAaJSrBNASMf
F2UmKwZUlYKevuSUwJaAOJA1RGMLcOymMOacBIaknoveEisUVYXlft7Ej53Lnvb0/nlODxihmAuk
5pr71koYqEIF94c2WyBOFXZN5U/gxJ68m2b1tWrG/mLrDSFl2IBC4dI1Tr15fi40xSgzSixPeBnt
16j2S5/UPgptboGwwnRmSXQmowon9F6QLH8gD5bwXdu8/vExpfAtLqlm+7S7APf37utELPvNjgLA
2QFJ0X+94v0gMBfMilzGVnPGcbSp4XmhrBlQ8csfoVzs+pDFmNrNSvTTNPC5t7WYx4vpNX9/AxxT
t2+57+pOlTH2WcIu90P5V23mwcDNd6OKwoxGvtiVxaNWW7WN892iH3QYPfIkPK8lyDAH69Jfp4eJ
X3PmHYBZkm9YbZDLs1eZuTIBoN3YqWpPz2GxR5Ry1VAIbcFTNAcdCE+Qccwnan/Xl/k9ImRGJryo
ucy7q5iIpG0cK++glMtscTMca3U+wtn4wfyUCBjtSdg8YP4S/4HPvY9bzYdodh8AbVeTcJD0IjSE
sK0lv4WYy/MItg0l2zNT2BF9PGenlDlkVZYsSdbq/z45J6YXohwLF3saM2iaOG9cJHajTWim5Mzl
+Tf43k+L47TFNGfj8o+kpg0I/gyQKRZzPYkYJYwHHHD3sd4n51UE6zWpW3eMHFiwpfieXp3bXcWk
blXa/htg2OsLS4w/j/rvVAQ+nsp7hqm/AJ+hxHQ/a/28ua5v+2rrXUBJpHygnr7hk3YdU77xSsL6
dtW25rX/QZVr01Z5vFRf5Y6v8/425eB7gTQUnCcMzlH4e/2dfTOjS18m3xYM6cJkgu0+vvHzokiN
iI72VbZbdGvQiggzJlV/dEjHp7zzVXwQPsU3wjS0QId/8j6X6/4zwnCPTXEL96u1lWIRp5KXlkLb
9KsZTeSSTTNAf62K1ZqE9OxYQLV8+JD6DtojHSXmS+ZRe3WxuBg/9tZQ0JdZp0hUtzHQFsTyJg3V
iqv52ejwEGm2tsyC3pmMiQfCoMe3hBzVmP/GJ1Q2FA/KuF60DMwbet9FE4TVVUiiXTepn+dvyfv3
Gh1BwOdX8uwOwrd/ATaW6Cn9lI0V6m4pdzPcr/VO95ghXnAVi1c7O844NvH5b32IIEwJp0fWHVy6
TrUe7WXi4DaKSE3BXV0kNZiArhTznY2jgnUKSWHKRl5SVqUqK+qIPPoopte33+AapgM5SKYsBaO9
Vgs9jLPM8uMo0KgPScEhpTTbiZ1moWkv4gwiz/5xImUTCnhk8TxOwb8xHsJOYZHWWZNq3k848axw
pzpIg6ASKnvXzjPZXhMIE7+EV73BIjaqVO0nR/O87Vct8+iWsJCk6p1Y1ffUILomS/OsnpaQ6pf+
ryA/k2N5Bx13fbD2kDe5SsFhHJiJ0bFza98N8iV2FRzxGeW4ioMWHDeA78h5D7aOg6/nJ8+W0a3I
mtjs4+QicNT/NjmAEgMbqI6tDyTUuNWDQEFDjWNUAvD/5XlgEYULKcn+P72pPbb5fvZxLz8Vukji
Eo6HyPQxFl27p+UUieOuA6UGDYdAAQk2ten4DpYkoT306z8aayaSsTz+UVyGBU6vXFs1OASz1g2Z
Cgvjiqa01n2UPpuiG8mIJod2CExBCLZwFe+GVCdMacZup00a/yoWDk85/L0kNWwrIhyuIh+vpzeq
u82FZ+Q6YYG+jkPBk0ZLAcf52EOe8DwMPwxpomLhvBTQKbuuelBqUlYv4J52E6Dy4Z3goy0PGOgt
JCxNmNyQO4MKlYD9rkSEEx/h6I9tB/u6rnyyLuAtavLVeXVBsSfWcYN31Yits3tz5nJetMlACMmE
iKzkeVUri6ZzXISqw+K6b6o2tUcHDCovOQNXUtitbWdOHsfAtEHyOfY73jkxwePXfHCeDHmVP3r3
xaVJ0BRueY/cr7KqMUHZal69OuD6vjS37bbYLO+1j+H4LqE/rT/wV1VLgijWXwk1+KHcC8nnnmk+
BEt9AU/K9Ifn5S+pqsS3AKu3F6SiJJK8K4xqginaMc2jc1JxtwQUYRVKE6cFijGRZcW51kVss0IF
mLVzbh5x+FPMUHtElt6mb46slv8XHUAojht9L3vhdASOJqexqPmK5uk6HT3SBOU2Cw/gOyoVRtWk
cgTGGERgtfHgdDDXE9R5kTUN9GjYjU7HnB+EzZYxYltYQcO5sR6jgtpGHEEdg6vpdaw44lCSASBk
JfTTtZvms/KbIBkNua3j7DZO4xw7ht1aSCfWPQL0z7Q/6OJ2wAh2KuUZFs+LAX7joSTzUFo2+a0Q
p4YrmV40T9NC6oZg2fiqjQBAMqk2+bwpmPGnzGQspsOZ/vpJ7RmlKU7/8FQQ3bR6VmgaPwHiEihj
i0vLVvkvFBVgZcnhEhEMAsI0WjU7kgXaFAa/72DqNkugiiOJRLq0jx7ys1+IDa0az7QELeH2DzRO
yzYjqLEFHhftjsLP4VC8zStQg1NkfEtD1QPNGHXicAxYUUl6YbDr3MabeVyMORYlsXjKsM8fPztU
roordAoXIRszaE6/wMjizSQSIW6+alTWsjhxHn6EXl+LmkfIWhL6H5za7hD+tknbo5P59+JqEFN2
6FmAoQElkv4dBO8MrEaQY5QWx4PIsvk+2PiEC9/U0jv7eaQfbqb6H779g7dlx7rHZjoD8d2alhKa
LwG7T4DMdzJjcG3qCV5amXfEZBYzmoxq8Neyd9eDjGd+CA+blHTKHk8WtRSfeor2eAFHju6aCE1K
c6w3EmtrYXtXgrCAqJJePO1XhkjcARWz0Oc3RILQdzImxIvDSqL6IXAj+CK2TG74Fgl3kkUgNr9s
GMrbjLPEG2kgnEoSBlaJ8rO+pCQzWdemdr/e4o80Rdjoac6u4ulDLbV07/S4ac/ppkDv7TWg3Z7L
h4FEaDnjsJk1FEbun7C70eT0aIve7ko2CaLhxJkXetRtrnNsK88k8F/qhTQ+Wh/es/ZbaySOQE3b
Z83l0P+aLEIKMzjKF8WoYa3atlOd9H3fvmYBPesCmcXnm+nnCiZclKjjbHY7LvYNfDeNDpcxlbWt
KOZdjjlahm1wtLxboOKQxBk/SOhQL5aXFanKPDro9VHELqm+rMnUrF9OmO1PgJzaq+104fTNkbXV
gtO1bf7A9fsAxEWAPg6l3pXYIBEDc/T9qA3zHVD3AoUIgKO4t/5S9aO853bf0cCtoRXSEQ3QiiV3
Mf/JTF6wvGmruTAXRjjoq+sTyyUGr2ier7d7kOZNg1i78bvkaFapYCR/SoshEI8fSt8TYkCjHUsW
85LTTueZGK6B+Fs0AjhRtGSDGjy/RrG2APgSAqzXVwgwaKo5klZOfkGHfjGlZK+77Fv1R7eT58TM
g/LqNF2U7JukLDx54ajfmWDwIn/5pG90Z7R40nBv7schB7WrcRYlybrCtAAJKm0btwp4WKkLYznT
OP+85pbecsKrBbjyyjVtlPB8zRCg5rG/XYMNCLa4X2iBNSSy22dW/bv7UN3PhAVju1cLGGWeIHIn
u3NO3NXRU981+PvK2gGy22Oq7fRpjRhUmChXtriieTjsbXicEa5CFIZXgrvFq+v2uKyh/LE7HpGX
9cTnlGYKko/K79KfW2eYuKlF3ysSeNlEbsfnpRPar5+fKzf9KUlzGs+tn/0GQ71SQl3EcQwo30R/
D0ZHDIy0oxjjU82lqPoTIHz88OCXjbJzGmEp7zfVSzqr+4wyDe3r6uRL98leqVppbyTphhhVIa6D
dLqPrsQ5cEILQnB0Q4fFZCuu0BdflO/PO2uWQNSIeeoxsCHfs3MSmA3KtoP7eAmz66H4wpFPZQ/0
97YQXbClrdWNVpCOSjBiGk9JlvGWgxf8a5Bq8EX9q8s8EKjlLNHQJsoDtQyLNAXypAL08Pgg5b2m
nbn/gzz2eGFVc86ODUFy+aDweOR3Lxp/Sy4r8mQmFKkGPDGwyBIjhVykFqV8R9ySkWhhD8xPToGt
enLWAJv/85u6fJGWSsjNH4kp0iJp8FxJuFB7mC6Ape38Q+g3OIV7/pV4vsD294IUbmpaORi8VqJV
aK7ahk98OoDj+2IrXSw2+46gwqJimxziPrlKo6IZr8bm3GevN04dSM4r7EXPRRqiYO8uiSZLNgm8
k4FWrO6lJ4zdGV+KaejDexyoNyuRyXsLlKWaCJMlkrDP/WAONsH8Dmsr1W4BRdUySVa9W/hwQpJf
xnTwfL/qe/tf5DlGmvBwgVh97XT23fNeq9vtFoCPMzWO+wIgq4/sAQadUso5fK8qcOrzHCkTtaDI
Poc9SM/5l2LwET3kOqALBysm0F+ZU+V58dUsiEya8oKBSsKJYdTjIHtSXlHWOGUT30G31cfI8lHW
8bkYZ05dZ/gTAjfiJ0QkN/AxZn7FLlqv1c075rcvWDQM9HcWW6fxL87oHaFRL7SLgQqPNSIbJ6f2
LzdrDNKYvfeEoHEDeepT/IgJ92i3ZDDFELFOLssTH0NvW8vY4O0o3ahVTzFxIQP/58rif1laeAi4
LDfiXf0be5ctWoLWKFsF8BFWfw98hF3J3W9G+MIyUrq1zUD1f2fFinj4ez9EuMQHmj3acauG0HOh
xv4hZDbHYq4H/eb0G9HAj9XW9jjj+3yv5TkTBb6RPzpQyhvOqusdxON4LouPy4bzmVKg633raiKe
gorU86gUu/9Ub3gZ0KvPB9/aU+nksQv+/uBFlGt8gsj2BItsnhHTNJhNLAlYb1mVUr5I6GRP9jv2
1mivzmHFolL7C8V2FrAKbb2PuGuGo/J9BrNEhnsRTxsXIgWXVw1p5tajHDAEsYnUoaD+9mcaRDQt
UGDBhIKuZcrgk3XQpcyyTKK79P6X0M2iFSXXnntDRyHCqJvYDsD06BuWXh9/GYifqj3Awh9EZDZI
6VZlGi20AkWd7Cl6agMOcx18FefQyuTqvJBy6gWfaHPlySZLyQ9iObujuMmikE+BuhMlHqWXf2T3
Rku0GwKII2SNOYtehiK3k7UhnA7wMTgorQYUG8E+boOaBJqDVDYsvKNbjzrQ6MkPXsy1WwW5mwLS
+lQfBqj9lB6VHtocBU8Nazm+r9Dip4S3XcxHWCIp8rlIBTafcx0dU4jR4DtuGEQIsukZKlONFpzo
084gT9Rvi3xBhOuUMKr1TjvqkDzwOA8qhpnHTTbBehRD98IXImbTeVN9CA0cec94lbL7WkzVYGCj
D6t9txMebkLbPCbu/dYADOBrgpXH9V93kesvFUVuYKMBNN5vcPQK6plGZEgLX7CNrZmc1Aldkfu8
o5ZHgk6WM9B8pbcfaVEDVml/PLJwF1YXeds06HYWfHsHjk3WmzY1m5nSWI4Ewz9KugT1alYIuLC8
w7vT6GuCCSlTBDQm5GchtvegrXbZvcoo4HzQ4axSKcNWG6r1ifLSdyWDqAK7sHmOlp+l40HdNQ5d
m0r34eKi+v0GruqNXkuqtgZRJhNReVosNji3Zj1BZZGUeBiBQYb9DlOvhFohXKA2QO29/z/aPj7q
JJwKBuLAqoRbRE/edj/sffiNKVxNq0Ul2HZ/U9zVfZ0hKDctHbFUAjprwwAAzVyz/Nn6AI/vscp4
z6v3dQgiiMZazXz97Zt6xYbgrZTr0Y/J5E1jwWTbBcyZ31XF+Mx0HhURaO4PtoWr3L0vtVJf4Jo8
ENeEFS8pV6dV7CuEjjZ6stqr9YxCmhWt5zeoyvqXKPpJ50EGfM0USeP+tMNPLuTxkGITZx4bTH4j
fCKN+V+8GX8LeHYqZHpWmYAGkj/KvtO3TQgtE+gHC1fIRxHxDEi0aet55H5hukW/jDlVK8JcjC+w
jsFFcKc9nxWVRabtflTeLh2U2fX+4EG8DYdUs2RDNig2R2pNQJjeYql0mZQJqoEakM8Owf+rI5Wv
vdPUJNE7by8eZqe9OwwBhEIr0gPMmCBHs5z/rf40OhDg4X5a7R0J9FYJd3iGntUVjEtokwn4YtbS
YlBGWSe/tEk/D9v+Q2l84DP3bC6nvNRK8XhRDv6mHc2093UeaigItjl4b0rG+d1NdZcLPjClDAuC
XLe6qdlr94KBwJgSb4ZoaePDO7yHxYHYsYkT781gzc96E40EL81SvMpULkj/Lg/u1tJhXMejyJtl
/UX5s+HCC8wj5lcQv9SrP8+yNfx6Xzx/zHUz8NmSMadwzyCSVqHZ+i7qWn2Hid02Z1njTW5SuVvc
EFWJMRBOrRH0rGQm1WuxrWqqrG55ijB+WOt+Ws+NHZ97esXYm+Ddp97x7qPbtL2RZMNKvmapECWB
p7DTcCc0dDAr3ULSe8g/QYulq1KQ0tnAeIJJ1Kdpj2PMTi7aDeR/ez4kCMbKc750mmCp9pTz50Jm
smr5ZB+7Fk0DAqiMYhhVa2eIw0P2wDcGF5NnfMYB3C/NEk0ZHreuzZD7oQDdzDaMaw29wuXw2LOU
vSz5tPlhhQ2dr1lnIPQ16uqQrGY5HRCIkOlhKtFOq3UNrgyKDogZXqA6a1d9DPupHAg8LKgOgjE6
1FiknlxqXQq1786wse4Uc4ZdC6HjefvwyViIX51rRHVfYzJT7iFkDnUFdhYIRr1kmlMECAMAgCD8
jt12t09AJoC70o5KQtfzJ9ptI3YzBdda3RAjc1gfr9SK2y/vkUaoxtxHIE3DK+CqhEwk3a1gVaCD
tQTBRpQQurroE46SWjhaJJcOusETuJQZroT7pkFLV6vEPqv9ogSOCF9FC0j+HZyfmUbgB91yaLj4
cWt4M8IJcp6jrH8neu2Ahu6uuEFhUFLy9d2e5I/Lhf8nZ8KmHjf4/DUDVqUcvxfvX1crys993QPV
AKBE1cAO9SZpGB8BLMgnW73aOFRcCt9xnEuCjAnKM6Gb6ZWSZall4HDjvjq9pH/5CqT0sELaL7Og
14DmbDcBgsq/SaPZwV6s9ic5NqZ9lXzBWY/I5DCiJ4VN+tImY4xjVnx/ApWdnPb6PuxnSUx/hAIO
B4VryPRvXDivz5wy/KpyVW3/4MFdsWtIjC6jZ4z6mjV+kOCweFp8H/KTciZFf0CR65YAp0OQmEGm
moTjJdg/LaiW8A64P9wz0hMkNiSryMjhCHbyU4NqYjsuw3pr8CSdU9ufy0UeAzlROqU471GJar8t
fRvWEbWpF7HBo3iFNcPEIJqn2IgTYWQCYsDJ6g5mCg14VMCMduwB7ZUAYNaUHYGi7bOjMtdp32iD
A3O/1SMkbewhyE8ofiw/w+/MmvBJo/5jY2EWACLmBT2qK9Hmu7hDbw9Xo0QLKDNH7oo+zaP6WUSR
9JQTJ+d7e0FX8LDXPyTJuSEJMkJ0ZQeXL0b3hpHI9Oc6aR6o1yXT80yvOyxY6pcUyyMvjtDUgWxV
lMnJNHoH9Lk7AF0495A/xMmL908TKPospdW8+u036dnZvM/eWA1SoDPBQ6gXQ/JeCj2d+VOe8m9J
kcJk6+Sj+yug6UiYo7cnFCz3sApKUo95OZb5svcYmGT5QqnGR1eYSjduVIdTuPqUp4H2zUGp+B9k
sMrkuvF8lkY39YeAaYBM8zxSV/5iRKdAd8140hgBYQ0y9cwdZzZDf+Q3KAn8iZw/R3A8dXnbNOmt
vgkD4MbTunmNiTG42ti62bP+ZpsImXQ4zZJjeacrj4dn9pXtPskyDm+7FqY59IIZu+t2xRmzD/Pn
rzCh2XyB5GOaJxl+0EWjcDOpv8T67eFZSg9FtVNFl9ujJ22wSPAWDYIkwsx1wheVsDWbJFcuysjc
IyaoVEEMXTXKoxgGs1ZHyxMZjmls+6zdjnzelGg67CVdtPYKikDOCzFWMDZ85ddOSEYmBy1CiCY5
fhfQgbD1cumfCUBF16H9Das7D69MvZnnfAGSCrSpdG2W3gz2P4dJv4KdlkzGElcnbEMicVZ5WiNs
Tq+uwECfPakt2fdhzp0mbHX8YylbaaDnVoYuAGVpsz+DomwYSrijpuhyTs0sb2EkNFas9bqPYCbx
cyznerhpGB8hsL00KaSEoGiRybnE/fewcmkRx5nt/0pVvkKcycFx0DcVkIw8lmcadgddiHwutYEi
DhUT6znYoCzqyG9c7S309MGYn4tWZqZnCl5Kh25METf+2giKRgPRJWWJHhDZeFHVV1cBnCE6PS2P
US2Xd4dWQk7j/KwCL5Lv80WU6lYwrMyk4gsoxyLECM1tzvYStWmiiYBrfNeHbpd4fEYjaziP2e52
S+tNXl7VrEG0IA/Yc3cId5r5pJ8LQ3yIEWRsFmXtKG0UpWpxnaN9StKh63ky+Xp/1HutLmVmMxDp
2d2ilke4JbihPPKm8mRg8Jvkz3YIOHyvVmf1DPMQPiNBOhassHAoQVBENTYzMnxPWt17CJFibwzM
GbLSMYnKTnu8TchkT9XNGFQUp1NfkC+G9VhaeK4QXhZx0oUqRxmZ6JYBzKlAUtVsP/Vqo7CKwmjW
jPTZfxaC1ZHh64RkVzVU4/UYa0pt8tXlRrh1OfOybBP0Lr/w6QKlPOn69/WiZt24pC3quSPWYefv
SHPXpSQ6wOZJz4OkqMYFz96EuRnQed+f+ywbvkAQn+Uio4F99+PY9XXtpeKjPMrDWvtr0ZwQfyZy
QwS+fVbaEo6pmF07HCeXb7MWAgubhjvQiV68S7hxlYFTyV87kW6ZDwy1ssiNx5Ooq0dgK5vzX2mX
agDaIz9nPfingsZnSLTKNB2b4b52ydG77+2nesHzPdus9NSH2R8e8dBuj/CkTPJbI02zkW5YFSwg
3qZAeSHt8auE7XOvdQYpIbKj/JR04YoH9b3bUy05EFIB1u9nuX8qTwZoyxKVlG68xdBq247SSdEg
MOhYnjiCo/d5hd05stZDpn2SNqHui9BaBBFxTdYWofNbott60t0ZZ7po3EEck/LBvSrVqbaTXtuc
KwS11xeCx7vtgSz74u0DfSMLsJADCDeO9o3csLFNB/9VlJqEri1gpLEav3Hk421274P5mqsjNcfY
fHVT2SZLdb/JTUmbGHvWXZaqgVjPiW4eK9N2+53GkuDqsrQPvpXLAfRGMZo4WXz5mK0hz4QHzsX7
WdZW/cMLv92DcSxYDsZomtqW957Dh+9YDibCzuw6aiJFg9PlP4cqjnJuc+5EsfADifeXGtF3tk0X
C121RDh36OARJgF1EsYcLn1vjBEGU3iOiCl3l0cw9gbJ/h6NMEPjsNXDsyxsuhT+xv5KkGHzOGHQ
madsZrQGCXxPuH48JhTDhSkHcxJoW9j7opPBYCampHgd/puwPUXADXfKZNd+Mx/iZjjVZgT7KJPU
baJ/1nvvsY2wHkSSqfYqBYKmTp0fdXQBsdtxNoAi049dSZGW8h8B85OPegNiDltgXz+qoCQ71a5R
oocm5lsSrCWn40kjkrkVL2qgyOR13L+RJ5iWvZcD2sY8O8CRiPYYdotN5OqeS70Tbcj+uL/jbbow
6IeVR7ah29PyqOOolcbW5Z9ioX/k3HXEnU3/DysrVPB57wmDVt/6iX/hCH+v2mL7KMGgTYhfgXwl
tQ/Po4m7NNRRk6PiVxrqcEYOAYwR+cM2t42cj0Pfx4rFrL8u5cS34//di/XAQsK+7E5//5iH0Vkt
hJYpbWawSRrv1MoCRB86VZCpaRKJYgXix2jDqKkbq59tUSKBmCEpgiSeaVlzEAY0R5LKbrGz1wzU
hmf/tUCU2kCKOG9XsX6dwEt05Xu8RHsSqEo06go7Lu3aKd8CW02g6mYugG7kiwGGz6/ooEzz62UK
Euf4kl/KAmEOm5m2y/jvzjdDFSOff+8RNOHwHnjWBlGwhdVFPSL0hY1SQ+dg6jzmL1FvnmQzPZVp
hYNsNQhMSXnheUlmtKMRo2oArV8o8AVv6FaIBEik7ISpLFdEil3Yljw18dxG+C8/EJiDzANLPLSG
nD8IweiGJcvPyHWXwrH0MJvre2csJCuxNFKsj8PxwgUA
`protect end_protected

