

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
U7hExZJod/vUi3z5N4RSr1wa48P7uP/A8O0jgaKOZBD7WNfzo6GmQd7doggkH00XJgs7nLyNvPm0
0zWCfXninQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
k253ey4kkVql4FDzRxE0SZp0nnUl5fXV3ls/4mgbh/6ghGRjfZ71MsiTZ71s3tpy77tZHD0rpNoh
xUysBr1hFwWkTjAISVTsWyokKm82DELzMzaI0lqt04f7kevY+q4XugjttAECZCOOrrnUQb5ODPuL
TN/5/7rekkgE3das7WY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WoA52aV8kh0bkIXA7aISXPgNn7kpio3O4wNzPv7z4wZK/v9qsQ4Fa+1FXV0tZ0D+Si1URd5Yt8PQ
TB8Mp2LGBm7aAfzTAAqLpPZr3KRYlBsnuQptgQwkquHJi1BcDR3dhZHYw2oUKeYXBoZJ80Dg1iyE
mKNc2EAX8dBe7hH745fnWjhDqr0z4schwVFz8IHUPGI/WDdrXtDdyYzuiWdux2vjC9Gao0MkqalL
zCFAkEPTT0xtWcvaccmMU2ICHf+NVjiwhEmFT/vt1jXBw7quncqpEDMuzTHteQFztMFqsgBfXXAR
/Q4rfhaHiuQ7xUCcTEngpAsL2ypgKweMgL0LDw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Yb4xLqu3x9ghRLjHN7QkYl0tDMsZMeJQgGEQuxDwwPb+acIMCaRAm0LVh6gbF0arOSlfOKBs+X6I
1sCY01AUXvqPtXEUt+RvllN5odbTYkY9f5RujZ5aQ9olezUe3+JLEML7oIeJ23v82E3q5lEn2hpd
Yirga3+XXZGIeEC2Q5F3LdU1PK/hOr/QQAn7r3cfSPSRAYJBv2q0KFRrpHEdaRVBAVRTnMADnWqM
+83djfdVuwjO+GhXELQ+rhNH9dkL0cqvHYfgIcRG0rYfPORpbXH4Uiizi44H6tpqRpTeCgmUfW/1
kW3FxovGX7M2+iedny4BJan5eJXy8iA1/NmnQw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pj6m4D23BtF6RtOvVlnmIzux1ocpf3A3ahzdQxUHuwpW9nlstiQd0oSmGGaiF66UD31sHUT6dfQd
yKhb6vxivgHto8LAAEiyTiUmNTH/c41wB3zGzcZFasAPOJZMvUysBGURofn88ip4eLF52/qIKVON
l8AKPEa6atmUOWXPGRix1yyvpjUnvxZ+wFAbBvP0ZsReS6AW7b6zRE+vUOJaMz0EaWEMMRdw3vLT
W/hp9Ruis3IsgHsdn6M611ZJnxSa2tuwXuWdXURUJzFjnTsi2R7EoD0bDJINDuh7T6iiDjBFdO8L
a4ER9/C3EG6IOxU+oP2sYgSHnI7dLthCIjJ+rw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
B2bb9hbJCVaDRqGS393PhTqcBLIIS3eowUvDjLX1RVvD9vYwfdlG9rjfAUVzitJwz5TOhOabACyb
mMpxy7hxgVO56ex26Ce3uZlntRRrSfXZFQT0ENioLNV+BxEHrr7uipCant7HxRFrLFt9nR5wi4m9
ZZq5zS207DucLy0jTX0=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eqzUQVv3z3gvc1IAF6D1gFpnG3jJXG9SSewyb0B7YFlkq+2WoV55oUnb7Smo54ZcwqBR15BnF2xS
jlkL+wI6xvjzAFZaDFixez8MkTdRnrNZscyGLFWOHz7RNKwEpAxAm7RSsBEcZUaS6x+lEu8Fai/i
gBi8OQLkjYbSnKt8sfNmpRhCWxhkRR0QylraXCBqvJVR8s/2S9YSm3zj5TqvYxlJahDh9O3V0iE2
aVTZ//VjzAQrgKQboTMB5R+3O0GmOfi7O8vgrOvK/PiOq6kVyAYEvce5/1FU9VRi8AQk3Hi7BRZM
1pWTxx+bC6qDX+NQvgu8HPGpHmqeqS/CQlftQw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 506800)
`protect data_block
VTOXDTDViUV1uJ5hV2DDsostj/MYTc+f4zmx1KVA8eXZIabywhGjvWffc068+JDT4sGdOH60T74t
rkLGaDhDIeKsJ/chSR6r3Jmnjz2VQyt7UhDMVe+mM8bjoDWNlwbd0Gyf/gssZRCa9661EiJbF2pj
bG1zJYJv+j8YePwBZRT/m5YlYKhcadTjf8ptCjuTwspMO+vK6oQ4BecnL4TD2DU3GPXmD8RWMK/n
qG5BKI8XNrJxGR8XyhYzGx8oxiX49oQ67b6SFaMDnFnPYFLwo6ujzyOiTGQdCHRGcojKsoiKwolw
F+9Wae5kMWX+Ek1j7jTlsBGgu94TMOLZ8Of2BjwQSE8tZKNdokLaAxAeFkxUwsAQmjzVnXtfa0oT
+JXKw2W8nmj2KgasANif4g8/tsjb1WE+gEHbbJkAyLFy9rDz8ieqKj8tvCfRutX8Rwm2UmbD/7vU
4RVBxaTgHErt4muT2UJfKS8wZLXOxVqZd20udObNhoiaWA3Sz+NQ914sFV/SKwLPj05yGomyZFfP
ywl1UZxFvkxQkY5vAbs/ZJSJMd3Nn9thDcEbUUbGufZ8kie7ceel4s1vv9waLMVgIjmnhZzNr4JF
O4njY7xnG+SwZ4Zb3NluNdZIJg1lk6eyBuszjADnDrCLQpqz7P4XCGn+cB0TEy0JaAoVRmIgiZ3I
3sQ9rT7bs1dYI7xfI2me+OX3FDNqkeQfIlNSoD3MhWFMsKRcRuqOIltC8nb3IoOH2T49VS4fCYEj
a4mrjjXQCrWPfEhZw92FzOQZlPjXiPU/QPAtsgqr3JYDPjXktri3W61DzsfgRnrFWWx1/nMeJq1m
bx9IqwiKmeEGNKi4Y/vfg4J03FNkj0iPLTpcPaBfSAOY3h83Y33AgXta4K56eWy3etyIwcbWb2ry
GTGTsyCT6yPeS54zqqfRVgF/Fkoq8PAms89kS/v++cE9fEaVKTODLMt2uPisWIwABk2Ik9tK1DtO
PXHEMSsJHUl9kUe0bv58ZDpkdU94TQ5NLyafGHR1LqnoCqx1vu1fC3WxBWOSKHqXJL4Gg2CSxEWe
np80E56fgRH/4rkyJj+Hx4L4pALZYD/vtLsv5X8VNKOU6WAjScbclxkQW9HzuuD+WMjQAy3qbeXr
JV8fmWyfYZ+1+Tvw2p81TDMSYIKgh8jYQ1BASTgz4+FzAy+csCfYp3sDNxyTTIKrxx3X1H5EPVXN
Ipn2OhzQU7jFIpRB2Sq2unkOevE1baqgRX0XBBZWaSH1dPfyPtXFtED/N9wdew3efXMj02yqVMOh
lawPV1kbULpXGUqz9M0Ng4hk1z2OS5knYYcvd2QLp/WnEVYJdETbetBFkG4EJbvs8HPQQ4L6Ha2v
WzhvF7rkGxY+KNaOs+N/8cVEsPEich8KETEIHt7Ra70cycNthyMMSGtYIaWu+O4WpywYcfObNU4I
Rac3yE5OTDlcPpZvnOLVR1avzEEhdAkNWN28Mi9ov/LW4O3pEd30L/3kbNDOLulvplWiuikUzM7n
XA6SOzYjJn8lLyFme1eBAcf78d+Auq14lsSqvdPCfDeiKS2DbcWTiqjVG+38Rb9MTkTyYZapnUL7
orBlHlMMsd9SbD7eYmkOWrQbuHti61YUxIhnB85oUaexQ2PBbWC/JEoa4wAsohQVzQsUs9ZoT0bu
vQhgdeuGvZW1agc2ZN9WHM9JuxRKDpXqC6QUXhGJK5e38uaLvBZYM/Y/zJBqR/zvwl5aRurkq3HS
cu0/0r4jTVR0DBCzmxj1VEk0a686V8wtJC+JTW+2PlIWO2bIrikdFyvi3k2DaYVS4lK3JkTgAzfr
TUNP0z4cWubD5xVStEDknaZnCSu24lOa0r/qEgXUFMyTr2IysoZ4JHR2p9YLC6xyB084huSi7Euf
46YwbkNp9spv6qSzH3kxHoTedSc9yjWz5/FaOCg+lElYuW40LT3aL0wzmza/BGuwY6QF5GctIdqa
k8HFT433D/Fmy2Tj4+n3+CZYI5pfvfBPDBs+eWf+TpOjUKahfzjEI4juFCM8c7HUZeMRoUrTFxR8
+CILNuzC2iDkuuKps+xtFdOeWoxRceakEg7sFPrrg9xoqD9NHpJvWUyTwXBrU44ipM4I2GmFLaGW
Df87B8wOPSogkqFCk1G1PY9BB4KoXUAxGU69W/k1b8D4X7NJSRCs9354pL55q10EzKfKV0F+oEoO
y/482Yopts4o92y7/u8I0z1EQmEk9kZukAmXu7zjniLwohZ+ZiPoC8jdBN6PkvCZSsRfJ0nyBSQ/
x29Ihjj8e3cJs0SFcHUdm8SCdQS3lJdj57kA4MpfiBa3boHvIP4TAewEAloozCPnJPK1AZzTz0bh
1xgSidCyB4dYxv+t+xKGaTBkvNGWzhnmPyPPNO1v7WLVFrInSPiSa7j8hiJeeX6IehTWwCdW4qdz
aZPoOusL1pZh4kiK6pS58IlHXYgdTcUAtcmvcy42Ln/n+C7lD2rHOxSbkVmlTPOOv8uFZu+UCPqT
p5PgTOiVIF+osZ+LPKReNLkLVGfYoMn+NeiRMEskOk5MsM16GVYyKqdqlZ5bp228bhSxXUK08hfj
Nl5SpiKNinJ6lt9rldXlKviA+sNnT2o48xzu7/wEI2qJZsp7ofVEKja/rHfJMLi9ko+tLtxLiVS/
7NXBu7H8+9JaVWvHqELP1ZPHL8ge4pb+RbHLwQS9aisvLVXDjd6XU1shSMmnFgLKKFSof1Hd0E9V
x2h3Cmlf3fU/IsrAthnk1LJOJL3ivUtu9cNJeng7pgn1QYkLQCJibc3AH/HgwB5YyELAhE29/ZJM
6E+EGMSo3jn3Q4DdK90Viqi/927HMsTgXim61k9mGF98meQPn9QT02p/QHeYDrn5wU5G//4UetBC
7IpHhDO1gjP7cYUDe6COeD0FZM1k344IRaF7yQsa5Y4B63IpjJv8yGL3qUCulObGDkPRmRB4h8i/
Ia/SqOq0RcQ/A1X7u0IavpZ1ZWFtx3Yoa4uYXcN7rmK/juYlbLxvehtEfydj+8lQA7/TmsL54Xaq
PFfisfAbZw4NIBSoobFR/zom4mVds/OSkljUtV5oVcQ+578rj85w1GsO7Jf+Zieisy97eSBoaCUT
7TKhWs+8nAxc6GJavFHW92xrWIC88XSxkkgk5KuIaAkzCt5V/TsEEEBfhBDGXEIP7A6GFCnjjjfX
A2A6DilS3+eTfI0ydPQdqlnI88/nMZao6ibTWbvKkgIvrJLQ1x4ubw/OYaydfJ1ABfdHkMWSQWLT
FH6n31pZ/U4ZbOxK51z1T/3fBZ24u3BJv6zpvXYlt7JwApvzphW8YMXxILmK6yINRxkp8MkAv9YD
sn8vv8iI8mZBQTrC9IlZQ8OmIsMACniMqh6HD/UQT0zoz0dZVR9v0Fgy84hbVLKT72d6BvNp9RRk
xciQ75YqtU1wOuzV+UX8btCNBaRvYViN5IxWudW4Gr/iLJ6oCuthsYp7rm50SN3f+4cpwKc3hIr1
edI4MVv4ioPYYFDN7+98V5xJTFWkDXMyW5iDw+BCDt7YadiXkCCxzCoVYZZ5DdtdWdErI/Iq6kBN
nyrfNBzjThNHFZxnwOx3Mdq47EQZvdgy/9imbRlqcBeZ3ccXc8gZdaBOd4gyH2N7OMOaso2JOqu9
lkgMJ4IgTdle0XYQeKQd5OidgwRXj3Q9qqQ0KK9VD6x1P84d95CeIDoopX+2+fuCpwhjGIUBiLF1
Vwyl3JLCM9begwUdz5LXnbBawgErW3H42ua5T7bMNzSKrXFNFaSswJQrxnI0bQVhcpJWWTTiDeG3
fV+1m4esBRDA78M+99Jy9H6uDglRIyGKYMEB3ihyHJidd0ReVDi87Ph36App7ACCfyeNbaiKIaGd
//9+OEmt/Rb8Xm/zGbeCGohbqV3n/8QdkLpg6DzREQxyqabAXAUUo4TFyQ+D2rtX8Bj1uhxGAsUs
dN0P5orMPMUjlwDSTrXZiS92r3YeGTBzQswKbB9B9zzt2rmiThYYmQSCT6IrbzLRNcZ/9sRbOseH
P38Eb1PUPuTld0yrFXd2ZHlTSVZwvXnSZvXgxfHAou1G1JELLBgfGRdULMHYg42J7q2udtH5/KKu
E+If58P40Lkcv87EXEuCL0H2ws/smzaSLMrQ9Spk+RbTXPg3LTgFwnd2JyNA8drPhxeD3dBBsyJM
syOZ+tzgbxCfErN/hmz+iX2r7V+6rzs1b2jdKMI0BRqJWHRufSg3QgvXK8TsYFoweCh91DLUUKJc
WjGT8YBx6wzrqzKsljkkdpPW8ZyYWd15UgSxckqB4Pl/G5ODOu+Mw38LHf2dQyIu6ELqMOgYagCi
VpDPpXf8LS3QOyO/NCtY87bcM+UaO/AyQhTEMFoQOYuFZcT30Ev2nZoEjUd0JVaUcIe8uOQ1QzJq
0hB2EfI1+3tAGAEsdZLMGkluMWrQYPDedgOjpZB5l4JGrL3teS5BkVVDAFKnN6L89m2jjtvAzUl8
e/fhbqIJ1GdTTA5tiDmYzBOXNhF4UvCdfYAqJrSHDxFEnPH/8pyYsJYhiLmfQs+srvPU5l0eISzq
rXmXpFEvdt5ZrUvIRD2YClfC7NrjSav0rycOijB5R4W9Nwyq7Zk/ZbMUvepwIv7561u7Wl/vqR8i
c2LFm6BI2SZlEFJ0acKx3R/Wlmam5Xv3l0fMrfcyelYNCdXA9xNjykh2WCYqw2yP4r7qdthJHxqZ
rBuyIELTRDchub/nDE3O0p/UEesgdL3oPoZ17rvWeqYGIA6qgcidsF6a3BwrIz76SyUCC2WZ4V24
CHG1pC+zoZd4mCnC3hwjgKBoRypuRTZfcRiT4EpSNAJOKrvQ1OwwIQ89Y22aXalJQlam+fDg8qZW
mgULhgwHHaYCtvJNzOsDED5p3B37T0UUqXt3hB9D4Ldd9mUuqVJI9dKXeRUGzn8gFP5OWKUG5OTm
ZZIqozJcSAvnehKh4xVTTNbc9MP6mXFf4QmnHYabiysize1g4UT0dSdM/E93m59e83fNjUXDPxny
yvp40em79b2WHipjatwVggVOTrpIeRE0rHEGYZxzk2aiz8VGmeTjbaQAQkSZLBpDu55/n6VxbdUg
NG/XBXmRkZYVzwywVQ7FK3VD5jNaeA/abKc+NHK0Ao8lS+skJkbWkxkIP+Qfgr4mql19RboLeFpN
LhWSdO6+W9u5Ua+bR0OSXRzjRULGTWFUWsik7/BcgpiqK437tzIY6JLboRaZzDwjxfdsq5cgFVj5
WIGdtzEppZB1uK4HwnXVg8jRthwraJIzHjwI1vLqedBeMDh5wZ0rP+0T87+F3Efbwu5GkkEz2X/9
0gP1JKE2hktcVIKib2PKxmU7ahZr1b+EHKtLkghokAvQLelYUxvPrfY35/vSO/1PKVOT056VdFPq
ao8LLPxhR6G52S7BKlh6ueUoiEiUK+HptxbWcHf7mhZeAUK16yvj66YnHz5xbeu7geDazQSGnwCG
WqT/nHCcNPnGGADWw0zHNHy/cO5E91G5n9DclBdVE7Yb5qzH4nKyZ9SfyCXSIG/EouPpaXt1kbnz
6m77yU7bhESFZR+XTOBmUfxKtncilhHZyAhjtygzmHwyRjf4xTsMIugRSBs+KJ9LwQP1xR2lrjo9
DQfMxB6BZ81R9Vj0/hHkeZOfSgvITMyYq0ep5JUxsr3cbO/ytfQlimkBfKvQTtmcxItR9KU3hMXk
1PVK3/cWx9LSUl1bvdAg7OoGHQxX3tLBSvaGuwAEi41xw5/MFPM3SvajhZFYvrAlEdsstYTyYx7D
h6OeunhNUxZgVpKZ9T4bMXlhp4mVhpST3SP2EFujxoLbTBXOqsoBcikAS1BER3CJS8LZRzBTxtc0
/X9qf80U6K+XbOnzNefKWlJqZe7ZDZaic+D26757kyMr0kVR+dGYievIPEJ5G2yP77lbCtC2XtbR
IvzykRwJVMvSKaS4AbUabpo9a6bHBCo8nKqYOLBi7Gcdz5PaR/iLSfObswve4wdtI7ztQPvjMDfe
9MCqRpzYZiRCBB+mhpRi107odM8lsQzmJMmgNRdYn9yarqoCfYiDK01nwERi8w0QeksLeG+4agDr
dvAdhluwmMAUewCA3ql7b7xVKS+dxwq91SD9Zw2NAg32MMmL2HiZOGNEqlPkju+cKyJLDkVJTHa9
SgF0C7KAwG+0MN7fBlsze7E6xJPzoYWhP36Wm8dRRWeko111zD0GlopoAjfejb5NLXilUYCETulG
03lF5AndKPADFCLhG3eLShnzunygeawb+NjasI9hoG2U6R4yllvdEr4Q7PzOn6NQamSHFHSmwLEE
s/lTBomwn/Bh4ntNeCHa2BEhq7ESMWu4JNgNbIo6X71eodt0s8/vYHZg50ihLZM85WOvH4U+ZFiJ
KHQ1GPPz0E8zk01IDULr9SRwbbrCnYy4Ne+ZqHP2Sg6uS4oaZbRSYgUf8vHFsjj/BE+GgQQIdkIQ
IL28vASCoii0wuXIGXvP3A3365YfLcT3cV9LvTpj3o5NZiqVAVeiFlZpDz7HqFzOAfOBLQvSjplI
DEAIL4dwmCabrLr33wNKptDg5b9FCt6T3G50k588S+01ClHCEwLCGgByLingoRxjadz+/YPSNDBS
RtyZGVNSEcPy5pYWkWNE785WebHK2kmBYHouTgNnNe1WmucBaoyhH9aOhoXUkS+3ZzwyuxFSDU6H
JQ956ROQHQLQNtzQUyK2ZIVE09JYIQ4++Dv1MX2OFc53QuEFrEfVTSnh52gDYBtRjUS0S3O62ZuR
MOaI/axIUzKU6hyW1eNf85RdrbP8k+IyQTfCvT2WPbzs1bhXDwGjZtwAu//F+nD+kNM+PAVG0KMr
Boi5++05zRqUSkutKwpY4uS4E1VhAKqcrPnqY1yPotJejzf5bDIgmE8VFkwLMlU0RA7Na1bxQJIw
X1xg8dc0N7P9AiK5iXPJylace6qDKJFE6bdaFmPBKTvhs5fWSSY7TUnTBtV0oWY5aFZhB0m1+VXV
aOpOLHnGqTjK/LngHjNYYZewkhFPTRXTdGBjbbaU5w7gJim9Tp+z2/tdaDRdeR0cXinvRUMp8bjg
cwj5Wd3GFtPWUhbgg9wZrX6uQV9sf6yuQJhySiCGuIt0NHToiXOJYKOjrYhtwdI24sLxdogAjvKm
ScdYgdgmZRiafV6r37TePAiNqZykliCwBYNQ5TfltCqxZXkX825tl29xB5kL3DbO4N7wFnsZ9Siy
Bz2sOuZfQ4kWYDPzxDcIUO36Fk2CSxNC55h1Je3c96wzNSpgczx1mSjPM4xRMYiQUHF8XyKU4hz+
x3O2163+Tlf+Pm0c4CY9Rid6HiLi1xZdXxFm5duSAOOmKJZLTNB6R0PdWMnEyQsSKhbyQCV+e88U
v3/JPOwNXMl1E4a2fi8JxSPYWMbUX7M46uNpiCxrvdT0FTByGw+RY0IrUztRUU8gzjmqs3D1+Myl
ft3eI3/bpyxORLDjOWQJkcH7qnBEHh2S/vs2GF1/DH8hg99tC1uLDw1QRYWRzR4ptmiUkEPAtIcY
/WIIJST/06xOdizzQOgyLvAtOC3RqeG+Ym9Ldn1FRlcpOHICxl4IpTJo/yHt7tfwFXrBq8U43dJx
lkDsRzBHEsZyTk9CF1L5ESA9vNj4tPagHi+ipVy1zR32S2HSCF1Y1Ge5T9AyI9pmU6WhIrFziEuH
GcBVPyNVh2/2/FI91AEaqRWyy7qJ+0XQL9smNxQ6TTOKHZLf1DAfDzgGZ7Yd1naePOeW8+um96Hd
i2P6/EUnSWBEEmVubSdWTGkGgWAJ3RS7jAOhz+epc1SxW4gn4p7+llXGb/uqn6HDsG7GKv21drL6
rxka7jW0/chvS6xnHT4X44PmygbTx/a9wYP9rDyP3PwnGwdsC9akoHYe5kjx+fXvEJZUzcumHkeH
wGtRmzZH+gCNqmjRYFIdMpg3egCzwPcn/2aPrGmhqR3sc5uHz805qkubf1wlwnUDvQooY+k1GVgu
PmNcmZFpFsbA6BqRfu8nH0Wb79oLfaeO05w1XO5Pt8+rzCLITfhYuyUVZ+7TvCXj6rvrvA1AV3+w
yIH958M5who3RQzy5IsRofKvzmeMT829Jr/zFGG7foi3hGWeTkfHN0p0DnxOFunVQe8TkfWpWhS9
WBkOSlEzkwmJueO6WgqH5nFx3ABctFpIocK7lDXJ3/VQXZGJWtSdTatBPod0HhefJpW3J538y8jW
GE/Au8VxOAVdaplFf49oJwS39pqgAW+44hjWlOEyAupC8WtJSyxcdePX1IBpZ458RJusrw5U4VQ8
bYULQv+fSc1ZUBfkZ8Jy9+L/aI1WK0hO4EsIBwucDxwcdH5pxyqRgvF6NjzgCZsUvsI+VhSdBM5m
+cv7R2xD7J68lwMDG48pbBNMJhkmViqWbZK16KmJylJq3WWRgqSun9ToHlsBE76OcZ5ddTpxvH42
UsizIKx1bUL4ZZ/l9wcs5WLbbg3uaPVydpn46ulQw+L2oQsw4GFkezK5y6OVnzh+TijgBGVY4e4+
JhJ8L7Boq+AJN5VwK0RWzrsMPLAnXGr+zI1St1otcc4E2I9NZXtSNPAH4nVWK1PLZwg0+y5CGYxI
ysfNIYXlkAiCTXwlDck16YByWRv/LTefR0em9YgOPsKocAJYCSR62gf397tClrQt/OF/DjtWu8Em
n0WQUhaYLehh/wd+pg08VC9Be9ufBPoVc2ZW6GXLnUSyJMXQSrt3c9SNyRVu7/xR8Iqa2OTmLICx
JHqzRFaHxCShObeuloNpdqduckep0+W6uYqBDKWMr6L8maJM+hNvJ3gSdaNvWEzw54CCuG3aW4ZW
IzC68ClHcsJApVcubqrXe1yGRokBeyw3M1bKVy0AvWJpZcJU5b0LCcdxAHwTYY3l8RTkTkF0Wg9P
0feoIuFujBl7fVpKWebqfRG6tK2gqAxcGsYYwWwrrcW1VjXqJ4Ugx2wp394aEruOJ5FK3Qdau4oY
kYLQRFzOzWJ5YH0NwUUVxJEFFr3Skq1xSM88AFEkcxFA2ARR6/8LM8r+7SkW1rXMFmfXe23Zs53p
zZXk/nbb47Fye1l7jBk+txkD56qCm/xvM8ST4arwUf7ffvuu+jHWvQgErIRu8slMntlbXx9ag/V5
7MgTRhUZ/49Q5demmO1FLORJnlR3Jcb3iz547lU8cd/S6PxMRTiPD8OALPtdkBvcg4U+/JBdlhuQ
IxqpWDmkY8PBWu7nxKMtUHQSl0LE25G/SRQpvTHGKVOUBH+71PCpw+ARjCxxQ4sKceh4Qn64EMBd
oEZ2ILHsbiOJbt8WO9anvTcZb/dSjhmqbIAstFnO3LOsDFN67nbU9uRJ6HYGLrBlpEx4rKIJGGxV
t3tcz52X5TYklYwgkX51IFmAOEhHFnp9/Z2fhDY0wBmE7DwtwVYmbz0iMgAj3/smq6AMqtvvOM6G
pOxPDVqLXsyxmtdhx8N0PaugYA7URJbuoforQQD1xtv127FEt2O6kKxHEcjc6WPiPOGOaOmQ7dcl
d+74RByMI0OQr2PdrkN4mtZR8iGkjk0S/+cd06yyVaUQqkC4CCIDqZxy3VUVblGHXER9tyuiUyZo
sZ4f8hasbOZqfF2+AGABkf+UIteiPAaLl+2zUnhvI75695E+nRogik1NFHyt+Y5ZccbQO62l3HVO
NAoEU55aZDJ5WSsRoszHyj+evDdLfopCOw/teE9e2WwWmtFAQ1X5Cc1hqV2Xc6/zpQoYJ/LTAuZj
XSFD1hLdsS6p6u0k1VpSAgNcOrgVUapNdmVcUJpVzkLV2E0ux0+Ic5SD8frvVqbK0SGRviAvv9Gi
BzqSeEyC/LP8STK25A/YMUZBOvCLPajab4oPT5jN6JvxTs8inwIO3VkKcnqNM1FN3bv0uzGeVZ7V
aytId+CamsFEZSoYV8B5xaXwdaxGHSHFW69tIS52uJ1NSDsVk50j3PTRIKElVbnpyVrpuaHxgwIa
JPmlL53bCuiJ4940NPOCyqQ+yfnILzs6kZAcrzQwvIGAimOWBM97RPALKrNYMFYQf1j1EgJQx0fB
YvRIwspd3NdP4FMvOdn30kG/+Xiky3Ki9zXTTgMb20RTCKx/UMUcDhZjrYOpwhmyVPlwMK7GLcmI
vLy/vcwol5s55Uv+kRTuKuX7MyYKCJtESqu7g5bFIXtrKx8aeQuWwJqJxO2iID00T0AYh214VcyW
uGUJRVexKZgNk7ALllKEGso8pgYJdzWjmvt0w98NzOTkVJH1fMyDrzSsC0NU5f750KC6Sw3ZYQEA
K6VUSk2mwO2ogrM/QyZLjIyIsU0hALf6Sb4x2KG0d1euBGkStC5Lihy03p5sqTv7+YnFi8Gh4Tp+
xxXn2tsm5WEDaqY0+HKMkG9hWXAGTn00z2rLclyvIlymUocTKO0zQeocDrXwDg92zfQLueheGzpr
HhevVEhnERY/9xHCjDYJM53XJ5ChGwfbvc86HtUf5pU7k98yc7F7yhSN7hQYSsv03OuJcf9gRIzQ
kN212+IfI9bDHsYRmk4xyxrA9Kdd3WIimw47m/s+03IZNt5w+wBhRTI27fmkibQ9Rx3D6+IsiMkG
Pry6eNB/tj5feLK4yJelDSEA+e4ti4wN6PGFlUNE4aGSyL+hElEsIJD+uqRYtwvfTuEPfoS9PVZX
PZ6yQDQ7XVkt5iQoEJmUk/UovElWhpQ0QrCgDBjfMZ/fdLMmU2F0tQnhM5XM839Q3mBqBzjvLWAi
g8qe6aFcpQrHaJnMTFE+db5v9u5aKwMBxngRumgA+cKwguepS9oflRs4bXLrwp0cBwfH+a9GMabp
1tBayGO60vD4VFrx7EATTfGdIVWlIIvCeazokuac+HWT55tHH3q2CQvUCYBu+eOxSXYKXnI7adGr
yT/Cnkq4IRWfDE/Fc2bGmK9eUbMahucdX6M/maYtbgu9gAB5Vpf6S8Zn9l/QeDwf+pU8CSHxTI1L
rIlaENdjy0T1GomRFpkBHZm+SXQt+OaVFUOSuiBQWtbxUtqGAtCyCegWxe1Sxg2Quay4qtbMwwsh
BFJBqERCybvmZoMV8ZZFbIIQR07oJmFOKrV4Zk721nQfWMoM2psE8JX9aKu7nmDS3Afs4cE+ond8
HnFQ3g72za773Xs2Ot+99IK0g4hIvDEp5cXiJjvYXZuAjoAUcD9dkW7U07OlVARglX0KlhXpheyA
XwNrnR9JVrgepMCRwO1Eh7E8mqjgQYW3dzfyrv7OSyJ92VQqIvpzSFffJ32YV4bNOk4c99ySLYlk
tL596EMLMOuTX/TAqbOzKCnXn0Dg2eNTv9S6CY/bo5QxrEnZwEg35gnpme6GrEGPOj+JpioXNbIF
S9J5h67I1tPhk0me4cZlRs4/GGBIGvtvTZprVUpam2wrVx7609DdSpShpwVn+MIMRcYsdyob77rx
lWL1TAWsXNpYmB0qrTbZoNDA7nlFg18dzE7BGnup8Rzt4DLrQot7ZzBXBpsgAD5H7UeKvE3y4qgL
VHfwhoIpZ2C6mVZennd4jZpmcAkIH44KMGnlbuGhBU8Nmm3sdD7/zetkeAzdSW/Z1VhTonjq8roB
/Rsd0XDk3MoOyib1QzN+s0s6t17eZ30D6PEEsc1fzWe8ttvOkbjgijnT6NZlni8q7owhxb0STOLV
OvxSDaqlez+HNitlWBGaEWk6njbufebGTy+FzJyPyI+k50kTPHmMRsPXv68Y1PZeFPXbghRoLxWV
XINlVSlj1CxUeEQLvjZwjktHeFTpAjnILKtMrt3A3H6jpCcRNP9loGjBVfeCtLnOUyUt724Qn5Dp
L+ut2ehMVZhlp0f3VakZfe9VU9HeaeCQd/eF1MMstnkorG6bTtxhvkwnggZNEXl80oUAQFxPRIs0
RUTVHM9f0gtdZXAYRJ76CXneQpd93wyW7zrYRDDhhK0BAsJUK4+iY7CtLgdrkSEDw8R4f0OB0CP9
pKdzsUpQJgXxEFloiPZAC4UhJxrih3tlOqmetjmBgvnkpCoBBIMDQmmBTCXWewphBcY2gmOKCMAo
/31+F2+c7qnO39uEBZqm6tavmbAXof9VeWWaid8XoS9aSewSzeUIicBklj2cbx2Q1Ra/4KJRyjoQ
9zgHLf5/Gb6pVgnB/j/Vl14wo67Oxp705YyCl0I/I+7klTyIn9BnzMKwtgDXuPmrfJccqJsxHx0C
/j8M9wvsP/kvZfi0TZ5QLVWfyclcC3UWdPK6tB3+ii7MpvuYSmI8Z3IfeoqHLaVra1lCdLEWccre
hqP88np1T5APUB0N+ISYacMeBQ6LRnGFcaexc0ABuXbf0GT+s/Fdu8IzEQl5TJ45IGWflefbodX1
vc9ihZbqUMDR5+h2m6Z5FmTqFvaA/LQ27sokIowYcGiYqBKPWsWfw+6nlv/Hb1Rw0hGQvsGe9KyL
hW174bjkGiz0b6kB8Q3Rr3Oab6jVlRXAvNOQ7k8kXJDWpaSWS/kUXzDa3GaxCvwaPiUxCBkMn2As
EPo9MyOdEMYmVDaAMfFKh4+1QtjpR9AWRUgVOKQiLLTR37ZdPb40xsQ6rgf3pYfjKIdNNlUcqkyH
FFAqZj1SJnIjSbdElYa86CDL/D7hR2aBQtdb0C0cZhNQwCcTnE10RvOw9hr9dy0SFlM3hLLSrF8m
AdiF6vebJ+5Zv6yDmUQYYgoKsdYmKFTJu9z8mWd1+p9aPu1qCkx/Gld2xuUx9Mu8F7bz2lJ+QZOQ
jnwqMtXAxa5eaFVpNzicA9UgS/J16Ap5luAi7ZEqpkwIdPM7ANhd23elrDOmeHwwFXgWiMUxkma2
L5X0/nIFlDa3aO0esvA0UsYNB8sjmt8X9OJR63rjMLC/FiUMEb1N/+qod4Luc5+lIgAEBRalPX36
OpwF901QfooLycOwVoog2dOMEVUN6tjQYhT9Vj2bGoxdvLZbXs5OlrS9vuZUbEg2cVjWorILIUau
2MU2i5EXr3pvH87eLcT8XaIl6i46sf+L/HWUpikmKsQ9oT8ebsucvNYG4HWjEyr1+OpkR7Z/YdPd
MfGBHRKJHD3wk6+yR5QvKGKuk1o9sUI683+H8hacvTUXxdduxcE1oDWwlqHFGgulL5cZKr2gUqNl
s5pJfnReDVO+Q8UpDBv3mhHgZyYGZqaK/x9ltU/50Q/oCIYGSl7Jtbfm8cZoP3K1A1tGDsVqh8bv
WiyijWUH852Hv3YtdKnR2ckxLW6XgbgJfh7wgf3FpaUQDGPziOFNsF2f9QPi44hMCWGe/jZEjOCF
s0fNQ7E77ZlIhYGPJ2RLeRVJZwt3+ecijwnbWhsG9iCBENJidH0ScUEvhWFD+klCl3LAyWp662r0
OzF3ajjSpfQLjZ/THQHanWlSOW+glpa+BjCBOmJ9FFP6VNKfT/PcRugObMz0+9kGamXJCbPjKHql
Nszb3pU+9H13FwfgiXc2+DU4qDFgJ7ppKO/6nQ9i/CFnrD7s8J0dslrm7L92KOLVO9khx9SKwBy1
4YfyMlcMjtDkuScauWdPkJxXhji7WrbZ3u3O9282SGyis0UBzIV6EUrm8wo8wNsVjynNGKSPziBF
gkBUEikHgFLWVTvAkVSUzq9MoXgDdYdTxqM3VkAwSqUKrezEYcsTqzYMvvuHe0B5an+hDrZA7kP2
IfldPjBKCei8TflCiw6he2QJq6MgYN+9SRQqYYuIa2vYfizQyWpOQT5u+hkoluDBdG/oZK2ss1nR
RQluol3qOu/wSuMB+ZKMOS45UPxdusqgRR3MfrYHjkigJz0EetecrufuLjpFp6pZL5VZJ4pCnj4d
kOz+MKyQEnSwQ9+/c/ySwbFcTigMYhFwcxENTMy7CiGZkFbfKDvhEnT6ajxEt965iCj7adEq8dk7
qghDqnIY4aJoD30yTCmDl3kVitYeb8zrvp8wVdbSYgDaRDpQK4pEf1LZW19rAYSFa7cDGnE4Jrx6
Al10CFroB+8aVgNSOgw50Fw1t6D6m0TjjuMuw+y3L3VsO21cCGRtc9HrG+BkI47sQD+ByxYkurOl
RfsJQfKxPrkOEdH8667hgec0+azBhiCbF5Nmvme6Gmrm6h43EbZ/PqDE0tfgMkQ2V/GrUHhZdllS
QoVtMFzfVvL86GlHd9YjdgHHUq1ZKahTTP7XYePf5enAu3W0YON46TxVIFEauEQBiQW88IklwU96
4iy+ooePitUTrdHA8U7SwrnBprxhIHrdkUd9EWbECCMz88Lvi6a6h2imvzF34Aokgfnc475gWdfE
XAthToIYkrjCevJgCanDeLAQUByPgQb3Ug36riC5+13dR+gJE/ybm9ls/DVvkmXz4DuzqmD4JmhA
s4qQ2MUF4ZU5zWzSeJpenQ7yvsCPk+2We6g8Fqp+FtQAAe2H/+rg+MLtVWOwntB3M3kPhlqiNNtx
oI2OokZV1SVW0K4u+6voJCcFD/9dmS9L8nXQDmn8hMb9z8ymHDg5BPFPe04DqL3Ggrfy0on5wfup
Mn62qx0imOREqcQ44dIGEIQjlfdcdpp9igaNaHc947Bvgp8b++0PaurbdbzRcgky+lyBQGBeDluS
QEtNhfCWVqqvU5uN7NCMf3Kq0FF0X5ED3obJWqll1LEQmaQVzLVaF2PzlcQqMJWXrcrt6FIEOU0R
6mED0EWfT2KIxX6YYN4y9ibHEAm2rx0YKNrsPSqhZkMh/7oMX8tROcDZn6hlnCwpgdoswjiWhZ4Z
QGGzXbsWq5+/AHc/e720ioPCM7DuteiAnaRCaX5y7HSiiBxiBc+2enR3T2KICpY3U2zVzW55SHZU
qW/tA+3dpEQhfkfXJuIV+Mnf64GtW2GvWtrbfn7aQ4IbKK/gJKTTsNprrwfAuJrRtdvqT/8d1GdP
fCHNaZH5reEXVg6lQlcXaRBihUZJT9FBfPrO6LfAM+ucO9q1MHJ+xz1yUvs2B+WDnn5WhUXJkYYb
ceaPuwXxFEBesbU+/koUbBnQC7RwB9+QH1OBSVzIlTpE3zWZXUNnTpPUhHhN2HAAvmHgCTD/MLI/
m/4jLWpmP9NFPXRnWLww/Xwzcm69nTy0QwPt8hy2imS+p97OsCkuZE1DQhZX8SPK0Kid5NCCxDSY
RZeYQGcQY+U23WPx0drZUPHdwWIG6QxdLiy1pFTTzJSgA67T4a8bk/2yiu6JX6k1EiASoQ2m5ev+
VxTIGUy4xDQiO2dlI7rnjzTciZphkmAKsXzZBPOu3gj9i8S4SSPoZSWFzzyZ0eqGLaoae05wJfaU
N6OUzinRq1n04J+Gjjmkr07MCpykWEoj3RG7tPlpJWv2n3e2wqrgsJ6LSIHGYrvNvZi6FkfSrFZS
RemYicU5oQpQMMzgohtQHkH4XHhEyPNHXB9j1cjrWE1xSVlmkggxFseUXNAYby7PJ9RgiBd9WndA
IyOVJNla1MT02Iw2zO7N1QWM7yOqorQgz5tWj1BweNPseNAV7F6NECRoiUvjWYXqdp/J6gJ8qKmB
qR1d5cjSNDINbWIPgWFSueduHZy+rduVtO9sDxHylTWUAOAWLBe89vMLEt3Mycx29Rz6JagTmMb/
L/BTIJciSnPq7LGHvdMAmRNUdnqb504fRV6Azs9xQPjst32mrJzsS1WyYHjCrwQe0DYh7YmBanpM
JYtmft280xglKhcsobO4iDWQWuyUoulxdZMdu0i1Uam3XbR3qFaijVFxbSyFpjPjyOwA7DAsvD3v
bUBEdbRQC8Xh6Shnfph0i8tgpN+yeiAYbIAc7OgWqP51ySC6yG8ajo65dbF0Ba2Q9g862pn28hvk
L4dldGQ/y6GXF1gTfkIW+J9t1xmiv8min/60CJPWYLadKyma/a1h8KrNnt4oqxVeGWgeWECh1ClM
9HACC+tLp0bEh7Iw/6z2vY8ILCzUdnzdjKdaNyteaebYlmAkBTkbnRv3Mk79/sNU+IP1dkIXkX1e
RuhCi/Qr4MjntBJFmvou5GjDPg/bf9AaV4BI8I0+Osj4EE4AJlrL2xI6GIidt8jb3x9bvvZE8eNH
PuP4K8t4/vwlPZByQXfCV/sZpve2ElDmFpXh4pdtKgnG2kzCt9PrfsLRoB6C716X2s8fwrM3qN8t
niVncsGdGVIfkxj5NzPWdWKWUe+Lqvnjv638R2ZnXOcs8S2GQktKciZR7/90+Fxpz6k0etDldpLc
AzOkzrtOTahwSldLm2DcxJSCe1SSOZX5qPuq2SZDc9DH+9DDUGco/3bxTkmwEIUTDd0Zay7/oZrH
83fk53C65iV0okKI0e0eWpEHgV9FFnlpsp1a3UuTQrxMwRhAShgGmZJUdK/i/zaBHxzkYt6VPzHH
U3OSg3Wb7a9y4Pz8HUW2ZgOAJ55Z0YpjTBgFNx/+xbasUV+nPmxoPhzFPZvYK7tEpnBvTFAyNFWj
oLMwPmG37UszFLUpyVdY5WTULUm1PHcN1ydzSWRKwyYnmsvDAQ9TYcgqGL0m4YyCoJwwOyCPuVWl
DG0+sJuD9rgKHepBLGv90KWQRCesPrJnXQXupVFdEhZNeVeZ4xowyKhu6PhqIkJeWe3s+vwHGc6p
p8YpzcDF521FzKRBWzg1Rfv8libLbr03hUomaMSgmp6iyolBGVoDDMMj6vikjVB4mh8igJTohas4
Lxq98IvxDLGbCYVFWq+JS4KjuTOtam0qNn7ADKT5DuRpStMoXxIRWKUHyQyCV5Hw8adk0CiER7LX
VcqTUXO2aAxdI/eq7OyALgMxPMJNoHVshkHnCCIC0k40nyLgcoDAOS9S8XKuaON00KALvkQsKyzm
JqTzAsxiDkq5sP3tiFPr6BEnELFaJYpB433FGfJLuVODP3M0OU3X4ROS3RY2Cz5X/cEJ2T6zfNBp
rUhGJtXknHUsaGJMT+6gyIWEXdsALUj7MLVYXedS1QGb4OK2L2XtQrOz2RdFqFgTPLj3AOSRKOTX
7QIWB6DSYIXj0s1mZ2wvn7a5NbRF9d0oCv+KjEFKTZsCxmnwAV0RWK4PuVVt+tgYnmE4xFaMowZJ
BvAL4kyd1Td4qq2kfGJHsJGMd0IxKk67v6J76oi23/qbdNTAbMJEaGrFQf0UQB/YBN5i4+AFuTE9
mWRdziEBAhbyYkbd2SWUbbYHxkTtc+rHC2nbrK0g7cNvnJameQeP7x4M3iYWr3jM0ylKt7sZQh1T
kADFcobeumKp6KJyGA2kvvVb4MOg8glmF2kI8QuL7elAETim/dTlOYIn3+lZHymjWMRYjLj6C58b
DGCgXBW+PIPjHkWsQMBEmAM5hc3dxEXn3Sa97BeWZ5qkTuFxdTTe1ODjUQisEK3oNUAPAXDpE9CK
F0gFw5qby5LkLP/dDlJ/S6Ju7q0NN9keoVeTr+QS0t5cwgXnivExOPWoyzD5okYsAdaFzrof1uvQ
qNf5ZKmrDmQ5HgZKXseE6RkMEIQqGpgA2nZAnWk45Q1bkiOt+V7BbDfkg9tN11P34ELqR6UMuK5U
H/eoXAW8cYCyraPSeeI3oirXoBmcSDGnbseK8tdMiKVFRobBDurTM7ZKw8Js6g+klcWHZZSv6We7
XjxzKrwmPNEyAE+JsyKkq+F5CFhf2p7KyuWB9HCCEy59EfwA3+zOxHD1JVrafI7u2j9Efbm8QBZN
PC0tRZQ1dFA5j225tGk03nbjLtuFO4N/N544ZIT1XYbmqhKDN6j+QqqEsQsINWcwhKeuPcTpP2Du
l8BP7Luyz9kDSUOdK7BIdV8LbDjtcBTJSHaHHp8iYMSqHussZ299VarfG3GScHzsPDhuF9EFb9ky
qt3MRywTgZKz8uAbufF72VOt3zgvymILEhDP04QPrc8d6zqAmXzkqHuZQy8XfdIbOdBzaSo8HCWB
yIFNvMX8KsqKwLlwegwObCvmDS/U3+4qWhusLAFogKM2nVc42+OtBfdKrTegQ3NeJlSayTiZqIEj
Gcw1FAVBDHZtcaUpLDGjD0s3zIkfuttGBQeAJps199gZtn551Ye9GaercO0Loe3AExZrCCqR0L2U
AEDMs18cPzwiL/gn24f6ODlRecjIx3cZGH2K271lP6Z/Mqxh9hgGAojs/UtzlL19K8NO59814Bya
JY4OFuRFVhtJybNlKwo0IhdP2ZdkkaqIIt5qigWiEsYlKXk1flq8h84vyCxv0G9ncZMWKLHZhtpZ
Ubia0XmOAE2dmgWqvRQ3w63UzTH/Uj/cy2XZEZvod08E2P79zHobcrAujKCSLu94eMcqncrCADPJ
WzbM/Y3Om2ZYikT8drNaUMmf+mkEHz9FK6jDfs5uIynZ4yWKEHrD/ZBlekIsWbn6MNJoad9tZEGI
musKSBU4x6e2MnRGTysJWer+3MYoFyQBXml4rNnnWx9fr2Nb4PHU84dQM1xn8qf1WWeMyTfoTHYS
qqYZbcDziRgnazH/iINqYzoE0lK1efPb+5Aw+vrmHN7//imV/qetdc+MWjvzTEjGd459V+C3FOUX
eK+G4XHsUXbzP+xlS1VewduTYC4UwzNBykyY6faA7tFTTxeVxMxXaScwvozb1Rs4DjZSv2j+0QnD
iXA+qf5xRdGOHsLRlsGPDI/jwVhy4wtxUiaIz5VSZTpI/WW4xT6aLYz1Ou+rzwR5oOXQ7RwqgM/O
vfvStTXqwTQMi8b4t4dK4LCjL9wx4bHqF7Y1TkSDNY+TK1VA7Icu6bXK3Uf23WMuYvibc2pYe2b7
eBHgb2gW+09bDm/IzdpQQOgRMQ3DomzVfl+xcVaYwfBgbZ3lMlguMnewxd1KLUPy0KDwfvxEwFyq
BtkBX0gOrokF5gX/FM0KvRz7oPG0Xl5EqueXMmPSHuHaOsOK1OuUjeRhIVBypcC7CdkXSQyM96a/
7cnWIFAXhtRD57IXeusO62Bm76khts1GCTw8yOQs7KVY/j4aiegoUVCk08RMLoNXx+eOF/mEQVXW
rlx3VlIRn7k8vBhesmQDZcT4VoqRacgblx3UEKWHfhIUsp3FbGkGDKCd+9Sh2FfifZu8luIeM87a
GkwTN4Quh6/4vzFeTgrqj9sn5l3NZheLUlXyZ2hmTmRCUtCO+BGH9fgXuyXAAOG3Jr+TwngN8okh
7g0CjaJkiESeyC9W9f5gikYpbP46FpwY7wJM7ETF46KymEKReEsccQefHWlOwhqPewRwcvO7UsvU
NbqjJX4MVF3FptCvU4qnuINqe7W8AzeNOzBUhJ1PrXwZDIcsz3CIC/hP8+4/iY+MTB4/MBGXBkqg
qhGBhlrdvCC9XEXhgGCp7LdQtZ1e49S5bRCWqsYRFKcT46SoDmIGgRpiDPvQeU997GMQo6jEYn7x
b7i4S2LG+yeaMbNu2SOUvJbNEj6IsRir/HjXPZixuA424lRdYYyOuuCTYdO5n2BMpKPPgVrno/Tc
EBL9cEWWjJTaFg2hcEizmEnqsxqPrG/Pvdd1/plIwQyR+Qa3xJgE8XVY8bB5STUBJZ3HIkNRTgeZ
YqHFQVQ7lznAIhv7pHq3GY8uXC7XDt+goXNf9lnrtA96ogggkNlKlKEPlHsNLwr7dEQNUumqhfRS
Oja0nbAvlsf87WW5Ce+3M1lQhXhlAxEzuwfaHJBfWw1nkmYNhGzO8W+CICCKTevXuqzmr4yc3CoY
ZJkE5ovePasbdDMdCxcw8LK42mgv4219+974/VroPmGAKaEIWAqoPZ90fgq00XruJ0+HwKdTQqf6
f5qN8urhvWv3IqXiJfnPaiAZCxDjwjlM37AXhuCn5HGDGCLois9j8iUKbA0fyBak1hBBwR1JKID3
VFFW93WQ8vMd7gMHjI6Wv8HBP+iIogOCrPnBt2vgoIYpAdcCcXcd5ZgYOY0D3NwnvwdG4F5F9uQL
jFHPUfHklUncmIXQxfyufZSDdzX+YB1445VuNPKXOKncG+1h3K05t0dvreteMCxr/2XJkfGX2a11
t61l42gXSw+U5ap8/OjXiWlAIDHnCDgbc8hLj+qsrYtTpZexEswsCQY1Zb3UCe4XR8npI5/Mj+O+
wgQfK81ku3BmU47gHUwpl9ndD4Oh7qiy9yjFWPj5E8QDMK45iloPfq7YY2B331RCR+ntP0oYpr4R
WUGoZevnk3nLhpKu8Znn2dtev6z42ChVdM4fELgqKjL9rh0y/sAhxCBCDWoG6+10VIVe8Ax5Y0KN
+467ZGnNmLPKwu6+e6PZeV1RcRPn6LSj6ZTHZ4R1xaI4KXk2IcY4BNtuYr+lLmLmcI6cO4KoR5Ki
r/CmZ21KB+a/xocd/fXDxNzj3nEvCSzjVMSB6pc7imoGUhIZzLRGiTEhXLLKULbTZn81EUsMtY9s
PUkSCceK7jgQ2g5A0GwR6VcNaf6c5qachDqrw0VMFE4AjvRndcylH30dg01MR26RmtzfRg3AP6IL
hlidVyTwc5n88cyD67Kt2+GFuXjFVNjD/4yGwWHYhsfhUX7j1QP3tQGE/ZdBkAOC1Wolsgal8mZz
LV/zPUwtxuGhBNz1KJiU+0onS+xnt7C++RFDvH7W0/s/wSYoF2qlnvIhxbI5TpNKcgfX1UK25zEt
TXNewIF006dfzs8soCbwC0tx+lg1FAKy3R5ugibAmoQRCQ43BqIanDqejxrodrpYSXknoFIJuFXn
+1dx9AEYWUjeuVAgB+4A8Bk+XHr6uuel8SXnD5vKklZ2c0wcHpYQIDYZAblZkSUD7sTBdPKOVxNs
wAlCG/v+EjYTjQdp+Siiq3wDJssmZYa/lf3rLkQPcfmSkPRwMa+vAI99nWo+9+G0aJNiD7pM2NX9
Swp6mVWIa369NzxpOLEoezr0eqHi+f1Em27HAkzUiv9xD8KiFWXFnCgKEr542Kgu9BD/y/Jzyb/E
Uu0V9w9VD1B9wCGpiMs9FC+emANB+Bwd6dSxHF4YPvQJkgaaCgnmlKxrWSQalqA3CiCRc+9QZKhm
c8gw0YK+2LE3+aWJcZvrUKNi7XgsgjUd7J/CTgoKqh2RZgdqHGCZHGkDD/xg1tp73tXz6hCHit6e
3XHaZs0SiIdLKYtUxZAuN/q78qhnL8NuU8Ev7AZrDKKmf/1W6sTnisZXPsnlnPxK/b2k6k8w0uGh
Pd6ROLguSZCEFksXBab1LKmUwNmWrUDqLc3O7cgkLpdiPYOUx+DipTwkkAS2Qn7Wb4PKJjdarbtd
+tLDgU4eR79jAC4wGBB4qWnc5bhGz0TbzA0wLkdJtO4oyW1zU3OkGawoLvyL28u0SwtOvmDgO8H9
NgHRoy3onxk8AbgzFp1tcbsihOMleUPm/yK4UzaIUs0NWy5c92nCP7Uh7PROSmL9KnN5rh/bt5hY
OkrI9axq80xeVTJypZw/RD6Twsprp0AgaZLo/PRHZVJAV8f3Pg2UOgVjwxZWgTV+TkzmOMaFBrf5
n9lIKDwPKYzx0xwC6m4dlLFYEgGU/+TUnu6KW8unjAiRcpuwPFGccUrq4OjYYT1VaW22Qbtw/xfo
xFurTzlx4vhZKLl9ID6sQlz3khSJN76YVysZlKncSGQc7HS8BrUt2rXcw17tmpg+4g7/gLO969JL
aGGaoqK92Fk1SJhcClF3OLuPk+y6xn0mlvA+zyUvVjqoD76etohudM4WqNvlBihjCsW3quSQshBG
VPKS3WRJhkrw8Ls/DnwA3auDkxNH9z7rKE1IxHpY3drj8i57562y94MdZ9L26MmlQO4MPh0AA92+
f9ndVPhFlio2KJXPWKDFIKA753jUABwYGU5o6+gOLUkRSY2lm56ljqEdATZT4n5j5kv9iKZPqzL0
+WyiI5a5JGeHhLPXncGd3zsVFxsofavTnvdFf95bYv6d77t0iZDgWmUqqLCcFTmuvl6niwCDvSJQ
T917R61F4gZTYxl3oMS015lYhyoTNds8ogcb9VzAf/P8FY/ML336wiwyObMzFe+UhDe4VFcnprhi
Ioousbht1EXdLr4f6EF7jQa5ckTPea/FooH/TeSSReXs+YoUp+E54BkI1HxQjRGQo37vZWhP6NnY
jBUZ16ynYefXN9G+rBhTHDNzmHaIp+9RUj8dAuKBdgTdsLxGgjsbi6Ff4S+MDJ5eDtbQHnU9re4/
SsqR8yCktSc77bP+pXOOKNqZRqndKGUaHE6mvp8q6KcTE2ix8EHT+dMO0tDN/1y99bp/Kcw2VcNx
LqkzbHET154HvgK6vgXHeTocW+dkNG1FTxpK8SLiCiDNz6fSpd+wCm3Zf42eGBl76AW+c/0gVu0y
Fl/dGNoY+psJX5kYKQsIfkJtJDxiYPcK1kKc2q4Hs8e907vUVyIe820voAe9AEOG38m0mUnCLDml
n96+dS46WJAt4giv75xVLHSIyg2Ek0nj9JbYn6/+qzvWzfuuAADjMmBbzxnJDsPVicEqMfuaSwtd
WJGMwuOmdFzK/isXttkg5C/A6GN9Nux3fMCCaZswZU4MCMLHY2pb+4RkM0vVhTiiYou3sX/xuxhy
IEdUaUBasX6C2aBh9PTrt0XjAS1JgR7n+q8UtP3zFtdi7oWC1OfdEBUSoFdlizw1IWmZAyU7iqm9
ZxUrCCOdMkQiUF5a8qhsXgKFhET+oKtFuKS9iVZeB/1iwuPYEWjfik0Y6/Rr30M2hhPI+LnpWADv
km3WIFRxzqs//iTwug/4BbgE0bBaKVCa9744QsHZAYRARwaOkgj71Pz/tbfRpwbAZTnhDwvQtXuI
gSZXCVI1b1hK3ieFKv61rL3HtxPwzAIMepyuBB22tH4A/agQukZiNLpWrDJwdOM+013itFu6gHNG
YEeyFwinORhNK+w2mfB/SK7i+3ZBQAjW5F41hEHRdwlGdwgbyNRayVe54qzH1n+chisRrKMR7eNG
OH5eLtfM17e+5cp2YKf/0OUCk8TEA17Nu96i9WBm55TwtEZuz8Xj1WvendYxs6XeLzrWkX0OlbPE
cKqwijhGL6xsFkdoH8GJKwAvU0bVuQIqn5cnDMfVeha+RWFDGJkngBUcAGE//VXokQX1CipXNcUb
PMVJWoTp4PCMg3jxN6Ln8TVT+zG2ndr4+AAUdde/1pAwg/x3fir2WXmZHzY38x4ClZReIKBTKAlM
mYS8zQywmg9HOsbOTSE/iPiCPGs6O7nIvsq5HnEycMN9UvAdu1M6bnorzMIEjqWozaVz5baJWjbz
LpOZN4Fgv59F45HD4QyrnJfd+8koIoeYkklGALMrUoqs3kxOIz7jrJqbWHm9286vOArhrh1thVow
etz4DnJxshMe3rWQ8IpWwfUci2JvNwe6nCQvAn2YBbesnmkTgoTy5OPCjNebB3VMTyuqtlvaSVjO
4lCpUTV9JGdTp8aEWT3f7A2f81LrNzHLgFqayv3Lo0x9Tbpr7rcMsu0Ak0aV8IoEJSyw5RUvFoDm
i4iR0mONMZRqg1NkMvm+4s69M2Hmi4mryZtcTGwOTAeg55+vnlu6s4C1nA845NJua7RJYAZ3+cda
MtfDeExVATyGbMyZhfpIpl4UcfiY2yrqjYxtyBSSKD6/h4OhkqAuVJL/6e/sjktJd6NniXy1n/BQ
/cehk9NAznLD/ZkymMCMblvlg4SR0jeev5thp9CQj9CoBMHIEH2UOVbx0bOyXijvcQ/FLplEA1Xe
6StLL5G6F75J8xwVXnClT9YGw0wvwh1iILCqdFyC4Wff1+aQLNOEEO9HkkSQLAdSh0JJucE/kgth
ub16kJfRKFyeUguoci4Yr8vr2WYoJPt4Z6jvEFFiyHSUSqrzs63eH+QfWlKIuRLFQWxrnVnxDVMK
ivX3niDcnFKFPuDyHbsIJ2nEq33V1RvHe7FcDlgaAewoAUK80SRUS0g/1ffIVGga8GXJK5iTApSv
jG+tTWJgbHdE/h7EfkYBpBDihhNHjh/Ic2Rhz+f7Okhz1WNcXKuwtpp9m92xHrC21fgYfZRd9KA5
yIXKbP7uH6QF13tA9pAV5mzujWomF9a0poHmkMyRUx7du++1/LbiY1W3Us4rXmSvPkwX774/l8Mg
Z+pdtDkJ1UCDJB6A7YkfTxnOs6L8dJ1dXmiAysA0kEeQyDPgNBfDQDA/aRGMNJfrPq5J+Er4zCbi
uckC2M8GFnq14IZ8I+nj3dILgKs86fBt556uBKB80xnNpTSvQZ4AhMrMURSt+0VGq7nDvDJMsRAv
IFbXBfdkxvNN6UjUydFq+Fs6DjNCycCm/vzG1Lfps4JtPEiIocNuezUy33nDUBWerOJOp62EgTnM
Gl4Im4KyhCsJvA04ZMapPubYnhzrkA/w90CBZpxyOifl2J1SYTTr4LqJkiPaKzRutPXXxOmApxO0
gjQN+425i6P3Wir0HMXs76LGFQZdlXGdEInVJKdElYlFpVvrASQj+bCQpy5yvd72YvAIMKN93f15
RJnNFPt76L4LBShVPWbPxsbrVoOPzuiwRWDPtR4diJTdBOGkRN1twTaBRL9w4kvnsKiOF5VojZVP
luv2r+g/9d0vKBTvBzfxlZEGCXTA2Jw0GGk8mxk6SxqDN4Ghql0AWE78POoVV7pjpPu/i2zIWsGk
6w/WrORDE/wEOmoGCh4/htZnOosyczPC3TAWCaEFJdeMC/r0EB6vC7K/9izNC9BQwaqCNuz0OScK
7DZNqOvFm//8+A2q9gXKSb2HcIGmNJ/IWUxsJkaKg98Oo5lYeYxitwNnbOoK4sptjAnesOaHBdvW
nZI8NWSs2Cb6jyUU/TG9MomhhMH25FQK5e/VLL6R9PLR22hw2/Fjf1gf1AccCULEVQFyYnWQeR9z
7IOrPX2SBO7mzkLiJLI2bql0hU3qLWLVqdjwXvf5GrodhmzqFBK63G+Cwv4MpamUWQUporh5964S
PxfwL6kUQ1dNMpGgMbIkcEipLKymyUvlh+s4j5F3Kt7fCs9npd/WZxYx2lGuxNz9a0VzaKNn4q4J
iq9UKBWY081njFgXtCN/yijl5FbCco6QNQUguIDWpNGwLBiARhM6Olp1wbxcNjn8J/0CUq8E9Jzv
n/B6JLoKOHLr47qFl4peyCDZjg499ERst75mVm3uayzOwaZzM57rk6opxl1l3gYE3+w+ufdFvoQA
/CepCjADoW6OJG269b799lbdGAxNZnF8BRuO3gmDvkm7FFA9/AJ9pew/XR/HEw+1U8catoPnKUMw
Z/cJ3sMxA4bNFRE4OEz+PD5OCvsOfl7L2RUBh+C6X9wAXPbeIfOjma6GKbotxLVWtIrMLmFjlWP5
GbkANihA7Ckkax93Fc6kvmL0jRMPygRsS2BRuGdk9qYhg3lP22rpjmr4daDPB0mLS/u5qdFiR7az
Ynpgj/yCRoh5rgfAy+A5u4QkF/weU4MUIcW2bqebKmm1hWEeN58+CaXPJDZnFAhfz0zzQKAIqUiC
m37tHUQjkol3gwiaosLzJmoCpGEsl7dK7bXLTcBxWybPOndYgLIfiCwytMlb8p3vJADErZfqJjIG
zPhPx5cmvS0v1Me6bptL9sAsZ33w+NgPjSPBOZ/lLfIl9iutFCDFGZ2RTMSCNtn32lVAVdaOO5Zm
3NlWcChIE6a6BvIikW8cSHMGd7fJHykUKmi6OsXKvu9Gjiy5y7w8pNyEczjKeaxIwGiXTnCllLBe
s5FJVdEOGtN9UIoD+V4Nw2vECTEQN8LnhPKmt4bGl2KjZ+Vm9nLadHSzNabjnWC/qaI6aQcDUFzM
gtK/a6o1rKNKxg8sXrqgH3blthi2/3irn9SgKTsGSF8vs6fd/7Qjms94JGE3xJvLqFmCYs76jmY5
qsMt3g6Qb0oXkbTXqwnxflCEmkyEpCM8hzxFH/y2xHTtDlLRUmFG5+Yxsz47o8qE1vi4ts1ZLXXd
OF/ts5SH4eECyq8y0ZF7T42UtwXHai01QampymfgZw9EeCgXJN3ldADgk2BOInjASslBRiDbQXww
9cdzy6Lu0IsYo7+MEo2cgNfrXdMTrSsNZ8Oe+bNbBZFz2r2qjq8Q6vdElsw28XTTA3SoVqMacpYD
q7cKFeOj8kBfOaVLu7xoFB1DsUgOKZujs2I/j3SEM09QE2YIiBAd9OfgJ6UJXZdsO+aH34LiZZ2e
XxMWzmCb0eahtYwDv5pj5kHUTGfHusmex6CCyX0oaNzCoa3dkQNjE2P56itd09b6Kcz8nM22hawj
279FvAykOuh6FGGUUoR+nqOAW44H35rj6KYcHEaaqr9ZlqTV3o7Pzk9ZBrP+nnrrNYyu3JYz1e39
20HWwABEE+xAB5Bj2VKTFPc0lLU693mqTlsekny1ncGNS7nQwDFYfI6KyCSdEUAEfyNCyGxeFZHb
K/2sfbLo0oo/9UmXEvg+z+DaZjDzQ8ZfV+IfpQFUM/AdmcPwz3z7ChLw2v2pmm5JU7RC+hHsMcjQ
umDOMi3KSTW0d7EcaHsS35d/Qvw0DMt+Tuf98kdA81Oc7ctq3SbK52sW2tObKAZdtTYiQfMwMfQY
zEFPE3z51sjZ623Eby2gceY6BvXt0eMwXCrg9ncqsnd8lYoulO/dbOmjhnGY0jOplhdspkbvwXih
o9xrNbgmpsa7rvuNXe8ohd8HW1x18UwXN/rlZTScWIx5ZYJKVQULa3oY6MlUQUsshmfTFeOHygvl
+HRV8DymBz4Y17HQeIRv9G1V1WHOuZOYaNbBtGgKjBsmpbhUxqLa1cpr222HrkIuzbO57O6ie2tR
p0bfdri1i/hp9t2ABePT0zKuih5bkjh/tvut8+CEVWg+7SMuYiJxh6WPDG0YAYAz9rkh5m4BbmlN
7a6KqGnCxbtL/NtD0YMDt0eFV/18ynTdBl/nyhYwyAqHd3C4W82TtHCWsWi+voKzAPhVysEaaZ6l
dg9/OQ8gfGkLF83GOqXYZ6IgpkkUZCFKT/rxOb4lbUv+TFmJ8Hg5ocs6+LroYt4EPl8+rUxfNl6/
i3cFF7lacLbAlwl0ewY0/4jFK5a3AGeGO8hE13Yr3ENrzG5g2xVAaou+jSYtPXzNUKTp510xHWcY
HKdXe+dx/H+QbWvEzFBW0MKok9IpnBW+bOZ+NiSC7bODwe0aq1/F5ruo0uXmLOi+KNSTe0kj6NXh
h3ygI2skOdgzoSrEzsnqrT3SC9a6iTqSQW0hx0IZe4lX7h8EQsB80b3xadNHwMuUC4gWzct6uHLQ
7H9JhlJOr6TQei9BLdJwfhk3023yPWIp7eV6syGwxK9eYAE58lk1cMXOrBJQMiXlBKZCsbcK/d9B
MEEC5D8pNE9D8YPaMYd84L6la1ZblIY+gVCw1HGVgcJ27J1R8yS9sYHSzn5QPeO5ngTu+BOXDDZY
XZCr0iEz7KosjT7K7DvjARptEMi5sPfUBkwdhn0Uhwl/JEkKzrHETX78cAg5hMSRmlWL4hMBrb7J
/g6E9NtUhFdhvznhrX2Ua0oHzBCPyDv3qvdMDIzKhc3tq69ETWk+kCETA0d3vMgEm+kRlGy6aDJY
JQFcXaPkU7XZjOXDb0TIZXY3oMxC3akeZ2p/i5YDF6YF9UyuLv4gNnZQxYEhWbLwDz9scHbHvCQK
LYxLKPUtiPou7LiLQ9ZLtlm0tDCkfFUPd+E+3RCAZ464Za+iEPtWXFQmF6pBrK1I5wxlK841/5ul
AFUyhzu0hsNY+V6k9XSOyIgsvGyLneiiNY8+xflCBFDFDPQOeVY/euk4QE1oeoVhPBWbYdNDJaQl
70IU68IfelN+kTJl1vGiVs/djEzUKK2oVS2rNmhonD7EPvRQN6LGcpVoFm1B0jxU/J4IVp93SeEw
yt7u449Jey+5/NVVvMDmH67w9kWPjrBz3d1ChQMdiP6T7mWXWJPh1omUYUeWGl/wFxgppHtb0XBu
NdsdP/r8F6LW2IU/DzvWDsTCOiwecwNLyXtb20MQMzAmSn1LTajM2WMuRIhapQPiuBjWlDSchsgR
XDv/TatPmwkREGRgE0guZVmhx9jPF3FVvtZGcW6sBTI0gzWKUtgwABrCcZ4zHQUuiTBtMH/YZPYL
oVc+awGcTSqxXGOxLv0LTIk8GZzl/TwQV49+qu/VB4l0VjRm7laE7ZF8kLTBQ6laFnTaMLrNM6Qr
5d6yeW7Nj6F/IZTnrX9lNTuWQB8ybG9bvEHhNPrQrE+dZbqBLUl5mJos3wBP5L3Oyl/ga9XmIjJN
+14g2k1FQ0lHDVKMNYZVwjSrLx4Jlkyn4fPHR+C+w/kHmIKzKK89MWDrlkNgxa6bfmopXndHL0N2
mtpeuHsaRmxg9g2V3lrjGJ6s6fGGmHgL8O9WhPqSxD3RS5W17TbaB9DiL+uFezKfRPDSAzYJpTTJ
+aVeH0r9P8CuSZw9HY9ytua7Bs2cx3XjxiXsoo4DbzEjkaAmuE1NLzVkF1dZ4nuh01hQ2YFXVuFS
C5u6DxeylcuUPJzbh3MEgj/vhqJ2ITNisDtntX6KdvXd7nBA3fZIovp7+xZwA4U5ojtqq/xTPLvr
NCYtqdQQlHZx9muSoYNM2eibN4kSvm1KTclqYw1GqB/L6a3mizy9w6QhPZkcfLfPSfpVo62BjSCK
lrZn/YgkmIeTixDMcZb9+g88gqt4fH+EKZ/TcEwFvxZ9ymPvtmAejgl24mZe/y20XyLdYBlKk+iD
7dDYQIyexkwDsvArshAWY6D1bP7+WwSB787aeAcas7JyIHgBDUQW56Z0DjNzPz4ZDwJmsw+zQ1wG
ouHZSvyUH3987gGPJEm+FKSOqx2N2R4VcvbuTW2lC6aKDaAHv+9Q0RbPFLq9cHjE5d9FPGKRW38m
wz/adqjc7lILDpeG2BnUSGdjuna1GKz64qRg0c83GFrIqja/V9s022KquM+1RQHn7i33jAHErkVE
GUxNupvs/yBp7z2RnLRBWba/8lK+GF1dctph+/UZ2JT92HrxwF1BZj4EOehAzQiFQg50L37Kkxbc
IusDMgKWxhRirln1jwVJ46Xj/5+cngLizCIABeRqIWBG/2VKrTp+/XpTQ51ez3nIaQWk5vU41P8G
d4hmm8x+h3cy4kGZrvO1q0adtsnRqK4TWv5lhNHC2SxfbV9Qdx9FAupGti95IlWxBRleYtIzvsvp
gdxy3yfvNHsLW5v1EE3osM9kKAd1HNivNFrJgWm91ntVz2rkmaBAXaitIQ5sPd0v4GQyGYlBU64m
qLpeyGbeL26VYyXh3nfnERmcvwk+oblCHQSIcZeCGPuA+/J8ZZeVIIyL0rRfEqa+fFphN/HUlEUa
wDDUrJfIeKDkh2UQ7cd9AjaRXdWjZkpVN9Wu2CN/eJkL10Z0pw7Fz/6/s77ygbTf3aMYvP71hyYh
dWrhfTbiF/im5GySFEEwkurezGFANCFa7FVifIBzf9dHjbBJTQ8Q3/1Vc9gv6YYub8qKdeLnQfVt
ZgG4xunLzABbHWAZc0zvUYCDQNpcXZqCf7zy65wpqW/K0E4iIL0bkpFI4XBJTHqEhLN4mzYuJLXs
j0TSuktbxPGQ50Rmcq3wq7V6GU7TMamCvW8Ft0fyLLwrn+i59jBa+QCPXySbaU2PeNySOz1dgKq4
zMMvmgEfQTV7zOvJYtg3Y+7A4xWyhAKc7sMEOhHNPp4WvU/4zLYK+BjnkL4HfSiCp1eftGGLtu9G
0vutnHDQEE73sy3vhWXNhvCaH9o5YgScAHYwVrI6EI36iBJ5ZCLvUa3LkM/dsRXfoqjPSBBBlrIv
dlMbQ0ioe+thOLXgToJH1N4niHPh8sIe8QfEk5oSNqnmSw3gCCEtbbthSzdgeslRPrmS0Mz9/pKx
Y2Y/i3+r6oQ5lT8SfPRKrEDBhrAn5iG/34OtiRQrQWCZmDCglnn17c9lA0GjyL3w9yAIkEcFqDkO
hb3CFqrC4+hxttYSmKp3gg6pMH7mpzDxWM/C73yG24J9nnh8Eg7AFvHnmYHol403CHMXE0oQ57wX
iAIIBOG6XGjvacQGOpK3FhxRHXX0j7cmOPC8Jx+Jm5gvb4LZD61r1+5/Rr8SxBQ3KK8wa/eHo9F5
T+eq1OYCDik0catDT9U+prCQ5XFvAq/tPxon20/GazhaflBE9JVHDnWVNLZcRfrYshg/hEe+X34r
3gBlYmp0Pr/UarB07wW8LpoCRzbmXDg3Yy4klZovRNe5qKoNqJWbQ8I9ZEh6JyBdHvq52baxWKpI
S0kpuJ1CbUlHJcGollXjFnSJ8lBU51VDYbMA/rts84Mr4H49Sfhu/7o4iLYcVHDHE06Os/mLyIXF
mLr7r1ONV/2kBzaat55Cq0aagngwazgC13dgZtOTufbihY4eD2cIbYxOhhG630HM+oTMORynSXdk
Lw43s81C91e26UuAwzFkrcKXnhOKZU0rCKYTFkWhxNXuVP01aJwIE2M850gvkH0X7M5fQb4Owtkm
pnduZS2HbZG8XFzsT/DhQDe7h3LzQ/aD3ryAmwZR3UBSVtLm6HZWq/wLjtye+dNu0QuCmgy2J74u
MtJ3rwiBps47Ie4lMWtXzRx6MYxYJOgmaIhbSrQ/l2Hls85/c38UdifjAlhIB6z09x7DMRwShuip
4AELY4jrfHj5F/sW9lzJR5oH8WQ69c7RFUV9Rk7lmFiig48GbNV7VUqYXID5wNxoIs59PUA+ZV8f
CGCLv6TQcVSZeKyTtmk6jxb+j8v6/2zyTjh5pLA8mT43PrCzbJZjxShFXY8DUaw5BxQX+pvOsjXT
Jd+eVgm3Rn/EGamC9GdluXAobcIcKomvS8TpAdu8+c6+sglsFhrPp8UlXAMoujAa5TWNrnSORjPd
umoB90vct3IxzxFreu+2p7oCYRC/4BGi6MmRvBtR41q5GB7yRk7XEN6MvFNCbzBGTTCDMA1yBzE+
5G6YZR/rJf5n7RAm9e8Z/wdx0hDL2S2JvjYZQRPbDV8IywVqgx1Mibo2o3efZh+u6DVkuUJq0bxr
PuqFfpZ3aJM+o1zjle4ZSaZpOvAk231g6QIC3idTF8+5Wv0b0De9+b1CqaVC1BKJ17w6ggHb3kSt
qxpVino2DsLIstAyEpmTKabxN7YQCXEXIdX3edan5d9seghG/tlWVsG2Bajq4a7llHy7QQoSFPwy
rEw/zRtf7grU9Mtp+PX4ggMdU/L8uJcns0lWbT/nk4LS8bGkRnvpVE5kK2lPJs9UMaziO2diD2Fm
F3vT4FKVFcAVvn4vUbbAteB2B1Gmr+60tDlgB+Du4kp66gewWFuxjZMd76SoMaPZ1/MEEM0U0F06
gWhcdaE3pjg3Uj+ohKPGC+4xwFotE2xLGAQ7w8VwcMKdnN1pFc31WQiDrOZwJvNbZpGmr9usRBWj
Sn2eehGSXXwjOn6BY3Jk3jmOHi0nBJ9BLO/2JeE1X/RRPhZ2OPDD8vYbc7Tfiuwo0/my25ULHgdX
u7EjhZLp7rSEd7QVq37q88yRAd/1VHEs/H3pRD8jSmu5DDNbxlDWxXZ3ZwwSkebLP6hNYWWIivw3
P5q4zlgSuAj3pQhIslFT3eyfTtTyir37zS2xC6awssOktpvSxM/yyhpJnV6S0gVFENTvROPUxDwj
bT73B2BT8u728UfXAwtRNA1KK5gnppVcE0EoFpsRiiRowLQ6oVUSqbw2ss7NIh1IL6KL7DAgvjni
d+bUMUVR5BFdNrz372aZH5TDpiCf8qGufarryLvBqYb4SLoMoIMl9Z+oWaISG0D36j/Y9j0Mjjed
8+Bhh92ZFghqJBZBpQQeT1f77/10zmRd8hcbWPOEF5bq3HHMXARLmhky9Sc9E0gWSjYqOQ4yBK3t
y+QVDK9pMtwm/6Pj9jRvTAIhgUeEjiXcxJBwEa0IW6bdve4spq3aAzFFCcihfxWNpDCCUuY+5BfM
avlt7CGdv+378OEclMPMnW31NY+lUaBC9J1UR88dITPWMgx+pvqUeq0e/AZVLU13G63jys7sDnwK
XVbB3Dx1dX3EgYmqZLyVh6pn2C41C+VisQWgC+G7B77w/bZ7v8iEf+I9LtAegay7yOQp1qrpkeCx
4nqQHsY3TJwaqnsPeX4693b+QUYIQpzu+8YoKzXBhv1bCusv/y0wFX/+Zvyjz+AI6BxpK3Z7LkTZ
xu14SopRrVMe/xLVJtpSt5WiqwSTJ16omDz2/wp7kxoHnRZsNoRkD6eHBg60fmLVM3eWvFBH7nRP
QSnhPHJMW6NWV5BJdGHM269toYMe9ioSRnfvm34KCsaFnJEHGaQ33/PJNMueA4/ytpgUIpPeCQzX
hVgCs4EvQIekI9eeIbGJSFLvpIfhw0WjV4OpLeeQEU0JSU4xIMPYKYh6nzb/XLQTi6Q1hswWgMxh
7HKd1VtlS2uPU+bEWDsMCBJNX7Iq86GKGMfRx9IyVpmHR+X/Gmxz4BpE+jAzc5O0rqY879ccgz8H
6iAP/8I5K8E43J4/VdNE7qS6rYXPw1s9MtSpjmBl+jQz+tOQGK12WREL5qX+W8odPigteTMaQ/Ys
qKuQWhng9Oc3F8f4JGM/C07gMxXfP08Epi/CXqJu2aqA1qy/QJYCtwP2gAZTVnWLgfrXqACTMaEo
4VagEA9LmJhEk/0jQuOYh2SNn2P2893H32szsuauRYU1zVJTIIRZwJO57f8eoaKMj5ijUBQWUzhd
82pmYaQ7xTEFPQlSqwDfyYVl8kgXxf6ftK//aCksjMZyprTFhxnjjLhSHcTqNmRRk0aa0JrG9eM8
02P1I0oHB8DKn6/al8shlFBIPZ5m4VJ1xisrr1C2WpIWx4nwiFM9+QdULIoYHzQqHFBvACyOsVS0
gHRd9Nf/us4XxFDxtkTgN+DGjDjLxV1M6jI43YfS+uIeJ+qkPc91r1m9dVxrkys1FwnNDiR9T3a9
gfiqgVqfQ7Z0qIgFOwyFL0XbfmuBE69HD1B/MjHq8VC/HtrK78d4wQ0Dz5MfWbjkYh434MdA7F2z
Ec3un8o8/lxYJW4ssplyTPo232saJU06Al4fdnTfhQCKfPH9MZqzIi1hhSorJYeXNxIhL9mNppty
PY3t0tRQ0bHFn8se8tyVgZYdLQMHgKaZdDkA1beq+LNw8pf0RGK/JjQKZsErDTT75IexQSV1Icnr
6qLtYGztdzAP3meHDrhUcCnlvxwE7w1UtVT4TTTiQV1hBXxPGOql5QNaTeAAIX9/HksyBJa3AgWk
0Zqqd3/3OzsTMpjpMvDsYc20db0NyOjpf6cPS/qhYo/p18vnRlw6YAJ9wQL6APJeBQE2MFro63Gy
aswVKLh6vMP26OnSbSd0LcK1eulXpUvwvV4luo/pGcE5bCKatijPTtRWGn40n9EvwYcOE6l91ISP
z8oXROsHjia72GRjRdmTYu+lA0e33WN8O2qXPtt1n2TyNJ0qHUi6U0tVR2WBgzLEcJxUgZChvRv6
Keb0vNsNJNJbawOci7qsuEY5wRHTDViHM5HHkHUZYp5jARf9oFbM7kU7WnOsK041nVW4iNmZElGL
e+87GGew/aVNbsH9BKKAVTuQJVOY3U9UjZPjG1uGCD0+kVMQYSgKD6xXitoXrOBBF1fA3V/zjz2N
CjaJUzLHI6qdrtVV3Efm4DDwe9x4mYLa8xu8sWTLkVU8bNyCOVvzwZjYlQP4YX4YCqFRmjURfeGy
9Z8md9K+NAbYNsWWQRF2cCTVABKcJkD5rcbATxRaUl9+598nk1l6IQpV/tzuXL3F2pduCx1IQ69z
HhMEroRcarbaf2xMUDzRAEgAItVAxQ42EvWXdhyD3tNJNIuAojyCzs0+h8q2oj1Jhh7zxjyUopVD
CtMg11hN0PiS+57hkEG4pB0gn7yH/PcBxazPIBZWwpoN9hQetyn510RD+PpwjTwPhaqqJbsuTFuw
2WCIE/gnZ3om5872Jd0pcDJ99B+XnxwHm5Coc1l+RinfquV+OiW8E8+3S5nhdIh08C9gjGwyQ4UN
0J93Llw1S2aw1XRO1L08bZF7+oi0wK4pL+g70UdJRmXTQHYgZVlI2UfUKOUyeZEDbYl7eKeGa3FN
8R1ltyOGiN6p09fNQwYsYajyXkWhozM7lj60Q+XCfRFM2FTbbfCGPRIKtAIwpl4RZm/SbRRXG6Kq
n+KUSMSIoc/W/vs8uIzq4FoHgJ0/lZ3XEueBrQDPCpZ45NZ2iYfR+HGjWsoZmhbCnqY+mUvPjaTd
s6szR+4zAnT7qk2vFKJx+h6hcfUbnVSmxi9DUWsm1inPOtiRZD8rusyOE+iz+Q4hnxJmXiXzL0+U
/rqGIk+wAufl3b3g/6VdyC3rLeExPcHI8HJ/eh0ZBjszx7pFJGs8Z2QyyYg0KGe7stFYEQjvh1Kz
9gP/1MsX6P7ZXzo0SnqIti5BaGNLVHCf5m4ULumasfK3IrwtwEuacqajTAHhlfKeK7HSVjb5mJvt
Lxx3rRRboZD15xgLpbxvVa3lGrUL3PA2r3dD+R5uAhV7JZvZgJpn0yhvjFcRvySjKcl5I+35di8x
VJj79rOwvs+V7F8g23FMqFsoIu7nou5PTV5aFqnCHai46yhIsS7SEWlOFqB9jPsHBc38GdrANyQC
YHwjKwe3W4Tg1qjGb8IwZEJXU+juWRz+TEZb0gcKo47kD8MsVF2uPu5zRuute3Tcu4dAjMNo+Om/
+uJ/PU+Gqg8VpEw1X99aKTo92rUyiXj13TKrfykYBhdzHdSw33zYbbuyv16Kb3UoHrrgnGa+U8gp
7wX3Abh13iCWS0YSU/JT/Ptuo9ExahRtyRPLaV2w3yjlD0i6YENwVBke9gl//FbTSfJHARnvHLV4
YBWuTPunOgixxPvv28mAmd+tmSgz5E+Zmh7nOlf333hUZITI/Gq5pIuJ5u0O0eDhqiYcym6Qmtl0
o/gXhQA8TWTOBaARIlQMp9DQyhh1HxGd9OHWLmnTLK9AvTHXq6l0Z7yN/mX7DeEKcSWcccyxcwXV
ZMjg/+6A5bWgfmiJ0mYl23jGfan394c2F01Orkd4YEyq8qeHRTDEy9QqXKBTqW9LAF6/LHhm679Q
Te+r/vhMFLaWnhVywJ4h/yJ+GE1QMhiU0iN/Y1IMyQNEj3oAyxsoFQSt4VosP6g2P2Grkwub4WM7
HGjPO7/62ofPdmB76UBV7hoXXAhYipGvswTxkmok6I5izqotX/vn5xmg+/NMrnZdepdbGn6H+G07
mDjFA5iQEnaTYaX30SYYvJLvpGwg3hw7G33T6r/VxZwbVfIz2aVrzEh3zvtKM9l+ROhXlnRCTyAV
ZVOpAxFskh783xfv0Lk698bsiGZym+x32sdHrB9CJHzwc5RC9rP/LD8LeW4+Far8tgWq1Gzs6f2d
oXLCZHHyGZ/9ioi4wHhK26ik6fthhYf8r0zTcmpWwJRJb1XAkbgz3f/HX2Txinojh0KlHIqJ9t2Z
ewMZGnIKihta5fwX1u922+cFDvr56DIKPP1x3WXIHaZc8ZPNUeNxFOVp2eZrtg6jwQbOYdNAi9Ib
PoW4lrtcn5/m52uG0PpUnDYEMGMU9SJRHMLuXO5oBTaNKco8W470nbaFpjNloKCDqfHas5if4var
/xTQ+w8IRP7goiUW9wuXeYbQsjB5q4M5ufWHybX9Xa9b2vQde/oUGVah1j9uzrhXK5NEz66NZ9ZO
kB8FjocHUljzb1CW4LgrDvieOZRUu3U22yvaFtTkYqS534LGV0OFYtEtrC68ckCwevvmFne9GN8i
MlJfSdWVxQWhoU9YCjBu7FcCCSb9KsrJWK+T3TZoWa3Dqte1wzgqqdTlNd/KuifUPufd9nA5sX3d
2JzriS69GgRhawbKhm/LtPDm/WfOI2ptqzQ5X107GcQzCHXG+czfQYcjnjC+86p+CObM9TJgqUWn
w403SOfAXUO1wEDHIPr7H6ZwIr+5bc+OnUAt4YN8POaWcZZGt8sKEAad3T9a7cyAZJCt4iD/xoLy
/LhJUsYrHgwTn0AkExtwT/TBtVhtpRR3tVp8CUpBAUbhFklsm6F+0fb9ho7OCV650agNPVXGvgjy
m6bMeGqCrxxm/BI3BB17r+q0/jli55cZUCEJsKZ3mA4euQOBjczQzjwaDQiFL9Ye0l6CgLSkkN1X
qYvNDxQccbAgiZNpxYtFW/01wL7aggQqmqDP3lSzNyFSyuW2g6CGJrqgnNvOEfejwRnE1AvE+8LF
EB0d56zgsxcMLBuissrFrWOfrrVk6r4zhWFT7BmIdC/xqg488PEKxWeqpMp02YvuP5JzLe44hlG3
wYXsOqTPxCpWnOHX0SQwTgN3aapJj9z9FfLp1oioeDADlA3wi6zjDh2N2V+UaH1pOVKeW+N6Fziw
OVDMg+roeU73ZLgPToSTfOeky9vba30sLvYD4ViVLb8EnD5J25YghHjEWfXclRuUfFiCu+r7tBfp
OhqFJsfpbVyjlRdPu/5sHLpfX4eLSx196rqOJBR6E7B/WrqZg4or4qrVoKuCvmTrnsuCOM25Zg5Q
6eeRq32O5VEZnlNtg07Ig4ODCfFwR1cVkln1XSxVuPNGQKcG2cY7O6z+tBzMnUu49XCE8BvbW0NG
Dp565u8JBBBjZ4W2UTlfoiSCtYE7cdO0mt8FquV9kf9MI+nsRh2NCcAVVkQzMtdSarMx179kMXio
VMum/fYMK37aJVl5ANipa+AtibQH/aug7/pYk3ngnfcE8hkvbh1Nu806dvSYAZdQHKqI1hg9FCR7
5zurE/8DHYDHeWm/ATX3hvCmdmYGHqMTHL3+WKSzN/kWUbViyLyEMmFX5PUT8yrwyeutC6Fgk54Q
6FDMkDugg9Li2MrljGm7eyIZyQqusZ1wNiIwYBmvXmwauKJ6G7bN9yUhZN6fNmILayjCnPGXFhq3
8xB4CejeRTZlxvY7rNs25U3MhIisiG9YSZE9qDXD5hi6pl+a8dDpGWxramZgKSkpAFl6wBpTbxAR
J82RjaczN2YvZEQScxnUIkDCkz9jFEiqARQtpYjQqqVJuk4alMNRcCovOuMLhvscW56mJxANKeGV
8VLp1IkNoutNqp4YJdvaZCraxIEGx2QkXNA8eBhQZjxNXvwbFyAN5btJSQVf0Q8rF0PkWLihEeLc
eekab8r/ZCsT8I8PftpMkp4ZtS9vYdVBv46DtcYvXvd7S6Hg/6yW3PMC89AZEPS+v1PZLOC9DRFS
GYUJN5+ZUt4NkG5Ptf+Afegk/VUOnhScPt9DLi15+KkjeIIWRRacaDdQA33GKgC73MEiYEQzMMBp
TE3DMEVpV4g6iTekxTVj+Z53MKSbNJdPbBc8bp401HK7L9LX29bS9aD8S8tlfdWAg8WHORFxXQOL
6QAngrgqGO0UDjQqvTu4VxoRW90YS4X8LDN26nVB8T6eRJSnCfAtlMo3J/IARv3j12mhb7Ua75e8
RxeF2oI/N72KcUpaxdULlQ3cG5fz5ZH+FYnBj2JAmNiyefab+S55d53c9ZehuT0vE0Riq7qxVwO5
V7GV0iNKUN5cJ3GumBqkEDX9PIywIxTad8GMbFxN00g7GrZZooG4pnu0Xj2Z8t3FyWfOiJDDi7tE
l9Qs5LouRpaYGER3hJQTz2NqsZlzsLacFI1CLUOxtaY+AJz269ZVQOCP3YCzZw64w2xL0LR7HbJR
xGnzcEB4pYuIu2I68WpRvl3bG/CX8bwqZ372OxF5iouz2Md1MNpgCi1KqdXEm6iAIKR9GalVXKco
l5FNDtyTd5i5wVAZ9QH9tHZu/jjPvyLfZiB4g8R/D9irFxs8tUNSSKgmTvz0kfv5UxmHoO56YYK6
joASgPsl18pvsVqhY/d0V6Pa5SFyuQPpnkuKF7TmCMFgag+B2DjN+LHS6oTWpByEubtGEwR1AkeG
0qVtuuYiIE//jLduoultGIJUTLMMxzeoeSoCyMwmshCWZLqDLL8ai0pCVwM8wEXqJT5U93tg6ATY
xN9F30zaoxRmxl/xdnIkx1jg/PP0w/Bo1WR277VUue+nt+CEc3TYh8MWz6jAd9jDV3cQ2SShOqeE
bz5zWRioiQ7MC31gSTS6w8N8gu4ufiUWNIAvi+u9Xy1Ugi475wRmf+mU3JgHsZLEGtAupYuA7iLg
6sgtf3WYpzlmuG62fIEM3Fo02QBi9rgHlRjBjvUAbkX+Bl+foJC5+4KLcnAyzid8Xib0aeXbBpoU
jPXSWs8ggZUXUaH0fRn4t/eEQr8PH3ENnhbzVrv3WxRR3krVsjMDsu4r3K6lkVPxo0TKnsA/KQPt
mZGBy8qABKre3IZNbyGx7jLB5wpcPHicstDhw8lm0iTFddeZZ/DsrNhGDqB7B/HmBd8tGnRZRwwa
RckyOV4lXFcvR8kBwxkcMkTlNoTEd/cQ/RlnyWZIIVp6YI1H7eq0dTA2uY0uU+eYHSCPltGeCOvY
C4Aq3hwMP1MjMc8xGTBrVg3EEUPhVUL/OGVDkhiwxklnQ2tP8GO4BxMcl1XE6oN1A75KJepEuGUp
Hd+VUdwpaqnQ/ywbn8N+H5mZoHBqQPQEThrWOxlYsioKF6BlOFDDxJJ1a9+pmW9JwLb9cmER9sxv
+doMsLkRMYZ8hNBN/VacEP1cN6J9D8Cn0WqYom/1DuMPNFHHg3Xb6o4R6cIf+gsD2bH4Amj2d0HZ
ve0bSoLcuNqpiUAnu2aKsWcfhEhuUYwuw7CGrxSfAUIz3RABxC+oyC6IWPtU+ocGNNo0maqUOxWf
1isUqjBZY0dCEMqaZsWiaGZ3eiSh+LbgaQP+VZDSmMGX42O9yKn1Lqext9zY11xLuJfPR2vzZTpP
RSCS+W0MiP/cslkbIE4tp3dYSPsaHSj2IVf7vBxzHbuUPeR3LJ85oZdqRPYXKRhgaC7SlCDGZ9bj
8ZONEQJLg9ONGsCY5KdVKOaHf1hGB657ZsToKxXOZdGw7mROdfoX49d53eJ93aSLWROHo+8mnR5E
+bamkq9LYtrL6DIHqpAzCcpyUDbqd9fQdkClwUZ0GSmJQo0LypAnkxkgp4DAfRPdyZDmJxTsI0Kv
5mAbhNcrQCwoCezxktJiZWKkMSlHhGoBEIsTN057SIz4z77adsQTmTk0tfeBtu1L/tQfgLGdxGqK
zrYau3/cYk1IcHhmJX86rKlhYPCKqbClhvIisV9OfAS2vM9WKqjFd57rYK1WvVrKgy4IFu/JCRTu
5sXfcfIjV+8RZefTEVkv5jH0NoyRTK2JkCj86JMl8oYa5HT20c2ScIVLZqJ+E81ryxb8Gn/nLJAY
E1oMEvPlWGm5pdXzkO/U+a9kG4XHELJ88BS9mLMhSmxOUzDbEKQXDgb4fwSJAIjyVUBCj2260XAV
nIGuz7s/MqzN8ffCfOcYYW8u1hAaQq7eFhRcY68cRI1/jJn/JGdcOeA5KMmqMZ1dFDskTcrTya2B
NmAzUITSjfCi+5CIUD2fq10apGebN2stcZWRjuf6jNdc/N8BVH7ATwgPpFfL+vA2QIhAoZI+0eLv
P2mn1OA4Yph6pEns6n5lRnYly13zuTr5DA+qpuxLw/IVGf0qlvbVFCnJW0d8GvkRFveBGMflu1Fk
TYc3Vq04lXZhBNXtC1hd2QUxtJPv4bYX/k/wAleu2hwUMgjlnN+CceLlnCMkhMn/jlsCZi6HTrfn
+Sq7EL2zfRGEQyAtmMGh55N/7+CZF26EE9ACfnRgM2P6WTX6ihbLVGe32xahlBv6A7bDLboUGzN/
BvqXljiYJHyAPyWvR9xntTL5TOGD4TC/tbIiEQyxD62IlRg/YV2sKS9atViIVdF0wKBRaYqO9h4D
Z5+/81xQFUS7UFdhYQfHhBxwixAKVG26/fWTn+HsfglDgQvGiWYN2fBblJX8pV2k1W9QR9yKO0P0
CcQJQltCZyU9QZRuuN7gS0FzCsilAXlS0EzXM8cbFbF/pK75n7fCBTcgD3p92C1LxwyfXZ/eSDre
kW6pcc6P9AjEKkxiEzXe4ObpZgtQfyAqCAW9qO2HOwJsBmOI1trjbILxmSSXXs+ftVkDTEqGQvkF
avOePytsIFjOoXWMglNJdWQ35pgGYo+Az9/WFhcShqSGDilC4351wcVWbSWNE4nPTKP9L8WE9kfB
WOMSgOpY/5SHgEorz5dh3ngdZnni4YAEafcroB9UFZI/pINkudszbzHKHBEydWyvbr8OhMzcZOb+
6V0G1lV0TsjuL3QDeypmqKyuckuNuwDtVu9TOiQDlqIMMG/FvrdugrBLE76kmGfFzt26+I06h3Ng
R8L0cYExC56jSWqenLFVJqLItw9sYQEqE0JLBKmvGmeX6fO90ML5AomsALj2gYmdGdo7LxKPfLni
E3KU9rKw7SALGX6NHf94tVRNCQuWGfyOr3URXJdesh/CkQNFHndtLYoKZo09xUwrS7s24vRld4Yg
jL2Dd7wgKqZUSKJR9kNwg/TlvEWR3axRViVZXvnVYVGao2fu19H8l9ZmgDQXvTzjJzHKCpeD4DwB
b1GmbEIBXGk/drIdHIEDsW+n+w3A/2ybkXTYpwMBMY62ezPqyFhFSREebxSoNKq53v0bubOVNBEV
sguOQWPCdkP+7GWY9scRBuYDDOGFx20539LqyxJSLEuyWZHvILbwvKcTM4IfuD0WBIAmqZ8IjfRq
A/OuytX/QzSjfS4wXhJ0piJxvYVcRCDVcoG+dFvfKlLv3n/mELPjVZWoGd2MYjt/T50sE1p3MHTn
YbrndKK69lXeHscmO5/1WXaJ73zojVNKPUFuwSsreVGqafC80VAdcD3KVcpumlW3P928RxQmx9R4
SH9PxItZeUiPQuQL0+BoMcLdswDuTNnA6jQJKjEQkmF8bvTdrhTrbJDYfcX2E7KkIKi2opDoMbfC
fmBxtN/+nnSrafYsZOQeDjbWrGhR83MQYF1cpipEDpGeLUT5oCbDyoc139qaiz6pRQXdFbMXY4Il
+bJTpdK8ZQhkRVJmZDyMJVywno1nri4lYhXPteKNPq0y9vELoJ1kT0DKdX5x6c0pUqy0jG1xU30R
673kw3E16ee5t2YNgrWCxx62blCr0kHOpK9PTkQKNcA1ye/x7n8iWExZEnczd+vv1iuCy3vSNt9K
CkBTjBbGNcCTvsFnE4U3XnI14QrYUx+ODvWLfNZDflwvmzNWH1Az9A1tvjOymzRI2hsjVNiH7vM6
dvxAZnTSZMWY81fB4LSRKN2VGYJmIBuV64m6TV7bJ1LEEtz4wGZYVlPWIZ0o9nyIZIV21J6uNEQt
F9uMweh9qBipIBR9pRFgMMbYNlVHk8mn08oFBWuSjE9FVf7XrI4o9VSZWUYx3sLLVxbdqMpkoOtu
Xa3JnHOL1CBCXugJEOr0W80sDK5Iozk6T8mQswCxoGXAWK4p1tF4VgF4l+10J2sMvrhimhRwG0P8
76sBHpb45zOTnQVw707DDT6IZyI2FFMGwOZqZ8/H3JuguZkwEYOR6PvWdEUILYGB3vMHOCWghuzi
6TSmlnrBEeCwjqnGU+KlJtpvo2wMJ57PlPDNRcqE742Ykx/2Wwb9QfBC8YMOyrIxWg+rcNbBPHCz
GQPlPdS7XYy+pDvqv3FDVncJFwyiYoPVVrFBg4UR2hyW3WJ1JbnO6E+V0xab5NilGdq0D6VtoadA
5hzj7KQJDP0B6mJ5jU2rpmMF9z1dLx8y4Qtdhx1yVMRwaI5ysPJKu1v2Pv91oO7jtcXtxVOg8vQt
zhqQ0jzGs3m3ywIiR/9iPAiu92c4HKL41O8ByfupOphNGsCbldbdV0tmqDZaHDHHZbaUHGPkoxBm
Mj8woX8Y9I/B5w57TTyC4nfAwqG17YsXIT2WP7A8unpOxc+aVfGMChgmJ9VXPyV/Ty4tSu1fsq+0
1iWe7sXmvS3Cb1jPFVC7ZOZk9SKErQVeykx1frTaGtsDJJA0hbfdyryWn1qnqG/vWAhrG/dcquF1
ezlDxRnPANe1S8p74YAaoBtoqcojiaZpEMKhx8N2G2HYPLHe2z8dssSo3GZDjSOb4PuNY/qE7nyQ
QGrEGfoPvkGI8eOdq189eElYoxqdoXhSebejK6W1c0QaLkwYCYIbFEi+yv7WqWzmy11EX7MmpeMg
OxEGfyO4iemStehVBBmLWWbe5LEHWlxnILaAlUm9Fp174m0StbudXRGFhcR5bcO40KNvKD3Zd6So
kDrZywA1pqA9S9Warbr0HYgcQTLZTUteRFVIpOuO5uDWCdaaHQ+75Z9gp1ia60ScKvB9d8gRWywh
vLnO/EEv3AffA7VWx7PBQKRR21uDR5pyCzgr95wkmQdV9DYCBzZ/iH/ceooGGyCz8mQ8NobKJXpM
iCs8PfV3hk0ugmA4JMgIZEMTa/q6xzEEftgWHVQ/85+b345wzZ3LvvJHS8I8nXa7tqym9/ybdT/D
xRt47QKzeoPEIvD6AzY6xAlcBJ15W37VDEWzFH96B34Ez+FxbcADDiMduGWgbztl0tdOXYykx7iC
bfru1br3DRjJW7jwhD7dzg0kgYdkiMDf2IzsShZ/+iBPmjpRyK+R9GUH7x36iNCX0onsjLvpYWY/
pWYSUm8dLiMHdfpITCd8k5tKV0B0SgcgoNOZ7Hs2mPXkP5gBGKWiTt1R8gx3sjIDzL4sBOLsPTCH
RSk3atjZdB7lRnVGGSfgSxbiWgJ2QL/7h0y5cYCXNzj4lszBC7DBQdab1PHaFNOibDP5c48KoY/E
FYaNdAKhR99aLOOFlLD4WNHlU92rHSGdf8HdpmjUqx+6O2v6xtLCWT/sYQEdMsTutVc8ks6QotDF
85Zjt4zlCGKfUkDgUorOEtqLCAhyQ5gZHpsPKGAmAuajMtupiEOQJ6zjzFBZl4dFnz6026WJ6XBm
GkC3DqyLqwd+Q5jlwa6puv9utne1lNkxRsZ3W+Z6AitGcdEL5l+YQXCqQxDQhwsGn4Up/ZR63i+d
oKdBCBlT/niZhOTlsel3q/vAAx1KLnIaSXJ301JDKnkH41nkudRIt3F45+7jDf4M2F5gnaz4xL2d
7ZVF5eBZsolx/Y/8JBr0CPVWBaq2JRFfumvzAV60s37mRjgxjDvyg7lkJAwEet+8q2C1MRTZEpk1
pdSQCKaE0q4nsfon4pwwhOGFFIrs1unqPHrj+izhwZUwox4JAsj3Mh19k77xlqopxHkJQznfYXq6
Wo9NATpRqo4Xc8jKVr54x9xqmBVo/tuh97CPsseMUAwM7oHRxpN0ae+UWCyAZ6haKAzk2nPZMHUq
mpBvuMvxXJtyMuUygRWbdxSGMPqndelr65bpQy2S0opakoPxKM/owLzJrpF/foNLP+SQJh6KNemb
CsMljhtzyFm/jNGitx8Mvmts205Yex/2snlBD/WsJrTAVe0g0Bx0Y4n//8VrOibhKLZn5vtZ01R9
BNnLOfn8mNu8ptflC/M6J1D8PFOGB1fXjZOxwjLQtWChhOcX/6x+7kIdw/BVjl/zlnw9kq3VAMoO
+gIG83ZtZoyIQsCP7or6Y9rC1CLbcW6wml/JQSvn1IphdwU2O2gKOrCeiGgBAH+PZgTSMr26fO5z
2r2JyiuNGCe00/l6ebOKdH1mkaZqIfwk3mwaIBnxzwB7g4yb+rxlqsDJ4yN6zsmvnapEDwpE7GyY
7ADz1430vu8Ha7JtGhhrgRd7bDW3etIAVAchaVhRAsCNumLZ/I9WrYZQm3tIUAaxEpi9y6GxC9av
EDNWWq8MYE57jv8rDhku4kLp1SV2Z37I+0Ykd03TD7PC7umd+Vi7ZdirEN4GYJk2kYlGfaJ6Aoax
p2ogy8eOtND+Qt6n+9QbxjxPBjtj1n0SwV0FUYEgwg/VkoxCLPuoSdcRll+2lhzlUEVz1GObwrzd
OgS12FO2+nDd0mgupYnSsA0JmnJI1wBK2vwMuUlfrGVOyczg4VDFUgwbqw0IlcYSZ1KCbc4ZKWwY
Hhs+DbcobGG7dLkfU7JS5eL/CcOq5hjjPZALSCb+fzB6f90x5QquNWyS749XVEO59DkL8a9i8NjC
BNRz2Ewa6OYRsaEpdANgkrYROSUkNsvSblW+yPP5ryjg/JdCoNkRKIpyC8A8Re4KfC8/miH7YW6f
/4q1nr1oV6qbz3V3ymRTPrxzE2OVAqB7rnZjacqLD3CTyBWTTIRj9PAgNSeeWFSPznoWgJtO8mu5
T2epQnq56ehQTuZteH+nbwnt+fasM82jXdEAFTg/z4x5c4X6BXmVT3N3Qon5xLljIrk4NZ1H06AZ
30yRAT3IrsW9EO3kdnGsFnsWb/ADTw4O/JbiiRM3VHmUq3QcX/uzFP3HgZ7Tq0UILjtsArO5+qjH
izZjnSM1QcI5Xview9FGbglz9yLkNqKX6388+yGz1PZxLatlzbqYTEtI23f/NwEXwtMclSX5puXW
Q0wBsLuXHZwUKSTA22i6Hzxwlo7BSKCc1/LlkVRwmUFDL+qEzaEpAfvOSJwS11BPeCBmqCKlV0Gs
p75XdS+Diws8l9IDgVdzuMg14LXonj8gaAwbdCH/o74M9gpUKRKJcS0C5zP52o7Zx4S0Jf2GAhvd
acNO2bA3suaxWK8EE2Zq0Gdej3lVSmvedHqTReH8/NvEWbhRrdB5hwAvM07NyPF1cde/92by3ouq
n0NWG02PfuFnOtmeouUDwiHsrR9Cj2fPE5SiTPFb2uhSl6Yo6YVEhtptBHMPT32MnJR5ItaFB4HK
oNsohwnfI8u4OzaqJLJXzoQU2lYfFTfqLwRxhdKlNVnofCryrHYMCITabSrXimnWc5XpkOp7BYkw
5vjUiAR7GJx5GX9fdCxyW6ZDHJE6kmLFa7ubj4++dBZzvw9L3KhuEwjM8WD7ybODuiCp2aKeeCLz
VGY7mJtoxkz7/Bj9igbKytc6tIgQtb2NF+v4k6Qx08NCRc5Qcu5E6Unaa6y1N86wne8I0Q1Tnya4
YaIsftxKTi8Lu3gC2ji1EUYlgJC5tLjsQjRNlbgM1mS30kgwUAVUESyrt4rPhhkqKMjHfKKrK4LS
gMhIdW90slit5UNJ2qgtTmuLPmlRGm2b1+LXdsdtLwhbwi67FsJ/VKDm1EyaqhfQSa80BLk96pcE
pO1tz/WEoLmqOFRBPpXCfQD8bVpqpIcTjVeh2nV+O23qDqFC7nKj8x2RJDTVZNd33j/xxgRNEgKe
9eYHIU7apBdWn0bMPTz0pPJem3wlQf/goeQEhUhQa24pz57pY7waTX7oaIPFFPT6L8EwfNQSqFim
MW+rDLFPaJFsmTmTYib+9vWM2sREOqtHRH/mF9DjX6VBpgROntpEV4+sYelBVF0v6+fLaPWeuSXZ
dzlyTJHfgy3j4YhYFUsbW1cQWhYEVPAKkYIuKqOXrFnUwy2nZ1jwT0cUTGSHaQoTjGm68zgVF+VA
gW6PcNXsVU1JfwyTDGXwH/OGhczaGIxtgNlQPnZjk7XI2zoUiSRJZPs/YR/WJV9T0zDZ1Jl5v4mL
POdxuLKK1L4pohI+0QKiCJyu2b6A/MazsR91TQ408z/XS0waurZoKZrQ+wMM0oBadjO+9mSQET+P
OL8qR5T3SIiH15lkVH+QIJ2BZhS0vfZGYw9Vj5eZckxFK+Nr8NoqaVmy9g1107R9v+vzUFZOXoz4
wx5whOMlR7BHxPKntlM8eRrbvK+NIFG3Qf/q+QKbOakgtEq9Nh8tUJO/KU8vb+HGK/xonvvkVz++
xoNk/jQS7UhnqIwwKuM3hOQPl4d3fPDgtzPtrPu6mxyBWjzv6aPFruW5/XBufSKBunnP+TkFsJoE
4qZNV3EK5aJUcDuNiJOx4Wpj+IBC0MQ7Jg6e/gW0x2eoWsN06UQKgUjzbLooXaPNWgfJtuSOee81
kkcQI86spnNBAVyurHR4HuKYmGAzdQde+mpTKJcXwl85Txtzl06pWCjwChRLCkqbtpLEy4ka4gk2
9l6byCR782HzUeb8OjUirRYkc4vXSJ6VQ7HuPU1tPmKIfW9Jb3DyAtZo6XcCF9Q3kjNJtuK3WG6k
tfa1B8g7kdHY3qEEsChOnbaoYkJp2srwhIEu07gqpNULSiNohIK2IBe7QBb1xrFP5cMgw/YSNL5h
Q71sztqM+e6lviHDM4LisJ8SljKm/9Z8X1vKJP2uNHJd/w53hP+FGAFWV7mhN4QLcT6Z1PdZZJtf
csAXbWcIiqV54TfEEYhyxRpq0J5//DKnZ0i88t3yTbpoUu7COH0WlX1kQh49H0W/bBJ8XJ9dl5wo
5HIs2BveVO0pHwmJo4gFKdmpSHaxuxSAPkhF2KBudFBHJtAnztAA36kGvrB+1zeOeC/GBuZdvOXT
2OxAhdy36UcqxMMnsvrWOQkkdylOYwBNuAu7TsD/0gk5b7XoVQGY7uOF7ckrnq4hYazYVx7UACWJ
3UM6NOPnAmi2VJhOYptJmcEUQOtS0y/dQJFPeXMraKuYnY4z784h8sKFVh3yrls2x8YWDWaVTHrf
c0wlCujf2KCdWdCC5VguYGi3xH23nru4ILZ6Rf+reidvR0vgGxv8GuJEW7tBanl+M3DjE4RW3Gl/
nGrDc2fR/n2ivLmFxlek82zXMbfmadWbZEt0siQaC8jzhsTEgBFmyndv8UmFvT/Dt2vW+1kz26zo
ozCx9XVPbOlk18DM47P5tgX4j+5z5FhnMTrP9Za9QfdshqCqJvvjVzBWLFDRxT6ahppGeVixswk1
d0DavShAQFu12QWV6d11Iv8BLhQozvjaKAfeBQCSDvfauEOQIaMDxdV6kC/IdEmTenCN9+kisuR0
3ZMX3wBJRDzQOufXkXLh5qVlXur2HIhcj6Z7RYJ19kvtKXSvtYFmrFT0WryI5TxjIK025/RqtRAo
T0btDZTUldoCOX0LTLN7XTJLRW9jc0xhB+1QogdlFb7FTevA8qGon2DqdWtkK1Fi4BJBdIKKe6uT
DNg4kLnpTi5PfrAPuBX5k42FZdH4R35hEw5Pg4/GJQjFjOlm5qI7cuTYXn+EvZGNZhQehR7gBTkn
J58ho9R0+fylvptkL1SxysfGQbWFkLPV90D5WudnUKjMV2FJZ88GuB9buisUo8bIW010zFw1yAZ4
2rLhcwT/ByEDbpp+P8+JJ5M9+FIKplyUOtF48nBVc0R5kwBb9BU/l5gqFPKP23eE4qVMv2+3he6m
QRghXT83l7FQKpN9IaXSiH+fvJ8mTVk3s3UKQnobFpzhIx70lRGP127nNMFpRB74bUpco31FRHOh
pQHNMBBXPx/ennBUH2YKRj/gSXJGBzu8zpfpl8mT0zdzECBWa44PAMB9od1zrWaLhdg8EkUw4zuk
DeAHmqUlEWg8XvDMW2MPoAi0L2xMD1EHP3cJneyvSSzXC9OAUJV5zwLsVrwnCCQT6KzwPcJpuxNF
8KwKUBGtMxvxCblSqTFDbmxuLJ9icK1ja63TvNRvbKmeAr8hOlDJWCzSCmFA1PiFH5H6T6xDW5dk
dKgk4LKFXHJuLybhkHJCOOtJYAGU1qr4vwN2R3JdOt368wOpoaoUdDYn8NrM8HKJaS8vVXBvg2A2
NDORW7sEBKh9yHC6QKSnNvyn4+im7Y2gDQ3HxUhVmsGo26TGHHeH7o4F8QPra22hDq+LHFetwcFu
cYwM3Nmdtfxou5Ovcc0enuAr4SH/a2hDnA8bjs+Ed5jK/tE4Y4jEthvXgyc9tBoaWt1+nyjWoRqq
6Pvg4Gr/+LMkq0S38qojhEWmnXkY1q40juzrXBLLuoZPTx0jssAkdRabxFpaitCW80rpBpWReVDT
e9t6iYOKib8ogcR+hcNZ5bBoudVADm5ADg5zZnfuU4QFTgYE7KgutuEWe+ZdlzKwq0jYlCTqoyCy
eNG1byKaBI+pR576CzXx7qJ/JbPKBaNMyfEuHAD2J4Iof86xbi3uiAFnuX7QksICMbjYp32xQsxi
pvHoJM3Qcb8yMExePBeLUlw/Oo+aNCsIJm4ARYEJgtDUrw59kMuC1wnXxI+jfJRHXrHtWXaNEduV
idlD+8igUKWm9XmQtTOUJRNOy649Ec+JUJD7G9NK/+iBTvnasDLYUF0aemsgMIzAs1wDZCHHatmc
nLbnSF0JyfX7wT7oZcZxs9ZMjwY0TISF9g5hkeH+QDhS2DPKKGV/toT1adPdLbGc6tAjF0bp9T0G
uAExwXZ3ev5DVHoo8LwSulcjBJew5DZPPgzyei/Ew8rPAIf4JF2yGZKQdrPLNu+LquPxlnbWF4WW
wvY/7IyX0Dn5Ye8+gqSVIh8BMwWpniGKnPUXeUhKEthACtuIVFGLVkoFaNwgsoiysCxEUbd6a7la
POI8kI1PrcxxaKlxtWT2Mk4IXs/5BDu1tlRRGFfNacYxBBatA+547lUQNNcHI9Qy26diVmrojgaT
a/ozKVfUU19smq8OAJUf1nfneBvF+zk68k2RB2N28Ad3vQFYMf1rVDQbAxBy5PCsAyBcu1pXL2H0
eXX/cazkaKiIBhokH0iiIii5qBpasYYRSDIERK9w3l1nPkBQkHNxkmow69SMvuGVF1wv+hYR4un9
9Qq0wx/737cGHx291ID3QA/NmTy6ubBbE9WYmSluaIKHgjR9q+EbWpml8YeXJWLzlbSCQAYn6/fg
c393vEGFMCs5V5SxarUKG35W5dvHu+JZ7BdfnKbUq/R10XW9FH8pukpNW1WmtidLalrnBtXwX+ly
kl1YH2TqK9r0SfsJeMujsFXMuyQ7eRX+Jpx16z+arTcAZwGp7MnoHAuEdGgOOSPjJycH3ZOAH+HY
2uIfIDJIhK0e53OQlSE/YQ3kGtxItTGgfjJf/kt70b4bwPjOmhc6BDLY9WAn+PZczUjjfQ+JyaTL
F6PcimjkToqxIT9WUSZOHolkd9iXbp1ntkzDqkUXRBMtGFFAQ0r18EWk4/P9NPC8Lg4wfOZaUcqk
fMk5s5rCHTrC/W6XoReZOL8pTq9io9368TlnkUuZg4lX6cVt7QGre7jnSwE+pFIumKK/dIxvGGdv
qz1ED0tJJWRDUQqdzetMGGo256558XW6hjXzVuKJbYp7pisGerlQwevc++0c2mGXaIVjM4UeYsLi
jg9EU8LgCT2HncNyWG7Ev7SmrjsOGsO3LPXAbeqWtEng2wdu1oxk+OWOHiCGyEOYUdJdXsPsEU2h
3BC3Uo2WZh43GRRENoYLkC7QURwK/MYbz4j6HtB+DKanhcWVjOLvMAqP10pnjkR0otc1wEl1uq/3
eGlXspITvMACtqldDpx2Xp4YdD67INMM/XxIpOe9EMf5E93NtTnFacV1msSY3tbGMxsZ6PfKuMxj
SpRzKjIcbz+cm0w77hNaS7kUlrnR5EFxIJI7ivuuAnLw2Fesuf+X9xpdsch0Cb4YMcesEpQPC/qC
3pjZs1CiD7UeU4UD+vQ6YVbMF9WV30WrOVYDqeaBoZj84t7nPuis3p7ChSxBfQGZKg+1mKBHbK27
KF41TX5ezsMb1QCd7O4ma3ImC3+l0sL2ZD45CqrQoQUzBma1StBdIIV1wMwqnnNrath1d0hbqdXn
L7rjEQ6QC33/rY8bTp+kTxvV1RcMJksY4m1d5s+Zd+3v4ESFi3OylGo3nGh9HD39KrtJ1p9Ivzzk
BwTPfig2cB7YKv66CMm04hvlhve+87miAOkthXvff5TlkfctElYaSeJ9JULhF5myxqjDtSsgFE6Q
OHBzM95ZEAqd2HtgDSWaABfAPbQJcPi+IdjyuzlHmMWBIPwvevg1SzqWdxLX8fnqD2YsySJ0ry6h
rGEBRSUhlRDrK/fFUFrcuHZdoIuTTCIdEbBNgr3ceWo2ipd+SMmkz1agtXKwwecQPyASjHtSXvJt
HXt7VLcDn4fwCbvFfIi55qdRxQEkeYABC42oTEgnktSUmumAowP2n4nyqhHhLO+9ypb6BPmSx2UW
emiujDWoaPyo6I9x6ltXdNGbIuaYUj9jwVBy8Wqj1xPVJFqekV2+U9T4N1MOC8jN3KyN1DSb+dfh
wMi/aFklJp+hf4fOv0OsR4xUcE6c2hJjQ8PSdY+0I4woFyJUccM80v7UaUrP1RTI8kEuYlFRFXn9
Oyj5v6as8PinQ87DVD5mu3kQodg4+I7HOp93Q+qRG2rrB5fAC/smiM1rRuIPApci9dKV8PabV9a/
a5V52i6Psk3mVDCfs3mTkh7+jDsmJU3OFUHRPuAnKwfYjAKEtKRcagKX4ELjelPDvEVx1Bo0RIhW
WmFuNMzaK6x5iUS98J6GVRRscqa364+84f/semwHTQyPkzmQyeFV5yV12B37BV/rmZUHf10Fouxk
Ovh5+RKxaQBGFEayPwEtslPmVwsdK/5NjOxZa9cpC63S9Z+GGGWCUltpgD5DUN+diRcLoN3spS/b
Svn8uS0zgv9I79TG8XOM2pNMJLia5/yuNZqiACwk5rkdjToAO9ingzbQMKF9eVCE21jY7c42nrAI
eJUGkKMGjE/nYbmfBNTmXogv2pslgXj9E6Y+UkDR+5I2025JrtH14G2kbVwnf+fG/7+IzeO1cbY3
7zfFlPkrzlxbSSaTeHW/38hpx4lsPdJRgYfAVL2QytOSvnUIzWws6qIm2ddGA/nwbWPS9opTj6mg
+r2NMg0aV0RdGpZfKh+A/wwQFmz8fiwlhw9QKPoFkrwkzdDinWV6SQoPbeP6Sn8VdxP9N0gRHGPz
p6YykLVanYmhCOOSvOvr3R349xcz0aRiUJZZC6LjCohBGd5vnP8OZ0u+1eWbJjhaWMSS9bi+RP4N
NbwqjzSovtvfoLPZZ/bIY6sHhRNsN80jTufPoWHg7a6+RAdOKCOyPlr4FV7AR4LQvwK/fkADpPRD
O8X+4xvlRjgwSbQ4uTddw/JbXm/OKwpmWZD2wQRgwKKtEf3triyXcrHGO0209V1yfhxL0Xi3Pj4X
qOq3SZ3dfVZfU7J0jgjTh5ogT2wKhpHmEHBO49E0+p9X+mX35trAaTiFlAw/DntLS1VrQvqs++EL
qKGejI4FSyIapJXJe3ovwBtWIJ6NNx7HbFBlJ18DZXljdhuCBM+ZF7At20uK2v1mu1aXwIC9It4B
9m0+xYNmGpAzE3JHDLiPpIDHE7vYgDotO76PIciYn2YTevT2341Qj+11DhYquuqKqzBEnRP4cdJA
udvv5dWlwcg1GxQPWvw7ZUTKS0GoYd+TgWZn8jePHx0O/Vi9dBOatX8dmLsUZwqZoTcIZ/6VC/5l
kw9BUDpEnI+98SEP4EbpHC3GBlIEjQsHiSV8sc9LAG518yizlNcemJMmjVOXr2MVN/5fye1cKKZd
RzMO9GIEsCQ3wARxqQiaZ2pYH0vppRlb/Mu8eIP2eIsf1JhQvqkVhoBI6BAqwm/Q1CXx8OciGeyl
ppAD19PdVyqcKgrcuqjTLJjJG2YuZ4UiCDp8+UDD9CqMGtEZXZPxbbIjw6ntiSEw62TTnbmU4ODk
Dl52Om85KJvrH9IyVjMgvBUHjJbxH3iGddXW7I2d9ethdylt9X8qLBWciqCwQpIpdG88eFkgK5xp
AQG/R0CEvl6bh/8f28BPUT7/yKNLSVWBp1ah+R7EUgDtQ8zc/h+3677WJ68+B85Rw2UwFnEtTLmB
0eE96voICOFy4QNwNGGuw8pWPzXT6f4XrZFu8tnK5TCXNAbg04UKCC9hBrAKR/xQudK7zHav+alM
rljzmsBolKdsX+tlV2mTDWQRpxJyOccs0dlTAYSytLtgfMBdOYoHk2KEQ2RAI7cSodWIkw9PbIQe
cqdxfoCnmg5FSCozpyadbXFqIdHkTwCnKEMhicKrw5HMszgtvfuIAyL7XuroNO0kQNcZmVoJ5+gb
HThUXJotqshMq8sJhrw6e2w+xb6UpEXbLiGuNY73+IWQiphluDP6+BqPaM2upnu7/TDMsDaKO6xy
dz9W0hvqxRTwpRQcRuPg+6HppoBX5aw/BiJzSbz6kSSGGWhPfrbR5+/WswJBkPM49SgRoyqcbioo
KvUlANJKYyXopZABR39VuOhG4vE0wkrtd5fY129Kgl7gccrVaJNYe6NwEd0770PoeX1J9dbCjB3j
xasHb6eikSVjCa2GRurEY/OA/BnC0Z8xynIX+EZbyKvtv8rL1GfFZBmH2/oNVboLh1Gcl+Vq9QcP
GegvppDQMrX7GfQ5VDJebMZ/rpxIEXd7fgpVfLnDZmW6yWO1KjOouvX9f3FaFZ6FGRQjG3HHNsbs
i/y2KJ/1ehhBHz25/pz7CrnRd35W7UxDt619NuTBPkoIjcNljDljQbQEg6q0g7XdH9qoqAP7nuem
6MSiQB6eZFo95M1TMEg8OgQGZLWN4S+/6TdrJfxbcEqVsZh49bz4YVrzlpkpEJHj7xaaVbbkszL0
qdqSUiclkNINMpUXepIZ/S6haYlQlzg94bFvqDmCcPRsGfygisGYw03vYnhkU/n9eQY53pwMerf7
R1Xf6aVluS57mif/ltrqIcBr2q9S+6PudW1eNHgfrQAK+ieNW5wOWHpbGG/H52uMfGGv0gK/i6Wn
Ryl9znkkwgMDk8LrWwU5e2X4vaSZktBVPlTqg4QHsoeISqaMvwJZaxz/bbqKnCzoutVjitY72zif
p6hLpk5kXvWWmLgBYbijJ7U7jZK4/iiUJMpdxPzKBLqwS3raRcdZBGunp1ifYhArOjFdih+M8b4h
d/DB/bdw2adUKmIDk5U3xeB5dAnc+ybfx08hXu0kC9b3TGhAD+OCAf5Dcj54BfxaSuS9bjNc44QJ
U1HCJw0FrdUuezhtrhLt7WWi8Ze/r5KcUdiIYqz2qz0LjeO4v6H2KCTx/uC59C0bzNOVS/mAX8l2
AeE///9yD4lNqBQcXPBjG196YYFUX6dBhBYw7yrva5ZxSu9BRus7zDlhCZtcPV7jxsqYbmiV1itR
4adosE6tcpp5JJs5GJHMMW7FshEHcoUyuSJnYEJKfGC6u0dMfpWoTft2cyQ0xRnXnIjfx0XqILz2
VkBE0M31YQvx49ofqSwwzQPj/lBx3ONbSvzsPSowIeiSpz3n8gH452dCVuRubQebMcK068EZqvB3
7fJv+4ZPz7AjOQIGynXKBXDtPsXPxMt+PCbWrgDtoEf9S9ED4zwQWqnt7xQRVII905V/1kTIycGH
jqsKHOOyv1RKMzOSC/D3gl1PioI10eATVqE4tKUq2i3Ub9TG6Uwbdt3D88h84JWTBzPasv++5n61
az8eI4dq9jqY77K3F35QTXEHUIk2l8WbMLmLydzGpYGemJtPOO7gy+m8pEGPofcYAVYp6P0TUjx8
I6HoZVbbO9QFSDGTqt8vRUaNO1CYHj2CpO239Y1II9rS8ZV2T4rq5p3x0/Qi3nXJIrbx+YrtOfHZ
lfthO3jsutKum+UIyS+o/zCxN+DZbsdhYZ/WgCjvzs2CFfMNK5IA38e3ufk26381GQFJH8bLLMf0
TFzJvu866kdl9Qv2zR+Tbs1G3ixfuuQDVbQSyuhcPdzrEEHa4gSa7a/bA4TORWonSm4IsawPGDkJ
CzN4/8wTLNPoEgArtWyhQodmotex1t1CcxrKIVyfTSqQnLL3dcnubVivWXEHoRaPgka9BRY0oXl1
x7EpbTKAdmBgrgiXTjvSYvovjJmKzgv/ha1Hf+eLhbPYw4sQVt4BUah2mxkrxvZ9ZkyTlyEcKSUQ
5lZvZhh5osm1DUAqUCEC3NnzYXAhAIaOOBQDc3m4pzJW+dG8EMXm+KwPdueNOWlQ5WcrHpyiP33N
DVd2bkFFgtgNWYj6Q2anI5sQvz60/wMpj/roZTTpiejFFtqpPD9/pbfulRIIaVyz8bAyZ0bwW3m/
HxnlQPDUAOWSgTg3tThABgIMRGagfJb/cNj8/cvd5gLzB36dnNmMVa82WSweWX55o2UuyFHIup1V
DHTEhtX4wXySygB/4h1jGAMMoSwLjk0hqDuoLvGOOpjYDuxe1pzrVMK8JLocAJXzQHJI0v+O/x7I
b8nQf2d/O23OgizDlDPm1Sr9VeBfxO4tkS4geLP9z1lkDHmpqKkhyCJlH1s44TXREvyByq71RoZK
icYyZ9jRBddqXLwhy8YtBT3e2oVihgkZ31ECJozsHz7/NqW4kvxs6nZwtVhzoIPy6IgWCSpv4cnP
yavj0TwjawJfg3yK2CDFogh17mofaqNEgsYr7AXcriDlBPRMQZzgpdV/yG0U6kPJfnR77BYZJyJc
FbwdjLJx3noNgcDwK2gp+cBfhOYDzvcUBNgFo2AS+e6zpiy+gNg/DGlHw9jQS3LdNW/G8Wf/+g9M
/xjwEL82zYIbGuRQJI/Qcm+A0tObgYHPGQbwQ+HWAft4/aqRZyty/qzdsrNK65+g1F7WoJLngNXp
aOvCBc1B+eogsEFrhS5mrlDjiVmPjxAB/Y1RvS9xZa1gYr7rU9U42L67lsbKYMKlPd/a0vD1D2A8
zJdYak2pKZZ0I/UlqgW+etduppL+rq/PBY3ipevlWhnIGRrPm+59RyOWE8/CRZvGDOu1WYPU2o9P
o50xRmtst8sDhCACvCAYfuNNHhYMn95eJxLiXVa3OrVQAypo3y97TOCpMnG7OelbMH5F5dsHGyK6
T7aYJkZsal73ShhpxiG8r9N5oVaCvkBm/WO9l0EgfynoB6i0uaKXGAEYvIuSC29aWE0a0Zn+phoY
cqjQNX794pGDcCbb+wvqS3Kmm2aJ0XRMEDUyLhTIwE61G2w93vD//mTjktU4uCiibk9b+NJPHzYS
sjyd3UPIqlkM/kE16sYPxDQPeOJ+CDUx9tJPJPQudWtGW6+96iFOyvg/cecWLDFLhcRFQRjopAim
WWCV8pP+UwV9QRtV7YAW0TPk7frougx2Ev1anIF3rnuDWx6/a9fZ9QsK6nNxd19DkFmLyOBj3FSe
bBmwcDeTWK2YuX3cdjGNNT1Jt7zDDczQFxJNZe7dyw/SyHfpoahMGdtV9yh07NbNDg4L/Pf0K9Gm
TpII7BCAl59aVfh5V6ZQKDnzVdpZU5QyV0RrcVrBnYumbMsZQG5I7s8LERoZv/SzlVPCP2a6PrPx
rWSOOJKW8ZZ3Z0fKJ7RuEw7yap0dKdrWpRK3w1ms0NE2Mc4gAd7uqeYsEaeVzrz6oypAL2tn5TP7
5/C1maKF1C13DeOAoXPh00snfwHkg92aPTrXAc98sVsiP+kXtVkCGlUTIn3z76USWydW2GWgiu0z
peO2gzu/IabLlIaBRjJ9Boon2X5CKA3oOpnU9Z8cxZLsX20kr+yHaBK6mwXueyX+cZ+bkOMb4gTf
a7iplSjj7s4i1yndf7GIN+CscYTzGbYFYHOREbSAtVuZB4K39KWo+RzKyLe4zcTZzioFcUGNjiHZ
+dXgN/sgmofnirDHAY85mEyTR87gv9SLTmAK8Xi9h8NtCqg5xKnGdCAxT8PT21IOn9ZpZHQDouR0
0QeF6NkmLtw6kzaiBl4hU0GAdx+Hicxjl7NHTro4ZvAdFnhxz6ydTRaPevn013P7LoZ6LR8Ff98v
6yt9uHLvqebGss5TkKLdVnQN2WsjsNusRI19kAllY3UWPMhsdW2qWPsURyvtwQQDs6Iru5JaUjKE
+8LM2s+S6540aYQ7s17ChpLLfw+npJGivQr5vhxwhHTqwF0b6H1zaj5CGu7fvpPWxQG1ecMno3Zc
YVqeQ5XrM1/3SWYer0tNvcNBlLBgFLiZRLiqp3nV2QkEoOglCNBqqpTC33DCoOcX+pvACSm13Wpa
rT9svBOKgWDZHGfInuruw8/THKc65sNZaoBtWhiXa9SIdqkvezJQovaNarmaM/q+LTmhFc/Wo1y6
V37q9r43v0/37hapeJ0kiBlIE0aqN2WOwARxmjajBMFAfv3UjfVGYq+eBzab3xq3Mn2+c2stJ7mk
+rTkoP572PK+a52rDwQSFoIpMuErLZ14LLSDo2IGkhfz/II9+PFQROu5yUmHNYTR8oQabNvAWkr/
OXtO79uYc7pCvEGVIcUD5yeo+IAZmqkJ7J9ISaRr7BztDCHsxxw9wHDlc5K9c6hl8jdo8l+xCwI5
Mq+lb6EuwW8zyUydpv8QGDxO4jxK8ErQxWFTjZKo4i+Nixue/uAkkMIE7MskTPVM5dNrY1F3b/my
dGgtT7vEwoml+ZkdxaNqkFv9OOf1sNqcKjm6cs0EzkCyWDhUqUp6NWEcgta6NR5NsfPtPqLvYToW
ThMPrnFN7/dFUZRyhGMVQO0cf/GvNtbux1KMvHlsHxr2ZQe1NdmDvnoPLfQBqx5OHCJc9pZyLBS6
EDF9yE5au20gixPo/VUx4jlsK5qJZUwjU9WBGO9fzgs9dBKeBl5UvOAsSbVFv40d7I+M9g2Iswcn
CVzJbKpUuKNzvlxB2C51utfBjjUOA6qKjgaO1M7Lw7poHuojJ/8dGGtb9fvPU0jxyZFrFbTF7Bpb
RV/yWXIn9Nz/OLRUJKPNnH74JD/5FY1MK5uvx4NdiZv4tAuLFwp5aFBAmAKWCVNqOnIw8Sa4x8jE
MY/YF4CJDr6jKcdjF8CL+5Dfe7GTLAsJWtQ9N3ia8nb4KvDfgK6OXqpowhxA1wMVJVJc98SoobEw
7W9MCLRUkpa/JHRdjFy+UOqIENojHiLYH6F+P7BlqmlF/cIpX8SjFdN0DNT+2zj718JbfdDcNwaV
mA/m2yRX2sXVBbf0pWE/2kTpiXHU54IyoZiYcKxW1vwWszh9QESovn6Zq2Wiha9Nvh38Jf5CY2BQ
MivRwa86vwQHIZWG4GMXC2K0r0EaOxkxXr/xT563c6cUaqRP9YPcWgmU2nURtnIfuU/79o4abW8U
Xs48GFp8ukRU27T63vZdrxHjJBH6GET79sYiaRTmPRGVQO3EHeHobauaTzMWcxJAPx7uHM/2XAoe
EEXaU3MNkqA6b9z2mvOFvXgMETflDAmQDUmDm2WjZYtW/i0YgMQTUID7V7DhnxxL/rPi0v0uffhk
RNqMzmOoljXZ5X4Ak8TxCPeiaDQgxeLHMDfQpwr4f2Zh/TzbiMs/Msm2spB/pMUyC8nAVdR+IX09
Hgai1YM4f8th7M8E0uwBOxr7h7wJjLlyva2co+QH6UrJBj8Jp5zQuOYkF8L6m0Ivy9kNgivkP6rD
Bu/hFdZfVl8oBLd6y8aEFGjgcjkobnkFQI5wmVXyZASZwY1qjCW/6393kgg4kKoA+TdrhaVsOF20
gsdN3rSLYLkE8Vo9rueRy9Gnx/hfXWaSBCNFUs6GtRg0WkV6TsVAI38gtQJbwV+SWL+mXa9EQM+3
gTEH/C335IC0c7uhXwkCkrEnprxerBPd53BmS0cIdiXAEfQj+jMvEV5Yyco5NJnCC5BFxdz0kutX
K7iTqFbgoQwYNrm1mh2sGZhh4DcFz4vDM9yDFBhoeE2KpWpFKfNlf8d5k9623HwbvalX+vmM6TM8
nWf2B0nCwCwEDEUuXPSbIoKfpS1lrjFitMbawCMT1Tkp0XsqVpLOkUxxKrSOYJMGpjZXk6J4NTXy
RcGNhCVbYm3S2S9zIcq3K0uPHYOSpnOOOAuPKbT0FO0lxvU1tq0A9hsFJYvQJP3vlxLAQYeM7vw/
3kO8aKobnEwpuhwVGngJ9FzPsCJrq3liYO/A33A5WcwZsfamXaGCTfTZNe+GRMShl+B+xTR5AohW
iHw91cNkPDdj73dWGUq1OiHanNPuFrSZRID/MN5HS2fNj58Xt85HtXsg1sCaioj+LfY8Ne2kOex9
rCTs5jzx+w09B9LFeqj/okS4Lj4p7qjGjr4ogjXea+A7rPBV31HSgTKylVzaHom8eWwpNIZtQM7E
TUNlx7jCppp7W4WcS222aRQLgWzfNurZ/tokiLB0jL8+2Bhbguu+WD6IAIzdNtcUhGJ+cgCwpvFT
2YT1sArVbk/PH/1+IkEC7un8iScWkPWhqbiU+aqf0T45PFsnY2Pi5q4kmtduXIdX0wlF9BclBoNI
9sgOWDYH0BFz0so6tk8Kq+TwboDKAW7MrHlaGMjWMR2lbn+kLLMU/Tv99IaEdWJ6BDcdO7ziWvnU
rI5BRN0Bmfv5KLYqcxKgq0s8nNUwLmrqzTbmNYtYz3nCDbIKWCdBdhf0NwlrTE64aGAdNYxROuOk
/TrkjyGHMc9qNV7aWJX1nxzY8Y0+92q7n4OpZauK1Y78Zila0Czo1nEDuzRfH0qM7PKc/QlNqx3i
k0qX7uSXEbPmXK6fBXylNKi296BOUbQjfktynw0roKR5f56cJJnCQuHu3rWCDXjLx97I9zy2qVnX
5x62psMrxnSiBKTzVR00KtzpgYpfFwjUR709+va+uZhtSTV78C5w6APi9iljXdUxXSM16REWuMSn
Lo1bYq1guuyuwWYCD6CkHYvK2ffGEtShD5qqiyQR+sEowQULn604xRZLQz6lIQtsRZH3XyvhW0Ry
83OuOocTdbL5dPsFJr8v/ZhlwUPz3sGLREqF7p4hmGT/HkRtciuMzChFLOZH9eXHwrWRnzTXRay7
FSx4ACYb8SNfw1t9OAr8MD2J46MmjgHUrfYAn67XxfMTqQFjWjcXpA3B7GkF8rc5FYb7lI5h5MWJ
vAux8wu5I5XInOR6YH8TmeZa7UTZ2j6T5bGAF3cTiD2LwR8aPXessZzo2i8HVvSrRCRmgn3XkHnf
uSnRVL+RqpLkG3Ft9TQez1xPsXVCrwAWCiaDESGViat2k/RoRJZ/qUAjxrWLxWWh53fVx//kvd+f
Kb/7p1vGtJrGDZrNFuTSwwrBJZOohJX35LvkZ9DFHO73j/x2dCUaHM44dumqaJjija+k7aUtFJyn
0T9+naW+XD0Q/7rOV+jXt7P6xDTpSzBOoGQgJSFw6UJF3vxJrcNM9C6H03PKJTvm5n9BEHUznC7l
Nn+0hsb+YA4YbaVnm/gjfQNFYus8zhH8EktB2JZJ08Np1DsuxFw7CjhJpnxdIBOZ8YuLoY7aNFhM
557SB7botqkiUZXByInMMtHN8Td7FduaJvkoKYDYOteljukAWwqPWUlkivFr/Axm8qBGTRulH1D/
KMsVYtdC9lhZPQTrL7dKNwznay30qypdr0nIBatkl5eYvjqzIgsLq+CbEU5cOh+5i8aAZSd6ZBup
FISEJZJv8Iitu4mK6Oasuh+R/Gklny+c9G3JmdtDHievPmcs4MZsIsjvI5nub4X1wvEZOySOF9Sh
+mocyCH1KMfRWID2/be6CtB5SS8XF9AdYAlMS4Ikg1qR8vF9kf5Nq64lwhXvphTmnwDC3t7tirrK
U2FWPuD4SrNo9CjzwGraED0ulUr0Djim8iRFUZNMvhej5u8cEylwtw08DImuB12R83jFMOY99JPh
2081CEBM8Z3hBYGWfNalDmdOePjHg6VYX7dz5N+fGmEaCZdgh5jQlWH18v2/5aQgKac++rytvzIc
oC7DiT042jyoep9EKbmnkGQIcgwQBJeRS91dpK8cxhj9rDH+EgrVDO9M4wKKLadGzYUZRCC3IlGt
zD/ZksnGnahjQX+C9/2QeqPfK6GJkMZm26uIX7E3B99OL0ld6MLcrRWbo9XJCnVEOaGiiep+lMSO
hFZNji2o+na2uvLsqnMZfN53CA4eWaa+n+7D8Xc8KCfjmDF92xdG5RNuyKDfNf4buMCbtNl8mcmy
FQgqzZyKDYngFju8qmusQl8LbsU2kJTby8TIVd9eBNUAqT9GsNH+CbAbwr7qCfKJS24/Pkjcaq3g
DQY/kjsq90ii2ZUXaN6nzlFUo7KgaAoR8ZO4afk1p0GjdiX4SIrJskeT+mIM3bmNI3ziNFQmppQT
I66JIMrVLGlBWUolpi6/wXfEHe+OtfSrsVJqhNnlP/C6uBMDHAlFI1Pe/EdCpIyb5UGqX90D4SYq
NETI146NqNP4ECLYAOY0BgV2RuJfuY36UyAv+iN/o/kyFl0Fyt5NPK6vzOilC5GTumWngeELcRyW
i8emTvR1bWS0cUGOs5Ypj8apffmtetj3xYMhJcvYO5HuFA4AZTnBEOWv4wCoufUYpUXEcAki9lBP
OigYizs/DmHw4LB7zIb+D0JVI8ztK6qJk+5XeV3sqOuET43w49FE1rxrTJ+T5gPzUaTBLwvKOywY
6h/bAujFrsJ1Fmjq0oZ/qI7MIAbzN4UsdHTCUsm6t/DaUyRPqJJBJylrIN4btSzVHS+bBSgHeJfn
Ifhvp+aTeDvUWtJ2m6eEo+z8Xb7NZhGZezhn0XMV3pMO8XncudCabrofZcYHHvt3Gk9tHvQrSa0P
Dp/oBbQT66+mJlOnKNgfovml2R/Lr71W4tNqtFWJLOEbzWonXROYsWHGE5j22sAWiV5TnbrfOzxr
Um8GMYY337t2Q4hSluUwyxTvuirJO1b0R2AE6mYC0VMLIQXC1vj600jUMlNp2n+9SdncqVzNCMVx
97/i5n94cWkVZiMG0aT5dNabo4Qv0zasY2s0F6EhEyZ+xkoORB/l7ny2pS9KYidTlcSYvqLoIl1m
YY/Zl6opTGAMVQJEIFG4Z9pCBETV/mktU/gZVSJvSXDqDvXlRW6LmJiJ59AvIyTlk4WcZ+hL16Zt
6t/OS6eXgahgbDxgWjmicKqkrmZUIEnR11ZRiV9Lw7FbW7o4PbVfnBVY0615dIiGYWNv1I1ASg12
hWHtehOyS9U265gH9jzEJDa6q3dmdjpURxKhKoJvPwN/z9yjfrSP/BQkiAZuEzrxi6l6oby/umuG
k3J4fqrziWEhxCO/8FPPgMJHCce4VFpHHNbhuRG9/LKrx4DMe/czasTJ2GjJdhIx5X2vLO/dI728
rrPkK0h9UhXecADqE/r1gNtbCLXehRJRx7ZISlYONdD+ugJ4b25eUCoCcCAcDshwz4c9ixCnY4uw
KVkKtk4+enozNcwcJoYBABCbNiMmbAGyzprm8LbZVfxcyykjM++SFQStGJEtNVc6M+X5EOoTnzUF
M5ZgnabOJ/VQwgZkPzZ77sVaeoM6u8m/lRx4X6FydzGrJK8OTkvtqvWmlpN7+Ew3lAO3ybv/q9fd
JlqzMx7Fdfv3U1Z1+jnaYU3kmpuuH3+KQV+Zbe5OmfG2S4qf8h85O3ZHtzw8CIGJYySZoASsJqy9
4TF2e72ijXHljw4W5+qH2brAwS+Zx0VjvWik1j70TsHEzTxTsKc7QZWl9hdzvIz5mNg3lw6rHJTL
shr2wzw3yVZcHLuHeg7m658I0cL1UUPB8mJMPD7niEUyaZE/nYMHeOIH2bN7O5qSzf1yil9kY9HQ
6/g7RA5VbXL78BZrwtD80r5a/5IMK7G6FbqNzsj72zqHM7y2DI73P7b2Iuyr8+ShmfBbM9A6Vr/i
0Etj8ayFJBPa5i9NKyMsywmgJ8ox+pK/njzHpSWm0TZhFuZTF27+EQi4H8E2yoqCv31MmM7incPE
PUpxB2QoERCqMDJAwKaK1I8upB7EbKfmL/GSpprliXRnNFujyKDxnoI/fi2md//uBR8prNnX+6Nu
4dwKtCfx0NwZSZswfcXNaWsSkm1Md7cSvpk9asF09045yEUIHEvCeFDJiBCITrIXE2tdjY1696nY
v6J33+Hz5p/3XDvWknlzxphSPmTgLuSmBCfZnocxjHW5GmA0bs673Wl6MI+BF4T//x42DOqlRP5Z
PS1+oi7s286CXe/VnfCsjqma2uHSPFYNfX0ohiPtUesmEITS5pXkJnqCEHVHVUfW4rFtFzUZ4yQV
gX4bwpOrokhsUnL5QATZKFAbX+rCNB0gKOEYrsMF03X8vhO6L7ekT91kIzi4xy7p3jKnz9et68BL
49H8cHBFLoHR35zABBQgDWvcnlMU63bE7tx/WZyqTO1V8lAGvSVbH/QvhXWYGf7+9L3dvaUrukWN
SuYGELGaK0zGER+cWBE/8QpMbeakhBB9yf7eMSL5Ymj0IZF1qDzql5ZXC6b90U+y9Q4acrw9IL9+
+IQBsR4hsGbqCGGUfqFEdUJNxJG+vm2Qc6CcAC4IjsszYOLdmneNdK17mwYzjnvxLubAeQQyqLTD
1aqQ6nfEurE3V+uymTosYS1rZkYJw9DbMvhV3udgYgwIqV3DywhQP/9WcRXUHVki4c3KZoeAgkpQ
VUS+ligPrrVPvqYHXXydJpa61bQ04LALzLwm5hog2GKUmuRpG8u/aPqHJ7QB5BQtTMQEKDKbwnLT
qw8gQf2TR2kBxj79LDzyw0Cal5V4fAUrqKePbOu2C038pmKQF6gBipBULd5DIgZY9QGUtlopfyS2
/go0fFgL6UPEN/0UYd4M6KHLlv64419i4ab8VP+lVTxJtQH3p7V4VIUQ207RTFuh88OV4z2DCSsI
nl4EarzW/SzZB0TxO/95c+K5pajG3oRH4L0tNqz+yNJ88Ws6l0oEAN0/DGewSQIssK/Cmz686Yr+
/5Bg1NQS77YzaEs3KbtbK7PdgJht97xflcNZKXUClaQs6s4sAYbNMpnVvKWvVnCqeCAYVF1i5KZB
MrgCsPgKkEghcevuZlG/k4tiOBXdjAi8DEUbHle+6uoiY6t9CWD9UXzWa7VD9rwIQK6+IoGtfZYJ
48Xjpwq4FCEK12JieoL4OMhKpLDu6ufc3x5uOcZFMqE5Jd7dfqmgM9KuFJ3F3WYZbBYA7YSrCGcY
wbEppBQJ7q5rt6bd5Kt8Mo+STJ6XRTUszf9Y9GxiEThSynerq2WD/NUjPBoT7O+9jM3RPZUTLLS3
oHn7g6CnUJoF6zfSF8voPoif7aesLh5Q4sr2EMx08h7R44fSUOsNPfI896QhFwpjkVplQQZXrMv9
YRe1QRpelTopr+2mFOaRcM6TNllGVszaNMa1iPrhL1ppEwOe4fySFQKsJGT4lzrsc8ffSyjOpf9P
DnUTWNzxFvTSR18ha2uXPN2auMEAEkKnfO/Pl8ez/4Wep65d8BPv9bs4C7/Pt3whLsI+Eg31oqQ1
jxcYpsb17yxKi2kX57teszYmKdMnbaCXVuTLyRw4PClt11hK5Dul9kDCbGMlDPr9jE1hrIBzroSC
JPsWC/1eVn9A7l3qsoS/sOzida3JB5P6JJlOEwO1mZsAL1jrTbPSYhCPrdxoEat5ZkYWgkEGCQxx
Od1xzfXXUZP597xvoRRCLFaPNvaph/6qcLLVMXfOPXfvTo9/V/AlWhBNkrcmrqYEPO2N5rAJGdPX
3pEkCJdSL1rT/Fa+b80Z2/khXPOXO0KJETc98zUBqgSokmo85e/WKeok/rq9E5WkN7g+S1i43uv4
kzZncQ8qjKCNOyoY3tbdZ/ThbmGj4vBA6rqAwUR30WSCUPFWD2YjRGVdwmPcsz3tPZOxuJcxQWG8
qXok+DLAFGdotgKb0JmOdiEBGyrAyUwDMFZxI7Ur3EyaMMirQKRrjKRS+84eY0Y4EWqmkJifluYW
IfYsr3sHzKLVTcJX4j+n1vWMKYwg2W+gX4P3wpOJiLKzzTBcc/I+5q301IvI6RWJ49kuZ840U0/t
8oVSGRfpINk4LSDhsJYhxRRl6xbljmPbOwMotEfmLCQ1GMsdfGCcHTe82nBRhJAdO97WhRk+/TgV
hPg1Vldiu7HLACC4gHUzY54GtsZH2CM9qh5cwEapBo0UwF11hYcybFIavB9/VB3iCCHix/DmatBP
iFac/UEhoPsD1PVE+go/RlPGEd1aHyGRFajma56E7c5DkLGPvJ6Lm49JjDB63OUDEWjMx3ZQhYr4
3u4IoLK9RX8KOKiBEdMOZTt7Rb4TW0l4CjnIwd/+UFtSbuS3P1b6NJPGIABijusmbLOdgGfYM6AK
B9YxyalTJYDD6p67q1Hk7ry5VpG0dbLwZx3o/2+8jkLrxFh7lsKBoTOETMTX7GKfl0JzKUGRuYv/
M9LAS+9nCTgrmQwjlaprtaLHRTHRZbgB4WriwFh0YKqMddaNrtGlCL4IZcWn5ciNHODAp7i/QY/x
k7tc0cIdrPTrv8zvbbZ2Mt+VNcCK9VqaVc++tr34S6bpbnnbbv6Rxshc8MDc5FdpUTI7HdmdxG4d
COkq1cst6D5al1iPcVRfqGGEZe53K+XGWZhMwdJ8vJAT606laP93HDNrYtI7gjChJ0FeFN5jaWIa
2dA55KhwnxT0/uiaI6/I5cM4qmNJbHKgA0KWuoErtS5n2UvKuTQu2FXKEvlVcfjFFF0SLuiwzwsm
TsYyeDiKHJcKikUEymMCIYC7Na/S68Xylm2jlu8ncJSWPS5BQ0Y3emFS1R7D7DqXNKPyfR9uYqYR
Wd3Sk9mQ8YcmqNab7dQvu4FaCAI7Prg0E05vQEqxRfaYTHTYzVKXBcpNWJFyRSo/RNtHKdUcP1lR
zKfbYM3VUOGWwHQV2Xn71MIVQdiqlIzMi7/o1YFpNyqw9QMg519u0SZMF4Ayq0JXZS3fI3fk28vu
WwPZrfU7mPP/ANgdIXGiu+g3DTlfqziOOvK3K2WKm83BA+tlWKDzxSieNX+E54OJ1nD0ZRf6jm3J
nAKl970zptxAjn599ykeeFIKOhm7MV8XLJnIXnLGqMffW79sdvnYBksIlaiL54nl2olQLx6sTCLb
1qj2OrLt/vsORQX2aQATwup3MtLsd71RATLd7Ob4wtY2UCa9m+caDVxIAlbrJimtb5GqS1ahk0Yd
KVUw7IEXhKKtZptZWOtmTXzYgv5lKsnQ1CHj/zQ0PHBkmHQTCVwzUAVlfOzipvQkEgsFtzhuFKWK
L4DWr0x7rDCf+ftQG32x3GpiNpyh7lwyCRopbYqKY8r5t+Zy4iKd5LWxVFO1oq21EdBqF6euCbuV
fk5jrxl04rdBV+GjjbPYD6M+BvOlMUmVYOQsf7+DM9vQ2q0BNSsHaBTArK2cAO6s1AgXmWjpZ26w
mvjQdajP3dnq1Xmmhik4tNi9vYcF8WwerP2c+Hm1mYR4xjndonzw3JMru7zZJC3oirWR36Lik6Cz
/azyxApntcgJTQPR0S+dtnNzUwvwsBjyHbAQxPbjBMVpNwqV89LsurgMVJsmlDUmh2Ndjv2GvTHx
AyTc56CzPpdy0YqbtaN4na+jGi5repMTQoMsnUanUBEv0GJFoLvYfQDHjNH3acNNwE1O+LGzhvZ9
SVJHw0sPsYjFUC8oxJ41vUXXNTAOXDOokrRTlbNX/52mtxuv/S1BtygxRk2OfWix8X9bXp7QV8tC
DFJic7bhw6mQaHwCfLkx4WMbjRQfbQHwMQkJuN3DtbdA7lc3TtqrP+Yj0NkgJul60HmLrVZ4PBLw
C3tMYs6fqdWEQODY6lawNbLkURhHiWNK70X9pmgUSdW89G+JoTkHxnQ13ub21hYZyUo+0OXaXXk6
rzkZTCNwxeOiutf/0wH9GdhO05K5dsHPLcw0AX72NSVa1fN2vEJ+oAv+GZt25RSUPnRuFB7jlgeD
5Ca5qjkLUNNAHoFQBzkiUWYT3lQ2AnPffcNXAxgO02zHDQZTYT8SgDHcUs0wBhqdJvFbUO2upIIP
q0VeuVv3ciaGledQ2of5KH1kZVRYeZcvJM0ougZO3OAeYyeZ4sjgOZhb3/n8Z5JEReTEy6mTQq17
N5daC/zZYgMX6jZ2GG5l1/sFb+ifTsZG2voJKUJ1ZJuJskkjLttnFLv//VRhqgUpeUIezE3yztcZ
LFM2KMIeSSBjfsz6kB/hadBo5sMDdKfVeF9+byvVHLTvD8HZYiUOL3Yoj/TT3tVVhekj2iIvXQkH
nTr0+7oVaj3zBzBcFsjANmCXYJDAGwOL+7iRDB4r36yDgVWnvK3X64pMRmTi3wAtpPHDdGrYr+VA
/Zy0VE1DdOxz4n6P1o1g3vKP/niJFMu47FDacCwaqvsDqbjxKHwasAOPp5lm2wV5Iw0Yqu3DK7Gn
uq55drEIs3Vi6PhtEOfRgmnMkJYpRdS7c3vPUROZ9C85YilCxgAXOy3+xGntZ6JM7KrBQbITUvjJ
fjQfOZ+tbsAn36tPVlOfGHmwGTneKmGteropQQ2MvD3sTC7H9IsPn99MEybY2JLTESDTgA1XXcY5
/65EDAJ/8n454SWRkV0I8PqBd8p1TO1QfIZsW5CQdpa56Ksz7WDFXT5Ga5CAyf78Cruj7GCbVQ4G
R5WxTG/E6A8Kt611gY9cd/GdpqVI57w4KDe+GyOuQkYzXr9e2V1poRkBkCgLJFKJ8Ij+TmzPsf1r
jibbBObXe+fmtyTkJ5JUirO8Gay6RLJJVO6VEP3cC/TAsq507MrF1ePD/mAV0+5idrRfzRIK69LJ
efdcUD8VYDLCsP2xdPDwtzlsS/Aw+RS3NNx2/2poZu8QpylXPO/hKpQHU2H+PRAAP+mIBSuhRclt
hVx8YlQlXQAYXnPU9rrcQLts/jt2idt3oWnLytZXrAwGq/hZhOuctYj4qBmOCZwFhurOzv3nadcq
+jJR3HOT1PFh+Ac9X+fd4NoLvo5RBuOrKM4am6FyGeqWLw8iAKWSTPlBihXEzogRVJFcoSZo8y7N
ArJGnZ0eVuyjAOCbdbVzZcvVO9qUjpOX1s7hFeAq+Kym1FUKRSKWVtBIWS1iZTChKOgjy+CDWi8b
n1pQfwzozD5/mdGD4ReBabe+yFwT69L7GTi7BB8LhHH7avqx4g+xqJ5eejoc2S0djFGPeNY2YhjV
G03Kn9o1l4cJBVjfXVfH62HLSBM7BRWcw4v/W5ebxWZI1tIyTbaJYtMs6NvmAmrLFSh+i+TQ/c4j
Bmt98mD9fA6g0YjljkxZlb+i8EjCw5K2sV3nlO9M/qpGCZnae8ZDWw4SciW2i8u3jnsTuMJe46Lr
d7678t4H/KvVkIIgoyQMkAQPTfEdLlbQR2TzNuoTNHCbZbaCWRJNvg85Ecb3sL0mosck297OCZ/m
Tz0G3paCmWXIm4TUnabZ9/wh9P4Ar8+1oR4xyh44PG1+QxAdDlA/IoJqIm00Gk72UnRj+pLULZ9U
gJjR4nz1CBmw0WCFrsN1Y3EUmuvAVaAPsuu/Q7TTxFSnxdMb4Vv0CkpmI6GUOm/C+AO5O9BObTx1
dL0esiK9kkDr6FPDwcp7gViqaUjl/oRQgbAakYs/7GWwspVLjQgrb1hIt9AxBau75k03TqxRBPTZ
Ms/XEEL4emox3VoM5BfrlOF1dVV2FSscKTBss6WNtFSsF1/VBXufXWKXgSgVe8PaR8mKZ5CiyJhR
Bec8Ebk+G6fYvc0IpiZKwJet53MJT5fVDnYHjwR0Unl5jwAsVZ/3WVOrbvHmAYqcvUfOJnfFlTyx
X/Blgo/nI6E1rgaXlW/nZoJhZV2gOd3jjzyIYSo43LdlsSrK67H1hbzvyPDcf+8m53Lv4fxixGAk
F60iNPmrpic5tNDFG/UNMNUkyJlXfkuEkZm5l1y01YEygIgyjVUbNME/Wa/wkv/rt72weMd/wyMm
g/UVb+0I/E7Ki65Q/OC2iwAEmnchkf27t0IJ068K57zEEK3+fTzTb8brMeiP5UD9uxdbWBslugQK
YUSk/Qga+OzjKa6kavDZ9eWU6SC8J7L/iDYOLb3sm9VoMryrAQLCGDgH2hB10dTY2wRFxrzPjCay
tpw1TKmaYQQEIQy/lWKniyDscOaJpEo7eV3oPqGKN72Ls3lYcu1RSh3L2BwJYPy2Kp2G2gmq8nQY
XDteOGAmffOKGjCpNf8e+9mwnnwDlPHQDnYLFpKstWZDlR4vqwdG1N9SncFy9arnuDPvCungglTp
JMiY9++IaeUrreoFkufD+t0bkUhqIgz8l8C8E8fT8GlqljTPMxqVtUG6kiIJP8me0Yc6647Buobx
f7YBW1C7/lwTZeWahhfKc0Y7K8cJG8/9wEe3vp8eD3oOUkihkPkhMK/jaiLsrkHppITPGdSEK6so
7SLNrC2p/ncrmE9UI6GWxQ4Ow6HkoaUVq/QvIpKEYRdQteXjD1MjpwGSrfkE4pLrrcAIc3kMceYa
t2zjoEg62rxNaT1fPsun/wdsW3qWAOkl4mV17VBzph1qKJpvAaUpBnMNbYh/o6rAsNMKDhNJyLwy
qxwhFF2LeES0lmFgY0ju8+vhEBAKXkRkJYRGDmy+fHjqpcU66USegtfiZqzTslSGEsXe/jGwQ4vL
F8IJ7Xs11I0+FXjhwhNOBgthaUCifTJC1D4+SdJkf5c2Di6Jisq1eHV4PWgMZGOGGJMjURrG2kSG
3XkHyiKoFzj08uXiGOhe3IoiWOte5+2Ros1dHhDUo0pE9FMylvI2GkqBIbg+gJNB+0Bq8fzwIh7O
xx/EFJjmThNb12Kf9k4wgd8JKznnrKHIx4AA6Sv69L8hmmyKbVdb1udFKMnrO4W36EUDGyd34iX0
Q5UWw+9iiREYHcCbuxBTmeCyxukReNtLM1lHQkWwr+J5Q2T9qrZxx+tXpYY/K1WWqERwm9y4V7OF
GnkBZtzas7R+D2EoalnLoLG9XIOg0PpAnFLTWo3C0K251tUOvja+UW/zyOePX3VqYp7TXocffoHp
81837pdwrEYIU+Roib29Se0HH+svu4PcXxld2WJQnU7mWobJNEIAkjEU8//TBocFLTs6JmwJttuV
6DWfhjwokCM9rT+neVX+5OILYkRMBQKeMytH5WnmeJPiIWP4zMmDmTQz/YH3anG/Ud2cDUBxkFpo
4c+SK2DFjfR1kpvNqL9qZXCt6cTuk642dgCBqlu4m2HOQImXqV9c6g9neKhFYmxksbsqP1lva90c
Vpxq69Pac/IRkUn8VTxW7E0vzIxGhFpme7AWAs/O34VcsENcNNetx8o9YFHrEWjGwr84r8ImBj2F
t9IgAFyPfA668C/U9y+EF/DpxTJE1BvF2u5AAsVY8Q0FfTmjWKHM+7bA903HaVmFeRLPAU+jMGvo
H8EuISS66w8rPzVK54XTxiYYxBncVeGn5B9/YrPgM/GrLVET6tnrIw5ExkMCfgrdh94vPb/AWJgU
f+ifl36w5kexfxgP5YMj/rmFrMOwDOO+kQsdqbwouCP0Ok5/2ucxKzXFuEeUOFrDgaBdUqQvht9I
0i9gePDGcxQg52J1PuhxaaH2OTNDiPw5MRWn8qIogu/B9FBnHu+HrkhbiztEgjBc1XXINF59P/ty
LPZTJmBli4RrEjDW3e9ICxuWA0fYntS4Z5rGHwybtJ77fdfXNHkoiuQyRvrO1JIQI8iiSuk9dyd2
U0TP4vpVK40lr4jjX8Jl+es+CvtYADy6irZksU9Ofx6WDbYylVZKGLiNsZAXFTNP01p0pDWqj5nA
WAOsslGIZ0NUmB+/Ng6oqP82Mgi+SNnyq1in9FygJCS8zw5jqRbi+HM5YmLGW0vxcWF5zOObPEsH
qyjNsD7mN+JBcGgQ4+nY2G564h0TjYAeQIQUStF4H+omP8l4s3txEjafPGETw48rtPbbO96C/oD4
ZXjs39Q5xDgaMYXu1q6ZFKFp3qeytTfBgctAvQwkLD1jEyFk9m2Vl4I5OHKjEgJrQRiSVtdMogy0
gmHwH/kAKWd4p6WrjvZ9TxyPcbyHkNW+4cozeA86abjAUOHSQk/F0eeFE4SQ1nAG63QLL+MoaDqJ
lOlSAODnYTBcrrJIVSzEO2XcBfSDVCXAoqQWIyFS4RZNLUGDzqz8yEvCSyGHTGhZJ625OEDBGfbO
VGnGZYxV/UhKrKxj0PW5q8xwKQE6f65SbDo4fElALxIaGv9q4mhKNYjp7grfO7E0xAncbixeRMft
4uG2G1dzAKMfJTSoe1aGY4ugDdtRGCUtbnljoSzsjQLGTKe/H3GcNMDTHUHkZQQK3JaSNm1Vxj8D
v7yp3w7op2AxwXLaeNa2j+CAr3dJWCEwUsGW0pjH4R0bP5+jHBWgWSzeJ5iurJgoEAk1r95myds+
lDXyWm4P7/CtaJxJU9dd0brAtmHMcbWkssmzxhzKRnWGc+IeeslpfDCz4RSSUi+juwVygafsZ3nM
XhhNH9+jbRR8Vt7hjD1n1jnyL7BM5JXwBCRn9ItoDRFM2+QChZGuESJDnSMKqb09SqEJ0m1XCfYA
Fet+IMcLvgXJtJRcbH/w6dloVKb6yXqCjwhXgj7bdcbzL6iy3tEiL0ZfQcQlBtuv4NrYwPO1ATpE
dS/PfdQ/pU4Cgkkvl42NiHbgRzGgOM/ihhVFxom5ZpgNQI3PbzR6kEle1h5OZLnypJ/bqfsJ09Jn
fxAA4DD9gztlpeWeAbqvgPzwWib24cLpiz/n+pilL0RSGau6QRNI3BuSacmtY/j/276d/9JJk4Te
Zjb3W0L0/nkJSv0WvRsUCejuf8LXo2w+ApBOwbQc2l/yQvd+SfWOFYQkCfMm6QZTdhpU3RJHQGy7
Ka1XF01mdDKgkkgfLB+orx1LrAbu+4k98UAjMHr9PXSZXppx1wfsGO+MzAn/SMc4Mn+93bVwVq3J
YAWgsDWCiz2JbvkyzTPPhQ0O0333yYx81PwhcPJQZbSiUhElgDOOImPCg/f9LuPoZlNBUP0DlJBQ
QspjtInOXrodpbKlbhlInFsBe7C94OmA6LtY7lhuMB+jEX6Qb/EDQlMElrCZaj7frd7E8BNTDZw/
Hs+FqUL32yPgZMQjSICvjEV8v2As91EFQlhuowME7TU6euj3cdKAXmSocXjcKhzs37oLIPkQ94EI
fJv/CuZGcg8M0oEmJ7BHdqk2qHJvfCSxEuxP3XHu8Lyzfx+ivsYueEBTfEow01YfNOZ47yGcL2uw
dSnSlnKebAmJrIhfVHLkidtTlQr3jE8eP9RqxhAzvUTddXUSS4ZjWid99r0iC/WxHGenhxHgoyjA
EVifb+1cR/ofekt9f6D8W0VSYVC1ZglaSYpz2zLm3+IQQgzk+b8/me8jWlZ0CK4lGPszklp37q92
HWqkbT34heHKG2g/irWuf3CJOgKHf5eM+1/jqA5K5N2mCC5rB1p4x87fAVkRTkMDAayGJKrGf8yD
gv1zKtl7nhPLW8TSHHqgyk7w1n4j1R99MK9cVkGmA0usr9VIY7nc/mExHckCvNDl7Gj7H92IrYym
WRcCwMpsJKW8i7boCS1TW7n0CFwJ4UDjZ3quhbJ5u+Twl29Ezm6gErY9SSJdhVdyfzT4gXEG9PbU
KlT+LkQvtUoDEIamzQq0IGwztkxePASP311kwHy3kMc/Vvw+6ycprJ1ngjGduL9/ppvaVpHPWXMo
9Xk0lunPLeFX1RjFmZA2iDMfZ4CS3NMnmJZnlhxf1fcBwGDZFUqrPz3/0qCel7Gp9Hmj5tVGxIH7
A95SpOJC1UdSTWdYJfTSyoaGr2bLKXw3H+mlicT+gbX8Yh7kIbHxxaS1D7S71+z1Ae8jKiKtiEUJ
VSD9kEZ6K3b451iAaMRM7PYJ2u18W5EqGBCtQSt9cTX5lVg39qCLGdmySCLSD/fH3smj1JkDa8k1
BWFyaCH/9q5v4ghOlAyTOdK2s1I3bvfbs+RxYpopFejoxwaTCcx9CygvTgpxvW6vz+y8KoNdDp5+
qXO0SgxVyYRlcczWVK8gopPVJsZ51tGfG144b86jsAx+EuHpdOJYJ/rBso9lg/I1wA3ZOsUZWKdF
NiqqquNc0svvWLUhZO7s46j7UkYt3AKYWpBCcARW//zF3LbG5zbDZ6XUkB73exhxVT2WHKloCew2
YsgFxZ/l+7L8bwHDBvl3gQaOI8e5IhePyhqAC3jKPZz24dI20jNIz0vw/AS4xrRVjvMXR3bqC02P
gHCGA/ErT87jQPQs39wKUU9rxJSz95Jzl8LIGGmKPaYsg7XKEMCnFg9FH4SOvvdI+Xk/Sval7hLx
RYueTDjL/mVoMeENZ0AUEfRS3gNulK8TYSiN75k2CTDzdM7Gv/vs9VdmnokLUbCNDb7o5dWsnOiB
QDpjk8I3ijpNHN6d2eax64AOWiqh74NoyqXRtthjJ4I7kL/YJYs9ceT0kVxQEWFb1Liroz9HV5QA
PK5AayQbtsRG+ypgZvobREVM+/vin/lGUNwU97Ydpy6JVXS2lWWJ7mMKawd3j6ttqu/lJwbRUkl/
Qo+TTaRZcL9CPjoEvXSFqxvZFLoV3cKoop4zhYLzn5saUD0SWkx/Q5iBCBYZ2SqjKbV6g9rT0SYg
BT4XKyHdUfO5EhB5A95gmU7g8zDzYd2aC59YQeR4Od9PCae1qoyKcQqObOAHAnym1uuyuEjjq3PS
2poihlCqxB/6vPyUOyLBjsrpJmLws9upa50M4c9jbCOMDYYnhc12aqNEQqY//GbbeQfLt+dCQlG8
QoC0CXvUN6RAGxP5Ui+/cBdmRBUK8ps3OfkBJ5f6DIMSWKqqf9WM2y18VnLMIOlGddegmnLt98hb
kQU8nD4RzshLvOcXCm49iFKyoomN2botQtoijC3ZeqyIJngyXHf+rcFOel5rDieQWtcoJvZoNF0V
Q1supAW/qKITCWsKk2M0Akm89BfCfhHQPUP0t+WRKWs0j9CtkN5Q4UjmI58RABLQW8Sqt8FGNVBN
dreXv3Zkkz/KNVqeiGC56SZLdB3WtW6L4UTEwa0XAY6tDCZnRCsG/JLRT30jydg07H+/o2JAOGTx
GpGhEQJw+xPiMWHPS06ITMmEfyaOCWheWk+vVbNC1l56RUfrK3V0j70tc4ZY0LUBxAI0sTweIK0p
2FVBXuzPs0sDEecy9pmmHuYXVYQvjzvx1CKzY2OLOJ4wNHdKjSZEV5MwxsUCggyxhmyFZVR8A2qE
WXR5eVmoUnaDOCrs1/a1YNd09qN6X1RazmH+1Fw3eebZNSEU4zuxtYdBs30lY3GNg+Yb3tkbXVig
gcxfciG+mQDYd8vGaDIn07LFMeWckphJN5/5eLvYq/7nvkX/cshUUP0U3jlIAGOcmJF2b0apcElz
RhOU30gRy+Wl+i13hWjasryoH+nHjZPBVPLYGWKXLah23pAdg7LU7dhJuojoVsnxZveJEGngI8dD
Gq0qhYT7H5QNYaJ5Kk+IgagsnHEpyo8XDviOghrCPcFgwyzyaQl8XZkyOFXTXRKnaz992Ybceah9
5xwOvAX72oIoPJmDOFLgNpByt3tPNF2GaycRUcUnCrEZ6ns/EV7cby/iRP8YBoGyPJbmY06ekwL2
/IXiHwzmY5qunfE2r9HDtQQFazXRrvxUjatNwaRlDQqND1H3NtWi89s8n7RQ33y5cpP45NO/nlrK
kXO1Ihk2XlkWTNVBiY2R4Doz2sT9Ae3tghjymm/kytc0xHGa2ie1NALlnqDDS8h0qnFkneRFBgSs
FaZM71uJoKHGm2F41aYOM19VZyadRGbICrU9+uhU8BCOsK7t+Xw+UWyJszbJQTZyAOQUyQ+tIHTq
BGwxvb2uG4Js4VPOC6o0Xv58ThEEeJ5Fke12LUalLLAZv1lRuh6kX/kAiX5MUAnRU1uRq8IJ1Sp8
YhIwohjXAMmVFQRzK4mKCCsejFb/LawysB1Y/TyI7SAOA8m3JBSxlAugHs6ybHBq4UVsfaqtpph2
SCgiLZmPHQHIs9c8DnlZfx0yVtDaydZGNcW7b4+trKGyS0fMwgvtuefQwdQqBoO3lBkC/vl46Csu
JsgEnYzg9K9HUBzRXsYO9NC7/hGKBjavNo9v5q6ixb3VuYTb4YqOZtLDKBFYApxj+PydRFrQVeMz
zrHukVC83Di4XKijbZb42cmHadG7uKTnusjI1HGZ4yjx0w9sfWG78CIGmSLDAM4IScIhnAuYxU/e
Qz0vCf5UZDBcz0Xqy0V3200MdraJpvKXrPZK5erWV56fIonGkPXh0C19PlE0SP7ifnkoPY3i0JF1
c4ES4gBBlqbj5JPoVJQRcZhy5Tl37g3tGKi3BJazoIxfTcTI/aRWkCuzzHcwN7E5n7thoF4r2YAO
N39sOR86FW7cUcSwPjsAtFPA5QuHvtTMnhSN1fZ7YJ4nHqlIPPRkm2AE7E9hHRo5Q+ymmFnAHxbB
Kk13EZOmt6BoIWjwlluP+G1lXfhqRpIHNXO/6NAoovelafi3Haxq+xH/+QnFnyJmxyZ0kVv48Acx
3UJugcNMCmXAS6vmscAY22c1p6IahnItsmOjCGnWybjJo0PSv1knOLw8FxTc4rldNCR5345HbXnP
HTks6BWtoniebOF6F0U1pou8Tzp+WainumcQTIoO9RLsVgU414eHGIdS2HF8x35WAuAof7nAjU8W
Jt0gW1aD0BSTZ+wDWlhyYqdMaRGbg6E0wGRHNUyBp9cS5X7KjCtC6pxjSWQOaOBmidkjbyMvL9KU
5Z5kSjpEV3HdJxkMChQltuGRMoi72r6F/f3EWm9m4MMGWs4O/RR6c6FGWzkT7jsUHF4HQzBbEqWO
HPVVWnSculWJuVPiUyGlOO9RBqNJr3hX94d3gAhvqSDdJ0IhqRT1FdF2etezrmMqZlb5S9uiYdgq
fVTMejzmDfpeAx4dec17Y7VuUHt3b28pU2riNYdmTRkQ8+mByTiLk3DHi8vvcAvhHNuEXFlCayjg
vaLFZxgxY24ciK2rJRJG6Ujxb0Cv18KPcm7S4jZMqwmBMuZJ4lW7dsELU9pnhFFetLL/CjAbTx0Y
OCMuTB1oC4lFtxa9qYkUAfQbM2vv0fqcD3d7a1PX29F9OZJCqljHPPK+SLnR0+1VDqGMH+ZO/an7
Jmn+VavAjMz+huwjTlRa5OrbFJP2fZOF9eeEIY5ZHhxwhP060aadFr5wWYP8OiloKM3PTqKYmT0j
Y8OctR7oyzpLmk+HTBRsM/Qdldm1AyvDV6cyyS8hJMThW9Rvu0QDZAzZdE2xYHDYSc3D/4pCwwmE
1R5BwOo947YooBZYGBPYyIGH7lN0Lf6NSj5//Uwqd/6f18kjyiTuOpjz0O1l9W+exw5aOCR1dM/H
AZzuQhik7dKoHIZCs4UkCbjroyKsD7NukokN00gkdvHSTx91v3Inck+52VtRdjQqeWx8P2+8pJnP
2GRS6+Nr59S8UshJV+tNMaGTPjunopibpwZxEgVimwwh7sRLKgGAl220rGHIumhvtKSjVkRcD0R2
u4oEE60IzBNR1oh5B5oUD3X7gSh4j/spcD4wgyj3vNSFJ8Arlilr7cjhwt6kxawk7Li896f6Ymdl
08SSv1wXUDqfq6HtWM9RVbRRQxSleEamxTQPYhQl6vSffPjMZ9lyF57DDrHtHmWq2VJTgcw2x5Pj
Q3D2ZAlzsyH8OKWzs2dBJw0NRlxD4Apw1/7l75xn0hR4KRpY5vhuB1unVr7p6e4ZleReiKl6e1By
7Noq+qa9TpI8H5cSoPwozBxSOHIzpPU1D1NdbWsFByEwa1LkKtpES1R56xE6lQDORUBfOunMJuW7
mLAxpvlUK0pfB7piko24IbUGenrjgLjUwz6bu/obUWpL/eycyV5EA63xtCSnzsfyBBumu9xfSTWg
XutbwzlBZcvq9wau2UmH89e5XwzM/K5XOx1DktzU8JWbYaC9tPoPEy1zH0foPtLHEWM2eOcXFs4i
MWok5sSntOrz6wnoorqillYswJkg2aqq/Y39sIb9GEawKAuuie4rCK8cAQvul7LSn0FXeF95Q2Vg
idPufSY/O1AHPf8bOFMnNn6CWecubxQRmuAPpdGTAyXbP77p6YQ9+s4qZPMtJGwFiZqJpNEjyQVZ
mJrd45C3O6MRjzJrWM/s5feVx0Hr07nHctgwFXicz0eNf6R5Geq8GUDmk/ZBbKCLcfGOcZjJQCt+
v8LkYfIIG+YKCV7N2DqfzYLRxuSXG9RMg77YLaQFJzvt4czQS/ubm0UeeLG3sQMtCPp0yK611wkQ
ZIMZ41mrKftxueCsmiyW9rEz10QFGV5TFMVzen77olpdjIh+bElAHcXZDf1qcqwrExUrK7AzsCqB
lSNP9Z4V+EQHxpOjvthL9jD3RBxUtm//4c58mujyaKV3fwZVBXkIFarjuAnlPYTzsAqvDyqLo5TH
NRCDOutgq4fh8OmYzuI6QrT/jp2MayvJcViIysGyn3HKyX22O73Qr56/YCV2z8PTcfRqoDnX02dG
SQICqyglVCxeJRBqRJavozUS1E5cQtfAz35I4xVPrfanq1ooy531qzSsX+MtROYuoxDFDeqqmIB3
ILQewDL6RVuTDeIp7ksPhhDxi2jefgFNa06XMbrHvm2eCDG6E1CjOKgm8zyVCr+uIFwix3hBPdrd
hh7KQl4oPS9PF3jmAUZgTVCojeoC4AnL/ky0phsfZzu60NiQs3nI/i8xMUmNa/+b1GvnjXGGlo1v
YeKzGgrWrPFKWh04IhK090TPo/RsDvYtjIhIUwbA4kHmdDIFe357Tb3uiWTYM731A3IdoGR6/g/4
yKHKmP1jgYcmXxu1xdanU2UCxUImjU+EcpVBnojvJKYwzpZ+wSzeaLJy+s9J7o1K/k/Z9UiOig3M
MN/a8t0US/Stmz59kU/tcx3B+1RJHVonI0pKxU3zCPq4126DBzfh81rqmqroHxx0RRnrDIK4wlI2
kz1KjSc0b0hmsDccCOS0KuZh4jesJyWvlX9Vn9iHGqpPcXxpasUlv/tyY6fl9M8qOOueAKH8wlWn
Pr2g8C5YhaSUvPmaq9OrdWo/gGI4/KbkC3V9xIchDYIHtH90gQ49BytqonCKABYW2D+5lhU8MuwB
EgxIHAZj56zf4imn7nSDmBY2sh4FA2p8F98q2Vsxeo3AGrwWlkhKW1350TYzyj3CojrHQEKrHYqB
OP1K3Bn2Kdeens1jBsLaxX0tr7Lpx9id3R7nZcowuW+58Hg/gUAvGrH2M0Q2O+5TNpaCmtWGnMDL
N04S599ZmwqA3+UaNzvmqApIirjbqYq1eY4PhzXon8pA9Lq3t3vXDcHSGVLgZgiUXh/97YgfVlgw
Fol0ajp1tQwTSA5zyogwWcc8Kn6U/wF9GHpXb4ju0fMgJEk/Lf0QGC/ohvV7mf5sXpsKBcAJdykz
8tv12/74NtN5YUA6fiSIluDMaaZ7DakOShb2+ohj3fwTXP0I6lEo6UmtB8PCbdjcCCxLa3TLrgUq
uEjL1aN8b/tWPijxfcnKqUuMkh5m+J1ka8LHzRE3+OOaYrzT1J6OltupIwyyRXkCvlJo30RfCzor
hWtNC+C0Ve6BH751BwRut96OOs/nqXuH3zWmDQgU/4IpsiZhK0S8koNWcWvOMw96FKTFSlwM8c8o
316sCFlPkn/FIDrCsOYbwDXIR6rn1iYwbYdkThAkrM59tGty/goYC8omACDTYYAYdEgMDI1J3NGW
7HVmR5M8FZ24bOIrKevNDPj+i1ZZyaDXv/JT73Vm/0T+YKHDKsgQKsEEb6Dg7QbCgdu30I/jtzYS
Gtb0Nk2q76v5xu+hCoH6Bg1OeSzPZ2rBd7bIHZsP31/Jj0b0xc1FK4GhgA0gN7c8mlz+oAKmeupH
hGQesaaSlmRx9TOCeeOZUWxrAfo4qvUqX8SzLFrsE2kIjkBVga/YiHuNxgG07LvXfpC4/K1k3TRS
nlIN+1mbjAcqkeinvqNoAHOTvAtla/fodQooUubTf43el4gmB5loH8GTm0lcUyDtuHFZch0YLlv1
1cZUg7xp9SFu9Vr3caTEyprfiW9SedpyUZoPaTSqGger+0N1sP53WhVr8MkvSC3WpPt7GTtHdfwa
OcNx9wk3mRBap/IA+hxLWwrYspKDS9T9mZSHRjNdQJq2/ffNW+a85iYdtM8scS++18efzTvQ3Wd9
FANHw43g7hljtGUCkXdPP1l5qaaVYQM8GdIQd4MmyeujGxopKg0GfItkZ8dNb2Vx2bvjvNw8rGVL
R/UZKlfCVrQykOtIaxxsMS/dB2r6BfVWzd9Ljom3fcnUCqCFrz192Jhi8Ury89kXAFE8WFHAgkNc
87vvU6WSQj4pK8itJ9Z1bv/duigz3J1BfzOvDH+tww8pogJyhir97Jk8/U7AhHOiluwBJZ3Raw5c
9qANx3P7OTJ7ZKMKZE8jqPYMZKVE0z4s8/fpWeVVeJi+f7nxGhDBcEGC29aZLFP6UAmldlQ4V5tx
F+QPR3St9ZGuV870qE/mxBueuASIKGdvZ87r2R4buuthoe6IDVSp/ZAOqmDGvhiYfpyD5Grpf0XD
pfdMTMcnme1UgiZ4t90yo79zx6/vmNCodb3vB+f4SjeggC1iksFzmoC2He6PxE2iP5AoXHpAwBpC
8Cx6kdaHERjeCXsMc+wBjOokv1KO901OArf2MmfNZlCrLwpRgezBmdQH8e5RlQj4H2kiCf+Vnyd+
ARJsJIsg6yyy8JdNmiFYzZm6xtmzM1YMrdQOAkf21TN50lImdjhagjGG5FXM5HS9gabWiaf1MNRZ
Yn+cGQc7Jn6NehkTHkEm3oE7+y20kOUGGizNrpsEFpiXjruO4/CNIlhAOx4eb4F5IauiSdNlLoWm
a+nxmwSb1k/Y1v5gouAWlScmjJzmVKNSJsfHJclMz+GHzzQnCE1IvCDcHkm638oArxpGQZgHHN7G
FsvQGCFCRgnakORHub8SwioozwL8TAWK9ao56XuG1H4j+1cV6qbsHMGDbiHuSpVDZ48JHzVxUXks
AKIIAYHLbcvNJeALt9PC90CflLW3yx4aiiNE9ZNUkrr8KhJzkOTGyhhmHsN5QgndxXv5ZzEs0JXg
lNW+SzV3aF2eBGYBdf5CU+sjeFpqChskIfcBQJYB2BZ88BB0aTGTIs1MiaJBf1u7p2DAoELPMBo8
mZkSHDW4wK2zsBi3iLTO4rlJrVGhEPjPXNpsDKXGftYaiotbdU1KsN1+vh9c77GHgpiae4o3ksnZ
vcyeGhWMdQZBc8GdaZ8JHpAqzDmEZzVLI0/HN/KI4/1UF1gAgCH8E84zy+ItxsswhOwqppmMvYuB
w9oxiaE2zPWeLBFBM5n2T/hjdrD1U28aEUmv2zIyLYFoUQxAmIT+C3ql7LMyRWu7yeL71oppHKl9
pm6qZ2/u6py3i9D0ZB2NkPyNM0pVOYe3OXa7tJB/JCI7W8jwcYhETKjRoXuMhE3it3dnfvLduj/E
V7K2cjsjfVAQHfaEceUQ95na22chvu65VlrYWQmUibQXOn3vFuC2IvBkcwu6A11FgSnwJz90bW7X
c5d5l64iM6TQAFyvC5qhfP7C74vINPSt/pu56lpEonMiHRHIrVUycbqvwZuXHu7gjM9WkYQkfpfC
htrB+st9Guy4G92JA/BUTxgJ+DUNzTcF/RbmcE8IxIrDI3sVe6QsK4N13j0n4LgrkYjvSxMwHE/j
yxD++0amPVnLh7i1rSxWYCtpXW0Bh65lMbfDetpnNZtd7Qme/g59ysNJajMOEulTRT9Im28dx/4O
AA8z0eqMCIKiBgSN1vzBgnb4wATNkwCtUj36KpBQox04fhRTvARKHcfuwNGpePNruJ4lxVWpjmy2
sCfQGaM6ND0RCC7G/BW+2vAnIpKfYkTLLfgJS+SbvZnPD8mBOKNGgxBrWTn/ivsTRLSVRCrmkTsj
Suwjjq2uBClFotGeVpCrcUX9C4jQ1MwZ1KyZ0I9jeLfgNdUkUqJTgPrXjTJs04wrC7Z1S5dK8xLh
IKz+/91kmr3BU8l5eErwlECI8JMNmZotz4UVH5YRy62MP6nCmb4Ag4QRBX6FXl+0xSZtbwDHVuOY
goTtt5B/oW/QLWdQerO94C42iR6n3gzRWqry2K8jX5L4fvepAJZXPaHMxMORGiWeswX2sNN56ZzS
9E1rFsZLOcG0vJBwO7uRlcNaxtIReAe3CQMxYFCISRGUSODQV6hfxmUaU4nb53w/fgkeGLwDVzHr
vDFoiC1XDo03suq8XzXRQkeQm9B2TPR68ZEykEzkX76Y6N21UQgeP0O7SNXcriUhv6mO3RekRTy9
8+7azdFbKg03Qu2OdHoIIs50Y9OXpQWuccMVygYJ2g7wX4K8eI3zNAlVMDaVjSVvmNB1VgS3Our4
a+BuXQkHRDE1XcFiPsLUuQFuGRhZYjF1yeoVZVhM6LIRRAaT7WSCzINf2lnxrcHIBTp/6+zLIhGc
Kod3AcReB3YwomxZa/bReb+w/C4mNKp2rqxujCqK2s2c+WnMLgqVaHpm0D3wXHzCRPKnqKYz5qqv
2+H7AFfIpBcvPffawHLTwlhtvXZCVoZrIC7x8+jnzSTlM7TbSSA9iRITyh1QnfsWzCUK58u01GyD
S6iHokBj0M6093LtvwBKFTWW3D2l28R28Wc3uKlsMriSblLWl1qADbJIdprQnmSUTTM0p0Epf+bk
ddsofT7Q2oTOEc1OQkvUVxCWQnMTld7y6Y4IYa7GeyjoPPDcSgDHdFeuLAUSnPRUyNow8HT16S2k
HiNnIpxdAsM/RMrVVc4BWuA8H1cnbRC19ErPVltPha3C6Q2eEGhc4aXD9/2EXsPKUkjw6pK0j3xD
+qwBInUr5j8GijHCmPgzY5jRa23HcIExEfm624veuGgf9JvxDih4ZCSHlwpWaPIlBmGL3Uyvx6ax
ipHPfkvl6ZqhxpcuDpNIGNagk9v76bKWtwdzJU8rOQ5t/+/YTIp5UCB91Ny6rIMt4LrrxU1vHDMC
skVIV7SAIpxL3zj2R7NJRFSJRvgpNkllIh8C+9sB6dtYFLpvn5qhr3lCUpDRYWTvZazg9z7vQFTp
UqbNDmIyv/jlNGQn16Ij4jvjaqEmJ20dujuGDd5ikBYkfm+MDYb5vMcvF+uuXzblWe6KklJ3ANCx
t2xIX5ykp4cZ43AHhNeYj7QA2vxoD83OXC487P0kQYxAAY5CxI2lo1d9bp+ZBouTFQgYAMLgIjnX
MUL3E0c1O0NkIHU5A9aKOhRDaRZbJ+hTV2XQv99eSXFvir+oisbFj2Z5P6hCOqS+tjLZWogzRkEI
jabvuZdg/mYuAjeBcbm/+V5IjsYBUh8JJcQpMxtdXsgPSDFpbzbWHOBJlFAu6J/8EkSf9E4iR/m8
giB+ngu/UM4Q7h/V3KgpVHwrPEfE8u3iY+jKyXiIPmQjGvoU814ymR7eTLBX/AycchIS/ZkgzQRU
RFl/meoQNHbcXtfmFzgmKTMnL1Vf7TejhWrYCgQCrZnC9JIDcQmLvNYUcJH0ZMqDmFA2V7saxw2X
Zr2y/YWjabFzIbWIkqHQNUxfS3b/Sj1CM6Q+HZXTCXfwSmw1tBwqe/LsIVyEKlIY68am2Mp52qKa
t0thO9h/HMB49jBLObPOmT8X3NzL2kS10uovkWAjNXUmoTJkKxMNXAGyh1tWBl3j7yDqY/8tCf/z
+ZI1GRRPQbf8Jph9OWgea7aHciNg2pjW4K5BrozSTF0M1k1W8wiO2Q+RUP/NcyWxdS3/OWE69mYD
fqWOOBqvQrbAJgcCz1RcXS3ie5BlQ8xduTPp5NH1Qj+/a81+7vYdoXBIjimqwOrAuFR/afYCh6o8
EPdSkfgUa+Env3QGwI5QWeG9znqA+AfGaaGHquxDVGfUYIJ/33NhHRU4ITTs8CdI+yVdq13AsN2s
LQiTxw6h18DV8zjs/HkBASwD+DFL4ZOWCe9Le6CyifQgy1i57ub3I2yDAoGzCK7h2flybQL6UThJ
wjSfxvosVA2rf4P7FbatIKLe45uzea/Ka5ntKIvaFu3VrGUtpws7SiRXjTYfmdm2yzX5/ikZH5Vr
d9x5zH+WFiTovcHYVzOrxBmRt/+TkbqF4pWDmNmPH9WlFfT2goo3YqPgQi8PLJxfhFWcKNAPBdOy
h8+YA3jQFZifWJeoM6qeAn0u8ltGUzP0vFV+USdkT4EwtyscIvFI5Q8OhMFsFtxJlJNyh84YBMYm
I21y9T29FsyDnRkw0pwwuY7iPu7hmTIdok0bICYR7bS1KF9yuaS+fw7Qzaiyst0WgPflpRr1baL6
Ge1/ZeUG78BT/P+VJOfr9SrI0wePL9ZWb+x4zBa1+KY+IOHVUXyqBZcvP6rQBPzo+Wwu32+Tj6IE
/5K4DSWIkI4F6UGlEjwQRFxzgiZif6W01KVxu16o6jAYtl6iGdDafKAT21rJbBlGoj1gIvU6/ITj
7YREOTVMzVDjSYH7itEvoIM85WicTaYfmXc5HXPWTtwPiMvRQx4NLqJPo1tN2F6eB7COj+lIsdGf
tGfZyid3YAU613MrpJGoPXQ8kGGhRfrLQQH+bb4iHUNsBMWHvS3k66XGPzsTF3HvmdyBqWgipDQr
NRJRZxXDnSeyvm1d2fjanqdThbY0mXi0VbXTB9fclHi+5nfffRddd/c9CPPjoSa+3R++VEcMxSOP
dbGNWYikhkXleZbenC+7BugX24vQ9DuOpAsUnfV1YRrABgDI/EHJy7RBSuToYuyCmhlhBl4FjiIG
bj8Q2d5ttR9LCbnZAC7y0h1PIFOXlYoTtm/lQgiN38scTJvOVUCsWKFODYJiJgYske48g0pcKUg0
1kB+cQc3i9iNzM5JUSBcTCDKDjDnvNK8+kQFrydijpryLBuc/h+SdG3SRXj5yhFG2Yju3ZNGCfG5
haKbkVjR2yG3pGw+XAGnI6vDiuvWl0FlT5H62LOOzO7WcWg8dMaV/0Ap8VPcqNlbyJPDJMLDNpWA
IXdnMbDhwiCx+pKtYWPt8c+Q9+GmUskDVf66TPV6v5gBw6w1EK2oXlo5ibMaT4aFawEl401WY3xy
uuoHOs7bV7Vm3sWUFV4ihwG2LjHPmpBFGREXfFcYmTxXfUd7R/+UxKn/u0BGIvU5scXTy0IlL9PP
KFFHv/hxkcj8p2tbw2bv5P3uvHuwkmlGbxgiRNUB6V/NCG5pc36TPI7UTOm76xfeB+YOsA+/NexA
JgebbaJv0qyTQf58GVdK+OWIMiNBmXSOxKaDb10CS30DVRGp3E9l/6DeHLEXUvzWNMl3kVMzdjK9
VFm6cOxvQVXv9p97dxRQ+eBdqI/613TJ+ADcx8RuqzEqs35s4NoSHsL64R2qwV706bzutogEdYqu
9FBcs1NFkTNeaqsw1BGeaOn+KsXghheSUXcjICDtn7e/at2Xy9LoTIdhx9LV98LlOg5H+k9zDzJc
rbB8Xuo1U63wd+jcpLSB9vfYBjDrT3igNpnk7L1livKxWlc9SgJe9X7gz8WnZlX48Sp9ikM0h6rP
K3ow9VnYUpzrFQZqQpCKI7R1Runc6zxHG2RKCU6GstCl0PItkE3eKXU4qcTHYYIFD9gvLHRJ3WnK
nQ+9PSmGSuICA52nId3CiSjecAGcJDqFEmLy3TZKC0LELp7GGkC+qwvCPO0YoUh8DW107xmVrLo6
5/tPiChxJSjcBaMigOSSSvUff6X9cmRMONl6Y9YU4FQR98IbH8xyyepofhbdOr7Vz+rHhHJFg1WP
w0yuimJW2kfGxTjEOOqi/LVY7EHFFuyhCe4bPloqv6fIBouv+BYgtXKgdEmyu8kbOa2VBm5ZWMFf
bx/Qyk8C+b5DD78/4YV6lE2lvxI6jNN/vHBtE6M1p5gZQfJdP27ZNJwtf9CVRAnocewdZYH6OPqS
njB/znqDxzQkjJO+QsKZYI5mEdLjW87Y55brc6uiKiOlcLvBvgVV8BdoaLcyaYyIFoqF2XYLdQvj
AmY/YBN0QbUxQbUnHY/9ZR170EihdI4wnjSIuZogBiyQB1P0yaCghxXSv9vxMJ2rpB5Vt4fyUGdS
r4DOYQzftuSe37zLFslX/mkQJkAcAjOun0oAxDN/zO0Omxi3KTbcTjsfZNSkDlcq54SluH3x2wK5
OyI4vFy9i7xuqyRV0RsyoicOrenIfcrukGzx89WR4VCs4BtwhUNejRt9YZz8DGmskz+k2x9sBaW4
d6AdefQ2F7Dx8YP0WNUDDJyDdOXfViz0JAi1cmtrTWRMyd8bJzoJG0nyXDQGhi7Dp8evNXX/xnw/
g+/E3/mkj+1MJF5jrEp5Kf0gRJx4t/BfHX6TSzdvsfrC10kL0LLqrQL0VGn9Am5Lt688VuqUYosx
PSjCjghzGdtF6rWlg7LO+6Y6SXYEJtVYgP3xkU2h01Sl5byF9POh/08tT7Sjwp0Dx6Z/hN90PTMP
tq2aAhThuCwOJFL3PdGPw3d+gFQ3RIU4LV5u/d3Cbr7IYrIgdozZIe5LuSCYiweD81WJmTT3EARz
TkON++94WQA5U5KDnTzXSmTbuDIcKGtj4lQaIJ9A9Rlk7MBFkQQ8Q6x6WbH2b7lYhLPUGU9/5shY
U7RzFkPlkcY8lTponKHazfdj8xxQwXoVcp5Ex6phh2Pzz3iRNhoPykLOsZLBLlkJMy/YHUmL9LRe
2intzeU3M7adO08MikgumJD3st96tf7DcR2qMkLDsGor3FoX5FmCrJg6VfZKKFjbjy2gx1O4W/R8
GAEBmawK1veDTUnyVHlmpq7+ZiWcXfaelcPdawLV3E8Mdbw6lVSv0f12gikp+drqkaRDE2iOJ8SW
GYAST2j0ni98m1bVtyO9Deu7YJN9DD7VY3tiSb8jp9bwGMTnnI+xVJLwJoHU5po2LAQoL3WDjGSG
WBoaQvlXmQ3+QFhreQqOozzqrMV9MgPWjqwNPvftl9v80nEQEvegd8MNQsOEDwk1foZEokknbOpv
1U8Zym1hD3w/w5eG4E1QM6tO+bk2U2ry7FxWAhvm+uKmDoQn+65O4ciGKUP6gu1WFerfsJUsDqoz
k/f9D6gaZzjxz430q8caYiTE4HhMu2jmzf17BchAuGGwRT+5WEIA4wltmRW3Xu/AcH0GZybJAgZO
aeiJYUQnHBTN3559XeTRNF3u7d12u/rtaLRlDqozIICLeSmNYULwn5ABezTfAJfbnByWeSp4VXqp
Tqs5vXxDOjJHsWrxSvwfpM/pZwsqCIpZz+ZZmbTvplAf9qYDTrUelI3d4MeNvm95OpryfTXyk6jP
eN3+ISEwrL+CXcoD5RcuRGY2XRG/0N5kYYH3Q3czhq/qnXl/haC1t/aLjBIuzZCgGjZ/GZzi0zl8
gVSjRoY2zwU7w0x3qygszD2dfxCbdMGRiaa8LCmcJMsV8wKMHw+bR1cJ9Eu1T4OKIvEUebYd7YoA
8JICuZcVlZY74BjBV5MEQJjJVJVrgNHveYxeTlf7kr+BYf7wywKV+85rPCLVYspbHaI7fCvl4gRW
Xb1oe8L07w7VUQ7a5bYGGX+hTQZ4S2POHdnzNBSoWnLImEyCB3WedAXDCpAwYNEAxE4QvX79RCtN
hxbBpmOgPO4QWD7L7JaDRHi05i3p2fwupizQ4cUTlstZMDOPYiQII5o8/mhhLsP798ZOVMX0Ul/U
WGOnRrZtSYnghEMlXpf/4N2Lo5uDXKDgc6GZd/vHRzGPVW3tUvOfdZq2xDFAR6yIXhZ7fJYsyot0
4M4CY/H+ptl8JRS0o7cYTR/CVz+QZzyUH0v0RRVYS4BvChfRNmGv5gSVLeGfzZOhAmTS/Dyxb8sS
6KvHG1k/TfgcLO419M/B1CJo4Zc389Z24akg5s8HeCvN1qnvM6yT14xuzVw0HRwFEvKT4g1ako+5
YSFmNaWltoydNpFZDuXSH1wj916ASwxgDOm59ZcdBfwjXfC9YuZU0iKbOU3HpMMECh4HCTB+n5Po
ioalA85rzesyk2jR104zK/NrDy7uT/1Tk2ryTf19jyBS573mu0JDHO8l1NBk+vu4hcGVJZ1eZljO
GUfEjpZKzjy3FDk+YZCSssLivzn/Me4rhnmNMOHmkHaufR8++JpHkDRmsAJu7MzCM2V0tWGWsjrz
HuKEMzOAQBxLa96ynT6S/DMuudxKF+NMjKQYXwc8eZ6ssOV+MTKHEJPIxKEAWGIfkC3ZJp/nzWl6
WpX5mCdCp374vQcBF2OjIyqFnrfDLSqysagm8IHFOOdbh7pBBjbft0i9X4sgqlz0+rNEJrugQyiq
fI9qzgAJ5127gX9NLs6+4fCYm7VPmELxrbr0TjD0LcOd+yErwdWfRps/A82Kq/ZK0lOXnxQajM0y
/3Q3VMQx98zk1GIXoCZTyBFoqcYrqltuGo6TPydQ11AZg1l3jwE8u8p5y/yEiyAnF2HOfF+9O5Au
lVBzltEyVOMFaiFUEoASzAF+Z1inSALWlaU86nQr3regba0zGfirrGJ0VWPiBXW3cwg0FIUJI9VK
b2Dh1qN3xt3N18hP1juMHj+fxs1Wh++Gdg5Bstc93mkX5omx727NedtyexKKqiJQvbFpyXEVeEmj
x0JFlcgIJOzzBYsCwQ2+/mxcrxBEQhvtKJ3R0hPId8Cu3mmMvLhRXZsXk+/YL46iyqzCGnaM7nNb
bi/hsra4NBbWqFCFDTGW+S6Xf43Wve3FwsCQc2Ct04ExBlDXTJgQOtNitMB6pST3SQHCXNy5gEWp
T2Q52N0f5M9z4Etbm5u/EDcfq++WkRJZE4hXio0ct+1NcASUA7omVqSPUB6uxGbUcVamtsJeYiaR
KfWkItRknw5nS4I9U2KJTjkxAepI9DbsRqJ05f2iR7yDBtMhCOx7vgGsxq1qNv8dUm3xGsSm7u9/
CaCK5FyuxMNmfZQ0drWRlMN7mrXVDNhu/jIPombkodwqQeGL0eb7eMhFu3WanbjPxm8dG68kvBWP
Tjuqq9XOe4gjQ4f+g6OM+1UWhoA1dwvBzLpy0bVVZMr8ZBqdhHr/F5FEHpN+gxsdagWGIoZeq87F
TgVE9L/YgHwT3wIFZ0IPd8Fvt0nlMWyPbfnkQ8BKhrlupro8jCFsIGgPb6J5rgwdm3RU20xTIaXh
TAI2kRCRvSJW/fBqIUpO5rhi2ZX+h/S3iNGKJJ1Yi4nL7VTku+CM3xvcbL7ID0J24bXoaf1FqL91
QsXPMQVmtGKnQu+IBi1fMDJWg5qQyVmDVB+t320cajalVHWA4tsobR4wZv8KT5H4hnIwvWaBSgPq
DPfV+PCa7djcdHd+El8SDLfgJsjwG5gUfJ6VsHmVbtdbfkfXGwaoBimQgSnaYTK1BZGKS9qhDVTv
G2xP1OKh1NAKE89KOrO8PwIK84fVTjp/ORG6E7fxptwZlrap3HEf1K6t9KJ0xHfgSMcqdXWv8kLp
aw951H2uNxwAaqtIzc/eqCPmxx22jWYRfXw0YS6V+pYGrGr8CVDXjuQa33HcrIOYkQ0Si7qbLKji
/zufcdmAV3EbUY3IwAputQw1K9SyeJzf1waHhKYPvkohUa7SE3gm8S1OjDGI0HVUOz7/dVsk082C
RFrd6VQrJKa5Cm6+oXYoJE2v4Pl+uX+SgWeYba3SwR6czioWiUcg2SJP9KZXuOukj5Y3OT1putRY
e29aRjR5ZrSkBc1YldKuQvwRTz5CIPgafz/ItbvHO52gpRgzYMhfrgaUXyYAmx/cU7fH+rUzizmu
T85AwxbLusK/6Q20W/SYYa+VGjDE9NnGnenunOwhzi3VZxu7QuNpPlIeYkisyrdVfhfTFcEBz5sM
Jwh1oUDrL5/5cN/fXZzdW16inbpCRWOhXVz/2BUhMJ2Tk2fWqWxkhR2lZpgAb8WMQAd/PYJWEoz3
rtugFrV1UWLJGf5+KR9wT1e82VV0uE0gkUbUAUeDcZu9NnFFxzVULdS88xoB0LaDZK+WOTo4JKT6
XHsR5PdN7dlReN3KjF/Gfqn5hvgHVuyfXPuBmt9+ttzAwJIp2QHAYQDMkeGNQ9lHX3ZTZHqu2RX6
u1RkUN5QMTs0Yz84UoWvKyhJS+KJEAKpCjNSyhvlZWltFYfObpNjAoyAEW+HXjYNZzpUnnbB2jkY
hTjPorpr15t3PSFXKUyuADXJ5SHrlDY2ySlK0jJF/NaBD2PQGPTVnUbfdxWhYXzevpDgSJfGMluW
KyjaO6BN6YPgntGjrO99iv45+7+yFwFknzTOixcB9iGZyC/j1IIE5BMD++CfvJXVj+YDipueUsvu
JxdmpmCD6N9/+Dz/Q1jOm/80nSlC1AOtl4xtelX/CWV7AKNVOlQJOPUpIMU9fqi5lkVeHVOlssKX
G5j0nnI84Ixpj8Ktsylc1dCYxVWSCikqFxrAMt2AaBIQIcRBZQA1zCm6/Y1/d38eXYg6WjES0waK
nOvYID+6dG6RjVlmBidBE5dIOn0jbaL8LUeZL4uhXvtJ9I2Fp3JD/ZDXcA0PxtZRVjKi8lLM++ve
MwjDDS0riuDqG1xvTHPnjxqo84BixLAS89HW3GQ6k5P4wYmLm6NwJLYj1brMwLSnsoNQgvbJbqDU
tltn9cBS8FzgfZglbW1E61gC5KkO38eZxAKH96mA+f8Q2YRtp8bHCwfxEuiu3lXR5Lr1OWrTsBD7
TOQubdh+W5BgUkblA978Hal25Dquy3Iun5ePJPOxL76h0mmXhQKzd60JtxHqEkt1pTxCTwN/BxKP
k+ia/xN2fpWe05cxei69IEchZqgf9nXd/rWYA6TXyMxsELZxdpVjATA6UmHvKagDO7pP7xKBOw1F
QS8P00Q0I7c1JpNaWZ8gd5HqaGKTnbdMrmLib68gnvUxgSdCMBvgktwNuvzAOPfFNwexuAaAY3iM
NBaf/YHLzBfkfMyEvFzk9moT/ZW8vou/ZJp+b8VY0EwuCx/rsBRAkncEhAyULa+DYKNTBJAtaC2R
9yA7gEcsebsxMon2HSw/AEDCPJ7Kx6py0nWS2qQefyvSFVvGh2zPg2uCTDHMrvRGE0LkWBukXuzC
SjoVIUzMml1NRkSrCpOSXj2qE7icHxa1ChnVXCiLb31oBqoQK3169wyGpTvpoCVTwHp6PqI7ReWZ
DqS5+hGqAkmrYVcFKbMz4yDQO2UA/EZcAEVa88Iuh97buctHjgU54WzYbhOwruacgNVpbDt79WH8
7EjM9ZFJ+e89uGqxecC87zSHlwc4tkjaypNQVvnnAE3k6ZCsJQbwaDGOHUUiQbYVv6DKSqHkujML
qld+KYKXLTJQEpeWmyjoonaO7iFz19Fm1QXywJ8JS7iTJSbG73R+rsfQJpT8rlc2ZMDfN+U8M6bT
GGJxncV5+tRVCUHVmz0yWvjk4gcwM5IelmiguYrwmzNhVU9ujYbxIgQwO0soPl/an5xsXh8NR1eE
kLvaNs58T0f8c1pMVXh+m3cy0QYI5B+ZpBhvfwVzFuWQX74XDY3pIPDlVZJFkXYCJYaQewt1UsnB
2mlnRNDTPY6BDEM/RpIxcfcVR9QrM0yXNacTdQtiLo7CxkPGy8gszUSKHBBFHCNGLZPQ/FW7tL1t
5hdT20i9Ic2+s/0cPckwT7cO7gA5ECauAXfh5WhKFhqJSULk01LHbIQNOmvzSlUaeohPgjcahsBn
1NxMTXWA7KmvgRf1kA3oMSwHIn2ycuMwFJ1GRCFwwWZ37j2Z+V1h7LfBl8bnT3cxQj7Toat3a9Nr
PXAigl0kj2lRts2hNa0ZPgHwDQxZzrV/JOCFcI3WOUJAH2bDriPI8SVeFMTSakJphX5v1MpfSuld
6+VWtDoAQoNzsdU1FsV3aN+Atp/56wll524JAJsrFpyAA0XflH5EIR7gZKvoqphbpzJCG4YqZ1sT
9xLTo7rr1A+UDxG4NfqR279SqxlTB2HDiP8LLWm/eRLlW5jrjO9IENro9l4hWyp4iTFun/ySupAn
cMEp3e/t5KBuR1Tzg4LAJhj8F4LiW23S4iwJQw9uXvVT0XBQviLCrU7m38tdZ5edQEq+e2qseUir
7LKsgeZSyrhOL1jsyL16Aj98I8IuawLADyR0joPvd+ExkjikWo9/0GxvB1n3V6nPyiIkuEf3VEdG
jMsVcf6MhNSW0DRt2lep1Vx5GTP1KEIQTariCFEKisNbwrRFOQfmXaGqzhGhLpAy3ZrhkLPT+viq
tOe4E4+HiPdD2siXushx3Oa/wPYy1A1JjRNR3MWkBVIeDqq1sinSCo2CRKrW7ikcNpmdonXbvIFc
mgHfLLLNT27WxuxiBVsdID8Vn/F5g1BG5vfgPOWEfOaHLEcy+Qxe5jPrdrSGZdxLtVOYPDjoFJRV
wx+rKQMtjVRF9MCboA5uO3dcvbc+8Qe8/WxBTAr8mMJcJnNRHqGifLKehDjwqNnfg64shEZo2WyK
qmnemvM9ldVUdajg9PksgfMcuPUD/2RvDEWANvFjK1QRX6STxWtjwr/cx1fw0dtMwpGCq5X43mBM
/shnU2Wh6TIXTKlzbxAKc31ikG0TSE+dPxrswQ3k1C3kIyKR4+Z6UNMfPJSTUIwScex6KtrApj3C
rPokJNec+QCQLnwwROZNeTa2G4qbzU04PEj3YUNCH53pkydeKCtILJNj52aYJDpB0g0KSLCCczMN
o3y64DF2HV2RhqyEYpF5x7ePO2YxGjpNFulTaPTmJDtDEcJZHvC6RwgIwvMuLpFfSvdDYsjDfns8
BaSV8rbIWhhxJWuAxGLBJVvRX9dmNCmKsmggKQbe3i5z5cYt4B2KVbNf9n7tX1slu1rVmwhNl/N4
N/xB+nWIlATsIVStvZsUhkO7X/8FM2h9woUUITPzpwykDSTE40SK3UDTWEzqLyV6TQR4xtlNhLPm
AQMZwEdvu2dg1vtyNw5bf9JzYSK66unXjhwSESEiLu2nr7eg1e2gKo3CYTwQScal/tiHm/zd1N6u
dh3vZIydi6HHDFySJN6ufdJDUZGxjA83Zm+LpTnlQNG0OJPWzO9xrskAEOjteQ7GdyIQ8yt8t34P
EDVMXPnTFF71xFPxawYsZxcNDaonZ68NaZQ0+NCiSWO3OxXzq/yD8P6O/a6lA186rVH6FpE0HYtK
GvCoh99hcUMgP4zl3a4tP9Uee3I/jFnkXY3cjinpiYL0w6SXiGYThNutjk9GHqKruQz3YlrgLM6N
OURTy4erdrjQKDsfFa42pSgaiYKW9gib4FGJ8gGm1HAa95wGV/ovEMolg8RXNkmVvFrc9qCmCV2S
7pep5ToVTj/Zc4W0JwXw6o2Xx4HJBvMGYLQia63Apb/KOIYunZTCf8PKpZP0Ix3dAMKn0LmdKGps
Kud7VQ+QJPOIlmKqQ4XsoJbeOuX3v2QQq2kJUB8KDKm9Rs/+CfZ8F/zGwGcj9g4+zBCET3oSwR3u
jIsC49DMxM0qk5pLBZkv4x/2g7lGxwW37Jk/GhwILVY1+u4drpLjyr5r+yEATpuku/ff5T9XKEMI
B9veFvySB7cE5ieuNvob1BjGVRq6OPX42q/2UiScLbMGnLH2lkiE6eee+Yue3xAVfwBZCWEd4a6f
HD5vtDX+WQvVaM0kK5VIc5AUzFoyg3i3msRB7Bvcf03Tt9ShcWPZCSf9iJCnadNOAalkl8rcsVCQ
daRJ1ekN9HzGdGHsCX63CiOxQgh9VBzdFQ66NHAHT3IKFkMNRDJHyKjrSSzvtddD08XASeZwpe7p
8CkYBcu1pD6Louc+iCPUCxy0ayaXpA4GDXSqtK1O3xpaaSTvEmkrqQfD4MkYCtwzJvrusyb358Qv
QDejzqXXbcoi2R/CYAer8JQ0IeGzm6UZRw2TM4QSQ36SX0Vk25aS508sj3mINJuhzABi3RkGAc4M
nwUOX9D+dEOpxR8I5KN88/uW3T912Tqw+0kIiIGl46U8TlHJoh79iVsuuyxjirjaJDo7FaKe/jxo
wd6amNw9VYHzT0QRQVX055pjHACrxXWJzlNfhl0zINcXUnm/5Y/fguNVtEEiiiUTiPd6QQtxHDCx
nH0fYgUGKgzTMZle9Zz//ynpKaxWyKiHLtjHf5cQA6OYe6ers9G2q2WkeayHpsHzLFUY35BY93XH
shwhXW32WlD5w/aazpXRYviwL23X4eGTeyL0ynibmkmlTo1Ms/zhp9tCRBgwVVItmY8CDbGrOOQ6
kJS256xYOcxvVgyAgX1mZH1swujVI0+/wZMDe0+ixcaLGPirCLuMrDDNN9PudAo75VQR0EqBuq2m
xU/9jtAQprW/jR6hMocmPfh0zVmiCiq4JKGr1bMSxgb2C0a+Y47tkdAmnLowwPYQADEJG9JXhpEO
Z1+5uHM8FgKhqmRqLP1zM8kPSjPBtOkzMpq9VVPqUwXO9lLfhDGCznr5FbtADv6kr1R/lAt7k7Uc
DQVMeq5EypfqELKgq0PnUuvBqITXFuIjq7fewdr18i/C7+bywdlD01SM+hPUypjAKF+iPDhV5yx/
D3qU3n7+iUikJCN7ciZmQ1cxNfzWjjlBPgpcWe4/iZkrRjlyuUg6zQ1qFKgqNKsa4n+jwxaJOmb4
+jK5xo74Kd9pC94jbbO5VESlrGdPrbislWjj/tDZRcp11kKUj0kIvwdLkyLCsIowOUlSHYAjYrjk
jqlSbDVPKDE0sLV/UAfXWalZRT8ROfpP5bhwlxX9xVRe8y02yqwRHovsrKFE5K47Umjs/KarKKxr
0tWUNkAurJa305lpZbONuvn6nPopgMCoXpz4ajM5sI1Puy+VIo9iuFDOemE/yGpMLhF13Sbyn0FZ
m2/urTJzVoget8Xws4lS+WKOOqUYh1JyPOjO30T/QAq1OpOTNpW54iixkEoLd/uKU+beXY2+J1aH
KTyMBLyqgrRQjGmC/Caxt9XCUjqPrW8st1xyfjkjYAWcDmS8p75DxFcv+Mqxn5LIe5Qd9ygAI1xy
y08GXwLO8HoCIXQNee9i7TZ5UUHxiUkx5rjayI/7EX/PS1fSn8HMhHPzjJMGnWsjHaezHcw3OIK2
rNjhNT92BX0Qk0UTSl45BJZ9rXbekFKyz/swsWBi3MKXZJl+J1aqX2yFNYtq2BPG5i04aaVAW/Hp
2Mm5EiUQ9urOC4EEaxo1p//LY/NNHxg4MXW9Xcf++4izDyKSynhURt80l4u3J2kvSL+uzdx7yplB
OKA3hK90llb7M6cGxBGcxaJcygBqPRjbSx/Tkj3UZch+09biDA0bWLP5rTvrwYeGc4ZFPpARl/Ne
jpWG5dLsDguF+4kQCRO1JXUBSwbTBKZlnlV/JCKDeRwYInjb+sw2v8CBJabxv0y746gmlqk8JjCz
VSohfqX1wvQgbp5DuvaTbKSy0Wn6/BtQiCNRcid3Z8CrS2o/VFbQt3MYhfJgvHlYI/Vwt27E6EFS
gQpHUanpyebWT2ULLd/atFvL2vO4I08QM9iTJnd3uvyAp3YOXWQWeZZVr5/sa8kA779pidjFPBsJ
xtB4DrBlSnlsxF8DZ4VoaFc4LWmQgfkLoQpZzAMDfhS6YoPKiFxzuK/y2ZDtkvbjcMVTQ3LQbl5H
jFXlPvlOAabQpX9Yekw5oaf1992C57lINz1rhu59ukLLXwszR+eOivnavsWX6uNZwtFtKW7oQ/7z
MNgQtrUtRBsFQPdudSQBgGS/sKbKwUHj9upEVjdY3jlUi0eA6p/M9vFxuGpRBu0YKX//jp2cEJW3
rS+SIs0CBnCtPGEF9otQ8hzlYRJ4RC+Olxs5ovRuqr+BtX/RS2r6R7oLptAnaVjTZXkAaUSqUNgm
Q/bufreNZ+IRITa997aeAREuBtlVp6jgS+NZ7Bq2Tx81LsyqQ/aj/Fb/SbVqLkbHfbV3mQHT51zb
nPKkZWICAUSGXVMeYmMtx0Mcww4VJw/FDfCfcJ4tI5JkWC4tGgJ+JHsi5ZdTO7J5eb/G5tGRUKRT
2IwnDnSh6yp8yIHM69PDcDLkNOmiRcl3Zmdc2ToOQC2jeImfcfvuM/N5xMM9FdQZY0TNRFqbSwXY
kjaG0nygZA9lpA8eaYkMuiaz3uuNPd13RUlePrApbQMJb2uPa+LGFLSlqmE11Wjht6V0HLsVEiyG
6w3jZbWSBFbM8/hdDGU+YGUJV7rN6Y4QYKOn91MqAqqrdx3+Hao5dwuCBONQDRoHtSU3IEIdPDjW
R/zDk7+KOmv4aUYnNQzdaurVy9nwTCYWN7uaCS9xFDBvab0fpXh2zMdubvhlnBHRvvbwisV5wwDI
ubdd4XJZNndhu7MUMmyf+SthbQN/EcY//lU/Bm7u5WctobcQFGd1QmLaECwABlZooLN0hwtZwr/H
4hrnrOCTtlUc2aNqEIISft0j2f9bOTgD6Zr9cWnZ/aycNy5PutteHDRohLOZ/tiWQcNQFUVsshC3
Idu2qwDNQGFZ7XF1FS1FPVONpS0rxsVSHPUWSnipRmVTriJaJVxrJT3a0SYIQg/peDGSOSeFs1UI
jSbgdGoaBIv1Vh8loWOXUZ4cA3Z/cUy8TBTY7u0lJB3mpIq6L0c01ExuF+R6n4STuQ6AoNshElA0
K2QQrxY1ox0pHEX5XHdyoBmuOfJcpax15x1C2tOyoxO/dI0nwpiWIBwdkxb5NFLv/Mn8JWkPr0Ld
dxeS3Ro5vZOrcUY74NS00hO6GIn5aiG1DjYGrG+pgTJzVpaEwV9ic2dbDouGPdzPbEQ5weUt0vqC
aH08ek7b6jwuAW1yXkGKnmj7W2hhfpsZldt9C1qG3tyt71dVkS1vPCxU8vDE31TxO5dC0ibWdT9U
qb9ktc32F+bFs/zUyQgtDALGYp7sQygTBDwuc0QdEJxZqpUHn0XxnwbLvRNU7Ix34dIxN5t4hckU
+FzCwjxbu3DmLNX/2pLWLPYGAamzcSH0YwHNiDfjlayAmnHhBUBrlKSjd+H9c/TqPnqHSu/A4pfY
LLKHtCm7Xaw4VSxNQJVgJVjGO2xhhYdkcLPaESNjyTcFkX2CcFI9xgyimsc1zcUwadmrUH2AINTd
ILSE0UQGssb6V02zpX6a/10OgiU0jPuRRVWee4Zq7MsuI/nbiUoiLW6CrrSCgg5zrJSWJcrxerQI
59iRpl9dyCcGfU4enRS6Cs+ByX02UohjUhQq3jMNn4EY+cuurP7NwC38SpW5ZFZQ00P6yIoFVnOO
sk9FgP+IflNtmLlB2UQz4/0nmPPqEWPvb/mgYsOoLkWkYojdYIz1jmjsicIvS6U2koG8bA++Jp1S
BXoD1z5rsWC5d0UZAMkQRQSXopqralaBwLOrHaav/oafonhgi75DzAsZkddObHtKqTLTyl/IPOfz
A5SWDNhR3I8/Cga45CW6W345m+m6nPJcAmYhT6KWmAZx/NJl7d87lD4d1rDJYYxc2m54d5Hbpibb
fvkm504oag3d89TV8AgDWH04g8UIjqL8sRwvyk1wN00ppZg/mvJVXqqSrUMpgeSa3Wr8CZlvUrtV
qife5oaYjgxxwFRaJxjgOno/3miHhFaRAlvo7s20qlqvsfVrlqkGgbEi80Dj7U9GtJq+AgtT9doZ
fJgogrJQ8FvcUHRqj5AP1gquQmAVeezAXD8vsgEbrjaMyg/l3e2NUGCmtdL5qtTAA5UkBDIWy2Za
qFjnmOP0u5lruPEIQNH+//0j6E5Cq9HFusR4EHP77JwCUrjn5KELLReyW0zGSDyS1BYUm94oRH69
lnw1bAWn9wmy/udQqUY77ci321llCwcbGbXQlHTovqIrJshoBNYTJZpiMSKWgW3asgLKep9jz2lJ
gMXdWFdUL+i++PH1M2ZLqa7OcmpJXbeGCp3S1ODpEi0v50a6oE5s2JEjElJiOgqDiq5r/Mn58Jev
1pwpAVqnuo3rSzzNemXpsA7wU9lJzKTo2s+95Sujb3884fqe5sb3leYPjQy4/fduGIeNQnWI9UXe
eaSof1jbAgGiisGzlDOM4/YXvyEgTVPSz2gSIuGsL+ivT/hb6uWDdSrZIWRfzQN7wsRI6nZ3OCLJ
QVQvs8W3C6vMxGqyT1ANCInmg/oN5Dvv7SrzsZDN5wpnU/o7IepiMTZ77nysEmEBH+THb+qTZ16l
yJtUXlSTOn5p0+BJvH3aXfluhCVDrz2h0oG44N+nVIHseD+dUFMhHmrg6XGh+IU8FftcTwj5YVSQ
807rLA91pSLWsQDtR+Ofl8et+aaOELBUTYWMpVryWRaArA0/6CEpak8ONQ/MLh21BwFRp8dQAEpa
LLQeP12luA14uWdWhdi3ndnaV6Z+H5fedK/PZy1Igl5a3WuxuHu5HnD31qG3f4i5iHBwbo0NfMwt
of6liynwzk43/zRk21yXjicDNNVz4XZwuoX0WUWcG2NmyEX5knMKh7rtTObNLw5yge6pfTthHerD
bGNsclKUZ6/DAhxX0s6z7UZfNTY/WyM8LIIdSN+GV+Oj8Wp0rhL4Oahn2ME8DYuB8Sjuaw9uVZkB
BHz21tr0q49V6TWe8cmNllw3lwW7t1mrsCI64eYapkKzGTNt01WD+MoU+fCI6nfcRGi1+a3rqOgZ
muUY00Gc6DoCCZTerVG0VX04Z84KwhlU5QOroNtcFzOvNQ+Kwh0DMiEnHVAVdX+it9aNE9jH22RU
2gsKxnhXzQjCbmcFV4VRzc+aXUHXX8eab47hAS/I+9YNaaTFZaPXPxs1lkbOxGySxzSX7iC+jnUd
WeTrUs+cwi5+QxAthZzmQyyg0GjUSOcH9BHcMGQrOyBA6pB4pZwRkSocINccBzDGEq3WtItfZ6bC
VwA7ZMqFjaiHSznJ/W7nCFtWbtY+lSt6fVDsRmSjCIc5EAnk8JB5+LXPBl7VZ1WLlH88U5Z+h6fW
vg51L33QNqukntZkMdwRY1VfWn5UD0QUHljTFJm724ME03segSHZf3M55wVQGh6ucbiF5Rq3h28W
NmXz4tuISxNPUEgy73tINNa3eOspaaNhZfjrAyoqr6mLDM2rfJuY3QTGRY9D8XvO8JpIHLCS80VX
xEhRATazYsl2j00UpQlJQphyj45QqjKpYKypszmYESUTApIZNxAWjmVviO5V1akl9650XBOqMWNJ
+nyjb/ZP0lbH3s3Zg6lDeR/GTER1N0mm/2DScqMttJP0yrl3iCDuLjWAoHgbbj/n02/xGzJx7pAL
BWOUPGMvoEFPAtj9eRzcrsTYsde6sVMusLkamDOc3baw1hJrRkcA/I9RwoDy156uHGXXoU9ZJ89H
l4OO4h7bunwh/Td6OGbG5/rGn4O+S3UGgvyyTRoAABJaxRmRxYn+yweUPLlslRJtK9XxfLgDs1TM
YYd/1Bl2NQxpk/XLx3ZNo5lyB5z7ynk35oCsdE/3pW6NZWPV8ScTzDtQeV9zXtFoOsZWS4GljC5l
cveCNrkrFo9iLHSKug7sZL/WuxgATTW7sYAM1J5c0eVKKVM+4KQyhw1OAH31USBdO8E23Qysg5+E
0MVjLWF9yFyFXALLL95MIEqgFL/RQkz1+Ij9iOX5AmnwQuwAaZzEA2FeLTvXGy54ugBhfo7sw+KW
hX8a43tSPiiBCjzbKu7Hm6o5ASasI1aGw4//PQweSyVqky3Xvkd9UHlCEHX8DWLmQltbxaYsHp/w
ctJhIIrFRIcAmKGXJk6uqKRKnOY+gb7hAT1chjtEYc/RU/HkiFSqWJ41rPljKzSGrYKV07PlF6yQ
dxBJsFblmMzT+Fvrlmjv/Y2R2GKC6sjTm3ADb/9gp0sYzqzKMgukaaHRwL7oYkU6ihOoD6PJiz0R
8o1hmJNgKxqyyIb1WG0Bt7F+H4AAClEciVCZfq+iXRRT4rFGmUPEuGIYwxKyR7XvBt0IlM5Q8US7
JMNT2Fk2k0A3/wVhH3WK9X/yhxa2QFf3/2/IIiH2ru4bzDuJNxqM42UDCHetreBRy3OdOq8KHY4Q
XzlSn5TMF+kVAjmOiEAq0X+u4VgtYHZR2RvlggBn4egMwhbJz9bs4sanWHH0uQsaCOOGKLDwxSlG
kpSy3lIq+7ZIE8CwlC5IQGTc/N3g1XtgeBzwd8C/fyqSkXzypJldT5Kuqa64BfXql7pIqzUQ9bn+
4SzoyVPnZYUZtzoeoyDW2YvLbyrOvrWYitsYcfVm1QgwECtp5YvkgvbirRYWdpTsMSeFuy5KAOvU
FbfwEGBY3r5mNIQUQuzRgeZsXsxfc0f3L+ah1dnCxpDtNyCUJUBjpb0APjx4Gx1LEDytx9BDxiFy
yidiillf0UXzpx7sGTVGkr6zfTIcn6ebybM9alIOmMsm+X/4YNYJey2FHGJQdxcYhMdzWJX+bY3I
PzZmmofnMKuyjBhB2swTV1nxTbVBUbNkrjPEetgxDmoexfjNbgqB65QPtUNtvRMGSGfYtx/MvYxI
yX6oBX9GLPWN6UDNqd/+HEhMbGsm7TejW1bgikFglC5W5OUfJHn90FGy99+ompN2hF8/4jh8ZFhs
h3S9RfuYYZDOTZnDayO8FvtX3gNq8tudMHD8xDrFD0axOnQhVyMoMx8oril6dAkDoNK+PgBUmIbL
g+28ac/rmW3zayj4HSsfvMVWzklGv4mUDHFL/FmEBfAiGG8F3XwlO2ykJD0ydvFZV89BDHp5w36T
yCmxHtJTAzXIPoh+ISIYOUlie5QeKvCgBSAm7HMxiNMbOk9ppmEgv69lDOTFBy/E2XRmT0VORB+C
ysigBx+43OIO5L0mtk/Cs4df4xTqTHS1SKuN/f+Rl/ZzK0GJGR8CULvI6mA0mURlquNQO7YZ5We0
Tdbtsn+FrVGGE8z8T4ndFXG89xAsy/IeFKtaXoFT1ICvRc3XpIPc/kwCFbAPqf939BIaUrELr4MY
ei/yl3M8GVTEK0KRqW2yaqKd2ZlNRX5dXtAoaM/VoilrgxAKdGUtjtWgctH3+q887ciScKi4tkT4
qqxzGDgDF3NVhihDDCysgY0FJUMCczKCv0wOwXpInmKZDqIGk+8FrOc0X5cNsFkjQe/7z2DBFRj+
eBpcGot3Vp6bjL7fJZmpoi1I+fhin5CuTFU4LcjRZ5vtAOMxmFBcp7Cqk/yRKeLsew21MP4jp4Ct
8idwk4S0p2i8pVRd/Ggnw82vER64KA2kRXoJjiszfsqgmZqdTYvcvJgqELWo4tF0Fxyfo2aazdv7
fgnAD8fC9fVKZGakDgRmrxO3jEomIZPyhN1ouyXbHYMbsaD1ai0TR3+AIi/ZLxzC58NxnFPhgTMh
uM17Hrp9ylFJMlCL8dc5nC5lxV1AGo7JFXzZu0S2848PzR4fPhL6oTLCfQtcstH+eOl7BjaiWjnx
fPXD4QQCSJMf771mMT5VhS72vnRBOblsXpCUaIkp7NQd8+96fk1UQq2bTrWVwgeh6uMmTDkUNNTy
l2kbOMi3m40UiGBfJ+EtBAmO1P2jOg+qSGQhnuqkcbTjNmxXGw35YOucWQQH+CvulG1ElOX+jzSa
4lzHOLc1RicEVuUJlq1HSddQIoTAVl1/t0Me2frz/rwR1ZBIZnAWyCuZ3NJK6IFHMszDuW/uoxJx
ZIfdtCcETp5vbDsZzpsci1hRxjoX/j1KoToFQ+rheg+xM4e5Rf7tjz2awRwP937ydhkOcyonyM68
h84NlX18RyEfk4fi7Yi/yKL68RjqTIgaMGWRH44ZhRc9kYZvSKt7HA0GM9AcPddKqB8ibH9yM0FN
il+02c3TB4zBYZ386Y58yHWeOKsFsXZX9hGxnri0/XxzX3CFGoX7mY7xBNU5gF7GUmSz1eG7XlUh
6dqelCx7fUQyBqecMmOmp87NC2LloIEVDYxQULO1e1fQcHAbIyJjGAYYMjZG4tAGqRvHYJxKxRlO
bwDjSkzt81EIGGq9Pq+RiK66OfWhgRCfSegMu03/9s/zd/CYURlwWxRV4Kd3IYilTpLOl326Gy/Q
D44qcygMV445M6xW8MtWBawQl6yUeV5pZkeKPhBIYnYrQX3NudHVP+x80QRq6bSVDL4PQZbH64AV
b+Y+jYTlWq841fAWnE120VxMDTQ32xtccsam1c8d2R5xSChYFhRCR2UJO1UG8shTrACcxCuuBJ5d
4FvaZ6ayDNe+LINgoFkUvSsL7YAOYt3WbAlWit7tv4KPSUno9WXQWnPGRUk0ggqMnoR0FwDTeRZc
EgV2mfXvuZSI7kHRGvJJ84DGFVxTS+0lcIMdELtnqxoq6iUJd5Xu3GRVZojHvATLMd0NBFykjALS
VcVoWgWKtAxfkOUPvLhT9MrtRnE9inGB/WSdo+GUKjZvZBHzpbUMRdoiFyhF8EvaWOA75cFTvA5J
ALTdxTf/gnePoMjTStxZmFVDmoK2SNWrql0aZ/LCvk0iNrfBMETUCW9O6TSHuUd90HKiT/QdqvPC
00vEfGEYPsnd9WPYsVPwg1Z+gGYSPqqw0VTCLPENPdBtZZp+tTWCQb0zySk1o7rIsX9yjETJrhHQ
jzkgl1io4Fc01wr/g3S86IM3DPVSXjFxFk0YAu0X5V99Ab/08V8Agf+9OvuBV4oVOEl1mN9UgtPP
Nn8FDs3njIrKT2i1e4Xy24mVjOnXBnI0icIdkTdeiXvDhwpt1eB3tZ7Mt4QrnEh9yYmZBGJUnzFT
OJx1nFIW67RwWpiDX/y6kp6ZdckkYauS1vp8J7yEQGNMciiRqRRCddoeM4amh494m+0qX8cFvM66
JtWdxkcnGYpcVqio9qrK97kWsLZVevJ/14JBgGTn3e1n9Wdg24uU628w/8nBwclrGgAkaQ0j+MH3
I6MkG2eXv2Wfu/vb9mn20LEMZ+QuIlWA7GIg7HcbwBHE2OpGiXuYvHkFXUUP/V8E+QxUMBCngE/s
9b4iaTkFisDU37JbIX3rViV5fPKKx5A8g4kr97it0UuVtoCUh7n87XgDLIUtICQBEWj9ftXEzreq
4xnmyFYqDsrOCFVGFwbmlDhTOBAAWI+Svp4LeGk7REtFAqxpxFV/+N5ODgw1QQt4Ku9NN8V8BO3l
gjdB2bT0s058T4Eg+okKAfAOCgLoler9hAJFm5XGcsU+NP1hMv0x2qyoVASnJIjhxLYsoD5PzdlI
3s+kspY/WmQH4yO2eTgveGtl18cKBotbZ1Ze7Qn43atx/Af1F1RKg9y5PNR/BQgkRLkd9WJvbViX
72AlSKRoS8HJsUA7PRkyza6oK/mvqblJXykffgUYPuNADteE/HmLv9devHvLo/FN+S+Nat5jR80d
LTFUnIwWEe3w8wYzMPYsnciJv0PqagCf5rZYmWtcgQRit5RffAou/VfV6kqFtLLMuVfPYsNyU6KI
2URMfCkhgSotwO7nkiCHX9asbRJF7FItxdHZDUcLLlpdY+rEVJQpO8VKoZ1gcEkWh75qDols9ICF
dg4pzSwPLsXuZmJf4BUl5tZ6ccpeyOnQyv1JlAtGdg+P2kQZqKyFSDpRBfMKqkObcs5/cIWsUVgM
OiCCnXixi3VKGWTi7L/6yI1BcCnuPoGTtcq4Ijvc4nWJ6PWYiGKwYS5/tk/IRy1rO9GCRBe0WbbD
XFNVOf0C8MxCxfDBB4vD+ksprbboYXvoeyjAVj/4VgZ+UugeMMT5ilNy5zOJ04X4hcY1Odf5mUts
KzFt+GmuwNC2iCx1V0D0mA5GhaIXQCwbEMdVnb7r0JcFAzojZqCCPN6M/jRiwW9W869RM+jL9epl
K2k1b4eLPy7Pvzi10z7SIz9NbG0dM0FuNEW74HmygO6h/TW2Do1Gmdx4CYE6c8s+03m3IykveF0B
1e1snAo/DLw9SEboQQKTCEs/rQ7tcvYg9MtPwgmDnHBwu/sDbdlRXCHhOFvwgXgcLfd7w4Gkm2ye
IhapYZoDQRToNMgVif0UHgv5Qsv61fpBOCf164HOucw53yXbPzj5FdJF8AQzfHS6zq0+3Kkhd05T
Utg6WX/Hqf/oiRRdMQtydNmOQrc9MC7CW0SMawoIX3Lx0GBvKqLGsFbnZmfPt1uVGDSaxxLVBjsB
eVHSlwpnq261FebMHV2+PMH7Y05Q64Q5ZhxPinlllHsjqDqzkTiIEIpgTSZiCFqZxfe1P9OOkI5u
PafiPOVUJ9zLQmLWE98a/UpFxpgBz8YJNvX5El5/oSRkPBbqj0DZFS6k5Lkkdjsh58UZLkl9oaVM
cd5XmEbsIHqbTJanRmyCkzw3j1YE4NhtJB5oZIwBYl132grOBRRER7LEIZLWS2OTr+Cq1y3Wn9KS
JNKsfShHDMmOmOwOa0P7ZJYpbHCibfmQKkm7cnFc0KAaDxCBYH29YK2Q3YfVK/zXe6+vtG0Y7gNR
DtNupTyz7Rk4QoYd76dZggv862QcEx1HHNKx1532F+z+Vfq+vIqwgoDvmMSfQLivy0dsWqtBbPEB
7pG6sY8cpo9oQoEqtTrz3jcHWssmDV8K4AD3TL1MXjddm7dgxhquqgMxFl5jj9S2bG5f4f81Qzx6
dmT4A/8JGdg5rTAkHcgdfbeApHicFkhHzY5Bho8GrvXFbKHWXFcLFgXnxv9/CO6t6N2nzaYKmICV
wnzU8xf/c1/tRYgofI1ZutCEWBd0i5LWvwkEBjkTglVs3zP6RQeoY0cl4H6LeuadmObN7ZAepuIr
GgC8E9sU7q42gAnHBAb9e67vzHHKPfgrb+UppUFVDQfu3qd6iaGtR5M+myrw4FeUHQCA3aNflj0a
8S1FUmzKVFieWklq27cJiYJTQgjhz0nqp5QqPb9KSPug6691aZP23BUTZT+BSyS9eVIDHLwF1sGS
WMu3SXaJGH55an3NkSSDCkbiOpQxgzB9TV6LJh5Z7RNjGwDwN68Q22nAMk69FXDXWnC0rGgHkT3A
6M1JjJZPN/guhmPPSEHf4Jze0HaqgdyCiL1j6DVCYMzDpGsV6b5rqCArWtEZck5+Z/y3a1+5hsG1
nbjxzdejhgAfhdp13+CSk6IN79k/ZKhqj/WZhNx+xIl9N5xs2BQx2z5rD3K60ltY63dW3JmVXKY0
5RWaU1wWLGtmn1nM8UUMgIt19FJvaNCFGm2OwrrYw9drhH2llLOWRlz5XJwUv8H8m4ZkW1o96r2o
HCHelIxBuweX/eLrZsQEB5o8Pim84EFi4GMnhGcQwcPm6b7mvIkBS99HmfGj1i80cwePrJ+XHnLr
RacoEMEMGc1DC1Xd1AtJWWPD95/czFAthhJO3J3QvTgXXoH+S0PY5L1xCG5COfjRvYj7yu1b1INr
FgCs5VKHHQv3OdajlSQzPckZaZjANIj7h+52x0fnwQJfTjmcVGtGLTTH1IrSfKGgiccxqOsQPqXc
Ys1N07saP/SZdDXnU/WN55o8JSVFfKKasbIL3gLj2y7ggfFWM9iFEnGBdE21iE+gG/zJUD78bPos
iE+T2r4Sl+VHWgorffWtDc+/b3GolawgTKnRaCQX3ktG+yvs+Asn/GTWKlSC+Y5KkgCQKNFBPGVN
ePsBi4XZtKkiVkHYupwoIZFSbU6+757sgXgxyyxHu5dDYIq5iXMgQkdNcL04VWajqtSLaYLN3ENr
rfS2xD+s91tQZNoylILVYHk7m/gXhM45P+vaeGzB8kfBoUJy5rHi+1DcoyNA70CdM9ifQfwQaaHJ
MN6zCoNrgRKbEcmX0YtghqEHVVvj7RfHJvqE95D3XZEAmyFqofDVQzWx4lG4hCDumzvy8BQM07mm
oo8sg675yNc1QnXLxBX2GwjZ4nReyUGtz4+GysW0+gA8C9yhGPDdVfUnjsF6xVuCVWYkMWpzqvN/
AI8t1Z+zudLi59nkN6KFsY+JtV/6eF8evKqLY4HnkQoAcGTw2R4O+S7mvOIhPp4DtYQUCDMxJ2YT
fSgMyLpBboVV5lgr8/zdazbdnShrnUSn13c5DWZiO2CyQvq22vVEgGetJLTmjCZm/w35JtiuPQJI
nPHzCfUgqEPQchpoX8scWtdL/THGbCK+VYNTVTm0Kp/muOZXCEY/mDME0u9s5V1/tzO9OOFi7cNd
ELrCxb3rnfN8UuxhZCNnp2c/58JXVU1u1t3I9tX+kdKOx+B9WKCAVdFUaNA8mGcH8/EWcjL4YbNr
TsGl3juqPadSUoUEs5GPqRhYPXqOu7+1zxBR7mGL0Ye687rvbrggXmyEBlor5qwHbOT7FuFPUhsO
z2o2+xWDZgiSZI3sMummQFEjJoni2rZg3+D2czA9OMauKDjMqu3otPc0cDkxotMg3dKQkNDOZhDw
BatS35f6Dr6llHMYD+I12XiowhOAfNbD3rYuPFR4vY/94ENzDRrAUhimWhSdH5daGMHdXkXbFAtE
PUpDebGzzdBWSdUmq27b1iP2ELezQYLqmFce4cg7TutwrdgRUQ/u9zxC3ye+Th4kX5ppUdI+5A4Y
nFUrY9Pm84max3ZoiCvw3g4NiIB7tYJy7FtE+aP4tVdI32EI7bPZOzpENWK5BdKG6JQ0lASqk7FQ
orOQVxGrQebvvPMEZoR+6KOWLQg1GFueMHMF8YLgTtxlkWx0PChY2N8dACP+qSMpTQCtDKBc9fum
dFf2FBXiPaUp7voXbYdKnweeI+WktLwjSkRP4yQhFqnJhZGb/UfyJlEHxygqunBBbfAtEN7hb/MK
fkJCn9r0eyQDE8JBV9i4O9AVGVdntPIQx7+AK5/sepUnTSyF9vxqpj/YofhluXfGDcLPrW1KsROE
3yw0rXI6d/lV/nqNcIb1KzlVW/7jfynBidew6EId53XhKw4vn4lYNj6/JldgSPmCb2uNAmvT/Has
QSVwTOGov9mkC8ruDvjxea8t1L0G0g/rBLQWAeZkkcGR3Em6v9h8BnMi6xPDgBTktTTgtHtvrTsu
tfgqpYIkiMx7i9gCRJlyUkBfi6ukMaxn0PB1tCtkVEyO4E+RgFrxZ6fEyc/x3mb2gRmE0LjWnWow
ah3lLfgs7jroKD6KLyuR6UAaPo1sQtBefZo5rS+pjzsZZsj23Uxq1koXGXNa1NtohYPyimP2wsSU
hMO5+ZlbAqMIzud2j2/G/Bv6p2C0Rgc2MgEnBm+9/0y9WzGfCMHocy0HO0YVi+Kj60KT/ZOS1D+0
pJ6agPklMIA5QCIjvVdiX/wKDyYqCFrKyRDe+Y3nImiW2lmH9/FFym9AjTGT0CjHT59oRTu+ong4
h6gWPcwHcC9N1yF8s3nJeSUts+16ahl4UUOP5GR7jHDSG6OsLjzFyqIC+kpZXeFQZAgLLQRBMHaP
ySLkTl7/4y60QGhjnfAcRCeHhkHEx/5dzmzwBekfpzr0BZgwsowsRccSTepH0KaPCBpnFx4evMb+
clEQBloTfD8S3Ip0Yghr65+wKGqvYLonNMz+VBQ+itUDSgjDkQOrq1//FShY0JVFyY4ICAE93QGX
5xwxOfUTja48a3fESHJPopW/+NlFKRr/g/X8j4P6lHMq8m2Ew0iPskkXNq4fQmUaSfTSO4FPMP5b
OXVi5HIgT4uc0Atus/XeRPv92a5R4i9/pg1bH3M7IqdAo1XYmNVh9xtBZa+F0C/fdNmNxV0VTCjV
0Q4dB4fxXzPWL7nn23bzJvHA4HomsQcP7RtbQsNXgQeXiSUAbsggdXdlOd/DNrHXNn+JY4wVhoy/
htLgr37IvRBoOY2HVAIgdyrcWhamVBWIILWxejYrU7OUQJsi/J0pbR9UkYZC6yARZ2NZf6eJRuAd
WpjOWVaXa2XHwEP/TbeaMDjcvb9mYrYPfNMUkAmPhBkRB09cj71Cj/cQTvAslF5bFamqmgWffwXH
s/M0SRcj2RyXNXp+fCBgyWgk7+t52lA+b7kd4mn+Y78a3PdduH10fxK//6gVznmRt4fol44961+o
efUX8Xwg4lW1fqMSrNful2MhTK4y+Qza6BuGSnowvJquZ+u9j245gz4WBG6KeD1obxWE2lpUviAm
3N8PC6HnD1PeqQPDRgPaxSNSCFfw6KwkQvX4O4+OvKqhGBnIm7OSG31NN+0nZYnDfMhb159ZNKLA
7lk/EWAfztz5W6jDedqxAekA31bMn/QcvAU7J9tNvjohAkjl9sERtnGDONNsHplI9vVdLuVjnSsS
1ckLvV1XOfBo0Ed22EJ2/GPNlc7C/hpljxmLI87X7JmHVh0Z4pQw6pCjCzryectOUK7o1G5qAZTN
3AuFM30lgMO1hKp9We1h7gb0CbmJTTv5xXp0lyux0eEA54YHbWVFqb04zilHGZptZU6DpJK5ln0V
demmEudzjpGwCF1mJmMY1Ly9iN1mQ7+n9k71HA5Z6AxWAZ6xD2jAXKez7LD5Mdsu+2BzphhjwBdu
N3K0q78FhQfWQGz+QpTgZX90W/4H2DS9LXShjQvVmnqMy6uidk4T6mubeIO1y8Sm+lF5+ue79nr2
Cvj5mDsT1jkUpmuywIFK4zfVpm3rErjb0M6PwulS+ySmqj7zlfILFQQZmSAXsRfPtFer+cPmmgu0
JiBuRdDftlas5Ju4SyoVwMiTbgRFeKjBnxBg7ghgI0t2KaW3jJYM/U06hN5m8HJJu4db2WQJxi7J
2xQ8UXOOvIcifAs9J9JOUy7O7UoQzdnvKLb5hQm/HbMJDi473bNYc6EMSYNhdbherz9lF0Ff88p8
41d42HUdEpvA2i5Y5lv6lObasoNzPkoP7oQwXpe1VzJqEJdR8dyW1ObhHxoXUiqAlWBnsveEzxdg
QlHl2W2Uowzih79Nou5eY4kELteDQz0m8Qa6NPKqgr2+mMcgJliNdPfP6igg9Dy9Lu1rur/jrWlK
OuxF70TyM42segXL4Ni8n9WvziEoGf9HBpbxXNlRf/CVv8/WEOTXMlB+Fq3vU4xzsOTwIxdAAJH+
2I5290aUpzlzie5bz0l9egQZW0uyiK5v2R9vMxkogWMvPHT2HSiws1zIx3T8P9J4pUbYwoB0eZIs
SaauW7+G4L1BDIcVxBLV5ocoUsn1wLA3Lc2ZTJBzbjxrxQtTAhR9z41TtI6zWDpOqJg8/RYCj3q3
Nt4d8u7HapnFXNqT10IBv6NKrc0AW4GkuyX1rhWfb2BYWK113nyDHQQFPOWddcIXQ7L3el3sGa/u
ju50rRLsolHCTlQ7g111/wIEy1PqTjR/8t++2+Rj/q4agiZfesET+5tTZQozcqp4DDkz8uGY+dD8
ar0E2o15zUn6esKIIPB2B1VS8PpWDEao43xjg5kV45flSPwsAJD7N9OrXx8n6gP24eOx0p7vW/ZY
54S9L8Nvp6im0cmM9z8hTpBRGuFZpRM0LgUOvkoyjoi1n09fLAYG8bB1E92DqraKNxxo5eWpJETp
QNFkKerE9BhtbN/A5RURw7sUP7lcWY8givT5n4o5ubWUsIawWcH/B6mNXMyCSNbSr1wFNTxqn86N
AqtfAt5qIebVe0pnQJFtzRuhFccGZC8U+7agFxlLjNCzXklJjm5T37u7zujv/ScTYNjbwtJGVzGQ
pQcHpzCIygg3ZtGI9COTate0H7O/pkM3keT3vgu3SQER8i6iIiFWHJoNZBaRI78vhf+INLswfXSN
UTi6fgVqQxurmYdq0NbPAueHMEHj4t2yOMBwBVvegkSGV/lblQTS0DVuH5ihlBQ1EXe1H5YVYJfr
KShAw05akkb9y+KFI3o0aTPkfFWpgGHN4HpQ8O+ZpiVuGRsyO21jCllkREM75a671OsaBzX+Tfkx
BhJPxa/Q5vS3ohASsC6+9zRU197m+xvcJlOnmVK78J5mN2PtFG8RQmEGsYN1RKjumikKPcrF1ahf
wbwek1Ouz27GYjT/GTBrVoT6mtPe0qAAyMkKupmjCjGCiRWGRUh+cmIogFoLjF03zR+UcWsqMT+O
bJ2jxzju50q2IRxa6RKImYRwvI9GKDcO2T4ksTJA1I15S1a8OsxjF+Lnp2BmF9baIiOQKLNK6xcL
FN/q/VhCZhlnxrOlJzev/n+mjaeGXZFfgiUdM3rX7qn+2XA+Gr38kodcWIkAN+ky8wxlM/zZix3n
iYG+ZvrF0g9pQ3u5uBXKO9oPdETDZc3ZdODtu2DNagX4Qd94f3aYUl+TjaQc47Ftg+MoZSG7zLhk
mrnN/Z1ihL2a6vT92+fdS+K0Gl9WbVcvXmipcj2tKt56dg1/RlMxDACqUmWVFIIy+XnWYUibHUz7
u5iJQ37Tv99M/v+YzHgdELjvYfVa/syYQdghjuddUIKc9rKJ2axTbf6EG29ytZPD+qh5Sa8iq5Ck
YbUizUzimSHRFnZIgkKXhev8L2ppmpyt/qVmclhbUJgdJHQnLJBZClIl6wWlmXioNzJxN8XWe9JU
KIl4mMxO7GVti7KTmJ9QeQUE4M5X16FPnreQUCGSkGibS+lhkeoJGEZJ5VL7JbD0zObfWJH3gJWx
eLwDbtrp8hNEDpmhXVCjMcmDXJtv95bD/bO3axJC52hFnBrjBn4vblSP8RGZZS+Hz6+Ktwbo/toV
sNgFGUzmLFMHRq6dDf/kbnykI+k6s3sQVRl5ly3UeGFVBQwYH/g1JUUEYgWozLR5dB3cU5hm6/Pj
zEvGLTzIkK+pVpe/g22lH7o+ok/AVo7azUNuvBWlVgN5yRI2mOPwAqHWMoJSdz5P/XuWiflX172k
fWgTOg0Q5rYe1OWaEVu/XaGMV6hn+XRUXoqXfS7ZF4AvyzPhVrwCx/TN3VxkAkegbL8sa6TeYK6W
mk/H5TtjlxE4juc+IBgjP8xXjriEwh7ORIPVrVXs0ocQf7HMoBsGmnG2ND4BQinknjSSJW8VFKMC
nB9OKAQSbwlhvUW7EE7bbDa5VlCxNtjtl1XELPDDl3xgYWeW+S/2NEg3ra1D3rU+GTgMzROX6LHt
rmbb/tlliXgKqXX8M5tiYmOF7iaIPDyrLimchpFJNl6QmbEti/8vI9gzWzyMxgJqfuCZ7v/mnHPf
J9KQnFHIQrwH9UtWeRIoOVD1xoUw+3aZp2hFj8uwWKKq9mLX9gilER4EPMZaG/81UCkpU4oSzk6x
9kTKFrA+ixcOUKZzRvhv9UOZYmpg2mnXwrWt6Bu7fp61DvK0Idb0GuhgidTY+Eha4ixxdzSE0sha
Di6WL4Yedp/+4UWG4EO5x8NerxIYgD1VdQgXED7ILyGEHLLZtGYi2+SFx5KTAXQvt7n8o8FMS6sw
RZvpSgn+6ihUzRtEf0M5sg7chfufiBDXM75akDtcOV5r3oh0flA18jWEf2ippFSV4jq5feu9ZjNo
7f8M+KzTn0ygFSsQvi80Deq+RLz7TrxT3RGNocDKQxYPA0eQvSnFNT74Zy8nuz7kCdmvKUxtwX81
3NmSfv2F/8S5Ne3XXm1D5ZHBcH8iTjh8usa2maG8WKV0ngMc4sQnMM/GfjtpmMH8eHHEm9iCciWu
p3E3a1WY3xuAwnBeVRp3+me6qFcPshtI2bRhYrg9KLMC+BtQc9TeHXckN4p/s2MSTQoOsMQCeF1z
d1HYmrvlguSRiA/LExPI54H5/QJYmSm4ojk/7E+ME6Io2HA8AhNmgO/9lavUQBOuieQ6YtVkTw/a
3i2J4VxRSrHq/AHpBnUsh/tAKVl2ldEGJTawZYb021NKUrndllXa3/5QYoBdreq0poe/fgvyI5+H
QlXUGET4wOuPagdHtZ56FkbEKt19Saj5CmEjC+v8C+qTL9kAXarorxOVCLxKdkYCimvwZJ9PrYtp
wlLcPK0ev8ImadQ33WOUdWmWwpAPv54P1laOzbYFh199boBiubI/0HpkN9cCHJejrLRsMIUn/al+
C60hS+OXLpixES1yI+ox6oQQAoI1SsSoOpb2ghfra7DmpdNPKJ50bFff8jo/T9xyRaR1IbX8Dq4L
dBN50q51LnUDgS6FD74tDZ3ex3DVZYFomCXiVHXK+nr27ebtDWhBf/Z67JSmMR0ddJx2q64UcrFl
og3hQkyx4d2d2ebvku2vvUg4DPpJl/624vGgX4BqlZzUlG+1rN71DlWTsbxnFMivcqI2i6x3y4og
5C60k2gh7HvrzMHILiNImqTywEcIcyLoTNd+TlDpTMQrYhWV9f1OJOxrH5T2Hs80xF9oG2FdxrG9
6Hq+nEEH1jQFV75K6dKuch5StiusarD5EcSiC7M4eFsucg8wprrXYKuzrRoYwYt6UrCa0xIRJ8TQ
XoTKGfP++6aMpJe3aG6oIQ53Uli/GZiUQ936mqCIQbYYLTarlX8Ky6BP6G5bVb4gfbg7QRmq4fuz
19YGK/zm+2mZX/G9BjB5RQw1QNboPOGhqsaDy+Om+UR1QoMAJCVKUGHFUkFlgy5MbCe7Q1Ouaa3O
aUWCjUwrpe3HcE5FDUcd2/ItVAohMmdEtA1YoAZKsAb3vUrCGGXKHJ55COA8d2GhChoospP14nrG
0Uc7sHSGnF2wk11dNyKNJmQTv8G7iSZhy8YwcqdawfFG4XqabtOD5bddSrso/XTVtHOyLTjVk2te
c80oAjdku+u8NU2y7UQxhp6U6Rpexukun3DAZleFNA9jWFfLgFkuGKgTyACRkisQFdQxOBXZJ0ET
V1czXJDuWLnkgCOmi3cewmGEmqhGLnjWQlClqbiF5pfmcE1Gfe4qES8pbKWs9kLJTjnwjg9nszTm
M5lXMPGmO6BpDkUQRhiyETaZylGAGBrMj8MNRQSLyopr0jJWlpaHcpGz/cydqd7RGyOfYI3PIC5m
o9YN/dmD5FyzzQyd5UkHHzZXF/v4CwQHM1dRpbve0mytMx8HhHjvBTOQoKTHakMGx14bxKoGrlpo
F08QNkrASRVit4n9nprXW4RcDqb76QRkTKizzUKXVS06XWsS27hKWzWMxZ6RVGY610dVyZZxQLy6
LBpaShhujpa0PQ3dldFdeeuy9Ab350q2+PYcac/DZ8O1VFHIgN5siGtqp4kqXRsNj5sz9OZiR0JS
C6Rc/wcsMQf+mU738w0navddQc0uX/n9apf2EITltFmeXnG06LUUGohIFe2iyZmpp3jZywr9ZANB
HK8b278PQBlN+5wi9tzkArEDdV1L5ZFbD2lY4uIzhZkmJv3Rcf+tTOfD1ltMmvJ72bCXP3rvpUIT
9erOy53AFS8mfJgxOdx4plLDapL7Ca6IQihA/o1xzgMtFELP6R1AdMzupgLaSTjTs0xpAoG4zumw
kfspL24GqNXeqaXYesfzrY1VD9CSAIpsZ92KJSRCihn5QO8yp50opRojapRZS/kNIfxZ6w+anRtr
rdZtb46KqqB6+/wXY1l6edp9H7/w1tEiC/duYIBiCJ1k1Piz1DED2xr2qR4t7fEYSzBiyA5zoj6v
SiaPvsbIdPva5j0gMR9gPEtyY7eGpARVZ+CdvhjFMMuZgI6ZsZkYwtqd1moYMYPWM8pdU2owdrXm
juTjcqsRtcjrG+rhPGlC2GJd6Wck2Js+XgiieNXP5BIDQuZhxQ3SWYM4jLx5anF94v4T5HogIcQv
cl/Py+41IAUu2yuLRkBX67SUHckJKi5E5yfeLmb1o4dtvWvV3TarVFQ3sL4H1/9SnbZPAsmtLfx9
sVmeaIYlSceYPWUMhkgly46tANERj4T/Q/yk8mOFoB0P7jG0mq5EZ1BqY+QuAWTmJFVaicrZLRJp
3IfSzrU9Yi1WVsb7h9N8Pf8rjAlzMonT+s2IpD9nI9WkGtUFbSijfnXHnoU2msUZGt4Ou7T1Otny
STHDP46U4zg20qmh6TGusGl094w2cbpTvx7Pk3mzX16LSAANFPaFGkeqeHJi+8Oi6YGsa9T4zLMM
GaxtFrGmsyPSu/TbQFJoI2j3LthGHovsID7Ci3br8AwreTGBLc3ai13PK0rjhEXsJQFd9pFHcETL
3NblR1j13siMyaWo43PFe26H0Ty+Gtu7UotbGoixMDk6ZpI/Ad8vEMUA2TSBLEE0NWW9hpQOJ5xM
SUWNMjRHM8Ob65qHmyxbnhBk0ZCnoiJoQMY1OqFSYqL3ustNCoNnZ4PLqL5SAsBrGlGFh/rGX4Sq
PXr3YZIcYV63r0eufzn6Ca5vBWs54urNSRypU1H3Ud4V0RGZ6YIhFFghfAXHGF9CkjUHhBprINRe
/oQ8SzJfwMxkA+6pieJuwhuEarBysWV02keBdkc4Yl201fXSJN+KfoIryFdlOpDm8IK5nvpcu+FE
Hc1ZVznTulBSbQ06vfeiebfDU//DQhJaC9lYlPKk3Cspqer3M8bW7tcSvB86frRvTETlm6dy1qBU
BkYF643vcpjAMmgy0DE6ZW/EUzpsieBi4DK2JUwdiCN7eeaBuK8F5FwEf/zVNxv6fMPWkxywL3pY
Pk9fAbcLDkB8VwCnRzxi9iYTqM62MgHVdqGw9FQcmS5C9+ZMSec7lY7K/bSsSNdcOOX33DLrRhCe
oGXl7reBzuXgAjJsnTBOuEt3yF1/53W/Q+Xo2zt5GDO7pc87XZURcWS1GPau9gRXgkQ6zmoeX9W0
J0VnMAK6cLTIgNTcoOS0Uq3ODcw368X7ZYerTVXzCJmZt7LWD9sJ+S+gqem4nA9LaIWJBx8GZCNo
8MQTNW7wIwfSq/Y/n8pj2Of6CXkc6DdUtwnCixAbTjYGRbdJ8HdUV7gfsxvVvBuw6ZZkeLL2dqku
Nf1IHAmwm4UII8rdO6JV2M9u/uO8LHBOS4VGbAxIvGqU8cxWNc3UfzbSWk3UY5i+OV4uA7bDYTBZ
ZFfSQy2P2yin3/HTPtSy4HXCufSpjAoLOADDWNCXTyoqUOcob19RBeCd97x2CH3LRn7Xp56QrDFM
r+MrMe7IS73g6jyN4HZzXYHyg4pkVbSVbhey2lluxAc8mComfi4kxwpkuri82GQFV5uW3G//tAWx
/kUSk/NIS3hai2a+XOEcyneEF1Z9uxcde+2d5WHuK9Yjanp+6AwFP3M1qMbRMP20K3Wt6wHfepwK
zJxxNIo1W/rxhJo/p21PfZzu1uIPMKSw0+Mu9czD9vmM9O1I0QlTzeLbtA+9wA/mikl6bb2AYYxo
angDlu6xuYb3C/KV78N4ybJ1MDGttEaOtNiayqei77MHojIkHwsvTFWmCGyVgh5L/aGOecW71KYY
XKWWK1hc/JszqgZCu4ZEln2YxqhqZhMWcJMmXqBCWt7Oykp0V9TDHj0SXGC6Aelj0eAW8lV++fZc
VKeKsIowMv19aLxCZ9JtDnveeCpSWDKbOKN9eR5xJU/xd0vhkq7yz+NrOZz+6dxPJPQJIxTODUu1
jislgsL/kMThRlbtzvg5SX44B8jIPCNjENk/Wx3kN9Fv0KtFL+XIRfAgl/SvHAjNpPQpJLF3WsvN
Td+7KVdIEUUhd2UjkCJ2bAl5gl3d3EazYko8RUcDPaz+GMENXcFVhwR7eAgPScCqa80jWQanNwJp
ioEyxidH2m4qvVHCU/qTeiXrY1DmqepTcZ9MSLjTvBubPh8GAiboGR+K0qphn7nVoeonl1Sd0tj0
l9yAh8E20iHYG8ABQY8d6iUWJPZEGDncWHXiAm2rb8Eswkp2Geder5Tvg3D6HQjZTfOu5cmGhH+8
eizCLjgNKK06Ewlfr8n0kQGep8QvgvKi7ZAefTd7qhwCB8S5Ov/jwv1tLacuojZWS3hBF/XQW9vQ
COJFT4/GKqsTe9RapgJcBcPf16hB0SLUpQrhdya2s873PfyG6zC5Rs4wS2S2lb+0nWuJIwIUNOyT
RYOfcAPcUvqFbCSL1/g7+PKPFoGLPw215Tlg+MNtH+6CVfOYtLPLj3s5uPV9YTb9lQCksLJamAE3
3/2qljjEhlC+6VnT9RdxHYhX91UtjQONqy0TB6iZFtbMGLfNiM2arZ8kO5DZbTVI3NnHHn593Q+P
eAtgT0kCPY2wR/obPS4PnrDQ/G6/XlaZzMqUwaaPEE/6ou6Oznpi7hkTeHJiYGOf4zxAycNPkB4c
1W1SaNnQF8aFsqE47icJQRPKr3gwebIve9tLJ3hOgGOh+TahMqKI2lOZrOv1uf8wHC+jxjw3vbHf
WFIofoTCt5PmlpA5ogs41McgTdN1i3qF3EOw+tcMr3H7CVqmtcZJ/HLI0x6RtyDqId9AiEQOiXYh
/tfeHrsp3xYem4+j7yO4oe/h6jgJ3wTRsJQiSznv+SpsfmVLYvqayonaLmaGq/kdbdd6Iq7kZuU8
1toJh8bxfZwvyU4N2GhJrstIuZXUvyff+pO84BfBf0v3kb1cGYg+ViNDeYv3uG1oM5NVAypeQAht
WnwniR4S1DpIVJdMtg1Su7xasBV1vtEIPi0c7sOdADLPNqR1QEv2NkZiTs/ChRPdxovAzJxkSRFF
bzdnHxy/6OlHS+p29ZZrMkKfTFAVCfFS+IUfI4fCUvrcL/8HMKS/lj3ssUXgKStNY0zuDxl/VULT
3Bf3QUqP0WFO9F+zS8eXenzPnyYLtKoVr/mwheirnnWjeCzvARWd3w+bi9oSQR12J1kzV1MoNZ/d
4f8RnAo0tArYE89ml6hieVRq5azT6N2gc8UlmFCCpvuReXuQnF3c4E1BDMdUrQeDoLf20Fn6oWqK
fiW5+qbv/OQt+MVTW6cjywH7sC/aKnmhuTp1qGRnH9eIoiWtKm741f1p1fxtXbM+vna4mYYkuJp0
dnawEuKA81/j32l09zQGD8HyuGRz2nTN9QAnuOekwwdi8V/msEt6P8J5CwMW/D98Kr0ibZmYGWJc
p9/HjHPIH+nx0EdW+S//rTFuMXAhBhPA7Th8rIKEI9c56xHuA3zSsMOqdY+r0ZF8F76jrM+rmQC+
cORd+NfX9swkV20S6RO7u+HGBoCLKbp9eIRiJTGm6scCQLx8cHpUQZARHGAarR9cK/9JvAZTJMux
Gr0B0io3knjA7XUxhhH4Qz1SdFqv7RAtQUZNIR8gaOLleEfMmZat4+fOaJshSnv2gBlJSpPiXOYw
YptApa/9W9JP577lGu2dc/NT7XoYVz01DeYd3yNtrTSfq7G/g4RNRGBPT/Ys4YAwI7wp/hGSUSjD
Di1ZHcf6hoWghfb26zK494AvRC+yBgzH5xc8cGQ2dEvGOkxbVFOVDPSmmlO2ljw+6lv7OYGTV0p+
lZN/a9Yu6D7GVCtWdDrdOaCUKpUXy88NvKMtTRxskx8RxzYPv46UZg2qnj4ZoKxIm54PhgyPlEoR
8yieUUaYZrBTCZKWFudN3yx8yONxpxzuhQLav42k31YCwvsHhO70ZypqhzUFqGmQtYE7lz33DXcA
ykVZy9wNNI6yAESqDJNQjzfhvsdSuElopx5frySjNhpf+tAUUB3MLy5dea98Atb1xhRus22fL0rr
tgoa7ol9iWUJ8KZVOU2xS8BJC7IaWDaEdke50j5Np2ju1/E5qlgZecnQl4S2LKPBuGxeaEQA7M77
XVpLrtxA9GTVMmbW1s82WcPKiZUHGLU5expGiX2DOf4tYjUucdWFFxgdlClMB5rH5dSl5AGIEBGA
k+3xil4PyAM/2VUFxomEqhklr/e31ZX8P9Vm/cnCiZo4SEIlqwHmS67GhU3CN+ddjw9uNvPECNLC
CULbGFBsTtt/rGd7/ZVEv1kemot5S1KzrrcWepKI0A8p1LsocK/xprX5F2gk9MRiXLBmN4fj+RxX
gw3aaSu9jmqB/w1IUQVBnQlkd9yhXx3Joayo34OCLN7Yr3Eo6Dals9umw1jdz0a6uqeKbGJp73Cp
3T2ivFb55XvFU6e9IJigoIRqWAGTArHizmJ2XHMGw94eqMnhLReDm6ilBdZAO/Bx2NI9IueqkASQ
ITIxgV4YRiKD5Igj9J1qcebOvPeICs62RczcScXjHSpEgejWhxcyKh8zwtXjLzWtOlrwTJ6G+xDJ
Bm4a9PknYubN5wEfIw/l5D8WTj8FhQpkFpTb4rXUG+6qsk82cfArFTM2GI0A0mEQPPmHIEFHfvyw
QaWj/Xr4nAC5uWg6+wS5djI2eKNXbpefAd8MdZTk0tbrCEBp+yHqVOl7hQ9gd+bmJ2CVsnByB8vy
N58p+VJRBM/RsZUpQvZOR3oGtrFKwwgHENIMpOO9p69Mzv4+iqjbx/0Y7nkEIItrZs2KUb46AiTE
tz2TJXaB126c47qNrHUZOj8smesK2hVnpvasonviVTAyBQQjdY6hKK7e/60ww79jIXpu6SSY8aQQ
eCUnWFJ3s9D47pkON6Olg1o+xaRLrzwe2SSfsemJ3FVkXc6KxTfxnLWx874ke6v8vuFn+8QiNvvR
sUuSpeAyESSopEzzozdcjujPtHLU2i/FhrrFjrIUZgf00FTAvfk8OiYQ+J6hGv8txLXK+ggqdziB
68Cx6FrSTDXmvOOKhtOKqYLzR0vNwIQVLw7OzH61k+JeZgbbVQiys0ktI39vDjtPLrkrr7ODOetA
ykhThMjR243k0Wxn8Iv2xjRDyYyrBjOfC/GD89jx4igH9KcMJli3opximHKypMvrhMMl1NpilhCR
ogNmZXQe1VAEdUN8PRh4LD9ECzRhcmTMGyZCc7DD/TFMd2enoMw8IX7quCJRrxm59b22htHXm+ti
CawBi0UdDz2JQHT7DlFLHqO1QNIk45A+nL3j9OAKgG8UtmsTQOAaOUDoUDGtc4sfJgxZ9qW9tm+c
AWnjuq4TWOkWUPn4Zp9fVyQfcGAp3k8uxT7rxLlejeeWqWkCI14TZGaP53xLfy8aXOnnE1usL8pj
z5ADuxEi48dO8t/vnXMsJByAzEiNJNM8DUWXzhXyyED1dTmPbddlB/dWL2V5Tc+ozSHwWIP5Fp87
1nv/RkstSIWI8uPxbiooBGeZL7XrX7HE/KsFo+GqBAEHKnSBPF09a3HcLNc2K0Yi2KWx8dJLjfoo
jELR650Fj1SeQw5TXEcOKWayHuxlgc8Xbpv212wbMrlTg+wuzgQAqZ49SEGJtPwW7P8+PwohlFrg
ghsBnoi6xK4tFql7l1YPprUf51S+Y22viNNdKj0l1XqcGbeEoBpyZwKSS9Ri8wKRyonnm6zq7HM7
06hxzEcMNHKpLgysOvZ5S5nsEyFen0K1LaD00LEaeu9CMBKcixZmZxJDGnt9D4nsyUgE+Bw9giTt
jclMbfZO4FJn8J9XsyhpmpRZ3IXupzDdnOJOQ7lQAb+q+FpQXxWSWs/M/1kxHfwIgWV8sIbeM4vL
fLuUy7Pa17WeP7Wflk7+QModaG475Ron/rPrWsT+S2AfKiMJRz55ae87uSAAqgvPezTV3GT2Vtgv
xvmPuVSYdDbgK6dBLMBkyd63lurN7pvOUwYpF0rjknvvJOjjE6iXZfFJLf6PH8q8hTJ5o8rPChuv
liHyeILnuRHl0AjTSd9+J8+e2gond74yTzCBmqzPlY5gZ9t4TF7DTHNmK3cJUR+W3kKDURihgfI0
Muy+d13QVLlo79CY2HQTMuLdJ3xQp27tDFGuJYJOacAHJBePfzEhlz8KTdxPtUVoEgV4d8JeWczT
xrT8a1FZpV2awCnLEVsoMzR+yEELSguYbzMG1id2uv0B8mA5r3TXM+bzhGzbqVRowrfDhs07+OZW
YX+NjhvX9HNZDYzPFmq2RTBclI8mkTfNTwgpuX3cJo9hgU36b7Wxb474P5JjsyFDwaPxOROYovvL
Kvw+dBz3iFfzj51WSwSxJmj+IgijjvFJtgMwd/v7dE/laYxy4gzNRXgCRLi5pepK5Ctour37M4Lr
G31xoP5iBAogV+bx/2I2F3BlK9EkyuM7fai1YIaM/aMmBzliSJHPuolEMKt3UZUtPp9KEIS4hNM1
+amYqwmagTdV8K10K3tZGOAo52gUpX+tnXnSp915ZKdYU54SKFYb1dLkqjxaIB7sDuvxIOBjolMB
YnKlw+qWdHlFBsJtSrjKSdMqWI4r0iMkv6ZWQqsx4yA5j4SH4/QnWp9/AYJlMS5dBVxRkGJGSHtf
mXIBl4L30yCqlY7llg58YbeRfPUlQD4sViSguNSdIFE6Ab+CTwB0PBRVYD7QcV4doQJzTF6tX10D
kNYSrQ4SMVZKWKWcR8V1z5SXzObMmsrkSXhFWGRD5rQ/Fjeb6/Yn0RrQj40y+GYESkA6I5bAqKCb
Cs+tLvl7j8h4IlAkVB5KrNYEcAVm9EIBx/n0QS26zjMt/jdXEkGJzEgRtOW1hqAIPusaKxfiEJmO
KJ1gfy6nLhmkkgMMTcsqvVfi5/6mdOBCVblK7PfTvnBqYpBF8hzYV5iuyRQlLV1Jj7Or2Tvkvf0w
OwVTl7IsuGDrWRiW8FG32CkMVenFYBhqvLfdtyFL6GkNzZ/zTl4gauo/0wrxWMdkjSQfswlNn94K
zN1nLk0TqKsvcPFp24zeY+nSLbJZINubudX6dpK330etNHWQ/XJClqTjy10iT65eekhr1DnvvkQ6
mpWLGX7spg0FNFzjiu8oiTa8/OPXMI4/nNnZo3HI/pv/Pyh7V0/zSmDgQBrhaSVDEyszEfY39w7C
3Flcd3V/GKxMZWQ2mjV1tMgWzm6hK+YUFOAw2FCOqa88wv8dKxAhTICz0WpVwol7Shn3BhlojgD8
Li5Mko0tiFKC4+964/MMLfB7qgnArfauzwgg7f7FAYBiVCseyrtPwAPH9mr9ZpA6VakNIRVczhp5
lXkrohD/nrqaWAPGuzC6fplIUv09cZevC1vCuXsldtE+ku9yLcYJTXBrsCXPDv/jTDe4jQgbojNX
C0ZDsgD8I0gZUr+44zWR5NTFliklj+yQ4w/O8m6gPuGVKPwO0lrW9IxNjrlkro7VQ0HzWQzlGAKU
wCmMKa3Gkgka/+g2P3zqBkUTfl4TCPa2q/z8cu3jf7jK8PCMtWPV0ItUhR5SShBVfGA4c3gSit3q
srmVa0OHbYzwR93d6UFC63gxNEiXreV14uk9syYIQ16M6bqgsW1WK/IYbjVUqnIv3XyuqBp8l4cJ
GGdLHFFEcUfnRMmvlvx+a6ZDwmY+0hwYsw7p6RPlgEtDrXjdJMO3gKiDgk2E6Yowe7FGxObPe+0Y
akksZmLeLNKi7XWjgQkxvYQGfgvjgwrR1BV32KJaTXjRzH4j5Z8libb0gs/SMeCGlvFG5K4Xmx4B
Pi3nEV3ijku04/uD8vLdoFhdM5bme+KMgy/lSbEv0hh90ihkVg0mn1GYdok8KOzwxXABgDoxz1sC
GSp3JBzwv3Zgaoaz2hMPOjbz2FDJfY6/GqyHW5DqP9sn+6+7skR5Ltfg0rx2BWdBZbkeC2JRs946
jXj6aRuFjb2LI+PfEViKC13JgV+LkpqWclH4dIKrmRxrIjjNmaOsCIlX/4OOsb0QpiOjfC+DTr1p
DFui+GmCfuA5mkCO4Gjggo2rJERrKgC4OuzL8dxxNEgt6x7jHc/0EJiM9n0N8MYjAYNIkIlPjY5C
QVsQFnmQiorDUzVOhNwHecfKWicD9hyBrkxXKjs71ucDHPpLK3KwVBGUArr+AAI/GBtr8TCiggzn
GT0MuOgE7ttpDICx/dV+wrgb2IhmDzDqfN8jdSuyOqK7oeBZeVU7mg3tsQ5uee9G77J6PBU0VWMO
JAOn5ojMT9wPMrYa6q06lLszss342K8T3+CCQgMqhqgHg6FC5TXLgTuDzNyCv40bzHvOcJ9MJmNH
JnsiZIAzYcczfBEWDG5ztM4Zb96FIoxZrI+cbx9M8JHjykUy6szdvGRvBG8bt7tcpHzD5g+XjKAY
Bg9lbAYBi0VZh6mY0wAZGptUHyqxVDtkJTS8kDbToVq0LcivQ42PI3YGViwZxgkfqQNkqEc9yGDV
vjDFaonmW5KMKLr4fXPZT8viYJ5r6GDjoEcjr6RaXKdKXI5SeCYkJmEqZGAFWP5pk0X9BqtXgMhi
sZ0h6hubZbOQNZWDmoWn6F02fZYgwApJ0EaokBYWMIa+wJvYPkv5tUlm3ifx4U77h0JkKFMYViPm
Q3ShVDY3ujZPwp8y/9+wWw9HXF+bq6adAmsUr8tbS5R6HUMisHHc/i0CGK4RcBP38mPX6Jyq7/0C
xQWFYvbV7KqHY+PgpEbNn2bzGpxpXMrXrA6CPY/hlABzarKzzOEDll5KA6+FNXEJ6qgELAYfIXw7
C/C7T+XvkBq7Fz4aet/O1YSMMjWes6djtzUqpVXMrbaguSgjwuDLfPDmj0kIbsFmkzG/F96EyUM2
Oj0oUFFMpTgqHjaU/KgrHtQ75u78REmjdtMg8Dm0kfOkC3HemqWeDnRvzDAJygiuBe19nlaVCsgj
LWYT7OzjggrZUvXHMNf0F0mr9NpT4KM7Fdhoil0dOKcc+Gy2fSk7J5rQ/Uyv2rCIlQ0gbkyawCW7
f+iFtYPfhAXQyPeo+wHkk2PCJaliYdQyqUYT63lQfTQqr8c6z9cVHqDdnrrELAKIKjXjVNVoCyaj
NOYKFEu5mniW4IrMrYYwaoY5Axwwhrl7oIEn+Ci+U0bx5caKn1CptkcpUlj1925o4NI02M2m6sDB
ATb8YIdQwlLy76g4w8YaBGXF6OLAuXuAgtnGyIMpTDAHxo07rLGZmmDTorJkXgxtn+fVUfJqI3h4
T4OBvJhGhGX3/uBW3Ltyv0c4eZcFkTzpsA1ZiMHLX0xFNzy/gG1b65RfoNOxdmFxC1i1fAHWA0xC
HDekmNOT3LPNyW5mcI/B+2bgq2Y/he8n9BAHe8Et5jhfH2ZVGtw9DAJ1VD/3pKDwwN5DK67AHql1
ND/biiLKIUwC+uC8yjYTBujJyyUXuP1bqsY/uFk3k+9Naqbr527CoXkFJm1dFY0oZQdia2bFr5vj
oHp+gUGWVYdLKk4CbAR7PNOfaa0t4tytpDtGtaCIOSSFLFvcq/AjOnpYnSyPj4TV3sjMcaCLclRR
0tpR0ZMr9Y/ETw6gKSQlqHPkfGlHlqzsa27b5sDejG8O7NHBMkPuZduJc08XkvrqYFAPzjvJwOqc
pR+MUvZRzr5JlLRr6+YCJKRmYgx+Fxc5lJRfir2NR+l3DTKODmxSwdPV4wLPBzt6HgskIO7gIHkT
ObcBCoSP+BCZWAer3Pqp0fjtQb/JdX02h7WoJHxQ9OryF/HNVUIZ2g7BlulBThKpxPB/jv8uub1o
Eug0h3MJhMAWoKxHN5tZ2MlJigeycLTGFl7nrsM2I0JOroGKX/ESDwrjTcxtR+8AZRf1uXsIoidy
E+2VBNlcA9BXXA9nx6DBbzWeVOIlq9Xot2HdPUztVOdun4M722bwKLDekpNRSzurSQC+vlowhJvt
BwaSq0Ex6Vs4LfRw334smn9oRjr/Q6g0oJEJ1ochBEavXUokC0+q8ig0Q8jZb0sZfbP3zxWpFlhw
f4unRlYh98G6nJ6MGiKQVVqugdSbkiY7x4F+j9ncs9DV0sn46amZrVH+fHfit5LV287bOGt96yrb
E1FcG8X/473mmF9ktOGapSYrF+by8hJYKGodR72BAca5Ci3dRljstcypfM2vAFrAS8WJzwKkjvF9
rmSfb2dSEcofqKohAElFcPPcDk5Nuq2M0NGv0YQPG8dANxZi2bSPutd+5X387DTRJ65Y2cNZu9w+
WQpF5uWcdDNBghh4DGgzX3toVj99j5H8H0yLqTdP1eqIBZw0KA1jk1OhIX+5s8BP6DywAuRC+Btn
7ncrBvDH2jQ/+itGkxIVUdJry3sNFMk9zVHo6FiRcr4A2CBO3vlVCbK7w2YonJHsS0zgJwWBvYr+
u9WVxjFPafs6wqSmEYvqLvRCRzOmmrsigzY/zXRSSn9rlnjx1B6tCKb9k89I1difYcN2tpftTD9/
93bIq2tRTu/NjF6XXntB0C1U7joi+xqDxCvo3Mkqhl6yluPC7BZUNv3MvNTRKUaisztF7nhYQ4kE
pGJkwemIHp3M6nCsYp7H9LqOZeSPO6sPivoc2Uk8ohtpXKFjal3CxTFmZsZkeYNvQAHwPnwb0N+k
h7h+GQtg83jYxiPn9+h0Mng2KR5O/luq0V1ETVsV70Y/KkL35eqEcNG8YD9mUrJJoaSqaN84q/Uz
RYhanwHJg7wOH8A5wjZjEdppi7E3Szf443A3OHxoIoDkEdlOXqm1HLnMLS4RyQ9cC09M5MbJlyn3
gDub+kaW+kKl/Ne67W8q85C+T9NXoEO3NVB/yoImLAQDWyY0Gphr8zf+4JGsgQ3fVAmsRolMvHRi
yC6X96AfOajbyyS8Kr0N8zyOTrjYxA/m77+laMxO78SktWuDs6a8b3otjlyKbw+poUvjjKBSPn8P
bupQRH9ByKr01TAU0azaa7l+EOBlvmzf5T9KCvvYr2fGp6zGKFMybxy098igoqKOoXaoIoxA+qAN
FZgyA51bK72glIZEAOhIvHXNigki60gk2esxoMHV8zZ+S1zp5dQKieIFWjqdFAy/F9VEM8fgNy4K
zGwtAqIBqN33+SJPOZO6NifNlKGu8UTfdqLssjZpN5c4/3jvVw9fzpgK7R5Fb7BI8DlmQVkbjsVq
93RzATzNPEWz4BMqTlDwLnLl58clIj1OFSlPvTsvzV0qy/2wFcVJEjInyxWWbw9SWvZGM3SVzJ32
S0zSEVYHM7gEaTaDIHrQxZgbVgwdHJQhW21uu0t2QhgwEyiiJMt9iuZezlwWhvGfc2co3zqIPgzI
rmc8IKiRhinTbPn9BquzSRWkxF3lRP1y3u3D7w89GNm6lS8lo+VdL0TPwZoP6KdK1kXRYTO1DBwe
Gfi4ylf4p3cydMXhZyy9ewPZgOQqwwDc6uN1AwAJiqngeeBralAJ5zCgr2m++uNZVdkLDs24jblz
C/enq40AWHK1IUhpsHUTCq215t4P98tfF5m4HFgTPgSc/6tgLbJZWUsFQcqZDlsEUqfBgvGPCuY+
slL34Ph7vhha7gTQu8lIEFw0Y4KOcAh/tIAa6gBy8CtbVcqQdqW9jMpsHi1Z+nd81Y51g7EWCQ16
Lm9kGA7JAsAnKg4ZLx0forc+g0/ijguk76LW2EBg0wfJyglCfY5q0PSoaoNk3od635YP6SStbeb5
07cKkhv/yTcBcNsp6tzhbMyjBd/yv0Vt6TC9AR7PgOcaAWf+nnpXgGl8Lr0tzGAV6yITHHATnecc
ht7inR3QKrbGm0W7ObGVUv8XoBoOniagXNNkfN8Zq4XuRuS42KqotJnlfioyo0dfcocXrBRa0BHE
axwCzqJTcWPjNHssinRxFXCNB+xFVqy/uWr1sLWuw7ibpIK14J3hxi9yNgiF8O4mT2qGE7uqA4/a
wEPHk9ePlZE+KjrPROGMKb9CH2h6t7tS1cQRKbRwQ+6DjqZK7MmPu7luAnKLF+TTG5lR3pgsgeR2
TmihQeIrhV+UnkE+fxsjQXI9Yd/XkIdEikpsbGT/GNYlIu/cuIc1gut0wTU86B2VqP7mRmFm4kBY
lq9puEUEiCscmkeuHwz5ZDRh7Rav9rcjIiT1Mm5zZdo1si8CbX0/5pLpKp+AR+krK8TnpYfsPQPO
F5FrJcq6R4SMk2OKjA+QyqtZEObIx+f/gkAivkw2JYzeK2e9rYC7n1ib/R0H8QyAtCLGve9L5rTw
rEmR1R+RMA9vUNfm3ZbiQzwW/YqjGrCa20KKuflKdfvpTCVjuyGjBUUib55pK0Az0Xv75JKTKJYO
OCjfAEGuAPSDw62eHuzyPUwuVIAgdpMk1FRs6UklDoQgbuzeQ6uYIAeuqtll6Tk05PnjYXwjrTYd
dtBCFXPW24gAxTh6dB/lraB0sgevWN7lvvi1QzmwlSYF4bfZzjUcyJX+4p8cxAYCzzxiPZno2ntj
5xrIocu+6JMtlvNop832ptm4G4RELtzNHyoUiKox7QIYvkd4DDxsCYphEUe/PGNXsmJDTbH6W0kE
U1lxvfrZ8GudYp3KnrZ4LU9VaR+wSE0ewvp0iycMZyo4G4pgiCCwtaZC0m4xhCTdIOA4ZCnGWnyD
F2Z7zLKK/lwSLpmPpiybwsVSRadAjP1i/+MOgYF0tGaPzQta6P9iY66/lTsRJWhzRQi7zK0JJROU
3a4uYlIftd2xavtSrPgMeEaxGmAX8j3tbTlioFE8CnA7i/jCoa+Y+7I9Hqi9xq8eBnixBnNk71TL
Yra0oP6Y1iwRS/qh+zxM2OCRwhAHnQcBFML7Te7atOVr54nToAzhe9xmc9fZRlW4TtDfhzOXndw2
RP+o7ckST75L1e10F54xoiZX8NyZUVHyYWGJfdhcza2G6bwg7ntXAkShoW5le4n47dRrq0XYlfqu
G5QsWyOKbeC7mQguJQVjfPyHM3wjrO4vnTPHKR0+WRpZYgP9BNds/s2Y9oTwxtYuhyYFCi6aWZqv
UcOfovrLhhTFDgmhf7RqQXct/ytccvfKpVz7Frnimlw8dGuS8BHvnx5LF611Jm/uZYJtymNZTYES
4cXcJMsvezJKBSOznGxDCR+E2D2ZKhJwOHzf+CO5u/H4Y/oBnaRgs73ScLKemEb4tqzETXtJwUFb
Zt5kSIC1oAx2WUnkosY3goJAtqjkMm+SpBFbfLrzTMpGzRZ5LNLjKl95I832+W5vbUYsxVbMSof0
3xVq8/m79HX/13gZVPrXZ1iVOvy3HRwC09FtyXTExDZMgBWAr8nrBMiPeH3dJDd8VU565mqFg1m7
AcmfuBtDmN5KfMLtDtUGhTLQFavR/dMX/otNAZyEGLWb4IxjyhmIera+kmWFBs8LcJRAhWdXLzIm
/TdCegLMjoS3m5b7l4QWcQ+qW5qvuBO95+2EWAvSPIkspboPzeMjqoYo3vvjGroVq/EaAvm2E7vQ
Y+obQ8lFyFGLFd1foY8ehUCKqfIXG4KjfjywkKE6AHn1u4VXPcTv77tC/+lUzO2aQdbIrAaY8PYK
g0fDqSoXxBfgtvdQgcaogd0yJgc03Cjrvo6sldd66OU22sB99nkMvPY4nicoc9ja7Zxg+nSY+Tn0
Phd6Ks5fMTUn+K6IUl1mWg/LjwwB06iL1S9XtYE58X8QxU/SRiqbu+dGecA/6rzXSTWjUxiaPBrn
zF/gse0+WJ9Vc2kXk74ZWArXlA/MuHm9ngC78cJNhO6gdp65OHgKAk9Ph/DzorULOaf2lQC+ILw4
ESz84A6yYoveUka3LvIk21F7S0bDycs+GD+ynvZoNwVbjiAEKCGSM8l6PuX0ju8VI23d38hW0HCb
a9p2q//C1wMMe+7G+VcDaLbrP+JhvcnLuKZPKGE/tFulPtKSr2AWEyfp2v+zoZqxpTTSkFJeZA1G
ZzXtjjQisJ7pimRFMUmTFtYJYSFk501+vK1j5ELaUab5hu/9CO2QMK+j+RQ8cBrzIeHZivFwJ/cx
Qrurs/ZQ78t11U89q1VXLeIh9pj8dNMiy8M9EcuFu3vlWV0H0Zy2mceEzXQ3M4vgx9zN0nASk/45
bbDV4IvaKych21OIY4urZvX7WmVzKLaYp5ZbVRZEKGfjuPdyTafFhtuhlTO/EN/2qLQ1OrzAWHRD
aiW9dSkHDXgvBcSCYIIvu/Wk52EUaHKwKoR8wfxzjf8WknWQO56kDL8V7Q+MCWHGnRPsQI9NbSlu
4EPcL4Fpop2C6vMmKgXqG6mYDWpW3fEuUdfsdEdYo7mDLkx6R5KRrRzZh7BV7BO7SiyFIACxi9kS
6cfSvrbphAmFVK6h7CR/IxHhJLbV+BJOvyAuABlVLcfgzooIaT7l+GaFWBEPxbbgX5BwHqrs9xt3
7KiIbnqG6I+A7vxLb5sxoxFc9SRxUAgK0Yomi4WQxYc+i9hhYuO+Q6GAU/HoTyyDoTsDHG9zgs24
t6mXxAQzq4K8MHW0A0Pjh9B7MjvDTttvYZIc275PowJZWrLN11Ud343EHNYj3qT+ZJCVwmMiTe0T
guEZ4qAku7kjB0ow7aVrE605qV+ehP+OqYtQgs8vhoAQYggA818NpqxNtVUJNPKbl1HHShbsWzHp
qtc3H2OEAwTQ2UxIL013wzDqv82JBLRpQefJSCaAli7AX6DDwtOt8T2YeeIBhO5KM/5zD36t5Ezs
W8evF4OqGEBN2qZZnLIbxRfYT0+rI8Gnqm5f3BXC/xdhiOLfUln+CSI+zqsZmaRuMhankyCRvCzg
YK+ZmLAHIZrYwM19lS2y29AcmS/Gq0hZI4yS2kdeJGL3Wu2opQ+XOoDzjn7kJuUh1bVaYq6HSKPR
nUuVLV9uBsplnyvfOaImysGKjWj9T7vFWt3JZ+M7TcjNCkCd3XANTkold08P8UfmaDHfrpT7Lc8D
xyreoUuk79GzFYj7YvG1K4XKLMN/e5OWZdu2xWaeOhRJ8yVJYEI0nAwI/plQ+pUdhhQFHy7+5U/C
ig9kBHdEfFJdNSqDm1XsYIXYruHiPqem+ST4BJZUa8hVST0F7ycPw8NKnAaWry4EkhDTIHgfQgUD
nNz1Fzwk+mZze/NGzOkt7mxtTEkfE3tOrVXzGG/8g+7VPE7CJYch4mOA5slUTh7uLgbAHlEi0/Ar
5kXl6grtMROWwecBwvDfAJJFOZ+lMGgYFS6gN8hUt1FPTuxl2943Ji9af7itPG++w6KvRZW2HP6s
Tc4luMSBHdiohAFo+vJV8RGs6aWsy+Qg1Vpcio3UqkWkmcwqoDoQySuNhawHgFjamGjlhX6CnyW3
ModrTqMj6MMaaFxG8cX0aryyjMDorPCSTAJc/wundpjSx2EnkzJYL8m0tZq1QmxPGRWRF/3J8WQp
kdp/sPahwxtd6pN3bWVoZAbUE7qeDdF0ZtQ2hLuNSuY4Kp31N/jqEMnJRv99kJ9/JLJw+HLpjnRT
OylA3ilpRu3as3//A3MVGcr9kLdFF69Xappku6iHvoveEyMiPU/ql2RsVDexYeCsLrcs3HuhbkaY
GvgZDZjzrbIw3n/8VO2IbIwX6TebPpXCsTooc608hsyC8Am5kF4ZlzN4HyZlOb2rGNbPPJt54kSa
qWqbyTdAzyJtLwSwhHA/ILBIL5bPe+SWZicWFJ07kiUY8aGgsWnOTO25XFckUvAcmhdDf3R5Guj3
RyyXONwL1CXc7vPEM4p7AOM95vfEHrgocJhX9TF9K50hBrbayBR0cVND5EUFrhomDNCTu85sU3E2
wA8PWpQQAblb2fi5N9cAFz/HaKNSvtdtyMhZ4mOg4J5K6olsg9+bBcHV8WED9le/jBoAWs+Xtu41
X+tw524jSI/gmOl6sM6QUu69Bqnb+bH2JsJP1UqDq1jJV4rJux7L9uIBjCxGWLxjqbAl8n10j5Fq
ip2Cu4etW5Nlr3n9jTJBr7Pk7TQgkadcS5tws1y+o3sucKhh1kgcami/xHmxWX4jJ1rvf5hY5lkR
7hGFoVtWICHKHmiQDmaZBDzDhEGfSvxb/r2LjZ8iTwKJBqKDnkKLy9j754sCJ58aGZbGXwl26BER
UAw5Iyx5VPJwMMxLVgFSnTIs70ZYIgSNxnRDpR/bwJDOJntiV9TjzmXGpTqC8Xt2E3JQpT/pTZA6
7vJv7p24H740MASZ4CA4sJwlA85+2nYCUWyYE27zxE8FawSAvkc0QHUlbUrHUJtUBkPvYNUisJ2M
PTSeEOVwdU0Ayv3YYdjsO6K3OrjTdMpdOC3Zwa126ifauolfXmdg0UP5L/PmY2LBKLms+bC4E9fn
vFOQrFr9qVsjPZVKTNB0zex+wkJJa+t4WHD0HPvLHVoza8y5eF7/aLz7+1ZjJSd31sEBs/7UByfD
5mcZGEq3QZjLIvq72nDxXe/C9Ca1TgCNXpfIsM8KlPSKucn/tYqaLWunlddKrW/WbuJ7hGRXXhB0
Nlm8+eFwKR/x3Q1Lib30XG4RxwfrF1+t2EiXcN2Ag7JBpjXNhseLQdOrKwsyAxPQ4OJYGPGGogsI
YAAltf1F6PP6e3RLyB6TLikQ5BLE9xdq6xm2wC+sgGGyhp2QeT9Qnj/+ixIbe5rPPHomq215yr82
bYqH29LouJmuGn51Nok2t5hP3UopiQnQKkjD9xOP8AUYtV0UrmCUdj6wviCCALpMNNEOKWjQDNnb
l+k/yBRpkjcZdAFOdx7L/CSA8jiqgG/H+4KFr/YAQviq+v0drTM6BzOybTyRJuIznYR4GuV2aC4X
CdtfE5RNVZEkzFBg5q1XJxyuQ7iyi7dwPnQVHdjRfVuPPA4UtROs8Eou18vuBwHECceKDwrxXFMR
DZwKZnSk0tK81ULQAgIXRb4I8GN+c4mmwwCpFL1Scu4MTqBQZOTQ0Sbz3RyO5jSKRbhq/y727oze
oIibqfff5gj7CoP0fpz2SoFGITI9/7O0AAO5nkfsvdKlDtmtixTMq/tEQRmVVAtrAHllt4spD+vL
Ygz/kB7E357kSUauJBiL9/HAr4Vd+YM1AT+nKuEqlSUOvmyx8cfdmIjTifaDKSC7vnZG0Qh0YneU
gSM1S48aYP4hM6r7rRLzE13LW6lEMZsWBxnsZ7gWQw3IXLmuW+t5mGwewK8f7IRhZVH2iLJErJnG
9bWQY4HHJ7G7nD5/kb+9UFxC0u3rKssvOjuSetyI9q+oifn5D9mcYLAGBbvTtX6FUEVSmOS3K8Vt
PcPclgPMXQWq1iqnOrQ6EjiIW/qjwdvZMOzsbOo/H9n9C2bsAjHZbQnvgbcL3kAGgZwVmHWGfh65
FIySVM8idwIds6Lo60+Ioz3eT92wpd8f2h2Z4HLth+6jpgj81U2rkf4KTE6wd6I7sM1W84QeOFQU
V/RKVXtzChzF2oO9LTG26xhw4DuT2y8b0hljjgV9zZobM02X1QanDQp4vUVksgm3Fdd/aA+x9aOC
oiR8N2K2K28Js/xM4wL+TL9ANbp6BPEVQUA33HvRQHkTwohxrtSbT7ACna5Lbxn+uQ+Y4d6C1Cii
BFnEHsK4qNNtuSYEFuW+BpxGx91c8SvjvqiIpurJktMZ4Nl3fszxqst1HCJ0vVSNGltftMPqLs4u
hn2+EGZ34HE6sYFZmdVgVvbXj2gsnA+iC83dLWjO3tf9f21zMPtc/vG+FZnjFFzKLR1sLXHgnD5n
oel+CmgLD1azSmjSg0Ov9lHcFLJSHZ3xmyZ6KrhpLuvynH9KkSr+wqHMzIG7mf0TlxR5VaqNWoAM
YRVM4og/GCrdbeF08Bys+LaPyqYMCuCSbqoTSPV6aCGqXB7YhsH9Hnp1XYU2k9B/b5FWuopBEFgI
FY4J6dqOWFllDiZX3vGmfR7a2js9M44q7HuXTKK2wguXENZQ3v9qM+j25dj2diP7gY3AO7kPbCa1
keojxgkNczOMx4ryiFyDGg0bfDE/usN3Dlcvjy4JbNQ+XGsWVhW2tf9v3Qg2QeCqjZvy0t2L96GT
ko0wbI+QZ0MAjS5uQAx26Owyay3c3usS3/BYwbQs7NERs6+BGyZBEbkB8pOTI/ozqrsZlXPBUWgQ
pLO84a0O/WKlBiZfMTNXJqDJ62MBeYHDAarSs3g7JVx9l4XC2fanxADdiXac8GLG5dKYtOor/KNt
I9qQuOIe0TFv6yydeka6O44yBRwLKdYCDijmh/Q+TSQrYPtEYRP45szYsidPLdm1EB9UV0GvX8ez
4P751ulRTnD0POaTiz9KY/fpzdCCf3oKgfLUXOA3G6rDkrhYqmIGrhBZ4PHkkHz8Gd+LiH7B4GIz
9wNLYOPWSoLJyn+O9xdsx25B4AVTEFZ8Fx0dP1nBi2pxMPxY71NnfZDu35qLseFfwMjkAjHGk30W
BiMsDQD1SJE9wOVYnjHLf1lsKDDCwrRPWvBCqAD2JRjNI0k6wlcGMoAczA1gI6TRrbcv5ES2RypD
svp0McwH0IRErxw4q84ybzmTG8O0wmIYCphx7PJPRNdKp6SOW+m5wc/P426kP4ET6T4FXu3jU2s7
sSR3BDl2bVlz0pKp6vtA7dV0uTCwjRWFMNKB7UGTkrcV7V1I9dphlsdRkkYHoTKfSBoWTr6ywbKe
brEOAUqS+Io+3rGktG9zLFs7KqwhiZGT1S8j3umxUejv22KBIWv+1t3k1ty/scbsMx1n6pQcq1Uv
ud47LCV7rZr2wlPrBdceSwMSH1CzqIDL1IEESjXc+A0g8ahHcBnrZisCiT0nSfgRREUUL3LD8N/s
cAKZ7gT8XxlOkttdueyswt6EaVpRq/nyaCi0wB4yy+TiEQk8PdOKVkXmelcOTrhOXvbK9+RB/hX7
uqKke9eyCZfqLTbKsTu70+oeqx64ZRYTlLA0PL+76QkbNFpPlf3M/ja+/NsPKRlpxaPqUaMldY3h
U1kDt8hLyKh3ltY/DAmlpnwW6pGxK+Hf37UdMIBRuk7vSly9G3ygKIdVSENb/8P7Fb6KVX9tM1h5
XV40lMPzco86VHEKlz8VSym/k/h2NVjeEnLSV3Za9xNGDyd2AExcgdJfM9YYlTg8Ecj0YECn9Oym
m8RAvXAG/OCJhzOo/u5KTDs0sV7MhL1terxBVmeRBRn94qBZE6u3nddDRHxvme4t6Dwfj3cTHkFJ
u2/Wj8gyW6XEHxg7C76mn+vtsJN8A+VNAhFn7KcxqRMBBOFLFoKR7H9I3YuoUT3mG4RPxkIijcQS
pP3Ws5pLu5lUI77kk2qyMcD7Nt3YMXM3PxVB2o7EaBgdajjpkhVPDmx7MDYM3nBIBRGKuqV5Wgna
zthhK5lN5ziMlmO4V5UZhR11eIKw9XY2Y1xFIzyvSA/jbC7pefJHsgjSZJr/75zFUgDeFXwKzF15
S2sLXs3RC8OOSs2IldyrMqfjMNgjgd/9D8riHNOAy9hsIA0f+SEXfvjV8iC652h79BFYtWx9w3HP
ouOENWL+1D7Q3+ez7YFUVpnQGWf+WlbIQ0aS7wezQlZzBwJjmc8qzf9P12z5r2EMbtTAxvdaKsr4
T1alSzFnR6fyJRbDaiP0A7Aykm3cQ+hRFhkCDeZIfYkrYDwAiG86Yu3oA1tze2KZ78ynftq9ySOM
eVISkSyJi0LtuUaRon8xW2ePLIRInRzIATtdnFGsPtiazX0ojw2R4URUkENT6HjIyxZR0bYVzjvb
IL4E4LoXzfh15UKHcNd/kwCKIoA3suOvzCs394Og7CnE01DaNtA+O2eCcfT5w+LfCNoE7qrYu2rq
jE1wZzNuhT+nsvWEdAv5Jjvj3eqY2Rj/s7vqSNsDc6njyUxoD4tU2kOcUFUfWZPbfPtMoBB+MBhO
y1yj/WXOehdNlWJExFq9zzwQTNhJbUl5gHddjCba2Z9Pnk1PIMtiyUW6mxnTVEhcIRaPiCJZlW1o
IX2UzOSesiIWWJQmA3d5lcmfz/o1yxc9MY4vInE4oUYXgAYHNN7RjMgxqEkLnf0Usmafp2ZM6HQh
UdO8E2REUKiS50nKqm59ZS2pHExZs8VQV7Q6ghi+AlQs4EBiXxjfF8yewy6TCek+1wJnVEPfyb7E
EEmG7+Sc9NZen8EZBUGt8dGfwi9EmK+32trr14keOoSsTrrCyF80I3UASfzf+aW+2U4j/CsqtCtX
K7pajRLEHe+z/7/fi0/xNOqF7DE5Zquv14VpiNJx+G74N6l5dtmFPiTTDm+4O17gCYN6/hUrn5ju
JEe3l8VUr4TkMr2JuqKeg2/8cKjAv3Z1HwZr9pbo68zZQhIySmTRjZU7I80+P370wE0RSw+moxdx
mAx2Uogn75QNlJVsKtNiLGhyVGIgbktiqWkSOBFLOLpkDbQEB5RJF5bT8g6dlFS+NEgaFRkrV0KH
G9r4eJD4RA0Sd/xEFy6hgI5GF15BlEnnFOxoIFsqfyIUzUppOT3/UQGH4VF9eyFbJ4QfECX8aeAJ
T8jOtUP/kw1QSSh4KxummUaxsGjZrh+XaGZGXuo5/pSjhUAH3sjZwN7wFmRviE4PMHEIS5Mu+P+a
05xDOTR+aR9wXJ+479KFk8B1wozoTO+lLpPTQQXSIja25yvSAUUGY7/v4Nme/KdVyYmnhKN+LAOb
6shDPZB65TUpjnwcAmetrsbpkcyFjuy2P3NziSN7wKcpbutkeJTgnyc7t99MVW2cjfn9DIxMfF5K
1e3eKEB7ggsq5ufJx4gBHPK7lHuEN/OlkfwSRRp0MVlIRCsCNTX01LT0eXnguHZ7I2JCqQSOvgS0
ptaPXNaMhq1JRZd4DRJTZ03qtt4xmxfIFUpQK82v3PMiV6HLNwanIzb7ta1Eryzy8Ycz1HuYhpj/
R4tI9c9xtdMCDX834OBU5r8eKoXHPc1kgwhVwvZy0phMM+LstchnsLyy5N1k4WXnBxZXFHIdcTrl
H+n4YOMl3zJ7sqZUB0twclAVAizIf81cVGmS4DXBW3dlCI/NW/JsjxxBRZbn4FOF7FB8pgiWFX9l
+FUd7MdiyifwpfyZgbDOaH896uXV32mC72uYEUHIm6mrapxz2lpNKAXwXVqmzraJCrJ/L1KjGb7P
Yl1yYyLiwstL84MFDrl4dLCfgSND++o+pC8WBTS7Iz1DnhuIMwgZox4uW/HH5r1XmNpC1wGMOrZ+
CtMkf9U9vyUdCFm4jSRO4CdpzvS5Du7ywS2reybcuWZttOFhm/1yeHcyzn5j1YMywiSyQA+dbKtA
E3CVLI0kIK7NsoKq3w2VDySfVI5xAevTdivOrNxaW6pgNFnIBD48VtS3RPZUOCsDFJpt/IYgz7CU
Sjs0Lq1bk9p7xw0IXHbqENInrQ7owpxJVdEooXgc3fKMXFRoVwz/SbEdyetn4TTybWRZH9zsfphh
QYwSysBlfMw6maJkHB5gOULoFmy9teimErjrIDLJdN5d8aDEKSPMus8DKS3EI0PV0v0ZotmlK7h/
L4Iq/DQxAQNgeA/DI3SBkio2tBYLe14H0OLzv31gMOMnmpmFxrCntwVIYa0dAa9LKRKug8QGmQtD
N5mj8n79EvP3KjjEoilK0H8YUyiSReXs/IVM1tvji4OzIUmTyWRXkQ8owrzPfn9oSUh5Llpii+Mx
0ad4BT6r5yISrfSjcmm710qznu791a6V7VxgT6XJ+fyHqS+5DpTrOubXbVLN5AXJ6/uR3hLPja3g
h53E4zrEgltdT9afAM30dI9SaAhrYxowx42DzjWBdxsh0poaaj47/zxgiP0rDdrEg/BpGsAyr1W6
+e8UcnyZT3PIKCNiwEArygygmQ8CAGJArMTq3NKQOv+o2oYkbBPxPjK4EUZ5HHJ0bvWWUJNzMnQH
AbcKAQ6xwRbqRC71sX9drPUotHp4sKP0mNY1JJV8HxUCW52cdNnvtjTGXpyRFvSlN+b2YNe1CQyg
5EMAm3eTsPsPNeYaQztzTR3pEwIuFvym3Gf4dxQPm0g7aPCz147wCHsNSROUqAlJ1qIFMSUwZtSc
LBPSLQ/v6aPdxhDc09PWvNxXmxpEy/Cl3RAa6ZspQcPZe+xJbC2yx0NpviJTkS64JWkSQofsRgSc
FQUyYnJAy2M5wkMiDceMkrrsS/wCtdvyVh8rXWzYvlpK+nvx19FFdQj/HWEHHXlt8NEpUgIl/NlL
+/2uea2IRR8Bb3lYgzqLAZ30UCUam/bIwutzG2T8eEKFMKk8id3Kq0h+rwxHLigbJiz2je8fVyNJ
lWgECEoVDBu0rdxWxsBdeEBraQmg23DkA8WU/Npwh06ZKot/oizGlSaXzA6s//b+A1rm2nRywx27
ekjSkdzU/oebrECAn7fvc7qlcI4NbUGzFDnpiuVhVrtDtBXEd3VPEvvpR0nLxOiywXJshD9VkAIv
Yv0o5ARQGDV0exbTQ1LDvNjIulXiXdXJOyXPynVfnOK51gojYmc/ZCs8izZNInOIjIAA4j3JAXoJ
hIAXFSaregkREkdAxmZWG+1BdM72kXxWoSeEzE4cYbo/oimdzxejdbHfx1D0A7ZnFXDy3xufZbFX
roHTvuxkul9oX8m1ZzmSrkD7o9XV+yymKzHoUzEWXbISth9vrJ3caY2nWX7j9Djq8imrXftsOaJ6
3KaF2wMvPFFM4FXfJcv9NYU8Kb40uvVGCHfiMxgAYs1uAaD828n+qoeiT4xn+ES7AH4eI4SV/2TV
pKSBds9CN0sPYyLjpuHiHELMYn46AcCQh8VQVEwse59NPQD84QXO+RKtcG3Y3l+WfaLQhMLWDb9L
xU6ZQx3Xxq1eq6JUcHIEG1pR4S9uvKk/8kwvVgqh5gjL4pJc5tkRTrh+8aEKdHJv1vfS7D1+5T9H
A8Hlq6S1Lw8rjDdKgvd6cKJpOPL92n3I6COdc9E/234n7NcgO6jgSIh2Y5yjBO1W4dV/yZ1ESy00
2EpbCXpxJs34jsYBhm38rSNmqf1l1obw0UmUZpLsiGpZoQwHapZIUuPQOQziYal0XuQsz0dgBpof
iKGvawWUf3Sa71aDTB4WrfTBLyNyghm+d5C1g4Awb9huiv9Ul9sgoAvkyCRXqfvfgJ4xnIELnCMM
6zNmFlI59Y1u/lVOjKxlal577oTIhHkZsCQC/iymOPiPs5s8UfEmPV21Q9YkjNR3Xb+yH58aFbXH
wNAVLOhLI+ZEFs+neUk8aEP3mbRCVCot7TD/H1vD8oUL4FZ15MGer8OcjodGK1SGg2U+DXihpB7x
JLhM163rdRLr+YhhcIGVi44ycxwr75cQV4U0+jCDxiPN8eUOWJb26cNGB1FZss5Uxv7bYmFsQ77S
Rjn6WMNxcXVBoEgJhGMYlfVwkThlb7OAMH7cDsH0kTxjXadbtUhGmxTInH1PXLO/yXr6E3y2UeTZ
TbbzgkjQQYByMkMYtmbw09pokn7/mLrOFgjzzuaWtypXfQaNYxxSGl3lo9KIvCMp7nr9eK+h4eT7
c+YdOyxHxxMYJHcFPkvgDwfwGBaX1vpUGgZrhqqFr5JkkwzTHrGm8jsddMu2Z83IOlVzeUp0t/Ag
/xyeQhl/pjTuhYYuKG7ijypbNkurjmVSuKLOGMr7GaVs+38ct1VGMgNELCayyxLnPsJF8zXUL8Hb
WMRUr/DTA4Jhtz5Fj1HE5zJhvgVg9WAv16GkN3nOZfAPRNg8Wl1yRBeb8nwxRMB0i3oSHXJ2MlWH
d2gnZhwXib2Cn3//x0omPvzS2gS0EOzaVJUVGdB0A3OUWXYuoVNNMcgiFNjDUvB5sOMtRSqgSk4T
A3B5E13DDZQfArSNep+bAySjdedsyGaSv51s+DNsc5VNSv5T/47Q9MJWWfu4hPbaGl7CLlVhlM4p
Y4Lj+PPQlUabg+7vrJ0ITVf3gUAfwWgXkGsOkzSvNvOM1NGyrejP6d42fQFjvP6zEdWrlttw1Uwq
2mKWkbkYCLXzycvCMm5aeD1WgZsPCfHEdJtdD5cqd7SIVEAhHp5K5TGXzu4e5jlHHTigeplktr6H
7twb6WzRDljzINh8mpnsuENTeNwlU9TVxYC0j4feRILME17hOlch77S4a1MoJ7+8hrEOcMRqKsMu
8alApaEJ4Kq6/hdZLORTEASLSCK2lXqC0r14BD9R8aSqQEZHaCP201bnZtABKOsrq6jhUX7IaCAN
o/7Q7lRSPLpPG6slemCgew0sf6FSrvjSPXYYC01rkJpF0A1pFJ2+fBg3GsblNZ1PeLvjXmozqsbz
8lo22yUCLbs0H/cUPFP8Vk+qiwPN87XYk+wrQD/eXUSuZRfKUL/+fi9b1h/xPScskUZDSpmTYJk1
1vbPgboqJxq1vYcOHJV/onK1FAuq4uK/Sj3NB4s555qncm+70hJpReDOFgaMxhOuqishnXnrEDEm
B/Bu19+nBfbEpuHwf4am9eHZCGLBRh8DkN8KUU6t7mYAVPQhBRuIfxkxSAE2pFwcN69Six1Zg50p
bwgUHmKvQswysbY0KEIq9j+Gy7GNT1lSgWBaMxVSbRkjL1k1WxUknlhqVfgBpG28uVCwdpv/+yKW
hkrhk+eZF6Oepn2jIGzqZIRjspgg80XxbZ2X4AmUTGLWPJXqJGENanci+oTNV5W8Vc9TOPf0ROmS
UbpttKE874vvFSR1wfzeoEQ9lP6+70X36tZLegUeC0lFPSVxgmIKQVJfFC9E6XwWsGOitE6Zw3Xw
tYxMOtB1ewjNELZffHXvxZXV8IS20wQ49Oy6q7jwJS/dgWomZJOJMPpMKpLa8141MNbNkEkb6p2W
RwJixzZvO3tKChDC0Cg/ifQV3nEdt0VnvRPZ2gV9qveIS94orKdTHpDAfmpxAHXFSZ1TtTZusvOB
gXmIkNOdtPl9VvzU0Inys+FxLCI0JSvRFv/MSZ1U1HYemDX7e9T3j0+tsGCPeUKTzBF27iUKaXib
hPY5uxz/irzz/4vCaJf1mA/pvNz09AJfn5RNQ3JTyfYoWpxzDfqMnDYwGxClJQqc3rbz0p4pTUYl
omrN3fJgmOKgrK028BRGVNlnGLfjXMOjCQvuLSVrdC6gQvXdLfExxFUiehKjJfKlN8zDRqeQmSTQ
uS2CuibJ8i6sEIaXqdrhX3u6mw888mlSMlAhaiMlJQIN4WvgcOZYeVULQ+r7oCtxI6QJIiHjt/TV
OuP69LDLyQh9SZHaTxxEeo1DW1leQ5FVicdkyjj4g5PLeHg2dH4KDVhe/IND2N/JgMj15lLO+/1s
AuvxwHpLZDwUCoSsDEE4jrz3k2QZ10gSHZFKKIr4aUA4to04GXjWYIWKm7RLVI62CwQ85yuqbAJv
8ObWMWE7aCbJW16ArHUxj+pgPK0vlI7QE+NMblD6+jn1paCa6WL+rTiTyw6OlUFpmte5dVSEt2Vz
kR73CTL6ysyx5/MCEu+2Uhg+5yj1MmdRyvWuzIMV7gojWnytBqwYMUKXvvM77U2U4KXn2AEBhV8A
CCQr3n5s363/xsTs3jh3goSZbYtJAUrh/BDZtn7dXwsbAkrGDvT+96rqDjG6vRMY13wUQ8BoNVcX
Aa6+BEoHSOwfsHNugfP3wO1EC4NZuD5r2XoNncj3S6Bc/o3ijsySPVZ5Hon1ILPa4bK8hEu9+rFY
epnOgGFq0+kwfPzeQRhTGxdkfk/wmeVpb3PEA5G1pZ/8Q6rYoyL2/6ZCG/eQnni6Wa/8lAgd4ziV
dehNGJ08LztckjRphfHfCZDm1WB0WQIIN/4Xm18OlJO61VsjgIoGoPmrZOX5PCNU/deEzGX9CsHf
6AWJrGWhUa0ZkqawNTA4WUc1VP86/EqkGljszBZdvEQBvhIcE5POS746rLYmxACDz2cK09SJe230
PjABIx3e8iGFuLTgX+vJo/Hs4w5tPZ5E7TxdrJJ9WjIG7v4UDhEr2n6u4dDEZKaZ452EF058AOvo
9kMU6arUPLEewG4+3A+tg91l2ZAFyk2cFvHPf9d3czrANcicYxh19CPfLoCwOXlEhIkRWUK+PL15
I1a8bbZ5uYasi+eSD2JV34UUlI/n1yNG/WfuGIbxQ5FrqwdGvnu6YrG5NXA+RcwymX2wlZvq4uBi
aj2r3Tc0VJoCyugvTEzkKb9LXI3Df/hzHOzTKQQa8+sbqyHRCZ8TqxfvZIhUe9xxAoXflk8lJ20r
AHkWSGe2yujXsQmgojQEj4vTNnOKU1Y5hh5qGWxGw/o7+MzI3JyIKpV+w0IsJuMx7r9OKWDZ32oq
WT3bpHOJeoZ1XMjBQFB6PphEgljuAyhNm21DIkc1otqF1D8IIBO2H0bbXEDtQWXKlQM4r/v7hfB4
q9FRb3eG8RPIniOVtdduWR+8B9BhT72gT4i7ojCY61W/bsFoV1MoC1GbvTqlLBIgGEK5gQWN1g3X
W091HjAtWCDyjwRCsNiuz/EoHBk5Sp3EollTK+lfBcHhydhB2PYgZ2Tl6eNB8ePqnt1ajLa92nsu
0xyW6fsUbvzbj5Y9fcTnrjMjOuWjF8GQjVsNBenqq7iSPWOSS/osharsbVazM4qbORve383vIrF/
PPxH2N3/Vn0TeG3nctWCU3QN6trN9zRl5tAX2J5mRPaWzaz9YVCtCPKzPTx5UcJBoug2xMQ9QMoS
eLrWQ4f76zlI5pzwuNCmE5QV/koKoBr/TSTj3uo4uWDozqYpv1r5O/W1OrkqQzpH6hmAjO64suOi
0iEJhgJ6rNfSweGuZpqtnZHnL8wfpjKca/QU7fauqN+Z1KwfOl+6Fr9MvYncLthEJQExdxNDpxG7
pl0R61QIUP21Anz3CR8AqkYsSCwgre1ccQqi0TYgyZ5P4OOtIsdp88Cm7A/CkwqDPM6aM/rYgmMk
/QWRHjSKGcb+v22SC2N8LL+KNHYk0W0XFCIzL0dATN0FioKaK7+wLfyycqP9xJrB0sTQx1D3CeNK
rX1ZU+GCR8b0YlKGTtGyReOk/W/lODoAK58bMBMMWdHHTsELZH1mwGcEjYE7dnU8IcFQqjLJ32Ek
iCitl54siiQg7yD+leIzr81E8qlhjihbbHQEEB7GVfbpWrZA+L6MDzpSJNYOWoXrBxWR0y0rve7A
a6enEnay73U1KqxhodCEO0Dr2CnCabYfyzHvlJPJpn4he+WrSQ3rYgXA8bK50ZNEKWylM/x2ywic
31kaS10JHkK6BHdbgo0vgAVRxfCXE3HUAqHRt2VQ551E79DDJwsrerXhA7k472KS66ykfZ7ehUoQ
uN5DzTVMbaao5G5xodRl07bGJf9/LycyK+qVYBjR6yX5Zg8JR0TmAcOJ9UBHk9NHD2tXasshfVEh
FdGSfC3vUislIPed5Sr3/wrVG2f/vbtqC9EI2980NhG7us2mcq22wVVHHg35HCYlK1udClXL+VaT
X6U68kenuL4PYt+7KOFo56snLdyRk6mhV+kbsxAou1u5nY/CtrvgODQ3OPFpsMcBnH9pku7MGZA1
bUyIsneUes4B1XxIlsN3N187ALaQsCHaWzn8Nb5lJSPvUQR1cyziIPbjKbtfWXA6f3ZCufle+O6P
NclPAQ3gSsFVvReK1or0YCh6opGkrRj7MTAbkdtSqjD/xN8zDBr72sfboTJNIi8aQzsSPL0/LA4w
5Hj4A4s/CrgIAbf9eX/AGJS4RnYHk2J0pXhWKj91xUrdmzyp4cvdhUSg9d3PlRz71ANWY1uFv+Qf
enukqw/8/8jvt/TK+6dueV2muY7z94fyi3ldAHEBiLOrUiPNStLjfhweukVEdk30JrvdM4duzBRN
+8ffn620Vv2DUJupvW7ITehgprjpxpTwraK8yRRlxdXJrOYP6RuTcXITzF3K05ptBuWaGfpCaArA
oYL5ku05Dir9pnU04srROchK/ZQnJXTTEd7DSrMVRtbtzRDT6Lrzpfka2eup+2OFQVjO/i3tkd3y
gBDV+I+XWWcutKFLuR0NcdHan3+Lm9A5jeuHpU5kITVwAqtrmNCMiRofaje3hoNo5tlyuxt+MTK+
1B6t/iqAwdgAmWOYyRBK/3yR5rV2Y79HfEJTsqHHIdRZboasRBlkh8Lc2VWrAUiRig4Yq/w70oYZ
N/mY8kGuOikbjEIMlaC9RsMZu7cdk0MWdP8tZylbzyfSCjbu7oIR9KLb5RKMxWeZL68v+pkwa5sY
zsoKyeo/zkV7xgUpQ3nFTMz6kRLQdgX2awqJmrLcPLgjp8dpecyGbxnnauMjUreCoVsdAX6nAQEz
1tCABHsa9TfYJZNhIXTPTZA993GCHSwcPv4pdIsEXOYn4ptQNhgbdu6s8aERfBgFWFM1unt9oXvi
XrhKykWGc+gAb7ihA1hga3UYfYFniWSRIAEa2Y95IOZv/JuZKCT+6G5xEXvz1CaqDn/2UZE5DORI
ztvJYPTwQGAglSiLtnrvxJMzth7t9eRF/jtZZlI9SKnV+8eEt9ivnKVbm+r/V1TsygdTjc5lwOvb
kG9/OtOZSYtdt34YfYL/Dh2V49ddboB4DI9Dcknqh2Aewi4hfM17TSjB77k5lL6YzcK6eJEd5ZKq
Azi19v5dvtkFe7ZrNZP5xHA912YGOM7IwEvIuL/5jCnVSf8wKs3QLDFaR67DUjcjwn46xJ9gNDbY
YfngYH1sZkQfVkjc0VL5sWardbcBAkfe6SZT0lgKIskk63C00KUHT9HvfWYHTT8UIrEzOWiWdga3
1kZEElWVBZYxh56nvScctNL/21zIqUkFzvfQQv6oyJeSjMW6YLU3OwLmw+MOruUlYJDe38n0Mgpp
Dmlr4cVrwGznoAoplqK0vWN2P4duzTkaEdsk4KWiCJsO5WEyU3d02WfB1+QAOxB+nAIn+Bo7oDJD
TvxryRrc49kVXlepVMvFH//Z0YFdRUN/rONrA4aB3YEvdCEP7ZTvmnODVa4g8VnwWvnn4XEo2w9y
nBma5rwHsd2QaEtv042VeLXHquS5FYOJ3f72SOZJ4Ex5y09v3q/njZcd3GC1xv3xtmuGFBiTJHMy
bplm2sH8NATHI3/f2/J+xJBPnByf3yhHcs5sWVnrvhZHOeD8g63bUEC7amtQva2NN4SpnvB2kQX9
Wlt/JInh3+QlzlUfc9ExGqdl19HAsFD20+65/+xnDqB1w7s+/bnivypeeFIMRFJMKvS2Lt9JmteX
HFdKIJXsJ36ByqgRlsmTN0N0eZg20Y/l1pUy4eUHdNI/oZXveKIaGTK1U+792H4qh5iAw9CGQM2o
+3Eaow1L6BQ0Tl831VfCXD2uCsggo0PcPhhwn6kX3523URd0RYdWFzrfk/fs0NLBQ/qTnThEq/PT
H46Rej6n3CkV9Z+SKTmKB/X0lpE909ooSfGZr3QG46k6rl3VyFV5uufzmFPpK8A6OmKBX3q54p2y
yfu/CvhTZP+Mx3pqyxRVQboIA4hBi6WxinuDn1lE+f7ILpHj3NvPNNS/dd9DgIuyDxHWYsytQXSt
q8BQddlqYxMugkF8EOYttUiWJulej99+BrCfhLuuDPZJq42OrTKzSd0UE2NzXqu7M0Pvz5s+yo2r
NK5Eg4hVHAAcV1LT61zAIIHpbomFNB2r/cn0HfttqyrD/Nx6b3I25M0bOR75iuhViCt6w9+7BH8M
Gy/RQGfaAtEYX1ojm+DhP4vhQ6DAHMcyXfkmiXjPuRG0HZTsfQmdAE80MR9oSLEH0zL/Y4DjXk8K
+DwaVBXQy5yBEmDqZ3S0simtgE0WY5KzwNC+4534GlyMMZEWn8NQNgitSXM7eO9zbX8HXu52tghU
4XRAk2ku0NbKv26ZVnQt7fUsgbBU92OJLvpsKDp7IMYNviE9V3Fp553rt4CF0AjcqIadIcMpoUUs
1uBDw8i8nuMa93EfdjwmdPPhfwo6xhOW/uqnKHq4V2Y5vNpKtORxnm1I6cSHu1tFaBrenos6Dv92
xO5dz7sxOGVTjtTwUsdqk6l/FpWDuM7Aiqoixj27hjfsnCkrSwa3zlu+MfkUWMLBViNQ6tl1dBfs
lFfBS6iu55uAnHfwo+yFazNXWADRJcH7DogBPuT6fNo/4hI91d+OH/uHy0leSDaCSZo3IXcCD+Um
KUX8ooZiYVA65Y2cWbSshZZ5ZzsCJ91Ur8y/oj+ZDD8G34kwNmexBGojoeNE16GEHsWaxKTZ/Kky
bBbJStLwptFIqI0VwmipWj9M0w/9jRYTVi33u5AD5ij36TjwviSdEntVRsNH3/kg+rz1Bd4ntgZs
7cuRig+CmXT4I25T24MPAT9wigVfcLL6krawucYfgKrf3mH7KRm8/IIP/m2xIagETQsB+tTPumsA
UWG7GgLtbvmfeRucHtYkO5ebNfBOn86C2Kf++zMz2+xwnGt+X/AGTnpJ8eNiUAcv6FrXABF0hSq5
gNGA07bgjoAS1n59PcWu0RA0dY9FJ6/nXntFdTj3LBJ0rVMCs/sfLMf377iF4vD9u11e+YR0x/c2
r6AVX7ZeqlICKDRLdtA4jXZkZp+Q+bLrQS8ol+tkqjVBLJS2SN/BWIBUd4g5gwtDpCxIz4lHqKYv
OZopmcpVpZGGy3F4N1MBTt2ZvhQbm3lmWnTo947pvEIg5BiMLyj/l3ra4IIbPGeOWXTy6vVRpuAE
PjhL9Rh+T8F8MQkwA87dluKb6a46F/AEjxXtnAXjoCe/aplwR8VqaEdeqBAQFQcK8S8uOBtUj2Yo
f2aAbN7HRWMLIqwUQlBRZTVFc9Uf7oLaSxgl+cf/4MqOzsYyG4wH65pCWLY7sIQCGkLLC09Bu1T3
dPZysHr9mBCd5JENNoEz96Tp4MrGzcx/HH6URsumbr/Owo2r2vpMe/spDEi5SW3go+ZkmwFdiKzA
bKxoX0cnfx0rX3iAkrr9UdC0ox+fgEPf6S8CsVjYlNOOLFtPa4zIucwIGSGF1gAqBXo3xG579Y/J
ndBirqxdwDJQ32UYlMO2BiKOob5F/Qd7z7tW0hfOM9K9wTEzfJs8sZWwpdhIBgp7IUer50EH1ms5
fXLYRY2DE954h52p1V7rpqmVMDnA3t/g1i7ygs3YKOajnGyUndAxPej/IlDYr/LiGon7/HHQEuWe
+g2YKWW4Etl+J0unJnAaqq+ilFg3GyVfCFDDJL5hTfm+JtTyOAlAfxWMjEvhoavWy8EiKtgkDp8I
51vTJoxCxxpftsRo91WV95pfPgDLAbjLK28iK08TzeD0sifsZBKN+JTgkLpFwZO5suaxglkclElr
1WJopBkuQS7KBy1Xi6z+3EkwcCc5A47HhjJ/LDW403BCDIFyl4MsLVwbRYuAs55K+gpM1GhuhqQs
YEYyQU1ozsvqqT3SGFM18cvKqgHc9Yr6jonIR6rtxqCK7j6+n5yw372paRGqh7UkYUTzq0p2eRvE
kv1GwkiHY9Epd/8qogzl89hvdtyeAh/sRuzLjzGkN+7W/zsIu032nlw7CDrKwZw+agl9hB2D1aX9
HDyFb6RrhKqf/itsRCSpuycIQf1mz72JucTK6Son4ZR3buLL7yIzaGvo1f4q0wWi+WDITm+t1Qf+
b84qaN5KY2AMGC9nVyKN4NaWnm8D0Ey0D9nKbPRDmTs7IGzZXlD5QI52xcxCVn+aRMRewA2s5Nlk
EX8qZ81xwvwGP3fVcqoozHxVs687RN3VXwVDdi7TTRrW3cilA5Bo8JWmV+YWR7jROcr/oKFSeQ8P
c7Vn91eir6ngpeiRle14D0B4CDIr6j4bN+/AnPkBNos+GyXOxtpHdEPWJEpAUgyHDozek0BtyGTq
0yQQu6lCxHvDxC7wb9Kd+pKTHYv7mohn27BPABPzHw3j8mdDgVM3K3Kww+H62m8byZhw0IB8PCA7
pS442J/ANFytuGKymNPWxd0L7cCDw4RIQKDTGCFYcEgrjHq5XBkepU6A3hhq0EZwOtKKujStuLz3
/Aj8bfkB73XcO5ac+oIGkI4IIBC6FSvwe5vEV1FS+sTZGaMdHq+C1dWcs3sxKO3Hs21Yv7I+0TMl
QfdTV5/Lk0GiWkze4D/W7hxWl/8eMspRWq1DJwXCY3Skpf5YaL5IjUPV+cAjBTMh8nOQuSeG29cF
vH+BM6zGHFXGYh2p0yBIF0tJ/iRZQYaL/ispQxE/0utkkLSwyFgVcQUo8eb1IQ6JLufolozc7nOn
xPIEdObK9QQZPfmYSMxg9gHohjKgrgqr09/vwu2xEaD4WMVXbYnRAvZ09Wp9ETSXUYY8iILjwJNA
+RLLqtq4roRRfWgvFcEV8yDv2x317qVOtfz+3WUU9GInI43Dk5XVEsLs5m1JKSLtP0PyGP4iVjkR
81STOUfm8y2NtEEdDpCy7gFi9x9mq9SlxMe16X3Y9OiN2Nu+wi4Z5pG89ELVXbw8V1KAK82nbSBV
qTnC4bY/WmOd+rmPlGQ4li3xB+YODMye/Fs0prsHwU818q66GboejPODLb11MmHg9GHrtOB1Nj6T
++Me7CGx96+inzgSNlaKyIgJknZ1xg9njxiYSNDH5YTwar7WRnCo15AJe58boe7O9gXTjPeIWjUy
1c1Y4uxcQsftOsB9fTj4udfLVHNPwKRGfyLMOvflrd08w0f98eeupaEA5HdEr/YufZXFpZ1IZ5u+
XFXfv/3zo1uoOjDqFLn8rag3CULuV3WSZpmSKIgoUmdVrJu4Oo2cu929uf9v3N6jgUq1uFdiUm55
sNvPtF1CthwoynuNn82wjrE40FTMf8QBiSNiIzAQmFZrK+G+Cq66yLEp0eAbw1qFarP+vTaJklYb
PtzRKzv2MWv1oVh0c5p/YDab+MgpiTIh+DFX99jpJVfyiTHARodBC81ZzP4Yl03pl/oYNUUU8J3T
zDEvksyllDLySDKu0nEXDgm+B5MWDafbpaz/Yaohz9RBffs6Ux/N6CsivLF1liLlUrc/XCHqzVyd
AfLjFQZ47z32exAZi4RCIw4AoyjMsZnAlkNj9nSKEq0/MfAWc4yI7jVToQvYLdczcfh6+Eb0/F9q
CZQlUebTlmoGQUzpKpcqbrxZaYpFkrqkB+7SWK7HKrTPyh1fchnx3f+oND5U7LFBHf+o66ZSJT2G
4fX/1OcDdsPbKJ6POIiGfXJOUaHvohcZAmHX6tuvpUjjE3pufluvQ1R+PQyKkhaOuKS9cY5lDtdG
kvs5ilC12GIkLFM6obf+DHUn2cU+lzW98nWEimPLIrhXnsG3Mjbd7ylFCoMiF5MtrTVHv1xJctF9
VZFd4oZpgCyTjryfC5oACXQImS59+hGbXixvHqBvPIUon9g878UIdw/16s3mWp0DnCiS6OOnfvLH
7AB5hkmhWnu7zmJ4ukm/wglk56kvNNz+7LOORLV3fSewhpPuXcPUMS6kR9ONcaZgF37vW03S9YsE
nYlFl2EDIEh5HSQyg630CHHv1z1Eaq2/3edb5h0GkF9juQ3sF/CrNhw7QUkh1LEIEc4V6Qi62M3q
0ylpcnSAFCfTttg9Vwqnok4QduDiE3s/NP46zJlFZl4J/g/wBotmyVcaa44+KpZ6aVcRfZoNV8rP
Yc7/WzgdO3/K2AbwOMPmcXpSxqMxLRwq2KfQke923V/Pap5fS20PbkEnCTkLPnVZ9/7SfvTHE3VJ
fiovdvRDflxY76+up03oxLq7Raeun28Qwkkslw1zXI76fcFz7Shs5C0TQcNihPKobcPNFFAUHHI0
t+9M4rMBMJBYQbKglwCweKgKH/gtWmJFHtkoq1sJKmVfnMjsPlW2ebMLlnJfTHJFas7LshKJR15L
cd+yJeSkE0QadRSPeQU2FOYgg5L7izKyWSOQnyCapAbkWcUQNzKQH90PVJxC0ZNqrTPgfIoibenJ
voT0kqx6bZ8vPfBKhTR5OkVU8PYYfjk61Bty/xccpghM5v+UBr0fLezu4+wWjgNgsuAtLp3+FYWk
TSuvim266NqT+vy1gwNwFIuniLK5bxUI9u34swmGjNXp0pfPuSssyK1G78VyiEVSbuhu7V+Q0Hvu
d+UlmVlZxIHkAkZGcDA4z1RzdNmF6R4WqNyItV6Swf2t+3VCpU2iMVedXXlFqAtZQm7mYligSnl/
u2yQLbknBAIfyc7WW7yvcD8CY37tvKEJgl6116Mr/TQ1j2OTQtd/khpZtRCPIZJOj1F7fifj0U6z
HA8522iHzDReX97dLDfhPyMzBYjwfHYH5fL21j+wrEJBKckBVW+xPmCs6+Z8Et9ts54/jqK3VVHj
35O/KVOgLnYHPrnOJjRUllCE7IBCYRU7REOfYdnkmW2w0l2TFZOMsikmN1QIzvNSWskVW5s3xcBG
bWol8Vv0pfwiYNuttIZimpUnSFVUdZ+QPNuoInolzYHbsCk7Gx4DBIIDV9E1quidrFFnuQq9mbPP
rrkdAHGeMOujhNySd2+LXAxQ/tjKg33lbPeJVuWK2onjShd4hGpABZQ5grF3HrMZC8YwYeEap4Kn
r4GiFRV9taFqAsriGKUmag3ifTD/WCybpjKCS3s3OWWqFYpCYmSRMl/z0Pm32SW8OolcXY/fzIS1
vJgzle6YjDzQPbkBdQcRUyzyTSe5AyKsvCfmrZ2zI+lkT/kyEEuRmNyA2hgSEbenwyLfpbx+3uGc
oNspMUm/QVvOBFvz/dacR/dtAgT6Q4+CD051OH60Qs7Ytc8FH8lNuGkfbV5bpgbBznb8lDSicSYb
5u0GUFNKm1uvE/YYVJ014dbVrGumZlhgBJsTeOVJUieoLroWbWR+iXBUSVQc6eKP5gZZwQsvK6J1
iP1vUHZ/5eGD8ndwq86zC+PJVFG2G2AzZFpPxIp+c7nlSjw2blpNZ0n7SE5GSKqcuQraK4lsOg1x
mmcDQWpv2kV5P1m3b0Kz3DDOFnLkNqKCxmiCSG5VpIIkwaHEAK/6Yv6P64F6eRMLhEY14azAN3Kb
kivFPjC4Txs7POHuDHcS0hKJEngnmDBuWL6Gz3rgBAH5fPylmwf5rtWOpLFv0+SHUj49n8UDlonu
jl3DMi12fDLCvtz0xDSDccngKwcRScU1oV0bzIkILGp9LHo+Qv8uPAxSgTiKIP4Crwp/DyFGprtO
1FzygnaqnlgKtr8vJFpEVTpmSjweg3xgFOx87IIOaefgzfxREIzvELSksWCoVnpH+FsKG7IG5cFB
5MwFbxVJzyb1Bzs90IQYm9Lnm6l4ikrA03ZbidiuomnW0P9PVtDk4V+8HAa3njFtDJPmiRVVKg0g
XEF+cbn1FwJkgCUOzL+l1NxTNI7yVGvwFsflYTtx5g6V/sSA9u8t35+W8dFnC8WFEOXwhyrE7Fh1
WY4RHJz7Md0HXOJ13YOR7BiDFI6IbyBBclyX/1o6hP/ecaG1OI1rZ/EpuRBWwHZR5906ZxFZ/QEB
0AA+Ay3PHEso+D+qViizyV1aYn3Lyur/vC2V0YU9Jtv2zW96eZjvwOs80BPmdGJZx7uEqvTFtpxD
i2JvU67+15bQanAdZdbmnomA4ui0KTf/XrJZoWOi/ajgOStAgQi6dAW45O9GtNShkQaMI0fNUvjf
0rBvhipammAxJSjCrJijIEYgMfWd/arrWupc6ERHbWKDlu7y7Bgy6rJ4hlPIlcQ6uJDlSfmSQTa7
7yDzX1uauHduR3F9kB3I4zIU2LwcO8RgQ50+8GGb3SZPHFX0PY6orjJW6FQjq1i5w77WP5MXrgEK
SETcYpvZ9gkSGoiXfoOy0knOvD8cQVZOPVvIzjh8orx/gEnY45uxCuC865T0UZOBLohAQvPmp/we
QRVgYORHMSDbWt+wiZUcxg9h2/1SqDAYVPHZyXnbLWvOHLSaJCwF+zyPG6bFTGakUNd/SA7moQPY
Eam/uWnLZ2Fd0X4frCFYILTZ6EsSVjY/3uCGg4qx59/zxfIbYICw0jQ+LRNwMJ7Csg2sHjPNRESc
lSz7ZlBml6/T1Is0YsWaKpvDVUCQwBurcRQQwBFYpcZN4+jXRU2RdVVs4YNFlH6EZn4E3W69Uctq
n99SV1h6Zr3VWWz8YJx1XDGlF1x0a2FzNZL7nrdpi8f5SfkpDMkPK0m/yI9gK14CJCcxRzmffVE0
c9MwJ25zAd+zvIyATYuMfaKpx4axzOFIjWfyO25xIPGIbBTy8teDfujqbu7a02fokWKUP5yR8aVP
444KfjNY02xtapH0/y6hxPRzctzb+WyuNrhTUIV/XMLHhWlt34P2unygLdiKuYTB4pjE5QuCJBbX
TANCzp8jW8wQBX339fRVqqK3VvWQhzpmzyFxK/8L2+QiZgZ0g/XFvKNn/QXIL8uCOLZAZXYzRtMi
FCMRzoFwSrItrlVKoQxMZ9+qS4fCPa9ojlFFWXp1kEMDnV3DhPEka7caM1JCIEGnIPcn+lpln+te
wpwFLwhVYUwDfB9r6+TpSCiWd6bymuvoDV80j2ORFheRBTHyX5DiSjM0i8lJ6IQb9DXeisaoeSYu
XSloCXfSWFPC0d26YKFXIH1u4+95cTAngyOJJNKMDJQQQXunX5BiYfSOPqoXxL550an3aXS3Pf6W
tdYfsXJe2mghiRqoZpDcEhBIvW/PTLIEWmk9m75q2SROOgWDeiJoP3iscewvaVIyxGNQS9LA6YnR
3gHLsvnQGINrJ6Jv7VHEP3qZP4KsflzVjq5l3gJQJlGvBeFfnXpvVVLVKBGh3zCbdSOuEA4a5TEM
8gsNIpn8Cy+sl4peuh6hAUi+3wVPfdbrY3rv26zY9KtcGBIGGE0zXC5qsCtMMyouBCIW0vxEP2vf
LQYuQMe8jrFYV/SNOdJ2vX6HBTrJHGctnHtu1wlG6+D3R7HdSo7GzcqLxBFdah5A59WWxhlH/udc
v9vvkSdTILPldC/zVxDjIZyS6j5kFw/4FQugHGJ/g1b0x0fS/R7xCIf++3TKQsf5B/6gOr019Cs9
ILjVRRePId4HPdX/bqDNgnYH05CE9rm0thWJrTUieyF1UD5l6mXdRSF839r/NgxMA1Gegw5/HLHy
qhBNTpqX4jzwhG5vwIpbyZWQlx8OqGVWKJ/8YK6pIoyoTXLOUcHlYEz69IBmsbU2LVGCwTfjAIX7
f/QgGnD+wkEpNjLLkOpKhNA7sKwXMqtGHizL7X6f3aX2YqS4Ep14fcqmnSoPxaJq6rhGOfZX6N7K
151Ps1FG/OFlrueq/BhIq8iCFmQmpPEZNDKCUN4huovT1bmUks9MLII4JK3fgW6NpQxlO0POolv5
pRadtgasVpaSfOaDnAzfUczgt2dr0SFN8XZa+VeElGt+7Au3ViRGKX4dsNWYrsyloWazQESIo6qJ
zscLCOsLza3IRtdxdhAgQcUIbJMuWXxcYdQN/XKdRgzFy3SRAHDnTj0BRF1igMWeUinOkLhZnuXn
Q3qQY1RlRGwURspNqDe48Mobc43NWYyk5GIGXKc1VAR+j0uJL6nWMW04NF/AMB/7jMVxQSmHpMVq
WpXaX1qCpbL1PMCrspT8CD0cMGe1AVRKn8amzeCkTyDmVZ56I4qB6bbv62GXI0mmCjNfrgyXGQRF
xTm74o+USKaSuLQHeykytpf+9qSBI0FhuwFoYosi0hr8lmX3DhAT5dzbbwgYXhrMZXiQv9rPy4gi
4NnBNJ9PdG7L0no88US3KyeQzLwsxPi+C9izCuOrqZHRc+asqucJI4eY7yrirujtQpjCE8whrwda
9ORGekzAcasWfIFYn/kcQv69cbgRcRxASV9sPoDTOJndNOxm5EzEgCdVxZeccolTdKOCSwXyezuh
DU3DGUHbw9mwJ+mJ9QE1nnGduQGqXUNHZf6myXeGk/vq+ECgwOhu43gulqgXWL6hrnsTUkvKrwOR
Vhh6MyfE9U7yrPQNIjpE9JNygqbrpQAkWzGkGtZnxuHgkpqZEQE8vVjXd+AW7i7nIWKKAg6XdjQ+
zC2ZLIG61Iw8usGm+Y5+c577QaMTIAFkLWZxiNqUnyCxIPl/6fxynPjlAcLx3qu/GC/AHyWlHtRi
1kFr1R/2QSVl9vjLusk02KTa+DtTsgviXC0kyNpJLXDZAHB6xQNs/5XXpDv8MEMIGirdeyNU0Ho5
n6dp1LGvyC4UZtInOlfg/vQ/Rihm92eJDbMKc0X/QjX3QyCR4vRD00T8mD+LYypqru1lsbg6AGNw
dxsEfuZtuNmBCVwbWJw48ynwQXrz0cbgZ2fVIlmkqSNV3otJxIGRloZhYboxexgCjj12TwFmRr5C
DXyUdxq6DfBOwCBOyAAil+9qToMAGJh0oKX7NMEhMPl5qkFUb3vWHrfEiwv5WDHbz0e+SAUF1NXN
u/kjOq/9FkAjbnTL/XJ9SHjaRGKa7UeySFawlrxTddbF1A0bVx5f1Pj9m6S+b9b8bKggeUuoLi1y
AeDE9xUgQ06l2kWsmMgpeMRFJ/YRbgZ401Mdw15s51S0SKJR8xRl2F+KhMpby+dV1C2Lr3wXGJER
ofjgt/OdKts3006WY5pjAnRkQKJxQQHkRHVc7o1XQPEMHOYu3QcL5WC876/q8AwlFd0Upeik2ySl
6odYU8cP8rJfxjZp3W3f6DkEgz5tj+gcHB7kbffGjHzZ11bzEK4iB6TVu7PNSszG1f79yGJiy0h/
41zDvukMfUWBdRBiWOoQ8MLYRDB3qugYXWLXx1Q/qgJeRryDZpZc7bTmQQtxf9FMvhrA8BQs36dm
Baj1ov7E3wG4wZ///r6ucjJMjJD5pGfne3mIh9xXB1KqwSXDpX6FZ3VRuuwNDUW0lyVC9xawcVlJ
xUDiSGyE5lQ3zmuOcnh9uta2LFOnBdgj6ut+WvadX7Ctovk96eWRi8pkdRzj/XjI93zIYOcpkEZh
iizKMZ05I/QPNrVRDtSdNasoue3nt7DMlkSzM/Lzl55qWaJ4ekne+v/wgJeKQT4EZYyt4eKwbI+J
QMH35h70JFu630EbRtF0VBHneMLc8A12zZBzj3K4FdBJWhTXp84YKthNGRwm1tE2JnjSTYGS0lKv
g6xtDF+rW4DvMbNiHORjjYk1RL1sUOAxBNv+J2U98oLi84kLv77QuJOuyx9M8rbFnfRZAq+85hT2
ZV35VR32PZTfLPmw+isM0xdGUKcxqOVMRgq1uQMmPj/sMrk43lLNqWypEVVmoiFYCulHkzJ8OBza
klstE+pEq7Vy5enawDHpILtaixxeU6r3KQa2i8yAqHVHM2eWhLh9TSGn71xCvhwB4qkGyr/gQL6K
ITZQnyVORFjvjAJuubgAuJodgwJAxRMVHi563Uru86lHPbK8ivX7Jd2LzXEzMjt06zQlVOD0H1gr
8+SbtUyu89HfXJR6lSQFMQqL7EHgNoTqAiSPX2pOPxvFioXgoDU/RvhcssGUmS1Exh3t906Vkn1B
HNPeKQJ0JZVF+TaHai91USSM63fU92ovYWTDcU9O7f+9gTjl07/KFYRL8YHHXg+eGbEzQQJi7YbF
On8EamIsSwmdh4KHm77lUHv45Mix2L8CYERaFHElI4QlJS7AdtH1CyWeCI2RDs0+TPniwXJUi94w
YL4aAkEPoibQW8EuszyFhbPN/LYg4nfeufscSqgu8QV+gOpq39WwqldoFIUAnGxyRJh/codO6MBe
qBVJEAxDYkF1AkjZAz8HE2kqYZMAoJ5xvDrSqWDgp1snDbNl7iDZnaYy58RNYgVJaMZ0d7BIcThQ
FQNFavUCTgRS4Ngam/E7TuwCafQ8yCGstoXWK9GsnDMpzoxft1GVFuV/IEG0+rO3A+O0bAoJdiaa
fTDczXFVV9SC6wHboZDLnPx+iadamqKHHMxGCCxQerMHsu+r62qKmBax/tO9j4FNkcyVzN+QxsUk
zoh4fVDE3jB84yiRzYZaxp0/B+Q66Ik10k+CICXamFyjVerV+D1c2odhCLMMMoONrh7ghWHQU2OS
4uwwbhdMnPDWDQ4qYt6drctL9xmwIIa05CeEPRoq5yoiMwGVcMbYQpYSTtL73fLg5SledGkys4Kh
oSllwSr9KK6GQkYrOhTuJ2i2Qt9kBAo7RCQZUNCfdIPkHlD9WgMpKpY/xGKdO3IdyK99irIWsEkU
KcRt2PwixNhpJJ2MGnTrkZoj1do0TBpa09zACRx1sS1drgpj4eQ2+4UqmvBRMJ9sb//zVIfZK/Oh
3w1wvL+u0gMv4UdmiWS+U2A+AYn0UWBZCSaenOJC4l2Na3pn3SCdLWTinS1ME7IXE8em+8wwpzou
8PlP8A27qdmPQvqqnYS36PETMITVMcsI7Vi0LFrmcUVZcqI6BojzuQAilboja+AzgE7193l4ukXw
nzU3jaN3d2JXwV3vBcUc/XrlPL7I3HpPivXePd6IMBu0hri8Sypd+srkz2J/AQIueRFj1sh3K56W
UwwZzZ8tZXWhtoVDO7iqthO6Z5rtLzd3DJXD0VXOkcVnpVaKp8poG5SZDgtdL7aJOPWX/cetbf2N
u/vhbGrIhUBvE4LR71cX1cBJiohMlDCA/NXjYhq73dHkfDPhVt4Bxsh8DCMf7dWD5M+CDa6G4IJP
kacNNl4+fMd3/wCkBStkiwwJ9Sd+aBdOXQFSij5VBOxKIGpj+OFjokaJE9d9mxNk+WCvTZtmB3lm
81CP4+gG9fUJihHn0rp2znDbPLTw2cGNwNv1XJS8cQ/+NgT7SnCHD9aNYcOzYmkDGi1mx+XfCLji
3jc8MhrMgMxKqAQwKlGRJkEM2XnDzpTu43XF2jwmWGtKd9hnZY3ZHQ6eEtOa4JA4f+TP2moPMeU/
/7qreUgxJkEG6MCg2nitHKk+FIueBBH61DcL1TvEm0DAl6Rn2JLzr1Q2T/EIQ1HhHAkWzrAMohcI
2IguYwb/ZCLPrTnGj4FbHng3Ifqwc9b3Thnej7cYv5pJp4fuXD4G5lxb2l87KblIQ4ZfEPVL2hlo
4fZOPglETI5Q70gQoWuE/gzRIccSqpnzEqg4FnGBnhxx8ED2lgdgxuu6di2t6LyIC35camXTUEUo
uQ4D0hoAegeUIhvURGmyM7aulTT8Q/t1XNz5+0tcUT4LLshZIQdIHkUftFARNntUmYIFriBC1mFz
nyZ+p5D6LRZmH7qWyiMfKjI+nQHEaePi+MrRB+h7IeEjr6zPLZzi6w1IBRE5TgqbklUQU3Mq3ZEi
P4La3mXp5yLewsqCrz60116xivmbJs9wh0h2t+c1HB5I6Y5GmfUYWqbIVwd/dF0mI4DF84w2HwiQ
RQ1PJYuTvJkanacULTHffL9MWh5CioD7hFwEtPyoeVufjfoFxLndklhgDWMqRnieIYorjc9cMjfv
OgTAgV6QxDxmxx8qnXhVekJWOa5v+ggmcVUiLWBQCVxHc8Apqr5PIWJnxRbCxLKe83JLV7EH/wbi
VyXEGyyMzuVYE0q0iLOCb3Z/4koGd/9F+aOlBQi5Ip5kroCPb+nH+9btrF6Lg7HNkk78+NxdPdkq
3ePhJciZsKe54Zx+/Bh67ZDvVFf/W+extGYZ1yWv4ZaEu2ThGNsuodK+SQt15RS/biI4zR/myHTL
8ub/NprFEHC1ktydNcXissH0H0I0+p/be68Q0/5shVxvWoIRZNYRZqW5DWunp95tuOAhmVfw9KUs
O+tljxFbKKwC35OeSRyfZFnd0PJ1kRlTXXx6SnGM5Su/+qOEE4HV70tedEM7TUqLjE+iD6BIt5zl
6I6S5XJUNsH1Tuc08m/4X57izwHfZWHWvjgz9bdI1Q+k6K88Pmk4n1sYGygWmzEeItDbuu78UzBD
o0r9v5ol6g5qcPYdbjqvbeIBr6yMjl9+bRDyrL8IaklS4dZ9DOoE5iPiji5le1SHgN8QwyvTgIe0
86zEZBy2OpuwqQUBRIEO0EtQlDiDbKsO27M4HcrJYRqaMzewDE4M5TeEWNLCXW1xS877wgovm+0Q
FU9oOn7DatnDAraF44mcnwcifaQtLQEkqqbCGrqD2LkImlROPKXWYcIMRAkc53+b/npHQ/eUIDRh
jcohD846sIPo6Qey923o2wE0V62EN+6fmHbIFssg45bsAl8m6EZOQVfEThWKJVnUHXEdUAFzcXVo
E27RwI2v0bNAKN/2iznco1fq8SLaHLqyEaTBQXQEosXTmWRNVhHHB9/c3s2Yo8UaC+N29zVO11TN
n1kU1rWkFyhL3rXJDSg8GnyTOpcK7Ipt6YtVce6yZ4VCOg5krCZ3HWwiGi7yWe4oWxshAr/125fY
whdt+jed+7hCm99omW/tNrTf3qtMhgnkgCIEo47+lXvgzPpJ7tpO9o8MkHwnuvwP36E8CZfGI89X
ETAVn9FS03SjyGxN4US1hrbIXc69BalvvCC0r+Ju6fJ1SmHzS07HQiZd1Rvz8CpbzidZQjQyDgkf
eUbekNwyswSyfEZP/WGQRc6SBSSWf3y5UKBULKzOdwi8vPdsa3BawKYCy0JCqZeHCDZpqC6RwPwd
WxSSJj5f0atB2io0grSB3YBrPKNqIErpCp45nnxOgx0n8R9sThHy5KgXUDZoPVUvzIzh+ZzWj6Jp
UlSdJAVtHCBl4fpGxOriwITN3s3NvRYjGwA+uVvhideOm56+9p/qSKwiN/4jcjOMBXWSuOSLNpzl
ds6XkEHE7NiJmAFdyW03RdBfcABd/LiyqpcmfmBoihu5PQPLYO3pYM+OgqdXytQvB27RojFRlnZr
slR0c3AuHcUZSc0udwj0JROZTb0JrC4IeaXtQ5KXSzKlxo9Qv0HvvdA1/lCPiSRKGjbiwKX03Zix
5VLAto+6bkt3HhXHa1KrokSD0tqUzvTMhgGveZEeK9+62jC8I0MNMg5qR299FcAYcDWIo9swZqHp
FBPnV5Nt3G51FB+DJ/p2DIsSWfIe8iR4pDOMt4lRRpwcniclCciOov1p0ooPRIT099uXBvcEKHNl
k6cVEWcagxbN08V6UAbm6f0Vu/9UQUzBUeq3OVqNFv/hDRPF3FCmXASpYs8a4DoXxq3BErncdCP7
klBp4U15kPna/3NrsI+YKc7uLFnFWNff0VrEtUixutLI61mN1PceBAzeGzULtK2qdK0pXB4eo68G
O/ZBaHQZuk1Ri9pdDdYIEjbiKBYHcV+j3Vs+i9kpAmDr1+kiKMI9trzC7i22DFeknHw+45ItmHqY
I89Pog+OtYNOsQEyhfckQVGLydNwqS8COcbGFdVI74gtBTlzzLjQhzTZ+l2Ld5EPJp15/2NBCO0I
QDirorf8JH88mKbcthpwBwXVck88Nh9TICcKI+FSDy6ZMJ3T4DJcy/+NvxXG369W0MWVwQTTWfk+
p7FYDiX5JTRmWSN9sSaIeq4lrqmUCYjowKdZpoRDUss5zffl37pW9LatZb0P0wUj/Rrj31zxsy5h
8nlwNQdyXkKy7cq1Xxl68GG0bgz2SWJKUBjWZgGibnrwzEsknVm6Gy0u4bA9CMLU7fENe9Nh7F4Z
6sI1RGWpTTZr8fxQJikPmQxXKotdwoh3oXa+PGCVmhHBsnRpFVOVhTyA/35gH6SGNNF9FmeG12CF
1eUKzrND0CnmPnETyZTTCe54S6c83s8GUwfxQk/FIgnRMCykrEkJQPnYUlFxKIqeaVNN+Us/GJxl
ZY9hyVgMWiArqHr8s4LbCvvG9nTOk4wuuv6AGv6iDVRSNkVpfgheYSxYphZm39bEFnQV4w7oE99W
8uO+yFSJ0XDZ352PClCuIlASHpx3gtK1GxdE78h22CouKZ9859kldSH9rMH6txWB8aAfIjjlR6Y3
VjMqpDlVM3DRezWOgXYOi55XXjrwZ5Rcf/jd1jdK3D0q3IQhKVllNv0xGPVLhuiHS7OhxnULcJkH
l3u80oZt07N4z6pjffQptGHnRxmgqSzaAiNXY+HfjmZ3dptau/VzLi6MeSho40K+CMx1wzkco16k
b8N4C1hPtBtSwQlKZq1ydAocVnO0malVF1+TALwXNRsOgP9IGZG/wRutnonsoyoRAQHzVobxbpcu
J7oOBmgq2WGyAhNSeLflESVbG7dGrmK9n64JPAymjfg8gvfD6rUPC1myapTpgGRsVTwNb2u72QK5
k37yYwcwZE+4VLRdUho+I/NBmIAANcW9TjNqv+SdbTUxVfb6U3W7sqZYR3sPwz5WAtNJ8QhYDAon
zTGB59tDV1b78ZtJZzImnss6o60K3ir3Q4MSlpsDDpcmkgCYZPZDu+YuSxK1FWl4edjG4qPFdvM7
loI/T36lWCn8RQFsmWr+SDFoEC1IwI6zV7IQ/YyBoKSCHe6B3JFcahimHLjh1eXf0neGqz7Z2aOm
h4kyMFO6ikC7o6IDBK2DBGhS2lzdHK3ZnAbFLNIwsVm+9CSRD+RLIl3n+gLt6WwbBJJdp/SlGZt2
Z9WuLCKiwwahM4nQjK24I3hHpJwjhzN0B2JBjomptjly0n+VFN0NnTkQteaAnv8i4bJrP34zrtp1
f3ia9zMlfpJo8rT7Lr/Jc9rEyFosjmSLXm0z9X8JqlttpZkPs/xUwj95lpd2ZWEBnTSKGgn0DIVQ
7yWHGMmsUCkIfmracONxym/TyJau4eknUxTYuCGfFRviCWHWXXtv1MHC4gRfkKIlPqss0lbDTBzK
+m+ZSlivf5Zo0FtvChHEt8Kfl0FFSiUdVOFKOVc1N1X6+/SLQp4drhTjbHFQA7eKke1fI0RaHQ2L
g+ORS+7tHYKov8dMLr2sDPqmD98E8AmNL9vb8cJGsBNJ4tDN+CvuE+xq4MOw2dxN3JTXOPaRuLn0
7BbuK0OFqGCb/EAh8PkjQsuxIBdwefOELj2Lha5ZpFJJ/BR5ynTGxiLfSJiaFY68CfOKS2DFAsC0
U0qE7/l8QKvfGmYdKNTOY/RqGfr4+I9Rpd+cUgx6wOwz+WJJmxBcKkygY5MIltcfvL2Dmspio4vd
/Zcqss4MfDnGcskJQBmLcevZvxHJcg6VhMktarHVUzOOmSlfUm1a3CsqGwzDgrp9KMt1X8BvZtrA
IfUKD5wevo3UBPzD6wLIFYHvGQ64Rx2b8HktfvL9t4kCFasAGnWFBEqYZBhFBsy1yX/POCyoNAAG
05jnUhK1EHuIqBitXgnEznRy2LdVOa07N/3pkPCE6mOTMyc2+x/TFeouIWpuEeyd+tCbF8XETXP9
QWWpIk9yt620M7csED7g/Vko6W9kE9hh1z2YzGO4aXiuzDWS23/hyp5v04w0NI53HpkbZYl2Mmzk
gDYrxTZcy0qt82oCcj8tFTKa6YhBPRw28reneeDMW5anrs1EQMDh9ygcqyz2L/uMWheqyvfucxzn
94QViGGB7fLPPPd2uxbIXXvMlYYWnVhMmgcMHTXhddvZMLZ1NTX3zV5ZwRoWz26D9B3ac2eS37kh
x3nHEStY2x4Gy8Qsd5LGSsgIm7y09ejyHK8pSw1M4g2exqaWmjNiDXdMyEgXILgQuaKKX3hJ69nb
MRNxWqjBhy4HBIESVevSiwnuBeHYjkgocLufgbVcxx0IDI8m5tgca3a7PReClLpMW9anOQOR+uCW
0ZH+4BpSalJJhguPEH9WJ4K69uWqrd5QECggQjz+n7uyqL1jeiEHCRoIDybuVD68IJOVftsSqCn+
8u7fBxIztuF0SICXqqRYvboDAlPcYXZ5U5x0486Wc0SXiqh33YaAbvdQJ2uFtlzRJUmriYqpmFaB
oURBZKP6MN25/0e2V9s0OenlUaxLWpF98mqm4WpcEdRnoUYtxO3rEVRsk1y9Q2pZXZwNdOEDpBFm
5Lk4tzq8VRnX/qfu/illXdnU/Qi6aUsQvNAVH5S4VA+1QBagZncVV61mX/BpbFxRyo15fA2Zds5D
QvXsZwaSMUpUwIeVuq3O2FTDR3BLieUliHHXsI0xsC7VmyAgeQiCU7Okg93mzZIxHbRX0iAz9NDd
RV2/TqgFyYOUAnTGVXqvJnXXoIEJ70U5dEF8oZYid1C/ug9YWLsRQ6sQUb3hhY6DNxjqWq5M4isz
Tb7fzY/6w6P7pPY2oExoEw5zjDgh972I81brBNbn6Ac1ebYL++4wfqZZINXP1PsqUx+QwgXYs5td
RP0+iB+JsKolaZmZP3bSB7RMkodsepVcCjbLFEKdcq+QQiSC+jBhsyHQh2ewta1zL2Z5M0vV4iaz
prYhr+a1LDVQfUKUSauSSNRupRC7D27rsXcNdsDszv7MDtsKV5tgTY0o8VgsEbEegLJWH4M2KQqV
9M271nj63B59rQXg7tOl9fJI33b5oQAvSe7+TOWJ0l5ElGNB/WrIL9Zs3P+Jik2uRz1WREidGnIx
T4njE1g+7qDWddssIJX/cskB4/9vvg6k7xwYhcTeZ4VQLqjEkokKXQmcjuLKumpgv+rOWSHEF9VN
xqFXbcI5Ik49bx7JQvDrfWJOQTeBTTPXiOpA3zTViHt/E/ETspvwbzybg912bWI5ZYzuaD4vV2gO
7K3G9Dj86OGpjIhZpfXjBtl6MmwXnHBiBLXW4Pgf3Y1/oHdhUH0KY72dF0zswqyGmptW6bmVuTf+
AWt2AON1jkTsmrQV7i5kJ1J1r8jcQrbYs5BAKnfjBukrKNdDvYyZpntl+Jlbqil2ABXmV2V8dS8k
2pGVjMkcurkdZ2EqLvO6Qk5RUx406ZHkY+e1BFJappHeHYoH2+Ie7VURJ3PZVE6C3RNB4rfahg1q
Iu5x15dKs2zxoQeZ63gfPwITtsS7nsKJeRZNe9sz03tBLXLbKCfS9mQH6TNa0+4cpwDGzBNSWOX7
RUoVo5XHq4P3pKxltixO0iCv/MCOVMtY1HxEvKCuNdH5SPMbhVD2zg+JuUSDgtXuSJ5KrcGz80Du
sBeB6iRiHEdRrZH7BgGQSGdK9b2GVQrDwO5sY4vc0E/DOfFO2rbTpQpi+Sf0vu45fGS2+mDYdOga
b8VCXOSAsk3LF8TaByhIgFCraUyMwbNUCHX4+MxgKkEovqgZIs3pWz1Y8VL7bNjS7bcIC/sLWNRA
5z4uZibHrVSV1KFuZ3yYsTA3vUy9gUq0n6yIdAU+S63IKrpX8OEcHnI+/JmFukXxDOiCtxp/2wsF
oSt+NOqLqXY+l5WC2B4T+qkcVrV4DpwlGPRtF1PwJRUPAxmYIzxfxvQDHAKpcxCo/2QCZZSW+uiF
/OfHDdzw/Xr+ToiL+0boFVVszacABLzETskCXOTjDnK65BMisRTQWLOr6l6QSV5lF7C21XRQcdPd
xyNsSo/9AhKmJycGOyV+R/mbYJmCTVnXxHiM8u11YCuCjis4Jhvbg2CRMxoQ44+Y2XXGNPA/po1o
JPz0Z5aaieO0FL1/XQpY1zxZPQJ+VT9YuVt94WH56V9l29dFzijVpfrl/W+R5LXKPmSXYY/daKIL
zdZO/pcw6ndlMKbDGuSU5FYtQnEUNujfZqJ+Se7DY2VTVcedvHn4zjxaFUF8Bn3Igg4nbrz6H6Jh
EJYymC6yUKHpwLpN/htjxrZf44tkkcLA4nuCwOLIfckyOPFDUj0RGxna3ahw1vJjewoNF/O4zelM
mHTS4z1cNra5yElrdqAap1SWPYSvqvJSgZnZ50RZ8JjK4mBcAeaWnjWG4FA+2Zf9+uwACiSsa3nz
DZdGVG61aMPqQhtXe8G0jizNABBX2aZPtKirXw7MVXpGh/ZrbNThu4QmYEjVIu01LhSloywn6e8e
XQEEhkwA7XMr95rerwidDsyvxiIX/SzuD5Vwmc+6I/RUhvEVvq0YtZU4f1wH/rZvlm4VIs2V5UiF
LN7lEYVUQmBVoLnRtrVMa5yFrAGq5j8lDdTz6nWZvn6Gw3k5fbLdx8Fi+Fyu7D9F9rnGlvUZ2Y0J
eU4pNWVIy8SwpzFW7jeA7Lr7fpAITquDF6gFyaWnnVtMpYjxOsEliyh0vYGcN5+iCRkR49olhtAy
QZq5TjjMOjlNG35tsxZBulwaIgp9biyPjyOV2hbshE7+1Wv8zPSIiRl9dubzGYkXH0+2qd3szfOh
M2q7F2Jzi53WQlUn6Wm5qWwXZWHG0NdiAA2H05GdMQTGmCNv7024ILahFiFPr/OBAXPJoKjqHL2u
AA2l8oMzuSRE07YPw8n87Um6PFL8luaBT4WVWXKkC7bdTZ3M/ifZjlITLBefhRni3V1G4HB1JF/O
7qAiePZOadcqkLDeLkGF/FS3e/gQLBgOK5YZWCskPJAq1NxrfAJQT0HJcXRu+pmtLAbyCNsIh3gw
ohhNlWQUBStLZzKe4iEI7F8wyntip28u7mITWJ1JPQsaYjx/p1+65lRy2MGEjlduPHsjLP1KkmBN
f6wQm0ShOnWsDpR1T/gtZiax8HLaNvHswUINsIuUg5v5ov1nnzSJST0qpo5S5haqF5iY3S8EQ8pf
Gu9u43D5EERGnZKyeYsOP4Bn60S4suO1lj1J/ct1SrWrA1qrQuP51Rx4yoaNGe3glsauyOqjqanV
naL13lUUfpUUneVtQ+1sat2WwtEofE9Fd1UfxAVQyJfZmUu7y0/wfen5jKlnoKSaDp5RiG4G5vU5
Xwti/0L+cdHd6Kpsti0hZ6Q5HnLjfer9EnMloZoHmvuyCdgOWyDjAxYj44si2JVHCLj6Iry8GQ5I
Z0T1u8MKIQGQXjuCunF6FSB0OitS29MqAZVqSMHvGsi8Grj0W0XXPrQvmVRgYsHSoLBKuno8oGqV
+mlszvw0Y2bswU/9qEi5mYlgJeBjl0M8V+XFTfZip9RHlSqff2Ia5WBIfQVbl0dWj0TsVX5OA2De
ep/rmbLGbhgEivEx8xHc0PHYGz1lQ5ogIVRWRsdvQmQtQMD82IUPlqJe6QplcF8WaYRWtHihOqgl
dmwEfaYicxd/E2kk/z1jG/CXjhb+PyjxUqxaw+agNEG7hzFOOnK16HbC8lg9hr89eBjjBABun/Qt
1TY4xaOOugoKjGu49Y0J3cd1ygDyzf/3FXpHwOodKEaB+c+Wq2B8LZBj3uRZRxYbQFAUkucsCPtt
ur8jz0U4nhoM7O9VwHiXb30+/cJGfYwRQIa/nnnQY5JExZu3I/rgnkMTrTu1/Sv4IeQwWVHv+z01
6D//n7hFOnbZaiH7s4Bk0lOtLse/2uru2e/+nuBX5EKPBshGxhf9HzeruTXt/3IZ73GyTv8kTuOX
6kZHUhm0JQcq7pVSO+D6GPLfksd2nMSz/7Q7ayFHpC+mGWZ6hW7KLbqRlx9TkrmiFe49nILTnzjg
qWsJO05PJR9hw556T5iOky31AopXcUDgfT2VUfdBOSlsOOXIh0Sebqcu9bHrNKrivKdiowStK4Gt
6T+7BUR8SmZF8MaA1+Hud1nT73Rzk972ho9yrbwZdLh/4D53fQ5Mnp4l5IpMu7RI5hubMmxlpdXr
wussF3RPqwaU81UOjr1NRxdMmqtepbX9N5cmKkF7dGxH1TQuK7u2EIKkjHwTn/whq2BpUdAKWfyK
Mytt4y5EOqVEKwbilsUY3di/zQ1nIxx1Wlz1GJM4Bk84/59q3ox7KBaDYUJ3gjrrR325oyBdD6yq
t+R8gwCTUUA29L9LvHtMFUhRalVO3yNByzv1MocHUqhbtYJMQNzyPLsTlaJKRjVj/jvUzycVUudH
SHg8Osspo+bhjtphhEmpHmlDTkslIx8QJJGQW3iUgU6OcWzdtr29ECHvOG/dZmGNTUtelhzV8awd
eIKnPBvXajlLv3YTszk/9Rdeu+hCsxWVvFODFh+4jwcKGKYJyAO9D/k2xkyicu4QwmlmEAon1U65
KPCQzb8+iIWNus17KaP2FSfY0EOzRSaLxWKqCZf+b5qqEXVVFJCFYFjV6y3dESQ8EmleOqCjEb8r
hU3gGQ6q4vGkfmUkpLr8l16zGceIY+2fHcnSBnfIcjBv/562AOvHHkBNkJ/lMuHGb2CE81Gt4mmM
AmbqMKGVa58EBbrT+FR3HMVRCZtspnZmChnvcPlRu6pBEsWa4kAvRhzBA8Ok3kX52U88a5SNInel
eTai4hI+l33aJE/bt6rfdxPBKbafCnApztMXEVTPGYn//3lrMXLFglTzstLxvZ2WBVFA3zVEX9N+
5310Xzsa8D0SRzm+iX5SkUjc1oJzGbiBRhhxVbPbGDkvEYYO7nm+Yvpt6NAWLkZnt7QGOizx1+oX
LAAtTZhXHCchZwj1XVFW3/6/hM0PrJ66KwBH/eh9ld26o+DJjm5Etneb6XbMTi8vrAT1uJrRVng1
+m4rUUSbADgydcZUEaxRzHXN3GFqWusKOQCSAAnTGH4qArYaS3uTrDugHDKnSePAegGnwhy33CMM
268rKekdEl9BR6NrOUP3Jsq4/Q9BAHxhf3+aPfvqbbr0UYUhtiV+c9ZCMZmoz1GSzNAGtKjRODam
FrwUgWz+U4n7uhecLKHdcUeQbw63o+YFCwL6w92YLtpvHl55ktqTSkbf7iHp8mYtaYdSRvtPKnRZ
pf/HKC25KL2swJHGpn88vXQoX6lhEGxYkqGSSklCVSrLDmUipP38Q+fRhEYG7E7edVSXjCI+2dbe
UTQbt3Kp3ER9psIdpPVf+1T13SoM0QwYB4nvgyhPvXKvqGcj65mfpZPxJxBJs5lk+/ZD5iMVQXQa
/7Q28fprTxipoxrsk0BP/uLKhKY+T9d4K62jMf/OACiN0d1GdR6zJfFLbFas8jnKS4P5zlMCbyVr
huIJLiXHQfm79G9+OaCI3SpOWJHvsXgJxFHdLNodp0hqpatCRGK9wWt5uQNbIYkKu4cwe5CqyTiF
JoBUE+guliqvazCVEaqzeXThMxAz3Ot12y9qEd/wq5aOlEJWEDBfnnIia8SDBTL21+5ahhcOG7Fp
3aXGlrE84oY4pu09lu4klGp2mH95GpCyjs6ERJh0wfFxuIxf2IkvPSSusI0oNNEUyVJcL2NaxlwB
B20ljft7t2R3Ams54e9f7Q/glEDNzr1i1WA+J9NX8S0HglKXJEKakBfJUAO3iZhdsnsTLzgnb3rm
DB5O9IpmnyBs6J56psw3GBfoNVoXXwvOISfQexT18nM3jKf4QBXzlMa1r7Dufk0Z2LqqR/silCU/
d2vr9RUqrVAcwkKZrjY/sayYMfbvLAdmLzz66UfClK2F61Is9Uihq1A2CgMh079JHEXIzHjGB8HH
nmulSBOV/ez1+TW4GP/t5a9ysJD4gH/iwMh+PERnOobX0xojlEBke3lNY6SyA5q222FW2Hk4Qk4x
934fFxTkDURRJRSHBE15DNDxIvGC+pMfUhN4PcDwdygMOS07vCSNHGyBYmN4cA1yua31Q+Kw+r2t
+80rz70tZlrVM4FnPVV8oBDYK2I7n2W+vU5fz2ltL3fA5YUtPop8fEoxKduOVlUR77ZJ6wDm8DCi
XX/FkOGJwRKbzMNxDNNf+Z0QUS/MzDvHGjFKJogU1jL6pKvfBAfpOUAivNKga6yIqidQUZaFCXDp
lPtDchCaqLohP1Um6kZFarXxMMcIomQ0N+yhmyAvkGjVZ5Da1f9KPDOXHzzvJIqABLWMElSn56hg
zpNBZojgqDENqBHzSi6hFpdogz6j/aP/Z2jTc4I7sT5vnEPMDKJuRbQ+AeA7kQbMO6EtWCdKUWrt
rWJ5naI9UeisQOiju+VPY88Tz+xJM27Z8n7ZrnMqvxCRFWuhhvSeBlRgEWYi7C7I8pTZjkmcwKR3
sfun84o7ACUZn/D7Pnh7LXmHXZsLf/4Yvj8Pysf70R+4q04CbNwyvoSbH5f/4VKsBrWA4ed5byOn
VJEeLdx09V/GxrK2sgJrq9q8Orr0eF9IiiQV7XKf9BTEV/6CJAaqc6ZGCk1Yera3NifQRXZ2wa5G
PzrdY4p/U9TWqJVxj0GMhUDCS0kBZFIiR9Ne11Ex8SRY7G4hu7fAs0TiAIsNaww/ZXJvLTWpmqOY
MThRUlwdvmscx4yHgR5VOGDhAQvZaix1MqWwP7KNoZYY0/tX9JKj09bnM7cwzMZMUUxxlLXuC3MK
vjuG3t0kN3JCDNZoU85tMn1MHSg0xf5s7rrFh9Bwri1n57FFTB/OPxL/TIlLYC0OwEN1D235DXZo
sFcM4l2ueFf5OIToWnbe+PdKvJigmw6oNG+7VWPoNhKket4SO22bsxxUMPc91Hte0RmvG9bQ/enu
vteGvS2uHGbFdWAOLCD6C8KVtDq3thDB+5i3h2FlwBkLcEajmpzOiwG6P47wS26I14PyMeew6zFr
A50meYqpJKTXvltbZdMYfGSw8gP2ejeqzryohm8moDtdO1XLEnpIH5yojzmCQYYZBW7e/7AFbXdS
FllD8P6A/7Z5N6LCeI4xZOWv/mFv7xpodEq/4VCKONpz5sAZom9qnMSQU3Pe/vY6rs0JqHxsyeqO
nGyr5p245DQu9w4j0lpcfctGLj547q9RYC2TryY6PHYPuhcXpLobCzqFTUS5tpeTERC+1rrZ8ID7
y6Ts4Jp0XaG+rqvlhGuxY3Az8SjrU2nLm5ognuMVJVvkjIx28E6CX2UEljYaiHgWoLhnrRbeEJFy
/WosLQ488pxLTxjU/PjP+Wmr3wPqr9DoK9AgtHJ81RZxMtkoSMtvvw5i3/UENNGgRkiTbGS1y9bw
hpu+ug6UVvczdewqCm/PP7Qed1nsmGHR1l6Zex9fKzzbHFcE6h0oScBH+StxRpfy4veU/9CqLhiO
5CyJJbItw/VLhbHZ4eJNOfU9fMaYAnlf7h3ekUMm0x8jXHHhyEYwf+Wj4xDg5Ja0Sg7Yma5ZCvGF
/X1jSraZfLLFiFeM8HccMVlaFuvacppcZiHxClzt/Jlnln0kMhDC9LlOG4xvknidjPqEbaFeiUVR
Tyn9gAmn2p6hahCeXDZ+CnZDezLat5XnL2Kg6AVTgJhnJUu7Sk0/Rm3UqEQiMvry+AMqd1S1k9n3
LFWJUK+EpJmUyRSv6QajExKh6wPeAKZQ6FYXEKY9HQbH9bJVFzdalXELmPD3Wdq8r9Y7a7tDwiqv
OeTgcf1vXpDB985AhDAZfYU7/PfMdgkfRx+i7+5tVNCjFzACaOoe86JUGjyBri3N6Z5284XgZlCs
WPFWJmU+4y9SQl10je8NxITi7eaMAmPJxOtbgzPHcoNm1EpM/4RgK4O9Wlse2zifj5M56ExP0GYT
d8m1MtKO8+VjjWxF2tDwGADWjfcWF/LdRhPyfLdBd6ena09FaS1MsRw/2UwG+PH+aEz4N8tusMOQ
H2PbXwnpJL2J896zkcXN2yggs+L8Aua5y/2pdWz9yFC4upjTS/SwHOQ6eVmZXjRBrYttPT0TOII1
tC4FJXWxKqgyx54sTdwpZlhbNr8IBhhR1SaNwoqPWezqhFhCz9az3TmQq6Ty/I9Cs8V27PLaHRi8
0Oo4BTR8QGGKrS707vneUE9+WwUwt/9TJwpC7SexK/q3DoP3wUNJfKjvcvFC1XNJzTyNIxgKAdT8
SfVXW8YO+p2yJVIBZTzqWpe9N1IalMuywDARN5A1Z/fS+f/lZVm2T7+7eRHDSqUXmCIKxr/Js7f1
yGNS6C9wNU1O0W+tOgNOXSny8HxXMCjOdkVR3CtVBlFU1M0whOmU3xVg/YgEOWhUEVX2a41DHcmK
6gFzQCBYWcN9Utz8FCtvwmuqS0UK+D2Mm/kfdmvj8slR9u+5BFRlwPtqnR7r/AL2bAc/RgV1YiQw
W9Ppopyd02SmQ5ihRkFr48DLcYAMDxwxA707gWW4eeLeCVfrPNGt7UuEpRe0RH/xyr8X9SrRBfO5
2OM1xE3ZD5mzcz6NTbbZnQBJQx1lxzBJ/gcWr/OwAbPiBn29gOxQ2HNXDiTC+uTnWJ8qh2c2I2qs
C8ZQSI9iA1GbaHD0VEJ4TELWF0XgpWatnBBXvGPFigzsZJ0CUOUZKyhJR4+Uw+8WtgCjQOZ2UcvH
5W2exI+S94IYktL+U8NVzTj7w8Db0DuPCz5i+r5/UJk3zjZ7ylq/QyNTpdwGccgNoVplEacLaGiW
J9IF9/2b60/V8ZESWUulGPtIya1N3QUvgleyTJFeKFK+Mcy3jM0J0S5yrAsTKye2y6KW9DsG6Rsl
XbBQXhdtnlG3xG+Dpz7TaDqO5LIdC1F1CarN/6k4aZn7GksWDdMXeDJnq+KnkXH0f931bclcf9qu
oP81ypc9kY1r5mJmSCiSIlkJLEZiEYwmUKebsGr222dyRqzJpQVRw7ivKvfuWy/xd+lL0/P3OUqt
RYixuUD2JbDyJ9iSkPGsUIU+Q11T89ouKbRshk0yHG7/SBSMaHGsnetUFLFdLItLB/d0gCnSi1Dc
KgkTfUMpkWu9+Kj7gIoTMKzmEgV8qfe6zc3udGoLFzF1BlqHRFfzqa4KWbouZTqYM8sd2bkO6E0o
7Umu03W+P9dsPYPKLkDrZIrTm6I0lCIbZubhKLwtmStG0bdzRON/0Gl4jA2cMNUNSxpw0Bt4guwE
vGkoOB06g+oGTM4AL9yXkLowX+tnn/KJNETQwv4jHYGLgPFfxUeP8n+VZEKOS2yjQEVT+gaKJuIh
QdZ0K2UZpoBmD7yp6gaQD22y9SqyKn8r7XCGvlW1zv2htZBIecwwKx4iZJ3sEqPrTLsQSHD/f7qH
yige3hQ51ukg0ZymNkv+o7dmz1qbu3hO/PEyOHGBWSFT8HY8xzlM2XGc/iXoK1M8O3DyjS7h1QEq
yXybrcVWJiei/rCUswEgsYzyGYVhWTI+O7lgyE75FcM9UhNL+9xd+XKR/FYrRN2I+d3V0irkwvTR
kax6JfeEDUkxSSDN2hrifXzN6vIPfmAQPkm/zltWlcrYDYPZnM4PF3VIJXdjieb6cJg8KxhsOgN9
sq5ur/b6F1JbroGJeojco3MiGDO6FMEXgalUM+reeZutzyzfCSqAadtfhjSFh63kXBnSbl22nouw
pDC0k86FKnZR8e1QZytNaDAnBFe7VW7+6AeeHRnDI74LluX7OyMvkOl2lzuaoI5fPZkDf9xggn9s
r0ZO2P2FCszkCUxfYtA6SV0UlWM7L3W3Js3BX/OlK6Xx9vEMESJU14oAqMccuZQPK3D8SAAQ8rAF
zsC6979AY7B4u0HCzNYM+DXKQ0qTIQFtvZS4GA5FuDMrBtUZQJISlXXiZrm0GupK2TENvIgD/krK
PLF8/SGMBXcuUYCxqPhIVTMttZwLrFUuWUc3eTq92uueqxli2JIoWv8TNx+/CihFqNTZol3kIUzu
fShYJv8YBFKapMLURtLRM2wsu3+vSAipI+6OwcmbQ4eO5ghgnUkxI/w8ABhFp6nBQ6HZRa0/DQaj
oTcOAF0/PTGjDsqIeCYPS584m59rIAqvyHyo/7Kte0SKdyiwKwInR6E44CUZF+4ZNhdoUMOYujeZ
DSbvUaRTz7BHvUf+P0/Kz5MOR7V6TcAbhEL/cwpygmXm2iNrQDXergQeF7rlG6SXj/MdIKC3eBrD
f0tPSw/BbapswaOdUiJv7LKnKOcXf6i+haAgXj6ZqaHqbwO1g0TlwWTswwmyryiMQ6ArlWxyijWn
GI8QS9lpcayIe9JIyUaT2ktIHoSPADBl3ClrwxH0Uulb7Y/JMbjM3aP7irtUpfOeXVJtnEOYGqFI
4P9pV+FTSO24F98jxBIWqW1GnJ16yPMuFSHpDLhwPlZTDBezt1v8VSSVs1seh0EFH1l8bJaJBkis
0Vrhgg4ZQdl4xnkjkj534Ap0JK0CA8/LT+FXA+8v3aaPmo3CqkypvvANV9/uRrhXBNQDOanRhjfG
1cD13rbpVBzLG9B2XVGwmBRST9DKLW8e9KfrYnzKr4Gz6j8pPHCzS10eSAv8Brc/LdRMwUIi1NPz
5XdDvnlGaI7NX6AMiE2qxAzP2hSX9FPb6Tus8v7s69l0DZeOn2/4ll6s98ahMnHWbpK/qoztX0wA
gQ8Iqvhg0/U4qC38AsrqOV8lPsx8kXwa62ORplwPRnVMALZKtRORTEqBET9ksi/q9BVJA3NiPc/8
d58GVahuLJrkWUlwYzxZEL7n9mS/bX0fQqi4TyQFuojS/uB+Qi+ujZ6KYS9kOoQY7HYDNIYcrxQd
iIH7m5JHNRX4W07BviLQgoGgmN9PzBUZAHjpDyFhMZdnK5AZ7H5XsmjupY3oa1jPBR1sy+uMe3QZ
FxmLfu//rSGWmbe+u15EPoR/dqIrGnjEzbRwvnMejaa4Cd0z/MLWlbmO2ZZ/HpGjojimmFLoPGZc
4+ugsBl3zcFFnE1Pm/tD0FkJnfCiOmR/qjfoJZnSR/m7EiQrK1C46AscsxGLzK5Loy1wmasCW+1e
pNO5t9L61+x6hzLDIwNnTNLeZVHsDrs+hNAqdRcsJ9fDZXMfXqHiiTtHGOD5O3gx808hmlEpbc2g
jVHWNGopJeDtR21ZXsDp0gjMiaVZPVh0Sx/fUi+SmdQAA3WzWZsugBzKw8g/YmGuIcq6cW0qNKYC
4gFslxQblG3vbZzgy0baicjDFrE+uS9ez6StJfow2gP6firKkGbbH6jFacXhXmLGktP7yBMw2Spg
RZUFaML8/h3R6gcGpK75FfVGEt6rmTZdtS5XE6I0X+MmBbE1ffDzO0zTDGnmIgQRL+pkF7OWJ7mj
dgNkveOOO12xuy2wjLs3pws0JFuUe1TUMD7uQ/jChVFH34l0Gfqwc495Xw+S0t99olhn61vGoOTw
qOb/8Yu0y4Ecev2HBo2dKxRZ8aKf4vHvwHG/WGnadp7QNMYgeCuUspMhG+87kt4uxJpgcX9v+02Y
57FP6XFeq4NY2wy/AQvu5U0waxFt2l0/3ES2OfhiTpyb9aExYODS+3dYXD5UZtmDbGppK7xZ3Ai/
mvaJjr3BM7QUpAYfqdiK1GKa4vTGEU9KaF1jVLLCNrc07MAIYqVb6WdLdsr/JOrwvjiAkkvBtkrC
B0D2lwa0ssKTpEc6Pu48Mzg/Clfe2jytQs7sahOUlFLv92WQL1l22TkI9Yw4Bdqtsr7zpeX4ZExG
qzqNSAH1toRekhg/+8Yb2tQAS+hOoU6R0sD35QiRaBmOiQ6MQKZIGWuDAxn+B36PqH4ApVXxlMBf
Mvz1ZQ3ckRvtjOza3i/8BjpkfrdZba4ip5jMYI2moY4oqCr847jnCTlLzzv9qLZCGxUiYOsgOBI9
UAQ6lINb/yJ8F96rz4t6TDRzCMmQNl9yP+0QHlPQcTIN3lHh65p3AC9U+DH9suCKoLENqwdAoTWA
NPbmSVEWPr5rUMOfNvfGNMGv+lgWyzWUiojnKpIEfBkBoDYwQbWi7XHDxqi/n8FOrLaiVHBKuYvo
ou7PSCpf8frnFnNk2A9zFDGms9SWBoj6iH09etxTaEfBggK0G0BLKa/cfuNZwLb9it2vxPihhmZz
krpnOXFWLWjCb/OgurklV356LZ6M+h5iCgQSOpVJ3waHSrRi34VNUbgCw3BRZVlRiwBRqzS0vrxX
w2mVe2UVDrm9CVW6iop2sbg31BUQodCHMSmZsiolekmO3OJUjGl410LPGCYXQ5SUB+o4xIELDK4d
pBJtukyn+7bWJEQ9Nqi9trHFSJdIvOWwW/iPkkpoi2IsRQlPDDHNXRv95cPzjxrohivQg8FnzzE6
ul2MfPe1eHD3/UspdutZfICW8I8S4k7dgbq7VP64w3Qxx/YZxceuFQyl0NGL/GEMScipd4U4EhJm
DSqLzP4vRZAkHsYliXbOh+Qw2QlvXNzL62hxLD7iw1fDWU9p5kA8eTxLCkXTizdv51NS6/Frz44W
+HaV4mlXshGsqtOsWwKTZWXKzWNvUQbIyuOzF4TMkEupe5EDDNNs047iPZbGrcS7Br40XHBj6afx
abqghqAljOi+AeDAyHiniYnUhTVN+HMpxtF0jm75nov16VWvkr656mSkXY3aNciM+s0qGd3gVq49
Meg/I9GDfgDFhw6I8DUByrrNtSSxd6Zcixg2c1a8uw3I2G8IfB/rURhQHxiiY9n1m/nJlm5bH+qU
L+sGYK/P5Rc1oqSFWJ8hlnIhMiDV7h6VyR3Hd3GN3fFdrAq8ZznRqtUNGPEZ5B1Q0bBS6RDKCuUP
lcrS5qCB3Jes4sqc8morfEcVnPG+x1YbTLNQxT13KcdGYvZRBvB4z6u/gZKoYP1u6k/3WMZ5iGeY
elCQTvBSvYvNFJAZy6i16+rFcd/6+EhH/K/ZCUgb9upPCHBHak5FtzW12Jw+ABjJIF6FCaXWnSq2
93N4lGds3NgF+nNa8Iy/naDdKKyh7NyHDGpJDfVOgy4rreFneM7oQqlWOv5DzK+pkCe+wQ07Q8FB
d3HLZ1h2kskna8tBrJ0IXuuV0aKfdXnIgJ6CrArI9nt81InsvUjqQG5oC4BIhl2mWrkc29GWZPk+
rp2JiSZJVvEsB2gzHNLp7nrMTwMfMhH2nl3m+mgsfz9YdrAz7XDKqkEqrjgYsb0FKTVuJzRzN76p
6+40uclldh/28+9Snu+74nhQH9oSuZ9iZC6EgSblCZRPvLf/2E5K4QeeAiB5RpoX3+Ar6nuX8azK
S7IqMmccvSy/hV6dvKsHy74MhX56CsMTcYRwcnIfaDabbfro2vt7AEZs5AUmoy1oHOJhSbx90dwT
HWE/rnV2QkrQgRFUkkFHgityXrJwpMjrxLIpKgdvdnMlVM1aa1ZKyGZ2ZaHmG2YzHjv32s1p5Dy7
I5mY29J9OodRP8OlfEFzifKkm42NnioF8Z1SRBXgPIzMsYMkWdVsdES8b3K1XplhdFHX81l3plhK
m1KSawAyKQT1KWtUKsFSu14HV/zbd80124yRRYjvvVnCkzftQJXr6R4e6cKxhIOkAKymPhjXctdg
bXSNHayrO3XGh7kR7oCG8txW58gKwbCX21ULXtr8enWr7FIKtLM3eiC5t7QLFnw1qw5EmgIAWVkD
rAop8OMg6Xjeh8bxBj1oPaOeWwb1iCu+ZOHy/VCohBLXSRKiy9tp6vOVc7AcuUXz0PpICOp3u/Kv
kRltrLlz0y42MKm6uSuJV3I9pBLSo5GPvxftuD4LqtwbV8X7KX8VoL/bFhcTWowsNoT9ujBuD3Ci
l76CVadeGjPhwgNpeJC42nWXnRJz7avepTMPOQv2RWxIY+5ruLqtbQnNMapyVCLs6jiAIxIEDUNh
kCh/VWoXut5ub5mRl7TJi8I0KgTa/0zTybYJQLEB8Zof5mxdnkqWcPsLPLDmQ86+0P8low0V8N/l
bZKP2sbKK5StOQy7Uw/2q1N9TD+IkZLQfUwFM1siE821YIa74w45peFTTxO+8WfAubHiicxi8fAM
OFytx7KwzVFhwwrs2WWm+mK+n4EiXw1SfOQ1YopDIjDEVCwwpRnE/EVNnZz+A1Y8OWu20lhS9H+Q
3g3FjBdF1avyhkwDI4MWXCkPNV8WrMEL3s5VpFW+Mco+yVB6TrdDdHEHVPbsRjyE/ITtuGe0cKku
s0mxdbp8LzOD33+TZu9rPt+ygdzDGcVB69qVJnh/hn3PVoPdMNwkNM5X9rQo+CcDMcPx/xL9iC0C
pUTj4+T9teDRHbOJHycqfz5n698GXUc6JQyHlVR59ZKLliWTBxbUK2rZHQrvPwQJXAxvMX1CtU9j
1XaIHT7UbOwRm+w0kNvIwuqgCe+J3WXZzxPLcGu1u6W14l3eem2RgrTRVaS60qU0Fa0njXi66XUx
1EFCAzquIAgKaouCZhzRLnZ0G3sRVQ1atT7COuhOzsefHxskdnAeR6MYQFdFQeBFdYZ93HTKKJFp
/NYacrmxnoQT6cxPHuQxlUwXvGarNsCzt0m/Yg8Y62Iuyi9BCVXayZeaKsS8qt8G2ZKB66HGQpp6
4WYjBgDcCkM6CVQekN1i61wv33jyvkZl/+ZGc6OesU85bB6O584bl5NRZ1cOnYLsf9QBew5aRvvs
xFyapFGn6CnCsqQtMQUQnbxfyuS+jDZ0UjyQMl+ky0595H0Bq8BByMnW2gGzgMg+h7yUUYyvF0fB
UjVKAui3LzRJjOcdW4Q+NQY/nMdTKmciXO99HG4b2STxA2fijwt7ofQKWVU43EmvVK9x5nQ+VaTx
cclnmeXE5NqVPkDDsQp0Z2joPqOurVFt8L2DWz2ddeKmq2LP+xM0+FseGC0mVyhjMOcI3+Qk9y9b
1dySMuE01KK95q3iM2pqvucD5VnefyeN/LBqweJtLsJx+p6o99kGTkG//UFT1r+i8PXexRauzVJi
SnRAy8tOXVPTIo8qiK8h3sJ2vqPIlfjMpcHqCSXt4Ulj39EUJhloCmMH6OmOcsM7WIOo2lmn2pow
pKRuxVH8PStsHAUWJtqEjg98+kQ7JmVFc+uIVJmZFuJcXSlw3Db0a37ZRZZpkVu8zhn11p5o1c3b
YqMejwOO62QHLHHGO2H7SxALC2IU3azjv11QYBXqu1qyrh71gqDOf4q/dCN2mSAObkn8yFrrBEg6
31obnW4z+qUKXsfY15aG8Chd94czTWWVUFiabumkvSXcCC9GXITefc0j5lR6F1iUwdU/BG1SfoXx
AsD8FiW0N+kpbxQvH0heNBIpExMA9PBVyul76meWJrQYNe3BFuA7cnxTnqYDwglNDfLfyO9lY4Z8
RoiJRpl0L1C6y+XJn6dDjvIZAE/xV8qGp9XPohotmu6wBF8NqUFHSoRBn+ieSOa9ilPsyIxioDWi
uED2iJiHbwLH4zgN2WvmVwgFm3e2BZP0F8mCKNIpvC33AAIUI84BnxI8cj/g+kW8di6+q/fYYV3c
ehlmZTCCJIVD1DfiV+lKORU+amoscuWXA27DuYFKbXUusxjHINsREWeaIomLMWY5Uk+TGCpjaMZu
9Xise4MLxUo4/iOYaUe1hYVZyXW6Kv4o2hmeBo7kT8CdsxC/QdJndxmGWP3MQEVaMqnpKbQce1Wu
sZAcsibMhbctg6sBu0wHOEtDzbiaEFvcK8RuUNVWBaaqVqWQ0sqZmMTCbeavNBw1RskpXFTXqwAy
u8+cahHLtHFTd/bQOjS0nzZHU61INVMZpk1mblLoSWXhk2WBSZNzDrEo6p0eC06Rcqav2Lcrh5pF
FfiX7pBPICLLy8ErKSKM/DcqkWxwZV6D/1CHdPnF4+MqetkMfw34Xcf9tlGFe/AYb0G4qZZddw2d
GfZI7Cq5CMBtdY85EOobqCuCSwvlm/vPZol/gmfUv9AQHTsR4RLFnrfr62kF2NNEijNVNdMqnJKM
BlcsKjYCbLG5HLQr88DkJPi3BC6dHDiQ4KF435rbD1BVZ72vGX4yAWQHx3UCfNU4aNO7Ps7jmxgV
WS91fHYcrPyFM/QhNgMX7sS4JH2cip6pvqof6QPq9vTycjLNPOAUiSSS/SjmPPQlwSeD0aKolPEU
YBsV+5vd2D2pdlIIRoqkpChvaXMpZQ9A2dPBOlA0Tlby8dhKacWD7K4nlnTGk1IrQrby3liuquW3
mJhA8Mqcjj6/v7oIlqy0k5uaAjVBSRW4o6Lb60l+K3o5n4r1DGE9rWJ130MMb9TNFvxgyzha2OKh
cjN1G4fuNloEcZhsNn5cW89wk2UN/+wIONK/iz29WLH4SCojzOsQjJoA8m2lxZ0qQXpY0lQjgeal
n2uEK3CYg4N2QnOH5yyFQLkG5lU/MUkfcgkoDUG/CCb/fYvlGIbEUfkPQ6roAAZ5FLzQoU5+NSMd
iUx/7Ra96d6Ja4khdpiKz3d7eQ6RBPGDrgz9DlRTtpUtQEzbdTz3opPYjenDNN34UAhWk5UGMezv
pzoVC4OCgwXes7O/R2R2AmJVybFrs53c5a67d8A5768kd5zcvdLBhlWfxfqHHErqsG4PLhZHqns4
UR7sPcqk4Q1scZ9eQc4WdTJtpPNgJq6Xj4/clfp3CttJcZSc4XPI5wRp12KiXFEV2Bc5/TqKaYIR
+H0z+CaFRNbV41PELS6qK2RXOLYqCBSROtbdhNRTVH7596ZZhk+bY3yLsplk+DYMwamxL1q6D6rC
DtmTiJ5Vl0PofnoUp4tjaUu63be+CKf9YN3bXqzxvVOInMcW3wYthSKYJS+bghUJCV1ySOiV0NHj
jCXsABmhEYy9bPF40ixQf0pTIxViFcU7ro5vfWRVzIJhA0wI0o7KtJO8WpTFAcf1XDT7bIu2K2h7
sQ/orWbz00vgiKu21ECOkkzqUbD6+D84dHFnOw+3/+yDh4RXupB1mUX9gRL6D9gsdvqAtEQx4Gja
Y7cCxgkv9O9Vo7ZvGgCED6g+4EN0Ay5K5rauvpQEPDeauMETjVuRfP1keUVD0aJRHGr4XSFxeeOk
/bVNOw5n3puERow4T779YrBKmcQsDvMZiYDqfpSFTF4I6qmX7crrG2/E6IcY5rOfCiLp3pvSP4qa
VcVXmQiPI481+Yo5CcTiHuPXFT4aSceCQI5+Zip6S4DZOtT0gq1yOpQF2525UWb4Uu1ky7xuCJnd
fZw/w6Btisj0U2RzOX98GK23mMCnBsvmp6natJgWEeoyrZW0B0Io1vWYZg9kUQolvgdGuQFc3J7M
Y/t/M0F9tV/oVwdIshPWDfDUdlqfgRK/yLFl/SoWpCodBolZ6E7o6A7faMMlrt7/wYS+2st2Cb+b
Xa8ahP5G8m5m0b+kRjI5X9CProXpBMmHqshmhnoqjD5nEpSU8uBcyNMfvi1/zGf2RLLcAXiEQr4I
bc00tOKgjSu0seknJZ6ANrkM4nOW7TEsR2H1xomahwWENReMw6Q0kWuMXqrF4qeqOJknxARBQtgR
hF4Jo9iaLq+7ae01xmGf+MWkgI6f5eyWWWb6tiKTq/Nnw6FJXXABNi46VcBDrxcAPuWyzykH3Jg4
gItpH3f982CeksoBdl2yo+dM1O7M9Rk0+4aCraBUpNr2VusLv+Nbpa4B33RDoo5MIpU6wjbEuQA0
f06STFQkFainW17Eqlmplqakd3xi6G4MYC1tVB83960hDUQeOwfk09ZVK6+jyQ2rNXjKZ+6FksO0
OXnSteZFRMt/ur4vs+NJxZotlM9PdoNA+VyiT+90STPQdYsQWiKlZfAgpEs8SEQm8GJBWA4/s2S/
piK3IR5Y3q0baP0DJF2KPcJkNdLtwR+n3szKkHZ/yiml0w90F7Hiz5XTPn5xJeCwxmYlNUesqqHn
XUVB+2xEyxvv+ay2bpg+vCq4FhB9gU6KqxY85iQ8nohV3DXuaCAxqu/ibg1rF7KB6neld8Xn6orA
uWdPfNJZLywFJhFG3cbTOJWItT75YD4edKbJEgg6OW0jZ52cgRSmCeuupdd65le0f3TJ62k7/clO
Oy+7oGtG0Q0IsJwA2BosyNhpXDFOiqMyN+X8avrH5yPl2OWObDDKHKF9/7ZLWthNsdGg1PwW0qeR
Dyx+xfA/HP093aRQ7f6d3Agy6Nr68FBlg/EG8tg/jRork40dChWibPGyupKfYaRJAf7oXWQbK09L
ei83beYlutFg9bf4Dqmpuc9xCQ5dKUkdgTYVEFDhtxiH6F5bkL/hA5wNbd1C7SldfFQfsWN6VB0R
bhyzVZ8LeYBcyLmTIUFHHeVBzTLIFi7jKH/6Ge11ILr70LsPtz409JiHzWM5iiGn2NYPWQqqNJJb
IvhTBXVL/++pUbs28dRpWWG3sZnhDoZVC5IllNfWbHNuJerH3wv0hXujw+UNXKAsTtquDJcLb0eZ
2hzR5Zfsvk8cEeettVEbjdsx48usm9zZ6WVwIm1X7idp4N2kQobk2/CQtop/xPSfCRU8eucMA3KW
I6uaDKeW+PB27pGhzW3tBz5Cu/40m8J7Z+Y1g/44tAcSJQIiiYdZcUQrGB5q8t/suZMJNsoBAblD
Dgt8IJ3AMChv3C/UBq/yFeQQMRpmYF4CLVIO+H89eq6dff6/Fvr9+xOLs+qVPWyVLBYGvfu0brGF
j22PlC08JN4frJirK6zY6UiYffCFSKBNGjb9fISvWKLeQ4+tv+Z1JiaYifdQuGI6FgwcX8qKydEt
G+sqppUGzxobfjTggzFU0vwP8Wmvkut/aD4mD0mIVKtsJe8RJo5aqBE7I2F1r/I6gfbR7/62fjT7
Tx2p45K0KqeINIFylrxrgEQwrObChpNvEnZjO2u8F/pOf5juCzCYZJXUZUlvn+7NCdVuH1T6Gmyf
S55jiXAmRB3QWbXBQrsfl0jgW2fDHClBg6BQwmU1IUtfXlB8a79oBqfM7FyAkShts2lUCNRyE+eG
4pZca6JgpL2xW3WeTMju9B8q4bDcMuVFNumG0dlhlK1tqDSZRPO2yU03ypoXfIEVwtCyGfFELgJw
FzG25ykCc+Bvy3RQIDf8F3GdbKvzY9jybxcPul33vOLHQv+YiB4hmHAUKMB9mZhcE0sVA9VQJAhV
eXMAIQgMVQdckCZGKbOi/nWX6ReURmTAVHWonVirwDn4KieGLfoMcaj5MIpTP4tEN/8oRwyVG5Q8
pBeka02fuxOIfRBIlwNo+OQ+FZxkJ2rQwqtNqlH2ExUwXsfDcF7UNUVVDrAPGdkjoi/nhr0w+Cjb
MnP3uM4GnIMnYmgkJXMYZnfIkv5pFJzT2SEx+ZxUOvly9bYLSOXzNmL/F3umGwQHwCBqo/q69Rhl
NXaP6jb+2+a+cYK4XH+8yAFaVka+IX2Lfh3cR3f3kBxA/ETYry5tl5X2WwYZud0F76AfH68D4i7A
zL/IOQV7KglLlJLcsPxidLfNhX7ulY9Lg3mTRi2EiUlZ8dieBUBx6vMx+Rig/XYcFZ1HoRI2zVDc
vuquiSee3zHkKe/ybeVtFiF0ogq6eFrqHKU76gH1YAtacZA2BJJ0hh1joyLoZjGiF/QkbD7Ztrrt
gGS+hio8gI7er7UbLU/vkau9UujQe8XIT64D1fs9ffMwLl8UP8+iIrBT6e49aB7SVM8JsVxEnaJL
P4O+NYclPXtiNhDwqOa0NMELm0jI8LrsEXj61q3LbBHieFbq3w+WZ+6J/aoG21kQvGC+0a7NJQ+7
mu3e4VnzAJP4LBTQTtCLHiQ4oGb27cXXURyriu0i8vjis+jnnrrU4TsXF9DavakcMQ4QMkBO6N3j
h7LyEATLsovxN/Weg6UkR4AzAF5Lhwi0JQweTtc6vxu3x1XHXY3QHIy5bwbcYBG/BX3F1H30TWQd
bUfeE86hWBL8R+PbNDYO/Vtd67NnN2HQokLQYpcbZiSnA10q/uKwhXXsDpgGHTrU22lqj8HFGygY
6ixGd7YDgOhffgUtwxBcAffrBhR1JZP6OtoUQonFtOg6P39dBgkZHGe1LPQdmjFHe5Zpwy36fzEq
R5CSWQ+sI3hx8N3TWQZtW11DEHXpDHF6cYtFINKcgGhRB4VTJPRGp+4f0qzRKYkGz+cAcS1+ECa1
yQgYu8QeocZhWLpY5j6d/VxwadqFKOtGdkA9b59Id5PE1Rc/xBH+pfSbN8Uv76AqarvHiqYlncKt
OIT8O9uqKtR514Bn06QEuAKxF3LYUrT/T7Q6wirZjcNvSzkixFPbjJFV0zSVi8sNWdAFK7bMAbXS
4gSa/ugUL2ZzNchJF4N+LvuLlSNmQuFwUngdS3w5mfESvYu1vtLE1HVPAa5V49GNr+PosMQHIMzc
ptrgF29DL76vaNcKyaKs9aYmfKf7YX1fC5Zkglz+9CnimezI7OC1XIeOVJ5OzIhUsaW3+9Pym3kG
aZm7pZC6aIC9uiFQso9HousxwnkRU2ioe7+VOOb/+ewp304oCAc6y2LPXC3MS2Yf1HZ0abwAJdpY
SyJPMFfTpKXjhQme37IYSA2/sa3OOgiC/ZbGx/2VZdNrOT7bu6oF21oRj+GznvDW1ss5qnzfgJoD
mw2Ml5e+WhZlHKXKA6YIVhUhXFY5jg+wjSLBemINRqx8P43uCNj6I6IFj2YCXspNMG79D7LyOQfX
+s8vBZiZotA8x20Ysmw62FwZ4Gdav7ypSZj186EQYRdUt2JkLfvrMiaqcLrWB95Sm+jpx+iKD5jP
10kZKSx9FykThbniviS3Fee48nXpIiW0MfFzcq90HnB8u43XjRjxqGkk3owSNPOZ3Ae7IX6qIuWM
CP6dKd/PGwC20zmjP5EcblJI/JUKDfbJDM6T02jV8MeII7qTdwape2ehua3nsw6gwOpGzxsBmtYU
U2ggUQgcgzXLdsr6H/GSXpsstieIcZHpVUEBZ39joXcp+eqepJVOWIVFzLURaus9weCUtQr+K8B4
Xi2drW5uaMdshL/ZtFRLecWWjFGNeQTUZcgAukxrFTyOyuptVfExFmoZKdY++7QHMJ+vcUotOCKR
/sbTFY0N2l2t9SDsIsh25fBXt22gaG9XMf9VLBKyCeogTmW1L6XvC6wkSk4QIKG1YiepqGvepAnK
kXvkWlL0pEDYMp9fddJQ4mUpnITjvb9hcsYIxqbxbvHm5wUI4lvXil2qQ7x0bDlSp5tM3KH0dJ3z
XsAwwwOfNdqhsP1Ds7dWuMgmPhPzGK4eKc9Ls038u46Ee2ZyqKndlUUrLaOmNNt7Ae9z2BgnfHJZ
0OtPwG8Obmr4A6mnKCqDVkcWA5mxOLpuB6wFMOq6tQUz3m7K69qMxsIjN8USUjjN7qCOBRSIqqax
/L1e3qAZYeV+LstMopIKhI8fh4h/eC+9Cvk93vlrO95qzdj4G0JpqL67SkRT6M61BbbB93h+w/N9
5uTaaYjVsf/jzhQJtptwAiFknzIYyBo3UP3hE9I+earJckN5ymPRIZi2L3F50lxNwDkCmtEHS1VT
RM4BXygeGQnn+1cOKt7JfsasVgHyqcBNUq/EBsQ0A5q0pUxqq/xxTgMdsK0hmK6UeD8lJVAX9Ts6
T/vtRSCfYPyUrfrlgs4rMgXPVH4+Ae4SnBzE7omhAWxqMTgEn/Y/Y9/TKJHSB+GsqOMJTigkwt/i
7Mu8YKZ3Cf6oOMawfgDkJzBFZzeRk7zYMSshIdSOQcGlic6EyZRsENvUJfHuqV2SfOSn8mOMmUZ+
6Ij+LCg5ZiOC9QwnGAnW5V2zyDvU4Zrj2JIZEfnhAK4C0Ov42fn92KNV6tgp3MMkF5Ub+bbliLa5
xAT0KEdjhMwdnFM0ztt1f+7VFgYgDnxaN0gy1OUc4MJM9GzDWjb5OQxaKT8MhLI34SaubOZlxiKW
eddeN3DzFqYCC1+1zCqo6mn6T23qfwaH2LE3z1IMV+XjjimDBSAhtCATBjDwnnDxoclHb64L+7qw
cvdusR0ErohHmmy1Zlkcgo/CJ7hjLiY5MCY5gEJC0UDHrwymLE71rzuih7LqnWnAUV30NBHe/n6A
a0Hqfmiih97/sLbZB010GqqtxxayJ7W5m0WoZyhvOqVBkhJ3wof1zNBO75qpzdkdugU7sAZxVC/a
cF4m7LxO2g5pCDmHBPh2DJaWCr86a9YL0zWyyrdwCCK83gtg6KtJH5YqPmae7T6L5C+/r2Tqypf1
+T7g2fdrESJ51j+y50iIe3UhXUVQ6uRQq75TODcWksLF3LjRJxtelXYFYc6FOVgiYYy8NN+81toT
TxCRNVkFqmlqMR6hswtaWTj3rRhB0/NhuefRiiTiCevTCt5/6ojnwpKKggCu1dXUYd3ekPCC1rkH
gMqZUhXR8zDcu8KpkBHfz/JBUaxKHKBkUWaJrfOX/iplc6xXbBZZMMW450AEg4CM9aLvwEDHfNjZ
7jMI6Hoe6pqAFD+Yb74REUGWTScTsB/ltZVhyWj7HYhwxnmPv2mS62e/jU9wMPFAOuULibXicwbU
JF7z/4KFBSDxewHspSo6+Ru/AhDun8g7WelMy2viQQdZ4pZHO7uDwj/iby3snEWAoJFvylmPMASj
nhNUVwuIf0j4pBTX3JJZup7mbtfkB/LOeYgrEFsptTec2dcU4C/3TAevNuy3DdgZgu9dYuKe2PjG
4B7N3jW1Aqkg6fASXdXmBMu2VzZkzAldERgS/1XzbRN/7YaSVIHe5wMfgXKlPOU5Pskl/Z7C/CCs
BIM3NRLOKMlV+vzmbvncp1Yb4/Kpqm1vzRHALrxkp2tENsYAF35ZaMYl4nn8ezONVG1LYTVl3FAn
fbDmk+PpFy0hRLWq9a0XPQv9ZH0R6zASbDXoK/vDavwlYy/SGHxBQArwXI8d4MOHYMQO+Zn6EQda
uQz9Ik2jg8iopE/fu28v4pGcNasNrLIcQMwYAl0Su2sJLEHiRjq1bQDGLsuxb2iPlS2i3HwlCplD
s6v3vR1YdIop1mJ+xO1spinS+iOzBDGUS9H5CJlENdpdAth/NE/ILzAnr0y7Ss9FRPgRmHHV+ieI
UhFEpYUY9ELPCyPfAWWJGojCwL5IqPk4hu0nCcOy3ZgFTV7PthXCbpkf8fpPU0yYHhfoj8ZVdCIu
68bZtH3BKCy+XIv3o692WKi3V50/Bp7PiS5hLfV0k9lh4cb98D5PZcz1jfjkJRTS2x4re5ujV3oB
0gOhvM6mMC/TsSwgVDf9cbM7kF1iefguYXgXrJ9fIo2WhsTHDF2PrcT3Ds0WOYtHy/vtemuoViUy
EofxxyYgLss7ZLXEr35GXyK+1V+ycpYKTqzOBbS+Sl5Y/zrqeM8xjEDUe25gcutkNTVSVYoOr4q4
jcQzv/JdLhI9y0Mqy/utkJa0JhgQAr17HrStvGIfAJrkNXeCg9KwmjSihANM3OsdO+q9bpqtzHBr
irj6LueIsBSO0YaVOp+IWBmY48zt3SWAb0aIsJ+VdJFpqgHTAkN7w5BOOqW+M4DC3wCTi4B8YKEV
Wd35kj6zvIQ1OU2o7DlVihzDpsGigLleUDhQXGVqMkObCVXYcJrYr7PTOHmng3xsMcXfk9nmhRcO
nWli2V9ANkYqWVGGASGjONsWyQPeB6PR9zkw4eG3UKL+V9hQRzKNKdVu+NyUfRxcFgt5CRfMnqg8
HIKdg8IQe2rGWnqvYgvUAABUaLrfh4Qkd0ewLnFjCyq2/MVbojYGfElJVjD2GkN1c/tb8CH67duH
ymYB5fJfwnEQ5mOYguMq1DXyzUvN0WEwYUZUtQi9UtkN9uN/4OsGrHpSonK/1aVCqqrvopiqWvSJ
/09pVqeMWNnXb8LfPGvIdCzikZAK6gdUZYW8cTDqpFZMZkzZjS6eP54nsAePjWTvn0uBmtFnv4bU
FGIUzhSFW+MOjGZoVFqsnfo1hClWx6V6cuzJqgUoaeM69V95BKV004difP3pH4T/fsFSCu8PhRwz
mQ63Uv4PyqDAzn9/vMgLIuJBUfRSSY/TTfrNulqeqjS8lKF2XTVubRbx+I4FyYIokiTx5ujhYusn
dyv5YTupJqyH3AEntdI15R4P0+BWSk5r0hRaUBfbl8awb/Z88kHnAm2/yIIIdpfF7ahbm2ugl+f2
MVNRBUpkUMrKuOrFsaJ2G3YDs7x8TwWWbZ+Lg3zsBrxSJSJmixO2ESJuagaitfkZcVlXSAA7szYc
WJQ6oxQS8yvY5cPoCpNvyTfjSvVdYO0SZ8YVItDun4sGhvf5EKExDa814xCTnuyqNtZ7+DCWmACt
5qm3o/7A/IG3tDmBoR0rYFZoI5eFE0PzjP2HOHWiXQlREg0qULgCsCbQjBT/788dZJ/lv2nVIrz8
Tyc7+R3N07Oe9ttRFqWRwXRmC4Jw0zMsCvVpliWtBDEmFYuFbINgvXQ0KIjLMRK5evlVaygTT3zq
e3vH5QqE7LrWS0JQVdgws+pdQKNptMyy25QmR23hq/HX6OH2xAt+LDwbzGq1kRmTIM1BucCoIOEs
TJMdLUu67Jl2j/zNItbCscepkwxDLY40G4CwJhkIC4Z3dogvU5UilFAkgDHpBwBikyBX8bTgYotT
6iAYO1RMOtQULfeCxH5OJ/R6nQLmdVk91HIwmnOcehgMP+vQoK68FhNNvgKWk/BMWfXqqeCueHE7
ywZBO73803Ayrq7prInbAcOWDirlDHx1AsAyJb0JEFF1nqBxFd4PJN6/Zf0dX3UyVwCvVFv2aH1d
/yLhm8kr513s+xpltvDaPb74xO1qh9QlbuEAe46ZQ8g98zti21o8EFMMYOJmJinEkxFUIchkpxG+
FhpJtHKt+BjM5dNyuy9Zt20utuPikSkwAG/k2YMfLiZIz5tNJAYOIdhXxkPncbwiFJgaeeh7M/Yf
3Bn6TZgl1J3WeY7NjuUkY29kiffFseo3lwu0ilk4daeYuYfWApEu0JPyVcZ4j1MIl1rAszaVBgR1
BEo7qXvMcjlHVDZTANxuJyFi3A4St5jfFuO6oWlZhLDLDhXTp11HNmJoqpQJxDu0pxoi76IHoVys
+CQy/whuGFDGK9aPat7FM4jm2JVluH5xjv3/iG6v2IO/f1oKwpDsKcq26KMEkyYPSDdf2aEUZKy/
V4NdylqCoIUgwWVTm5Q8vTCk1CN1Mto8PuNhiHJCli34gaEZNTsjPUgq2K7Fo25xzWEeparTyaax
jpRhErj5m+BjEgK1eNECzoeqf4MEhFbBrmCnv3Zhfw5WfF2qMZc7UT3wDzKBD4VoqM1vD74E7TrG
mSQI5I8CFf0Nb3LiZhFhW/I2hf3aGvEV/8XdloiAh63OAUWBsZjfxFQVcaxg8OjuTGfUfjewIPgr
YpUo90mVOVV+wvnrBzmXVKROig+CCIhOVEVYkN1PxvCqkkPRSLb5rhQmvOrN4am227rcuEUZE4sC
EiNtWyr+JxhrZHtwRxb2fID5/qFyNERWc+IVlicDvXAmIO3sORAR1wyeX40W5j6ew0f6/KyHDKzz
TTZWDkFKSrog9yB04R6nDuEVZahqZFSFn4E2DWEY4llqSwyTrPGzKu+P73IquzHKKu7pSECG9pg4
d1aNCcvIRzgX1adi+5WxAOtDj8CEG/35cVEX7ESZ1yqJuh50AJgyO1/DLh2tSpROz5m+Ys60y5o2
wy4xSxw24SQDdaXzqNV6UwDEU7TRoBZ3w+JQeBMxE19fc7QpYw3zSmkD77f/vwKZJF0Qb1uWJX1Z
TyxqlfoUEUUd9WxBAT7mLInamlts5r4B1oe/j3hndvoQ7dKaDRwk+/KOvDgNbRFUfTOM/brmt+hH
MP4xSz6UJQv0sHjBra+avkbq79unu4H/6NLBDiP+h9hJnLjCXHAZX5H4t3PlYxhWq3RPJOz6ueCR
Rt/5XgQngHARIuIyZ2mpOiIdvhSCY7WngfVQRo3Ys2fZsREN8AXBK5VznSZkXza/47M9QP2IKh9B
gHBS2pXz862nyRFjpqhq8fKIPHpR9VZKpzgqF/YoThbzo7xtH8JXgRrqKdQWmVn2B6pHjLdn3sTX
1ksz9LF/lZ0i33DMhMWITMVmGFX5BJqTBbQpX0OL5I3irLdp7V7+Cd1U6sUznHYc60afZdKGXrJF
LdF49PQrVg0w3Jmkx+OgyKGrvejUwEo6AwSOx4mgXR3QMPe+AScYibkpoIK4kjkbM2natl0pOsMu
evD0NblbzZ3wiqNXThyoHrCI5P1LbxlZRa2VQSJUHqYqYLABDgqDeB0zrxbKanRJyqkDKfQgsGRe
PTnMiGCjlQfh/YeAlKNP1R9riO/S3NQ5ECBbT4h5QsQkifzlOVcRau24ai37LPJg6+7iCmUlBAei
he+OLawCVKWvqcbY3DPS0uxgpQ4VvbqagCkne0T4OGt0Ws9FsIVlorPjUb3vE8UQnuG0UdDUFaLD
9oWY4/5STQbg8cuMjol3jDW+5C6o3vaF08Xm1LNHTM9NhBm5a16fxrUAW3UE60ed6nrcMpoQmV7n
iA/kXdZkz519+eS1MnUVKz9SxxabpjfgP2+Udi8B2RdoO9t76b/xkhedCWRpUJxjA7ggsTW2HuXf
go56XKdvam7McgukZBm5i+mbJzpAUn6jbeCARyefHIWT/RWCCP36eiiSkU+6Y42hgwW0BEgl38bK
Kukj1Q5slXdnGx7XLRdYuTqflij0/GCxvp5LJGVvJnLn2b/rD6C8Uj8QKCk58YraJHvh4VIWJ4OC
55BDxgf9+uNcsQpiiJUIpxpZStxhP27ehZBWoojd3QgwmNHdgUaUJDbvuvpxufslLwepQ1q6ApRp
cqs6zh1guOo3a2wmlP9MQNfiTjdw2EdTKRooPqLo1M/TMiUNCO/wS2zKfAJlwpFymJz13dv9v5y3
seEjp9ag1mkeJlOzfdkffFFtFjKM+gjDUr53eaVSohM54ZpKYq0JYpuo4/ZUkURji1qm04Hc/hE/
VjFTpbs0FOLGWF8BFaZb4vb6NUYf1Xl+q5GboVlWT8JMRb2TG2Gk12LskEg/DRHD/+kELG7DmVWR
V2i0QeSt0syRewijhK7ZdFRVviTC9hRysC8wAoA2eoLZpVQE2wJIj4l0JHrDHX8/L/9E/amn8tEp
zRuNeTorqE2yRc61XMEuvIBn1O/vV4K3Xhtb8H/br8ljyqJ1YGZ/t0D/DEq8bkaU/9JPIowVTFy1
+jvCXKXvR5Q1DIsTi05WDzxJzbaaD/qV1bNY4ceNFhDDBw8U5vCOPjjl2bKIzJQiZiKt9k0qLA3M
suAAbcawYt+5m1r0A6wepo7eWPWc7RVaJIqCtTLYAAURL3eyiowYE2nwABS5506aqFsYhma47vtE
9wSEQ+VFWi3o1EGh0nE31XooZcQrmctFRFreEiEsgbNC30IUSxLLoU1hc0PfyDiK6oKzJavIVX7a
l60AvfhxhCPuff7yiaRhd2IIjoIYvGbjdExgxmp+Ha72O8IpBkX2jfkyXfJsYeoHQrv9v/d4lMI/
/dYK8btNfqQqY1Hxo4eBNlv0BhmCjcvKdVZeIJwmR7b3CWYSuaUR+7/PLW8Zvj+OeP1Y9OuHb2NJ
66+WedKeL9KjiLbO2+LXBO8jmkx7+w+I3Zfk4qKbIg49lZsntbGcVO6CLuzY64HugO/CbrNhdvhl
vGDvqVKmQgkJYxdK00uCn90ZwqYqL9p9b+13VQI/a4nutNaB+Gk7skUBx1j7vvIomT3O3/d6z4Nz
wiB7gpzDPMrJiMm/XteAqOqfYiBZ3wwjZcQmvTltnAwHFwFmfBJJ6c0giNAbbg7H+ViTOz/u0lV9
+XvSM/yUT1IfObp+p7Fa+1h3yUpDf8bSQY8irNH8fDdCswcpT78iLWyL5pPzqwJgvwLLf2acoN54
i96Jm6oMkLnQOJa7KsZuS9XXC5A5F03nxvErck/MhIOQlUM5yWj9m8WoveejRYrt9mebYPJGJGus
8NOKMYv4onz6tNjAZ4OpmouV6A0ASrBVGveHn/23gUjQXht+Vq2/o6n2MsOjg+YnnkGb1l2IH9nI
zb4sw7lfT6HSoI6UdLcsh3M9UC13QLNmFOxeBVXJv3DAtOf/YtdHVBdGFMhpTwmv94onY0iX7tCK
RSbMs431f2YOWI9HnFQ62g5I2dghQKrWBsJmvHmMAaxptIsLR8gCq5cxq9a94L8FS4GX2C4jtV1L
1N4AymBK77++fFFAcj83XgGkiIJyeWK3W404qP7Nz2G9tCAdww1x26DVdxvuV1KzXgwNln5LZBHM
Yka/O9yUSajNefz6oqNh6hEzh6GimCCS1P6n2wv9sq3Gtme4c0BSmqAIzZsSYZfqEnhI+86mM6qJ
ZOEhuH3KUxItbNFcnVZ9yM2Rr+lbEyeomW03meGcJPaVWi6oV8Dxjfsmi3jCJWzff1LIZ/ZWUPcZ
pcs2ze0l7U3kcTEZ1S9b+U2jid37CDo81RIHqnQ7UOa6mmTDYcrxXPWRGoz1Vde1FyvoRqb6Eeih
DNG9wgn1Eb4194grz6YNs30gXCMiTGU6n6LEqyaMoPlNcz8mW6s6uQAzInbwu33w+wgqTgRINUsn
yQBuOd6iipIlba6q4qktBHBz0uTW2aljKyTstAboK2VXBU9GhmXtM9J/1DznElmd/65+iMVK4545
XAu6OGPttHb+M5m/pUFQMwkj7yrLJZgalZXMIFMxcPDaUJtgmgA/uIimOv0T6YAS9X1ORm7rq8R3
SY1W9/uJz7HT3fdZON3gavXZuNdOfQUQFgx8Lij5LJUWVmAhM4074XUSGkgACW3Zw/wJfDwmWa9j
yuSRwZWR3q68mCBpff8Pa2LI344igPN2HloPXqDeyGLMK6bVqSQmYoRvRJFTfpRHLC8d/1WsiTi0
5pyLJVvVZLH0B/83VUwz6fXUdlkUzASr1nwu2qLIr0MM7BKrOHE89Xsqa2+HRHfbtG8FclPkCRaL
trKkHV03Tbv6coB4WJ0JLlpiap4OvUBbsgZGnEdsSwfe+B4gDS8dJfRalKxpK7xMJvWJD3QI6VhX
cRAuAS6ECIxfc8vl7aQgZ/Qtty+6b1DkyKfzEbPgUEF3fh7YHY/HfgfBJqXftLk6Sv2+l9qsUnnw
Y25ecUNhQ0vfsVJMaRS+6Yq9RdzF9/TymJ1C9mKMFeQ0yewczhF1Kb2K6+IYFUc4ahKnJw5nM/AS
Xo9bnnZRaFf+dd53tIRjyPcNGQ39Kdv6oLeMmtOppBRxstOh6NUwp2BvPq4TYCozjTEjKuQW13Ui
lYDhFoqOTT9cv3At2JNtNFG/XRH3kJ41cH3nAfuXdCxI54GjgGKuGToFTdvNodN7pvwI4Ji7SGdz
ysD/100tuwPWSbKhJ1jwXS4kt8AewBWRvTYdekDf3kXsaED4ENDTnTjbBoU4Gs/D78tbUxLBfexm
XqjTW/OP/rd/OyivfD0aQZn/PchPTq16zL/yZAQhRieHmnbeVnEf/vEyil1WALUx0KntaiS7EZpr
yNNzxC6oUh31Z8HzY3tzkJBVXx+EBl2Vvp29JHQ68pOghg30Jz93w+wKJBwfd+l9LXZK+lESE/0o
+n8tQAub/tEkFvrO1smVMKCOYc5kEQtpHn+JepI6ZSJIEZbFh5fkug+VAszpwjHsNATyTVkAYWYj
lNQqE0RpM8l8kO0n7R+gf/NR0R7u4MHTGoNAgad0S+U7cEiMv5HYFgz1152yy6qyh6D4ZF3Tcb6m
0eBiz6Z27FNoQzbXUUt3tOh7qUIX58NznQZGbAYABDnkN5EK1qepRZQEEWlylZ1idp2n/gMPSZSu
Wz6ZGK7FsFpY6j2RqeEIBOA+0tidqH4YjWMJLNHxwpzL2CqxKG5cC6lZwlAAIoI6015ICZDyV5YF
2EkIax2brwJUdjQWl1asPXaqIdsNoHkyb++se6fC31avN/27dW6cU2OKZ3WixXJQjlNrMMHXj3zc
PANyQr6n78hxFB/Fj65/1Zj3PcD+EPPCq5eJDSFaP6fqILmvfGZZuIUIUoQa/KpxgUnFw+ho4dy7
HBmG6CEdp4zLtUXMbf+vUQ5iLL8r3s9PETDyQZ9e3IXuoAt7kJ7XBBV9Zzei3j4LaI2vvsdxe50T
zT23aDD1FxAcORWtZRXvSV54q54nZSB34NTjEHyMFdQZWhHh9RsMJD5fIYTZHmhnBL30HKT6eKIT
jHDAwt36XjvoWQAJ7bIIvEMYnz8Bn0Ey5pL/Ie8gwTLz0zDvw33HIUg7e2Vc4wWUujcJaFNtYDuN
mU84JBCvmLcMeGfQha48qd2T8zR8Qd5HO9fMZglMx8tSeDKv4etsVUM7fEk9xS2q2PijPGPVuuBs
F0pdMDpMZ0ZnFnd9ni4WLKlvulKUObjiUQsaBvbssM9PRfVYeI9giNVVbdEN4ZFvEZf6SN7RMoZU
O1blM9d8tiR0v841652YktiZS5GxMzpd9faOYeAQihn8yIZlIxR/HyBIOPJzZPzHEZ+V8jU0yU1Y
MuGGABh5FSWewueQzA5OzPuZ0Npydz5P0sPg2LXR12aAId1RBP/+H0MXrkW3SaJrAhWa9+Ur5Orp
xITVf22uk9fp6Nb2ScIPhYzaws30E2Tspa3GZ02/ndSnOD0CBZFICXTmOiYklD7B5CnEsGiMWoV8
0ge94iug8XkUuzdmlqmfK9qachVb5ytsAtaXb75TEiiRJh8bLjxsM8lTDOAIOA5HA+6W+rram8h+
mldz7sH0bO4gWYEyKt+E1hQralMEQFElTsrVR+7q2qUWG65MWn5EON/JZqKYVmpNEj8ld3EL2I7E
9/wMStAcGFV14+zXi+XlftQ0rMAV59090/7qgZO3YiiWK/nwHschO7mKcxEMS1Xo8GMM9HBK+atb
dbpQ/Vg1QU8ep82H2hEMVrQvbNFrHi+jqWRQqc7JVYeYJYrY6+DY12eXM29tuXKYuTr7omcvq9ej
331inU7eW27ZX3v87u9QarXeEWxKh3HuTAdZugVThfYBWoXU0KftUO+hQzLzzt6tGkvO9fbAjGhh
D0jLCn0BIdUaixCKyN8AXJx4qlc7zGjwd6dLC0Vn5AOzbWrvgscVZZgtRQzP11DKuN65f5+0TkgO
QU6mYl80B0gqNR//lhyI0lHWzXoeQYPs/VmjUIsfZ+k5tdnz7X2bpKlU6GsN+iEGVi6xELV3rJXo
kqXg2DxaDgy+/jhlCLWwZUZpNbcnB+ZvzT1Xp5vXTo3b8Zj/4SkSkPhvjp4VCX8RtnYg52OmvAH6
g2iLre5o0mVBNKMqkcqyN7hkm1B/A/QXLlJUnkYQ8D4/vFYjLWAJ4xDDm+tXCwAeWSZNNyvJq8cU
rTFJ+XRAbR0ib0BXvbeCXh6GmA8o/NWlFtp6Smw7NRqiIgKbmTGoYvnOSglvi6/Ow/KAjWrKl2b4
8LCBUg0FhMTuepSV6BIOzosKFV+1eCW9zxzY+oa0eNrVizp5dbAM+Mp1et25kcSdHdGGnkzVHwfd
9YBkPYjqNV9Q5d4Jmtsz2/joGQKBbFwVU/wwUcmjtNU4T8eUpOL0VdM/+i8cl4WpX0hyUULLAOAo
STWdPXPi8/2rkFjQz9KltX+l0daB7o7wF3+0n0e72Ssi6wIEO0uvJX0VEs2Xu2RtqBTDDDP4Rlkh
+6zwlov1f9xRqR+4MJ1w03/DznusPtaK9VQPm7u+rPnRZKJN8goAyFgJzNkfeiuunCw5kJu0GpJb
BhNwLyFSo3gV9NGetgh8EscpNnbIOdaMo6YIfG+B2BDuTeFSm1gUe8dzQQlMQUq1YF8Ac4rOk3ZE
OtGIJjeqVNbnB3OnTVvKnRuXLOz9w34c+RvMB8Zl6l0XHdTC8b4n7q1phfOjFGESKwbtxBYBYY0X
SLQxrdFTv5HiQ4iQmzBjUg/OQ8vyHg4kPHAtR0ghcROv/BAMbGJgI7tVX0auMXMaMhcMDpGBByS6
U12RZUZtefWT+7mnvxvQDNQNH6xhrjVOYTlxS8lkzOjO0wiXygSO6GYjZ0DX2KRRto0pDr9GI+Xg
BWARKkQa/7yZ65HKZj6LPKI7szgscl76ao+6K7ebOhIlMv34kfW6HHH0DADthHd+qcYsjBs33ePW
xvtsAUWSzeqxvENJBUJWKjYL32Ik0raEUYWu97k9x3Fg9v04IrAmT973mhpK8JpOcxb33OpNIYSi
aa/D/ibrbYvM7p+ia9rM1byWTZREVVGM4AHahvmcSiAkc9mk+inWDn2Ut54LN4egmMdx+g+EF8C3
9DnwAh8JLuxhdYIbZE7S2d9mmM7+roZ5oraMIgnagEVWvKGx9goNoS702rCVqAqAAzkkU0LtbZlA
DKUuEF3IqUpS1klSNYtzpWwhpZdSQWgOMddLOFPhuYY2XNsDngXJ8zuaheWoRStn2rJIm2B6pcxl
tTOKftzIP9TShBRXahWKcUXCJeE8o+bkieg300DTOtOxIdrjpdQQLvB/tzcINIkCT2jzWomotnNW
ACfuE37ErdAjx9OfEOjAHkfZZ5myG1NODNRXcwPg7ztNH/eDkQVL2Fh1TB/91zcywtYGd2/J8nmn
vjBXI2NabNq44Icv82oiScC/FWO7CKWtf9Rm3GR9yK4g9gD1IGYp5uwCYyaaRVi02wxumi/eXerw
tPu7K6RFb3WqD46LRcMd/L6mIP3GY0Ko5JuBbG74dAw5jWLwLGeJfGFf/C5ILeOfTIhu+fTzpNj0
F/X4FaErp5jfJTF3CywdD3VKTdSJNXvfFHbJqOuz82jRHpdye9JjuVs+WboaginOd2i/HBPfxdFc
Yg7Q/UMW1A/+yRlUm7sGwKxpIVXIasL4JcwcqlzghRjx2ymMsNmOroGHQVUllMcuJVkWo31uApBa
5AaTL8aE4ahqSMFoWqc1Oq6Y8d0rZM0M4HfId4EOC0KQA5ImorLgbTWR3b3lvsaZvjM7ZgGVQIix
vW96WnIKz/VGQO0cfWg6HEpBBW8Y1qbQGuvS09pIdo7GQokOqo8glK4lJoinAmu7CgFfwG4XXhcO
r0TI1zUahDDATMtP8VzZr97BXa7n4s4G4smdFAo55wsT1Tkn3baoLPWV2KRB/O2+fIZAEQv5bQOB
Mt8xnhUpsJpIgd7L5yvI0+I261SJUsKnhZJhXmyAlIwQVYQpfRfUh+jIXPS4KsnsSBI8IQVJ58fZ
xxrapTd+jkyqyH9bFTyfbbeO9E4iiXUXt4uLr5FBTKFhlKxFc9MLByU0VaX3WjTcguaw/p44Fo1w
k/I5dN/rE6w290CXKsIb+qXr8c7AORq77ZJDBdia5JBhpYz99N1jEpHetU+fJ3wO1Kef3eRCEg2S
pFeJEfEZldAMgo7+AFrwGj5qadA83fYZ7uR1sCbJ+a0Q82tWwwVlaPQQ8yM0PsajG0fLJmNhdKIA
+RyaKaieWLyav37cPGk54y+cFnQ+QGlBHBGkbwNDOA1i3l8IGYOqc7jB7wv40EgeKQ7deytsIYde
Vh50Xr6siBAuRMKg7tt1BKlzas4e/ZC8rf/C5Boxx/oOPhcGWZZ+lrLx68Igzdkst3JYjy/uDMgD
KWPH5cSWlRBhHMLyvz2y1Sj5T+Zhl5jKywU635LgyPlRiWST/bPkPcFv71ZKmA+HptXy7SXRfjlV
zK7ACHAjTB0a3qNINHvuaUDlAMVaFc6+IdBals/Hize0MAdrH0Rz9gZkiMiz3VlAlN1pkfx+OfXu
6ZGzJIdh9kBYKk5rdu5LqjQerJtDVdw3k4ZGA7nB/Bj6qfWwm8qCGy4QxmTauUabqlb4PaYzXx+c
HzwQL3npRmvyeDH9Jdohyyn7t31dUE9vAZXMGoapTmFAPutgPKfZVrPU1JqvxNbFrBVfE+Qcp+6T
GOem8PVykYTgZtUNKjb/YdcQqBMFC47ocnMX76+NjT1+xzeqHcDebYqaj9F0XSIua0XsFZpQ2zJv
ovnWUvL7xbNlFhNnPhaoMw3ZMM2mYh3S98a0FywIjdU70g7mwWowGOVtiRrbmWNyjZCMW4MdrVnj
FCed1ucIF36Jy0EmN2mxx+LalB1j/V03DtRWhX7yHKcpaQdWXpCWfK5L6FBfojg4g5GNH+j9B/Ff
Kec5rc02ZP3whNzP2LhoDd71tWdnWc80//UMbIMX7dgBKYWe624UusLrI0qS/9bi04FIhyeP/jLh
MBejEy/L1HNvmh8zSpTVwL1GxRg6F7ae01NRvZLCzCcLijojdI47LE6TuzIhOADlOjWYffpXrW9h
4RM49Zq428cMCVdPB1bmR9oWHFjBB48AmnHpfMw0W6xYiK9Xhe5NdCOLsRdqCmhlZCFLYDnR5Qp2
x/54GjNqMciximjCsF2gbBW3r/HqO2sJdZYmuyR3UJDOTy/9036tOj+34usbkwuQ49e4wbAAqrdZ
7CRzt0vsbb4XP6TsFLqnVoCdO5vF4XsBLXI0e9f7gT15e737mRlo3sYI19qRPPIsm1rsttfQZbix
l8z3vCGBG1ItB4z/Jb8Wvdiubumgon4Mw8Cwy0dOMycl2sA9lWYC598IHTWZME96+BeqG2OPaXHZ
13goNIKzrdytWWHDppUwUxCriSGFLqBWmsovNJOu4jG1h3QNYj457D5E6ZtKTk3OKgQkYsJWIaeE
8Icuk1rAsg0EL8e1NoxDMDiokmh1p8895FjD6tGHQ2tYmNr8oMts1cx4ePsAwgaaR0AS2E1DvGl7
gPb+OkPV/f0k75+Fr4buHN3Zj6Z85ZZeux7+RI9W1eYJ6WX8nkZljN4QRSXqFcZLk3AOJ3QWFC4s
kZsCDe+m4LudbvUuBxP/QsPhKh9Dn9wMmzBg3vdB4ClhQf5bn5gPjbcAa5ZIYpYuVgsyV8H+x02E
2AcrmkT9tseHLymf6iABEtk3KT/R8+4BVwn29/B9X/Cl/jWAT+hjOh2g2EQFWpseiKERUnolf9xE
jwRl055utwPCFkJjXqfySMfTHXWxTSa9g/cyO6r2GfVMARKYPO/zzzJ3ZDAPdaPo5Ry+vNb94wvv
CrrIkPh9qXlfAwjbsmQL4EsJOvogH1K2RZSuPnCVjWG10qNRhj1se8hm8+Gh4lnAtj+th6ALUmTk
mXog0HegCjjhBV+eWEON/Q8/gRjIkP0P9R6Tyfzru3+uoVnnthOaJyziL3sYyY+iaYTP34bJF/PU
JJEZDrYuOORUIohgYFP8W0GFYwO3tpjfmwbbQ3WQIC0osvtNAg8Jfh4FRtAEyoMyvJz2qrnP2GXV
RQxr0VTBNLBkqknWU4pksVLv/RLwZH6nGIAsU+0lgqPmqtDX2wLwGmGFf2m9Wx4dZQikstW3Tc0e
EzA/yvDBKcER2Ka3FQhzSI5x/FvB2g/ETCmDP24GXMd9qcjnlN4h0Ux2LgRjzDwSgGGFLLHY4i2L
ZWK9UKmeKqPQsJn4VoTyM5S+OT1dqQ2gXioXDDoE4apOjfepsvv3cmupdDnMw2mLAdiEcay21aez
6aW3wvchqX/qkjMX5o6dqa5Mj0TTGJ3S+kLAxA+MaMB0UJ4RdmiXdce+4D8utaUMTF8+VxJ75q9C
eF2LIpW9vhWTkXiMfJGJnlvJi9K/Cb79AOzjN14PEq/d7biK9ObG6HDkE+8jDG+TfqHKyOP7VUOw
5LF8u/A3TvILdV8TgoJGtmA3lQQLVHVtcI/eHdWJV5Oc0xyOvvu7hMXj0hXMDn+OEQkI0PYfEUl7
po8DPsgkXsz2w+xLjJSJ6dhghmk6KEsxNx6+fn83KTJhbT9GeXyzJkwun3zWiu0YPWUW8jan9YIn
IIEOenyAMUv7d3/VbBH1j/TuqMYlWSQpHhOAvuQ5tgvRWiCCg986MVi0Of4npm6Gpb3+lpFF3Cmk
DDOo7V9geiRQbrE7OLPOmYCX2Fv1hWRliHp53/jxr4luurkZ7b2CftnCY2/g56o6cdCDe3mxpH5q
M6IHzH0PLUNBWT3QI2Z2MAj+T70OiewdohK9OD7bAQnhD20/r/7DMqEP91XPtcXxOQ08gw41lvS6
2Ocql6TrVbRpf1ZTEsEyMd1GQ3YMxeCraznooovjjvKmkNZ+JNf8Xlrl8NzC4eqPmAcniNCMxJh7
eE/THIjS/44bzah4b9IsPWlX19gnM30K8MdypqudbDJFNo9zPfx7cAQEotjXeEKe0byyx99IeALO
jx78p0rCzOr3ctJyfe9QO3WUe44MQRuocgd0cTDjfFy8m0+QE/Roy0w47mX+JOYZGgXiMwmM/JO6
8REsZMMajZI4hylh769G1Dp6Fj7wecnN6LeuHTZ7IqCnI5BQ4AzzxiqXSEIaYnFjAuztc/tYEr5O
QdsnlBSL/vQEp5ItXkkGcawDrvu8EVxKWKDIIZzeonXk96DTSOuPZdT8cEDgKeCGvMM4wIqF2h9k
g3fFWBj0vmjpSlQdwmzgmV7gegETzpKz+94spJmj7boNWv8A/DZORKCdq6f4YA9F0EdxRk/l3IQn
RFe2kBAr6IIp6yg6ehryIG8bH4NfR496fFKaoZ61fXHX7lHdsBeD6zeWlw0WE1JyXXN7kX8RFZuB
j7XIeF7SdC3HKusxqybwAYzFotGA194dV2xXLHvtCoaTWHHvd00k/DvbsI2MQ5cVYwA7RYodNlML
17oXnihXkibZCr4JO0jzLWd2A81jR1cBG2MELjkXp2LvUlPLTI/bSBR9RN76wQSJmfkiogIdFDjv
q8qRgbzH7t4eD7ZbgDNctGdvvXFiH/KMFb2MIUFlVcSKVUMp+LDHt7G1zYHraJCpl2NFYt1HQ1Nc
VVnJPkuiTqyk3FUiH6vVHrwv9amZr+YfQayBuR4/tN1zRTrG1857i+Km2BFf3rs0TcRcwrujs9fI
V4oc5o6yNJ1tkXfgrU9yvGFrswmjKoRJf0fGqq8YfaVdwibrnXldVviD0A5waf5KhZlDk0240+LW
p6nidGxSIdtXYYc5mZVv10qZkRHMdywEc/Rk4dt0tlSB9JAgHhrxkCp9WsFGrWYHP08UCVU5Ptkf
rXno69X8e/CvGqptpC/MOduaifkr1jwhFhKUckVIEpWtPGCxEtYLWoRxnYz/6aghjBUWBR1z7KiI
cdFQu2BZnXO1+E/MMo2RtVA0ciQXYalpxh/RMEaiuoxEq5bV3LW6kDRy3nm6g2gB20ojzIwGx1sr
Oykf4soLFWQ4EsvJe0z1FNlKqrVGRPjrYPpux0DF6GxFXrqjipQxZD8zHQ3kEP3W+9cDTIDzjiks
z2SVcUoGP0jTARLbJm//SBnE2qfCBT/p8CLTlv+CTuXk45/tDKj6wZj7IGvDeOgpFIDfX3w5djAV
tL0LGhh5yQxgyzRqBeXXN59xBvHw8Y+iHBQSgxxxqdkBDWyFq+Jyu4k0mSSXvtUt8/WQ20AEDWbm
HPmM5n7H5KEgCcxYGXuIlXBA6SYKt/MryHDp2ijWAsP3DiZ/pvtWDjSvpSTxO7zwqrMWx/nFOrPv
nzovqyexSW+5anX1mbVRAv7FnboFlob9Q2DmzM+6CH7kfo8sOMr7oE9A0BXdBqJRVN8LShPw/UZC
pcRkZ65htMitAE4ijyDtm975I5k6CdbaK5eXnZFjRss1sf2NJZX+BFE0NDbonXiAHz5LjBVTH6le
u2e1DvtvIoOH6tcWrQa8XCIXt38v6jN77vnkM+u+hnEBZGaixe9xWy6P1hxdfLmVtPViUQU/cKX7
pzWGF9hVNSVCuE0gsK2fUv4inuvrVutW9OrwWEY9Ckf5rkCTBZot+mEhyO5kJ3lJERE+PLHVGqqk
L87vH67j3NuyYuvg/e3CShNGEs4mHaQHpWhL50cV+ODIc6PVdTPBJsRyDKumBA0bui99zGRjQ6br
u0jUqkl4YU1bZUJWg+XJ3xUfl/HlDAgtsvzJIogowWQ8KoaG2KmPB9uL/3/ggl1YAHsBjGELbtyG
k58K3fj7UAY6/ocRZUUbZGkVLBbyet2z85LTIKSq4A/xhtHCbQpTYmrT8hsAf9EE00oXNRVeMm9Z
qlD4J/NwgTqH6iCh7TtcGtr9Idy4rrEyO6BnP3Rj+8hxRgsZKv01eURzXiy3Ed4B8pVScHcQZwCN
kEaKppTfsb0daxHcwfLdYgTegfoQ8SdmKKoPtghTFFEsKodZ53kLMU5eKeIMV8dEoScCIv3gZueR
OzdRXRrp0REMJXApSffRvFm8Rzb8IS+C8ZKidm3zjuA6hmM+48whwVhf7WTMp1gMYmafa7RPpvrh
SMcwZwgzdz3j4PYE9ombQy+K+cTZytNWGUij6EKoC2BbEuQ5WS9Z9h1JBbnPtVGTzKabjE55gc8D
Aui1q0yDtsT9kgjtg599kmiuo8lFWnaOpYcd0yldeIZVbIUSxse9R/5vZuZ4yDSlaF85ARhk1CpB
Pl6syU0mDoniaO7czorZnGvB8ReUvzTXyGUrU/EOwJmAs0GEuQ5/uT3zB6Rx4IzO++3isxpMuWS5
iy9wXlO+B+XvODi0SlNZWXj8uR8yVL/a1hLp5PqvwEKJKwmip6J1CYYuS039qN4L5eadmC6eRjmK
BW6bHVRE0BwxJUIsARfJlOTLhHx5uJhiAHrIohYoz11huov/OJjD8R3UZX/QOfsk/zZE0fa0wSmH
o8IUeLnfH59KFlyRsoKEvYQwJV3tADkmrQK9Zd2Ra2jeAt/GNF46EAC2LgxEj9R82n+OQREbF5zy
wBoX2JbE1jH9zQuJp6BJVnz7XtLemoWHxExKGJYx3hBQeZTFEtrzN/1cLguN9lmL19HxO+Nxy/U6
2CIlQ8phfTC4ChHQ6HeJonVkoMJqm3V1+uUi5c3jSV5JuD6dFUzbF/CA8b6mKw5WgxnQpB7NJzUK
JeVc6k7Eas9hUaze8b8GMJyPT8f8ePyCfrbQVKXYgc+4OSiAQohA2070F8CsWMx2/SKCfInyvGqV
JRVxlHgQ2EPgd00akTuOWpB2IRhul77PY0D9YThwrTqlTvZfo6TVCzeO+j9i7m6+Y09O7OiK8EYp
hZrSBtQZPMH4GxH7QSixVN1nJAKBkQiwUe1FiOZrWD27FeD3vO9sLMl6MLiJV6QpMQRr8EVuZ2tm
NSLHoRuk7euhWb4M4RNxUULWN5ELsT//7HqYtOsoeW0WTGUBeRZ3jT2sCOtLLLm5Pc4yshrqaBCO
IbUUUq07LRnndzA4mJyBpF3AhOL3INFI69WqBMwE+BYgkkytUncKEzdJQ3uguHjzobP9jmiDSClk
MVBGln47T0x7bzuabXWXQ6VkAWKKj6cy7G3g/Z5ZdkQJ0qLRGgIWE6mMDfHxamdWE6Z8lHsfVNK7
y8uJUdTac4AQPpwjo5lB+dHXdkSQRjIIkETlAkqVRmhTVPxDkdzIl8QZfvrPnzKPz//NJhCyc4iq
8Ez5XqVhOjCtXlYgiDCyHHcWwDVQn0t3X0+PRwPMp/J/xcf21nYMWBdocIV3yEntxVljgmGrOa8n
aoD+4e2VB1xMji5yaF+W1MspPWDZWimHjq9a8xKYqM4qnAyzb0rarRvJVrdwmgDJAizVWzFCqNNS
l0OJaWRCWVRe9t1MK3tSkZkW4E74AP6tA4YhjIaQTtI6/uZB1FWxofaQo9H7AbQcFAxrR0jprMRD
gXyqPMfuVTz3mVgPWJ8CFpLS0XpBVUl4L07WlwozfYWt0KckYdjmjXmVXuUnRA7yK9zzgXXpQdfp
g9XlnKs4lve8SkxiyAMZO9NR97XWNnYJlV2C0w9V9Rh88WzmlVIbHdX/RcvlQpnV0NK3GKVHi45m
7fm0ztm0BlU6jRkiO9T2ScTtyCpyQ/79EVKv5cefCBwjSIto2MJONY6WqpH4rqg90OgeFm18HR/l
Fz6yyHqrMuez5b6u99bfQD6tKAu3jg/B8fk4FiFycAEDo2xYpcN/VXBd4finKJkIh12/DS7OG8Wx
XWbKkkSu/BFQCPXVMv56MgPSNTmhFokGMrMBW2s17U5AxbyZzQPcxFok8aVV6RBOs7XN9eaMIxcM
ORPnVF2J3SpZ22Pbq9cEzDbqmMv9nZqccsJE1PfyCKZC4LmK6qgI/ibqQxgyyTaqHwS0UV+Ww2K+
xyB3KQiMtsWqYulb1mZJbcx0o4hy4nzVB8gImX638um0ySvOvdDzhAqHDV8P7NivSkAGZGWZPtNU
cbA0PkbvFiiHjdnAkr631SSJsmxaR8eria0+sT+E6qzyihI3vrmt7QvPg1xKJhLK+i6hRtW1WjwC
ad0ms4conG09SHC7p2sHhEWE37I5KfBTGx5CBAs1MhrwHDZvxHrF5MR/SsDijGs52X/Abliyo4/Y
y1jQRLaCO7SYMmTyCEda1nEgYguASLIW0ctUc41BKpAnuEMcauE8avcOg1Ko+xVLsKaxwroFr4n5
yNJp/eqJeeuZyJnHMR+p2fUCQWbAG4KQ0NW7Bm5AVRN9mKZqFGDhNB8ICWrg/RQV98YCe/EkflFc
WNis0gMvmta8ZAhR7N2T7e0lIcFFGY8cHHag0i0xmAZqmUyg/nE/BBPRoJ5vxHIJvqMdxuTA88VI
ZgdrIiakLSyQnEYDu2m3bYwNez0kPeII2YoJM/g5SZAcgTOHtBpW+fMQRVolxEIC84ekh9tIQPp/
zC4FbSDMjseKMw2A6+Bv3V5gWZbe4OYdLEtUivqaNTqvFQ3O39UCdrHJ9cfT4YasOXcNR9+f8eHQ
BOTq80nqEpK2PF05igpyJKL6tgBZ6wAK+zZ9EPBfnLfNI5ZaB9XHwMu3V6i5HrX1qP2EsbUwuQOs
MADoecbggX1EdtRd6k90JM2eBLxMgY9G35n47w3dzSiLbBTMwzqhk2YygYFoKWsdGWbdbhAM0ddU
FHwJjLmmCMJZBl4Z6FZK5m5DnKQ/ztoR5ehoqo4vG02mSkE+3E0cJg6fV/pDvoL6HAEbUUEvF7Jv
91h5nYe0FHhxcamn2tNYbxtZe2Ou6ZbMa2vBbIU/LSkeR5zIC3O9H25lQOLq138azanw7E9akcwI
OLTBe6sKqfFYt9Knuif3JSovW3BD7FWA5j/BCOTOBGsKi0AopT+0z4Mq3JmYCTZZ9sdZ1GOYrmZ8
2KYNjQmAnOGfdTVgUYIOvTabq5OlUvqfa58EsNq3woBm4WTnR9f9scSz6rOsM5M+W5u8GeONnUL8
ITF3j2cslyQ08+AG2lYnvPymGMRAB0lqLBRBYELibNZ8HnLU3A7xlpqfZ181+FqSHOKR9BhtV4rt
Td4IarkX152rrV3euy66wwXpaGB9ljDFav7CQIwj/9hcduVt6BNZ+852rmWvILA684nHQjhELFB4
eM8ztRym7l6e0oOCxkUjIDxLOAWDNLvwx9RJHtUVFs406CmPg44CJfbFZYAJpatTtPxmI/jBT0gB
Rve5jIGJbxY0ohchE6sZG34Zb9oULIJZXjZNuyhMYDnxEEjoOIQx0F5oWbiHslP7deObq7sYdDyw
hHsgxgX3Pp/3e38+y0Qr3I6dqSCTsGmK6OzMVncvN3oHQFViLjn0znW3upVcLihd3eec9ylgR2bQ
wuuMgjhQbkzKINPIHhHE13Afuy7dc5yPdN0vCyKP8zJYnN58rXIgH4En7tPyGE4G1BCgwsMxJTCp
Erll/8Zk8xAhQOhiBO+UEYaJnk51TbGXUm0bBz95ChQt0sc+DhTvtYlH5FcgO+pTF41hU3q97ELp
0Uz8s6/sGBqD2dOjoybpcfYwSICljSHib3voLoJngsB0YLChwiU65Bp3zgzKWEC/iTbCXw/I6YQw
QvUC0ebIjMoWL3Nr0kuxzvmHL6rWr4WVM5nH4WsI5qI10MWjH0mOxufWTs5WDLRThhgMAX3QUgi3
t4rmtWEF89P+TRNQjGyUR5F7rLNmllyQJqXBLmlSY5uekrp+iIAVvEb+SLx96o4KaL9o/YcQLKis
SsqLT/83XWp/822OSAr8G7Z0lcBnIvmjOkuiQRvmuQ9lmKoIIHcFFdpd5soF0pLY09Tc5SCk/0pe
+T/oGTVZCGviD5GvsrbyQyIn6q5oYoIK1VSXv/FP5acBzijbEnX5LAWw6q0bZnbRJdqEKBxqlUtT
NlvU7Y6UKSnjkDAprwHYJHN64Tjz3AdHAGJ5xRgOB2w8MluxqYoOXo27yQ46dI7j2HslInnBRhON
MfeNIRrPZ9hgqjNMMYxyYbMLmFzL4JgLYbRvSoBwuZhyF+pZmT+Wc8ss0BN0omUHpamaMIk+IuXt
90YNb3l1XlDMKwyj+G29ZU1IZW8S2T68Q80+n7jeMYyLf7li4J0Zd5+suDjcIoDFmLVTtuun77xU
b3gBMDge2olbdbctDNtsb4hRlfiTwvrGhZJcTeUzgDAlN5NECAR/etEnjYu1Ha5uhKDQmhtQmghc
1dGRAy8CxOc9jpGTiBulN4RbHGyT6SFkWouk2R+M0unQrd4fu7bPZF60NOEfZO86nEE/lFYS3X+U
F+WJs3KGmIijAbzm9W4lBbKNl04Johw5V0CN2mAuyWFU0SCyW+yxdXKwDojGKE4HOp1OIrFanhsp
7ORd0t16msDWuy1LxKIZraGfUQ5flMZgJJZZKfeV4iPGFnVAjH4OZ6loDhWcd4aJR2BlLXSCRH7n
0m59S5NLzVw3VPxAExbFKczfeliMJBFC6f1zfs5KqkO4PPlPCDlAn4K+NQMZC6SNG6BJ8vVywmkY
P0aO3bhCk53YK0X4r9wzl+vXOUE09gsIIpXyJvxpcr/WV0RgWGpsFTzYmzw93gJDZxNeyiYhimcN
ldE/x2cLn0gNevTV1ULG/f9AfKERjUU30fqnbiSyPjfQuBtq23YRntcEHF6b+6ywPFwVXMWoSBAB
/gzvezi4MA6eoyKNjjtO1DSauR2HxSH4ChW3TAgdpxNpoRAU3R/Ir5PG4LqH/pOMadmFDCEzEfwT
jmreKN1QvAVLUvNHgE2/hquD2GhY7/EbZYtp9WsbeUudXf2xrOg7kQPK0GOhntbWVwzZda5DDsJW
iczMvXobBVpmMpVRKi6L5iBSjFM+3PrP6HFgjs0pdxZ8bEet/qJIk+J7bn26dY2MfI0aMZkBQlQo
JKujIq0rsu1O2dSsf9FL/EFeCAANnEL4Wj5zY2N760foJQoVuF0kCsbxl7sEaZr/kJA7/rtAaf/C
qg/kwa1n5fCSdfcdZplBJTDOXm/xqOf3shdavaIlzgCiHQSYdCb8m4N0W6uz3Z1/Be5uXx+3pgcr
7MY0f0+XHf1gtl7lEGtiz85YKtBUWFt1kJ5hWCErhIvSpkeeRvAvErb7ecjR1sDh8zk1AHWa+9X2
rqCDY3yOduYcew8shaPnwaNUE8AYG8+7sFdFi7582fvbIq3UV5/5ij2KYZkmMNSvXl+CCDKKq1fc
rNJcKtn348hZorqdQKP4IeKizOkZyBlSXLTDjslngFMzCQ6Ysez8FO17nX4Xka1OrxFlHeg4y0GC
fG1BjfVgwEOl9iAXt0nsdIkipMGAKPXyW2KOr8f5VNv1wIamvUUaPjm+mUF3rfjhmsQqb7plU9ab
scS0dc+NEYL2xlLsVGlY7JRau4adGM2oUU7jYSinYly1f0jyxpij2vE7+EaGDPAhm5HhHJqXa7rz
47FMustf3kotP+H2Yx7A7o/XvHhzwU8FqIHkLXuXqVLUT6Ct/Ewertcd3DLz3hWPO2Voxc0uSnDj
EdLv15o8w/wGT28asQp8CE9HWRtsfVToUopimWLbqJUVjFni+zk9VMRHx0bdVWqDdkeMUGniF2ex
sfCGaBp1j6zp92Bvq3jpMz0WFpHVoN4GYzE5w9zeAjP9Y5MnsSYos1d+kMZgtv6AWBu+dm3nEV0D
lvvdcItTvmy1EsGg7FiA2RDQ+TXnWhKcxDdQsUV2j90h6b3U2qu9kU6/APfTTo+PwPXuAzo4L2y8
7YOy0UWQNoeYkiwgfpwRaQeM95d6kVxx5cQDdleeJ1V8WrDQhLjXPiWLjOIShYrfB6RMqX14jYK6
THudIR2nhh5ImvoeeCPNv57pL3C+FOlo6Xj90nKkfFVwhnZeVdcBVI8Ixaz2WAP58lU3NRLCBcdJ
MOaf4VAdc+OITDJf+KzxYQiIxHcarDo66Fr8tzUEyeF1cp1UbZMOeDkLHVFStDqJRGdrq/bSrrmL
c3jYK2bezG0DE9ReE68QQT/KmuH19kfOojQpmknIH2RIkMkQ81ugC4vqnLnpnNTMECZLiQd4S0H9
XqMB6Yp2OEo4+BFfAoz7kxqfzQlyhBkb8hpylbPsFTpkAdftJ3bcwy+Q9Hr0yBHDH4htDPcHefFU
8/0HZPBLftTmLQZsrB1BZdSjRB07B8371H3nwvP3Br7I2JfvNFBBoxhXifQKBf3kDOMfWc9EZtod
HpoznoA1w/UXwqvuiFEfZXuMW43QeEVAxWivrAiGbbHKb5tUeawY1/rRiDqPnHfkwCAy//5ugAsR
mMaEDvdWHKaQeqVNMmC5nINVhacrQ7BsnoqP91rsvd9QS7eaQAmu/eslU+XakZQBueOOPpwU1q8n
+/VL4hihbVLV68g7Uk1tq1GPPL9KrW2MI+2yhgzCBVXvBkTKmImQTai/+0xK3y9XFlO5r+aX/rS0
jPXDsEjsq78qXc24prRZuQvGPaOfw7pRi7mwQu23vKCarVNVCMNB7R0QSwfAz9DS3tPH19dXLMDn
ictFkKf3c1/k8F/YzpqiUWbkjA2fZ7/rtcudRV2DiQwVvO8msCfVMwEmYA7otj/xM+YBSEtAuIhq
wj+wcwl0unUJxSXHY6UdBPhmqLv5GU10zBTVR+QCvFAT+RfTuFkWROAdRC2v7V8z/tUS2AjQtZlQ
iVrpKJBAZ/opFPiXuWt/lF2Re07Hadadh02BW66yrrT40qU8t2mRpzzznJsu85dk7Bp2iS3EqB7Z
8z06SXQrpOmZ9jrOkUL0UbYL0wi7d9FhdIcd+CWG+3/TDlVCn3GxqbgCE5xHHAKw+lF5Te7CYcTF
hFypFmVHJIgX+Qw3hDwB8b21PTVUO6H6aLLSVbGpjlQCQj1d/91MEJm3tCvr0L4SSuGnHZWCcaWW
lq4TXAjU+cbBLC9ysgMa/k/w3kQwzV3kKewqzkOeVTLkOFhD8J1qa7fWZy12c1PhNe1fzdgcJkbx
mljW2yot/AQy+bmchk18wWv4AH+cZFHDjyj1Zk7wgHeXp+vgDEp0zG6F4Rif7QKKEV+I+KM7VCzm
F+L/x0nujrsXJX19+jA3NP7rkrcArTwUJONoF3quCxn3oCOJmUqRTrHr2NOLpkrSY607/2PHwuyI
YQkT6j0xK5rzM1b+dA9cG5KwjY/2eG1OrtGMVUeWDNgBRfCAWHX/9Tr/eN83j8bDoK7u6Q0mDNRs
8r0izx5aL5wIvbFZDi0owh9zrtEza7rhoBbCSijUSZEt/shqdzHJQ1bMQ41bGFdHdtUENk8srdS4
lMDM5aO/aq9SK45+A1RRiiR/lKc34g++g2GZ7GEtrtwZjuQN5xBJ7jMC21qqdwMaC5rInJQ8lXZr
oVCGbhB1Sr/o4i6qpfRUkQwZsQH/PBNO8aFvPaAoprgMNL7tjrpZyJ4j/yovmLs7Qy5nQuGnM1/4
cMy/hYRvD8G4tyW+tI4uor0LBGzIBZVrpwWlA5eG2aHD9cZ4diItyUKof8HEA/OrEQ369g5N0LA3
wAQDMh57isiVCxg1cbcMxlyfaEqDuiFc4zuVY4Hn1wWsWx0v3lGPZ8pv5vHjTNVwhl4PwvY8NRNN
9FyawMmblkMWntfSHBCR7cruwH3q8xm0FBf9fpmHbRmNlmb7xA16MWmWN/nSuGWHcXo2g+LG2A3C
N/uYV9WMFN9/BbFqkVZQSLtDYa+yTra+OrAqSgShLNOurFTPAM5jBHORJ8Ku5XCVxdtzm0+vjVja
tmtNSxm0sZ5tE3ZWIjWFJmXSPYs3Cz+5SaR6wiHDYiE/Cy8HRfaSFchyvoPZJ89A+2oEDWD5wfuA
0fcyyC3U8xaI1HrGgRnEIQcHQR5Z2qibpPle0aOr8PplPhuBJ4j54gHBR2X6EJK8azcFJCtbSiSW
rbVyWuFxVSkJR+y4zeMtqYiA8OY6/gqrNReCk3yK5nrbNpyspBrY9Tg7di4yX0/Y8MTkrhQbNPzT
UBNw5iKgEZOClUTUkroSo1jG5DdXFKaeslmbmRNQW0boe9WsKCTdGLnnE/JVlNIsh+4Ugg+Bebhm
dbjl7RArxxulnd3xsudJkI1HpeKU+jJVVpkHbBcX/dHtC5mDy2amSFzPSuaqikrPGGBopJuEJk5n
v5yuV9Ojdv4qoGsSBTepJ+ZO8EMLxsrMDHaDMA7AUW6hleevCi02BF9m/nPc9hEW828hx4sgMP0W
+f6bhDz46pNhgRz60qNthxkJKtbf3dY0lUeoMWweebTQx9Eq2wYTJRSeWdi59cd/T6+6jWGrshEb
uWbd5i8Kpd9z9iOCLmyXvvJzjTa5DxBvAUxq9SSIgPmttOdpAgfBcpQfB3KAcXTf07o4KkcGURor
uOQoQcMN3+3XO2uPEJ4h5nRyDsJ1XDTnW+WN4Mi57glYCmIfhHrrsVVqEl+gnj+P/9cZhIrJEggm
1r2qzt67/U/KIELQTDRtR0LRr6kZ7m/DF8CawNBvsH1HbRs48laqOmf5tSV69xeNzZtebYEJKW1Y
jfcA/QroZIN4t8sTthJVi+aOAF4OIZ5KY4FmDJUQkWO3dxBxgvPqEfOOipAy8GWqsRFIU/trXzPp
JeiPCjZMNsLN6kdYguyzr+UVWM5oFrYkMrAfLmFXPA5vTi/SZRiNdi/Jy528KSbCHq2Z9VzX6DAD
zzRj3vfxJ2jfXLV9nxWHtBcgNSw58dTQlFYkl/eja5RZEhqImQinWWAYHIAthzb7wvvRZLV7QIRK
UnptHifyyw86u8RPqK2rxvlfbWo59+UDmOPfPpql0i9dXyzd0S32lat9sGLo1geYhRM3OafLyRhE
OC36pbTFY7KYQyBr/jC6m0PLCK5DOBf0dfzrdrhiamce+sbJBDAttrV6zV8k4vn4dyoUd1f84ENE
+LqrV/ZaWfexU4eq0xAzzLV5H8/pBYttyMjdkBoBYn0EZtkXBcIBucPjyJGTnSz/iuCM46fodqj4
NW2ugBPK1rUhgaaEvnZdk67pO6E2q7jKjRBLrr5LPpSo39CYyyoOBvTd60RA0+avGKGj72xY6mCS
kT7u4ZGBgY8Wn7nZKj19gNuncJJ1pnmQAiJgwDnthENY6Bk66POSMmfhh9vkTLpLJfTVwUZtjcny
OXjLBARKwk1jmS2h3kcHT657JCfUXU5LZIhJr0uosa79vmjKTRxMjktOHeuNs48GJS9v97ZH4NOF
ErhgoF38vc9BzcNfVomZslFIFrwJVWvZQM+2JT7S/pMb620+8irRTt5pr4x4Pl4GamKLmxHr4fzq
U5J4g74gLZ7XaevSUOKv1NtJumjWgpvLLw0qrXsXsE6eDIuacVtj7sCnuxrgqLf3FGF0IH+sFWky
VJ7ZvPKBgVTxtZ9HB3AiP4LGXSZcTD2iTuHqCfFqPo98QmnMd9iom777fSFFIUdkzgc2bMA7WGw3
G2qANWDWzfYIM2T9cv2aZWMW3PT9kEAuWPmBVXshzSlYfRgzNsfx5vkxq0hduYfkgFBUiqbZyN7y
u0cuLBU+Ejn/XrT/uoHz4YnJRczlbs9oU+C5zfNGrsB46eU7VrhmRoYFh5PsmRqpfryJ7VfqQjPP
MipGRGfQA40wWlvg7E6K0hsZxozXaNjrb5rvjCjTlsscQsGK5kEqwpy3ONixE29DGxMv0gGSb7rN
hDGA3VhIS+GKna5Gu1AbCibZ7ijWEem53O2xvLhGiulevbhl71z2SJqNGTjCPoSUHauAb5P62WED
PPNzKBd6tIowv74jD39lBoJkGeMO/pvHWZEY04TAoQ7rA+xWs9hJVBbbN0lx/FYzzr6gNgEDJkxw
2ZI0ZB1hTNb6DAg8bCTS2CbHNR04TD89VJBZmFui9BsUd7bcrng3ZVL9zfWNUZSe0/t+jYBuLFsl
CcBGBYjG8Ltt3UO0lDnI0THRzIomEJLkqYl6DvhJrLVy0DhkXQRmQeb84+FuERWox1H3fxRYqogK
y460q+TElBMkAYtXH4xqN3tyhFrSTmq6dMo3gJzztHdDvyVXZxO43xQzvhD70mnkVuDjwXkVAhYa
FBbwJeV1jBZFYdNMQBiNyDPHnvxx/n6flCeHwpTo7KUrzvVZ7KOXTld9q92sT0yOE35JIeeN8vjc
BUbrHIaA0trvW7FoUBMT4EIqpFtHIE5lzUIDxCmQoYd0iVUV4S9w9yicbpEy20D3+jiTKGj4gSYj
aIZfXEG6rZCv2YmgBak5a/G80iyDGReaa9pV47AS7MGL0+BZ4IBe9OUFzvbIK/r+/vwnctficJsp
nK/r4M6Pn9lGc1Njh3XbyNrmZMEYAK420yNM8Mr9uQ5nJuNjXG/Rqc0ACgRMnQzjsobtstIyJhqW
G96TTu4y6QD+repG3A1+noHBgLs4wwJpuNgLTxTb2pXx9RvbEVAU3fSSrdiPtQPjPdrv1+9Jwh0L
1e00nBs7WkjkmfbFpqDCM5sOBRE7OFHG0IGl0sT0VOjOnnMSQc9W5vy5Uz2U5FAxfVGxLc4Xet1L
19pVmOXWnfEXMA9rxGU95/LKzv87h817vq5/SoiYoRVo0D60tVol/K7kqimDZ5+OC8ur3zb+ep06
VdRprbuoGoZi/D9e/4pACsjaYTT2U0ndcgUmetWNUfhVlIdIDxgyF16/BrrGGX6ePsodjKUIU5NJ
yZktrfALyjabDp7/PhHjWKFoFKjk9ayJlxb9Li3gNyiXvTqBNDvlxeHAKJypHwE3JLUahL8IszWX
W6L+AOrgSoXvn+os+1JYeFkco1DBN0zWpV8k5SyahiWv9wzUMWU5YTiWtOu0LB/bChJUZUghI37Q
aS9wALstuRnuyT2L9KJPulWYAfaPZrilf/x9pqTbtq7t8UtoaIPgw/MV+YStzCX4EVNa+0/EoI78
2qY8YRncGLcX0JtexN2A8srzhkIKDHfiZL0gJA3Mannf/0AhmZqE9VMaAyDrxbNOXRTx4tIMsD8a
wFnFIANs5p5BjWt63Nz1JDoOAWxxMHTyrNGoGgrVxnEv/oE9ZEJKiE5jSLo348G6Cr09xXftaVkw
KgwxQhAmRkWBkD6a5giO+B9xRSr89LAttVOaeSjaLx6u24WAtUizbgQHp6NveqIkeY9ca3+c6bTE
i6dvwh+X5stcroLoVC+xDZtKYRIa7Msv3MOG6rWQTXB/zNDHCksAndYonw8Mxs3CsKgGQBjU5WBa
XY0fqWE6eU/PxKNDnlPEKX9IlsdbyjF0jXnh+Erk70cVZpGAGfGStqBh5gXcUvemk50yrmS9E75R
kT+AShy2iZvCXLgxXv4vDWxffB0JxqRv4Q0Wv+1tmlRyXisQV+Ww5fHbWrdYXWnFdJx6Vm2i1QE3
f5Za/lCM3gth7tKb+yletL/9c9LRqDvcBGlNwPhTXQ9ewEYoqx4P3uo/k8qs/l48LMmBcE2t0dVt
5hJCx6Kmbr5okX9NurQLVGWbbj5kNDIZuzXk67V8rnJXugbbQO1DoWYgkJ2yszZRTsgk3P8mC+bB
tTNjKrKHhMKrYWe5UgW9IytKmYcUG0M49Xu0UgZCvuY1IiRKWIMSD9SLaeegDlXAYARlEla2L4Du
UrORnT4Yf8EwnBswBWM+fvys8M6uT+DTmTAS/yNFU4YWgc88uHzk8FNYrqhZPcIjUIAirjyXOYWa
QrovUEuo0BAcx9RqtSF9Jp9D7xvJjLYqGulS76DIsaGUwVWJjPk2iG+180Mz2RqYNgMLlIA+wfuy
ghAcGF3Wk3nv6PYxWSVj/0G6G+DEM9HtRiOWxF2aWWffeDeg00vXphb+8sRVHM0NYXGf2njZy9wj
SXrqUgjvQb1nK4+3VaStqivfzQ3FkaPy8FlG4E+FxlCL2Ih8uzfoEOG3lwU/QjToFybOW5H2GUUm
gZ6HyP81wZe4kQaMO/FaZE2eWFlhUFGR9mREPLlHbTr4CFfq/WFYYVlBvAZ+gbDMSp5ebH9+MD72
Gq401/DIXq8JZnpZw98oUo8dkQnUvjkBy07HZf97D1oROFwDtvTyKBaaYVmlZB6yCu4dpmW4JNHb
N+Ec9ybR5PnI31pdgwySonqAgUVfQAKnk8Dp6roQXXBaQOAexjtqnmjOpypXLHKVg0FWK7IcwPki
n4na53ECvi+OU5YQn0u0X8SeBQCtO0/U7xSlkj4L2J7R3wsl/Fe1nbvoHfo7dBqKE3oJT6TS+z9o
zGKoYhuWVrirvw4sOoDYNsSvhg2vKAkLV4CzkwkSoQixdCTilwzNkWMQ59zM6y10kkYBhXwAEtLk
Lw03trRh3OMXDq+8JGdZl5Iy+D1qQz6vCaNnRWbX9l8v0SnTGmxPo03ZDsOABK2VZUGUko0+QQ4S
oFJaPatza0MxfCQGfCwneOLsgMnPl4RZU97zMdcxCRJrrDFgxJBsfKm1zGPsUnzbkaDc0AJZ+ecZ
4N8acpMMY9riGsiHv1DyY+BeJQ41ITp77Y7JLemVUGrjtcJk/vFBIprkhVWCIlWXglc812ngbPRB
HNBKWJ7r11P6clVDLpzD8dr5O2eH9El+/bHK9vX5OLRqPf+ULvMARCJeyxK/ZdKlSeEthqU5uYI3
WjCbrxX4+k05O5mwg+ybYQQ2y9vaGjHuwtqHLvBZQHsDs8XJs0Qk4IdU5wnQLwzyU0FN47JM6GWE
gNoHwcirGk7ojOajpxoKzq5M7AgKMy3Jjyt9sId2waTjzE16IIsl+UzD7F9DLAyi9BWbxZQVRgX9
Gsb7NkWEowZzKeh3wrMfEzyBXpw/6i6v3aThgdo6jVvEVQJr2lkM/Ig3vTuKRbGbzZhvw4+uU6Dr
YfMjoihoauQKGQ4LLr5cdujqcYZlSWjsTdjFxKPw7B8AbJOpkoV1kY4McWwTDvJTF1cK0AJRGHrt
aqCBp2MCUA7LhfsiTzoQPaPGFv7bDZi49ARMNySIfPZnRD8jNnvNvxdJGoUDpcLnbTRE5qZEeIax
QkonsoSZMeLkYLcAn4ECJ5WtIG0vKo9PVxlpNWW+7wApUa9dqD+2wqimdmzd0EVGmRTOVNEPm7eE
p7+gWlVCR9IhWaIV40x4Sxle47eHhKr42csQzI+bFRKC9wD0tcC7W/sxktPfBYl6ocRfHEXbIJyn
0p1XpFxF3FpHmc4qqmJYT9LTC60iRPfoCX0dV/J7G2MYfR7WduW80pml2YUchC9BLjBV9kGsFBSg
UW1wm1dde2sXs3VW2mXyyJroYNfUR1BIvZmJsIugA5G2mgsJ+7pMR+C0pnmF0m6hlwDV3gbfXJ4v
sp0En3sZQlynUZ4c9tfHU9kRASYpRQk4B8l14Dz5lcOFa/8HEX3MzXLBo6Uzkkc9l9CJcNro2BjU
m1dhk6IHuU7TrE30rY0n7jAD8cQXn4nCuAZoo/u8aHNrBRIlaqwfsmHrLajPsqSndZNPpd6V8REs
Tr1ELj52PJ37QYtKxVfrME8Ru45gJs81EsOTheMSeQXey9wv2d0Iu60uKYPQKbt3w2Vq0eD8R4uU
ziPvFc74mQiUGo8oDjyYyjdNxC21nk2QvK47yS759Z9a+7YRF1eR+PWeCeyhCLhLitwupz34Y75h
jvc0e5AXicmEwHd0B5gU9jhmt3+2/9t7TXGQKcftlmfzaO1bP44llogFd3kwg9nXNy0mbNFJRBYZ
6/UkcZnWIyKeJMra6u7AB+/ee3HWA2FY2AiTTcVEyiALB2ulOXTyaCmuZr/O6HwdZba8YWMwan7e
9mOT5Xxc94DYIpiXAoTEASBBoHsgzCygClUnUdKN4q8kQFudiqtaoiQYF0L5f2/Z5lsyAEdP9Yv7
65SIfqhHG3A1eePq0fAoT2c8iq2LVcggpYmKbZaJxHEkpnT6DUKCL6paJre+VkXPgIU7pSgFNmrb
bHjGQ4VmHwxhBXIY4b+emXeRrJrb2WHs4r0CwY/zqKT+JqR/68Bw9deYA5Y+fVO4hQplb3agQlGN
cO1xzFUwjxg5NapZJLPbD0O3WVqPoJP2mN379rYLIq6vBHSBjcEqg+f5VDV9EO+48LGtaNDpdt/5
KDM8rLRf6BdJn8JK7oJBeruJERPqUtKByX6jf/sRayHs0Jg0tXzKw+hayt0DQ3ZeSw0Of/j+4Aog
WxrVJja5V6ZoETM9gnK8V3tb9jG3mooFiiCmLpnS+9WhXyyr7zje25WTcIJs/UafoWnfnZ5gkS+H
klFYqXYiNPVKiFD6TM8ADMbYFKWSmvHGnYWOPSK1yhxwAHETN+A0qnElYjLfR8AYlMUBrR0BXcl3
eDgn/BlrzMlLaiuMYRvsLd25wtz92QSMh6XMiVSfsNrFJhoYJp4j5M+E7haCdnObDGX+zVrZTQdo
0G5fgAcdEygrIAUW5mWk5hcKREqN48BkAc6S6Iv59LgyxQ3RRQzcy+uciitujJwhqkZdJR3Vk3Ci
4HHFqexgc7mM/N0auS5DFLDzHOixI76XZTahFwsbWYuwf/ag1JEcAqS3p5Ib04uAnOgHB2Q+C5WK
Z8nJnfeA9OekcPJQX4vfDmiPg4ys2JM69eW/8oAoDIf5IcSg3sNvUcU4Fg06qflki4kPHugcaFYr
B34PdEQWWtk5/aJk4ITEuQwagmXawgB1ewiA+33WNxSBI4x+Gr19iAeo7JJloKLLS13w5Wntp2Xm
cIFMDqNO2QKPipyxyv1LTzWwBrJcVweOnhBGYTQi7jpBKlUXSVtf/j7+eVTXulfueFmZBQeSfyhx
3/bq7mzlQImB8bL/t/9blnbnkbjUnJA5Hd1l7TBRyVvts4ZMxBpGesh1/IYxWnVzVVaUU8QMOQnI
CIrmgGDQ0WtKzxJ1j4MZPmvk+K5B2hwHO3YENI8wogjdCHV+T+8jrB7zFAen/1WqmdJqX6FYZTVu
ol2PBbGxqLFz/EqQtzDJm+g6hnx6FXMT0B7xJcw7sQ08VRyBSlFDJCPFW1Tq6NHGBcnwef0dW2ht
WuTtBB0CWhhBih1639m1moDDvPh/jDtYjnOcvUyebltsoD1bSkl/daG0j2QPH0WlAgMICXiu5OXu
vCQK/ksw83BPX1IUy0GcTCnzIlpGiWGi0RQXpoJM8WQ8x6GeblFZwFfQrfhJIO6mrVKmoqkVZErf
OuEI4zw2PmJBxKZ/514wIg/0DJluk2WmVno3ydQdx1m1jnu+mBxqxfHc7IUtrrKzgFT3j9hE+KZA
bX8Ej3WL/x+5GeVv5HVu+l+pLxjBWf7kPweu0AfTwzxjc+s0+3A6akyBO01824x30oIE1bBBIY/c
zmOt79ZPAEGL76iTq7TNxkMp2ag0qGZU6aTAo7LX0i4L36VN126XaJxq60akQRhFPPpSPWYmtKOx
vVcfzUa3ALvmSnevt8lJ6JlI9r6wPgAE/D+4j8eqCf32V8Hqq37Xe0N49N9wDySpbgzEojYW6xqO
VM7A/5bYy/3dHnQDaSmUqXYNNmzleahw8Uog+/thA4orBIafNyV9n5WhUqwSbm3Zs5dsjWBii2fm
lm0sc17ObsVoyUzFHN9PyrnpK4o4jaa3owGzM7AhZK4dWnwc1pXgmrQ4ABfQPsbTRgM73KAhbtSf
kKjwYwJQJZdg7YXz80EUPMPsgEDf4Mlw/96bZS3THESEIxcZg3j7lrJmKIl/chX2EV02rsXZweAa
+P3zf0fLuQrQ7SKuEHiKaad1kG74lfeIFEJy3q7shnAGw0yDvAct+phuRGUMht5LkpB9ao7AtVFZ
0crymGfG6R8t44QTaOEyn3VPCi7QXCYs0F+NzH8loacUxleXfez7DSNSGS+MDlx45wphs2sdx0Sf
Lh5CC+MoCLGFPvNlIoZfpj8yEUpOsaLBA2+gsbmwUTeCx2KM3vOohMVWd0SAr/SuoOlie1qN5C9i
bM86LtyHXbQxsBH9jSmeH+GWewr03ZNgVS9SBtYxpqTfPbH++ugqcK9WwBcKvaNwOpn/gEz12q8O
Fbu15JhG65X9+jqIV8uxnXCa3fwFYYpE+zkCXkapFyQFlqCWv22U5lUQlNv/qYtBJBPahL5xLGyy
onC6ER9cisdDh05oiw0py1fPpMEagD5WYPM1xPy6aRqx7wYLGaj2G3P7puE4AX8B19b8q+39V7Xv
ykNa4ZxEXKio2PLo9owZJrJ5e8xF+FNC57E0Ir+KtXHNCY9I2KRg4PdpQpU98oY36TECwm6N90Ih
PgDI/8/eCp75qHVk7TaAXpMwGCOZxOLGYs3LxNAzHhPJceaU/R+LPFDlaPx3KGr9c9c3A49S3Qp/
Hi6eFxg2/pqf2oF6lkC6rpKD/opECHxQ83fBCR5vnXuhiy+5Zndu3G+3jTOqgD3Ia/SKMvC6hEHy
DJn354QUpWULRedloiizSXBxF9TBG1XyMNf7ggxTpVw4GcFwhBvs0VEnqYTPs33c62oCMcZx+ws7
8tCuJ7eeVwNOVdvrhA1biJalrE6+k8OnTOyoL3NU1OA6e8+rLnMbyidei0CN2cZbp769NgUgkB2P
849l0BldbUi38vJyJJIzGJ41t0lTuxqHDtSkQwm1dG53qs7Khs/yjBe1BW0rSj6T8NLzdsHVvxqU
aswmJLku6MFl8oQIc3o/ZbouxeXjKeckXgq2lzMevXFtvKZEntBMhyQ7Tj0JOYrxaBZ3jcoqILqA
40S4BTi39gd4ArAmLHfGYdcJ4WhZFnGnwcuNnH142dtDgGFvpkZPLMEvoWc+Mm4Xp89/xnjqHTtw
qSQikLfkC9rDorxHN2qq5FNPyC6ytyr+fpgpsqrnzZQLQ+xU6YFzADLacG35YVqEm82x9TBdN5G5
zUkd4iXyop83G6OsBOuxKBwOCFNWCIqQKqD9NTzhbe3V938ZRVv/hVfJg7miixkKhQUQ6kZZtdby
vpoLIgrBtrwXWxsQM2V/1NEI18kI8oYvcxkXQVW1gF6bGAHY7uUvuOs0sRrhk0B8bJFfawtwiIMF
12ijQIC2xnV3YlS4IyIJGwPX3+8GI/k/lKOQsDfEyMjc+j0P70oZSXwwzASjZaHlvDoTRFt+BnkJ
QaCo17/boKBzQI01ZEsTYCYd5RjLZyUQq/kYUK9GZtDTVDRfROJdOcyZzQwm0qT/U3c0GIiKWuqb
NZxXEIE9VSDNdxwVmEvvB44MJhMoDkmgWjxch5HkhVFDb5xRfZ5smO7v6QTAS6B6f8wKtMu8LdTd
V6THV+2H/lkkSpfRYAUHD0sWMDXV93/hA28SsOE38rHIcRResqqVU958KYVYNnP5tQbqc+cxi+v6
9+i/U9bH/jgaWyL66dxd5BReWdQhO7K3VQbAouTQcBi+Q+chRQuJ+HdKz+rPZjWxwfdBlw4yUZcM
4cKxjSgaabYGf7bzQxhldcIgzXaUHYuOOtLyOMfoFSWlu1aCw/OD7N1xoHe7CUc7Vml7Xx7t4gSi
Rv0sppgn8Y83CuZrW8IbfV0BmUe4Qz9dAGT/sLlUyqT95DRvsgOwc94R24UdtPqr9qFfL/xmowtv
Nxunfz3Xj0csMi6bBI7OmPWNRYYCV9FRcZQuiaffK8v13tLZ5cnIh9WUnP+s1GTRLKLoQ5f7zHJC
WDWef7CNVXR8aKgkSAvTIIKhObmmNM2aYItOWA+GTrjXlscpLpFXcxxfjzIjZDMoAR9KZEdu8s1X
EWNhAz+DF77+Ax0YLsrl4nUD5YKJKgsfG+UpG48X4eQBdy/pVjXIGHxZU8zPLPnYFxJ/bmAp7n0X
6YJcy1P1knbLWG4jU/qdL9snZuIWVqd29f7e2joD3SRfrUaJCtPpxmnGP2cryD5iSkyHDZM6NAXL
mYmSpROZxX/bGkD6ZWvTt2OiMLNIqXF+xiCdj1IgZBi+oB6UZlAVUsLUgNHoE8L46p2iKVgNzXhq
Kfy2Hs+oF4Z44wp/SjIL+p940i+b0ZRj2d8gS9BHcYZ/h9Xqr7zYK5vIyKrlA1OYybNa2dC47t7B
qTTg93E9kud0eFctaipZBUjiGgp6vB6K0qUoOHhEWb/XJ4ivWNesXrHSdcg7GwaRwdiMjJKEdB7S
SXs9JYj6/9LxJUUpqC/FFo7KB5lnhYirwffk5UEF+JjXIy47JU7MYZz/FEKVgspdxPEc2TNI3QIj
OtE0vA8g0GO+5KjXBTJ5na/gJlgAa9938X68TCrPAPH9oWH5+JIHXsD6yOBlTVmpExJGq4sA/VFy
3w8hXXOyKM/tGrQS+ljW3vcBQIH9e8G6X4Y+g30YoeJm0qJ0/ZLAS8a8GTSXK8ySWRy7trkB9s4s
4/Il3Br9yRqil/2zg8WcFs195sISbsOG4xLtjqGBkPzXoh27B/mHE+iS0fc3O37N5RSF/4Zj28xt
I/H4SP3fkBf01oTDStFu2UVEcbgj7R5S9YznFFJpJehOaDkcaauUT03LFM2HWOReESCIsadqx7rG
neFpFcyOvjUMWOKvG3JoYMRCZLg3JY/Z4hSmEoBAVvO+spLc0wKidJqQy+BkCbRQacjDl4cLsZ/D
BVGORO02AInJrQTgfC+djpCPUFA+wWd/XvH6SuHx5QsES9bdB+S5gXf94xKZuzFMloqxmaHNhWS5
viNdbDIFBFbPknVihn3Q2fvJZydlL2fVmcjtwaY5p8WynTewhgpKEWgUck0A5onKYwE07nsSHoQV
4c74FT2HhpqdQ9vckNlEFzKDGPCwY3bLExK1N2wXNUFoAE3zQT1P35AtWZuMfTX9ww943wjO9m8z
Fq4/ctg+/TVGZlS2Dz6fogiGjv4baI/SeOAGH+rpWrt+ZxM6JQKBJT9tX6ObVrUzRhVE8D9ig7eP
Qq1wpq8qBZacZD7tXU/pJLHImJ/Tf0Y+WCTnk2oXuuRTUG+6SLoEFvbFxYq6iqejuegArqlsN/Ss
u3K5Ut2bBKEYUHPcJpDAb+SznzIgjR4Rwp0dUYPi2m35qYgyXRcWB1rxtVIJbIPa98xtr9aE+KI+
adl/fsCDs/m6+i867hjJFC9Ng1XoWcDs7/QuVuQTRdz031HCiRrJntpwi+kHyctx+Bgq1To/liRB
5Nbc652vEmcNP6Sm8oa53sk+VWbKAET6IydnZnU604j9MSb+0fi3uSpNjoI3wEnnkoW8YfdwEvkC
N99D+zvJOWcLFTS+kQ1A+YnJcakxLMQGHOQXB32P5Jt1R71dPV7A/iluqiVy6v8qvmvjQkZ9Mmw7
PSoWxvhC4Jah20mUIpldCSyoieXAKUE9rifLxgqVC4LGNywjjcc//9nNdrwZJ/X66Wn1/BqKxns4
aQG9WhheYcJERhqbeJ7wxfQb7nDRrDFUhTmoeJDGBgGkkylU+r2NmHkZumR8CW0Nb3EupXdpzObG
jwYZqNfSOcWBsoxFRB0dxRXttQFF5GE1qdho/U8dk73rBfW1vJW9lyRsi7QnaiSB1JRoxJU3XULh
EoHwdWSczVK2DMRTukaCjY6GuiuwfZvYd06Wnzvrm3k2BXAYxK3QJnAclDcT6NyelG1iQROGryvT
QzhHqz3eaEl7hRkAMNGewZbhwZCrElEeY6xn7Ehaw1551D7vBe0tYbpM32fR81ecLyJA2qixmKDi
sh1dJvqSumn+1YgsJFJB05R6DqX5SmkpXMCDiAZTCcnJMooRuzpZW1BdPFHBj70BkgJRinmaDeUm
7HRt4ze82BGcKUxM01Xd6nNhf5mSYetCNs4TLX9AkwHAiqUb7zKE8wkOqbVwcxqdt1tIh0fprlnm
Tg+tQSLbrJQl/bB9ifSCBACbo3S/L0PLieko5lnFFClTIYCuNNJF5PRhCRtBSFabt37+zoqDkssi
1Jt9q+KZbIJwKx0jt0+CJ8gTiOfSwapcxjJavgNcCRuRJ3cTuwa0l3C752GdValvgo7m3ilc7E1e
FJYMELMIYcAndHEPy79PUf8KwADwAlo5guGxlMBwDxGHwYz8l/BU6fl0861Vg+w9AivSwnrRDKkl
R+FujNZMXTplwLUTbDuYqVllZhGJzfRiZ/AxyWYrV+dx6Qgf9az5yi6UUbpCmewCBwTU8USit2X4
ptNr3rSOtqOnzF6N1sv8uEt+MVar+ngR7L7yQQJJYJpM1rqS1bn40NBbt9Mo2B4ldmlfBxcO/+De
El+kbutg5yQBWPjX+M4FmYVt6hkGyWR/ALwTB6T/L/CkkqJ+R/8Woyy82k3pef1paeHuw16OXjLr
Q+vW+mFsvq+o15Np13uLcpLBOBdGu1Bia+7w3WWvC+4K0hq3SOjTkJ8zAAxlzYSfo5Ec5IPAOfrJ
TUhlNgN9hNDX1lFqpYEHol+Lm1OgPMnwEaG40cF5uBdMkYdacIrCsF2Z1e4i63tdFfozPsxosfPt
tlwxc6bZJqJCzJzo4lXV9Er3oZDsMBf3F5YNa4Jcw5JxUL7cxlSoeOFQe15CxRCMs7BECQDausQc
jeb+CNEiSp9neH01OObqzdwh/C03PyQNtrHlVFpYAvhDh2s7Gftk4OLtgsh+VG9ef2IlLCI+uOIj
fRM/2rS203iHqxcXWcb+SipP1ReTxskCPf1Cu6weHwg3z2HHGxv8yLHE+7vwSXKmkSsYC9uAJ6K4
NafoUhHopGLsGwTJpM1LsbTYI1k2xP1i9odGqLDIfQZaF3auX4YkZSEJcOJBl6gHfygnRzEZFX3Z
GZ6jRapBz2f8/lRv6dptOnYpwYLDIkI571DD3Xif3d3QFGGNX2lebXJbRO1cQUFZsC311S6fR0o6
elvaiTWUhvExD+3eZ9ndckxlP8PrDXNl8q0nC0gkYM1fmTFTDjcNIFpmlqtttqenkF2VcX4llSw7
dltnqxmpoUkrahW6W3jWevD/5wI19Msj1hG6UufqT5mPZ1rEh3sD+QDfC74waemiL+fgtuM0WlGz
WaveU29xS0a4BLeF10eGMrCQXi24m5q5GbFvEbgw9C5dZadRcM/e8SNhzi9QUG3lyAUTdMZvPKsk
nLndMlVyvu0LTdZDkrkhWgMSg1V57EHBTJXOFxGio5ge7Cr0boPZkS7masG0ywiZHa2HmQ9lgtEY
xJzOt7XvpHyCnLGsiILi73sIdXNoGzeIpoqfoUAmth6GETfIyLGLCghzSwIVt+FsmfAASsmc1kqm
wXFM41HCs0/NhkfqtM/8ZdYJg3aKLBfD5JCvj+KT7SjPTozg2Jt07QWO/9tEJicGKmKuVjSilfyX
qgz8QZ+tFs7Gmo+pjalpAYmF6d5bN6/R+uWPIW2dH4mAf+jjil82zqeHd20QucYw8GENrVVnVpec
D8oWrjz4YwqZOpFpye52EMGY5++eDexnTseGQc7TJeQKnKDtWq2Vb+2G3nU7FMwnBzMjf/+M2B7/
m0V16G0bA4HFdu9dX6YAkWaw5wFeXpYDH+i94vFF4pHD9UHoiwygfNjYrSVJNfnBYy4TVPQhppQ9
g/e/uC5D488R5MqsgxDc21bII8yUbGcwYcYujHBZyLg7ePpgu12DCa+4Fr+RKK5gARvLBsiBba+g
GgGzNV1ws/dcWYEjj0hQwXJQPyrDS0qESYOeseKRs3KXkHvin3fIjJUAAgbsWtn5zmNL0w+HKd/2
+2MOdEZz8g97DhJFwkXst9vq3hwe12qmKzJAteFpRof+PZ9exOXzDDUL/wcaqKOuVcrUXdnJeWt3
z3nvCzUBVz97RAeTTvcxYCYJ42xgF0mgxIjzaD//eh9kAad9FWtSzlZNKZDA/IC4yYpgedf/4VCT
p3xanjHOOJ2ojg2AwzX9pB27hwLs/X1sPG/3N4Lzs8ihjlBiKfLR2TGalEGP6gUCBv4XPs0sECAX
EMh5iHsTdbtOXgalXQf48K1UCFJ/3R+j7YdZqFnqi96cK2Ugmgr1IiLzmSP5MTz0oWSXpe++Srx5
hzw44B0mUEV+H9x+JOBrX37zyTSQlPDrd5YPsD++GBCmdKb7pc2zRmHH3tcFsSKFmlED2gwz+vHx
BjuHskup50CegWaZkSad/juVLkqI2fiGGaCJc+Od4Rt80lCTT6I61rwatsxmEIKyJqEblNfH7hHz
MpS7E52f6GtxdXDdhX5qn3Zixkmv62JuZq2C6NWxeGYQGLAdyhumlvZpjezN+0zA8Nlb2eOuHfNt
I1IwdEnoteRgXM8BDJqFfdjJMvkN9Gp4xblEUi/JemQ+tYJU9CXR3JUoC+Txhxtli6vG/OGDhleY
L91k05gJH34/WMgs1AKqz9CfYic+1qXnsGtjHzL4iNTxZwzhmeWrRkQAIxNMGFfbxZYPZmrFOf3f
0XovdqvrVUtBAn8Kb/jnyySEBSqQIAMwOJKzlEpkPU88nwvLHy2OHOLeR0/w5O9XiLnyKZ/Lv91S
gWy3yaHg/xkYID5XVwkRRvv3SgSRo2lx1uW8XeeG+ZrheC24neyUgchpQQp9uQF6dAIceMubiUBI
rZS9Ot4dMiWHwwnEmL3k9ODOxhEzihMTflyVNtGWeMIpQTLO9y9K8SqWEK0wYfg/vaxZhbWtB7fy
+BQYjOMZSeVBweSEkG4DA/y64HWL+RJx3c0xaMFue6HO3umkhfbtHQx1rIyPo8GPwDAPlO1qQkOM
cWokYdCjHEruksnwkGtLxljyrCXeoMpaxFJUXO6tSO9YUEh0UsyGFxRssdiUWws8nKCufu4QC/31
J0+caZIrM20BfwSzsMSaUqAv0gO0gJiHdzlslbcjBP+i+1a2yKReqS3T518G58KNPFsydrSmi/T5
4a3cJswkhXV1j250oqXc3rtha0UhFlQlve5jbUijkYSsM09GISEMkAQjPeff2frkbkNKmfIxtbSi
2PV4PZFhc+d0W4PTyq6dHUJgn3aeYPMPoxPc+pObEjlPyU7JrH7Y1SFth3rfnnIcTqwOs+1xi6r5
tkRF37FF+mBL73MxcNU/DbRCN4YOCeZglIZmhtooqBjYyFe4YM/UgVRDD7b2LH3pNj6ry2dalt2t
MabazRP3oTRzXWaARm+BF6TVsM2CZAeUVXsm1NdRG/wzaK452cMkD90OIMbPexrqGLrDm+q3Zvwv
rOnu3mbJsvTPYsrVBX4bnm/uQNX1SQnBu9S1q1h5PO4E7SwKQl8l5S3/1ghO76DkXD/QpV41kxXE
FHS0PZBF3SWGCs242NWpao0QbML7brVw+SzQ1GK6f+/kTnWjnHWplIMBAACDwQtOfsbvUFCI1Tt/
nNJxyEHcY1uq2uFSafVRej0LjiuvZQhvVOtUobsUuCGKb75lBTx+gNDRV0aMZ1gw3aWTt4vSh14h
OoPoGdoYSdZnAp49WYusD3xVS7QHDnrpS1rifTaP4cog1wwxbVBQ+jPrOuYOTgR1dXmNu0ES2lRS
1BmWUgDyT+Id7y2r3Ol6+iZvFqbmwBXIm0zzTW5ZkYgWprfTZfmvKOafEe6wmCga/OSB0U+eYA/d
3DiChLa1KXbXQU5MExnJsoEXrhXbh24djqSUV0+we+hA6Z+4jrDSn4irvbFLB8UdCNOH2ZUX/gQl
IRAiYV5ni7j3ezgJfiYUItfLSy2jwKT6USIlkcaaKFeXKF5+jIW0PBDdD88zeRFz4XLpH4a7y/Y2
w/rr+hSa+EkORHqPGnwqNfgKjLgsrlpxWSeFgCEno1a2sm7t5BZtAtkvXnxmcMXXP7Xs6qKLbIJv
zPcqLFS+t+r7w7mRBIGaYb0jS2c7q4W4P1QS6VPjdFEzk8TOLMnfUBCJb2LV5jznfZwX44TNLzgC
TmQX+ex7TygINcTCJeqNaAbjltbBBjCtUqn25TkLn0sISfxWynOUyscqEJMHZ/fe/2ji7Au5k389
1H8avN8f2koenTJnLLTnALevUX+otVzAehlIPwQUVH+gRDRqOepchGAvF3bkyq+rC2ZpDcbTQ2kX
MGGQ60ymliAwyZD2HkHnzBjafPaHEAwyqzpjVC/YSiUEfFmP1+Dr1vKDSSm8so85X8D0H8NOW10W
Lm3GcfkNMMQf/R5B2q/i9xT/RjP33t+KurGFD3hQAmMJNa9BS2pMFo5ksmv/V8vqkbbOCUB/OodG
zodoJ5KZHdCPX10h6o9JwLmhzsS8XMzcVJAM0hneSb4FgU4Nbx1iAGS+Rr4VlfYh2dMGs4k4TUBk
amffk1PNwn0J38mSnKR0C84HFdQHgbL++aT8WYcnEZj55oTHXKR8dkr8tWiIK11Ck4zz2HQAoU8c
whozZI5EeH2dfWi3RN8TYKwFaeVERBSIdlbO5aJtAlX4mXuTRL9A2cOWhLnyKVS3/3qfbcu0vpYF
MkMhkhunuPHLxSqiznWZBohWC49sfeh2azf7upHuTimxY5ONsiwnZp5/Kg6+sbSh7CwML/QzKw92
nejRhPbssKQKuXdZsN0ASOKbJ9GRUqJxCdg3rDo0eBcK72U6h7IB0x6tWPXmTMEOor7mBd/6Y5rG
EY9MnJNzF21ugY08W/9LCicQxmpizNBEnSMuE0VrJg5I+NJ3q+FxhfE8lLzHTyychklmyZvEfjDz
8awOO9xZms1mS9kyCS+zV4lhhFJwRI+6Au0pZqAVFFHn2lBbQbDgS8cE8txejpv3Zl8PTVr2H/3p
BcR0+SUKAD5HudQiaUt8xutfK6V2V2Zf2mipRaEyZem8X/cUODDSquLfqCMoK67ZLnMN3k7ht/7s
7JbwkHQZERRbbaICklhr1I8C2ycdQ6m6/iaud7Vvj7xA1SSajTIFnLGL9SQcEq//DHtHcoQiusWV
ZR3/x56A6M8UFqNGw3QQoFTPx8i9CVjFntf4c3t2y8/rNuiGEMp1qCxgGaeJxqwMswyGJk4biqwr
yyCj7PRC51oSuTdqS5hY7+POXtqKB/vKylKignmLGuWC05Gj0V7aQZQJtNLnsPBA+OLDbzxvhyGk
bgksYSZDoVO0spJ1Z/Rk4quLMInZE5YZgnBkX7pf0jPj/xD7n6Glt80N/tdGFrcTEW/BUIQhVmKB
bbtBYmD6cH7zEX2AZqorRRnjoNI1XBaVrvVWjtCi5YjPtedHKfkT9psHjo8T54WCouSBgk8F4Ds0
dgd1dLxUQmphbGOO7u73mx/p082AJGi13hIHI3jfah2WLtrPrIbQlVaXhg8uKrUDD5zrxKMMc+Fp
7RcRRktnjGyWnx93ISzFReCrE00jLac6Ueh3hrOHHDN6hRLTOB0YCsufvh7YncP2+k69EUr7JV4C
2uCFJ9lseFoLwbpXCvgxKgFb6TZ9BLh0XFCw13u+7LbSk/og/S7Qk+HcHJgeM7VVe6dJnkt5MUbB
vbkBIf42CthMMKQj5GaRoygygMcmU2Y3SWasG23fjZXblqZFDwbth0pcw0FGQjVUspZnJ7JjosCJ
EWJ1pST4vQtwaUupkhJ4M6DeMm2aWBnNFlJ+dP/c5d1JMROcFbIa8xaxkOSgWw255AD3pHU3Itvu
GCBZAQrbhREhFjzo0kWCGrHevzpRZg8TO4PxHTD9S7MDrE6pcZZDspRyx/nzbWikDd+j73W/6iHB
FUJvd1uclNPV2atVeAiZ3+uoVQK+RbWHCLQPX2XHagArfYT06IcfzZpJSUSSh2v/ZFrRSjDekL5+
ghhOm6sD8OOvDr/Ec59Z/8i0XJ1ulXK7JwTmwfsu7oegniUyDhSf+WQyz1BGH87O3gBjwQV8LZzH
bcWjUvQjmWYH8JsjPafOXwPeiH9J4gWyi83Ia6lKeykKhr3ly2T+x/euNfn75VN5hDABdoPoEA6A
dPkXEUF34SErkJqyeRn7+zpXFDl2fpvwtVFQqaxrlSAE/GOlHd+nzD3LrB4Alh/HmDAOWIqHWjAG
gWUIzeNilsEh3qKdOF8UKewM5G+NLwOMK6C3tUujz8v1hnR7R+zRwFjGejKFyyR32bP2IJbRgyK7
P9XawxPksX6S1jIMXv8GNBlIECerBpoeFeBdNqjTrv8DurwYU9zBRST3yzse+TlTyi0loILOaqMK
/rJBQGH6IQVX1gG+DhIZ+TIP5LWDR/MOQlw/ivx/IuWk/pADMOPmq5YouQFUEviVM6p5a4dTx5YL
B824D5lg7CRqeoxrjVMmA0osTzoxiGBl4yQ2xmSrTLbPWQVC9/CkNa+L3zad5XuFYvANKuNXE4GZ
rh3CzKeemFBEq6OjFwL3cHr2P5zVRY0pWJ/MozEVeLYi/1aJhEu1To0J7Bhq1ToydgXDK06TXomG
euPMbFXsBRmQs2UO+Qj5C0K4WlX+TCymBQxlwfVsQd+3BmE3xqNIdnRGREoa4tmlAIaNJhorlFDa
ly9OlWa1rzn9iv86Vkjps9QEfgGNWClxPKHBMJ8vkGmI45qfwR4tuPvQBFZbvA+FUZ8QTqWLLVVi
3SgNC03iCTRRYwxRKjaDn06CODXBVW7N/4eQoQTzYs60j0WbYcovDcgB5fYJ3srIeifUklQGl2qU
YofOW4TL5v0aPmgKZSG1RIzcKahEgy28o23p0n5Kt1E2qWJ3yfS4iwHEZQOJNuHgQBmiwE6i9uhc
Czz0IAxCj3t8Arce4EIw0FHCv/XB10EmKV0qrH7HIDIFsTX4fPFEfL/2VBMRvslMOMTHmHJ+EBsc
k6Jm5aSLMDu3Cnm6Kbf76hyaPNxKp4rjaSTRF39qyOMwuM6mAvJngWtqKfCsTwfVvWR5uI0vki8d
vdN9NL4qgv/v5zfD7V+Qk6djmxYG7VpN3NKiEfgPYmcz3XfvSc+/oftdD/vfsI4vjIY2V0D0+VeM
oGsWxRHuTgppZdw5v8dQOEV8sU0DGtlRls2j5WCvAF4jqcMcp5KyNhxH3ZU0p8tpOIrxd9+7Neic
xVQrUJI5leDk6YunZznhiY46/EJlCOuBIfll4cOLUBuQHRB5z2PqH3oA76qZi515db+2pmVkQ2mv
qQomm5O0cXD93YEiSnaUkH0LWaUCYbHy/eWv9QHIDMOD5k+p1qaJlR3GQ1ut4TitYElNUu8YwlUH
op+zE1KY08gI8rByNAj5FEtb6SUdhArypjsiwlbGqx0T/hJsAfqEi6OHCXKyBGbVIxvRKxVVT0HP
bE3MoKr5fViDLY2z2jDCoWRHP7ggfZoxjTETsrD1aEmGT8rWaScGl0QX9PZu8Qqs59zyX28ET+Lx
nBHYkqRXIvLxxKn8D+yqokANUpzBfpL+Nayre26TD2WNXPO+3X8cyGE/Poh7Ho4w/XqJQQLmqYAP
ol9Ul25jfMfjKFXNJp64lu7ohA4j9yxWAIZDCBCujM3RyD1e0nhpuWKdCcVYkB6lGggZuGlB9x0h
6NYp/fLJRkClPp7wLkpyNhudR3r2GoTsm6+g3X9tpovkh+81J6wEyJlemfheYnoAMnCL1KxFiCw5
zDV56UKR6jtI8kGZ8RosXOtAnj5Y3j43ihZggda6yrnbxD+HgRH5trM+dfjABMJEHVjvNkowvhEy
7nYQD3jaF1YdGqU1Be+W8GcSU5TE/n3OhO7H3kPvPmI6vavIizj+FFAjv3v3DtD44NkKtJI7Y29B
yynyRwn3eIzDBbzXp2CfQrD+qws0+iTtQsv6wRXmdZlGjM0o6Jsti6bQS12dKUAoM5LYTtbbGmgG
mUw12jUZtB4sJ5Lsi9AoZLK8f1RZdFUAsSDiAR2QuXJ+tT0/i6UvjG0EsP1HhtMO/jAQxgg/8Ya+
mxI4Gp/nU9f7uKFvzxmYY7M98noPtwLH4WgyS65vxKaCAN5dY2VlISSXKMiLymikzfmsj3B/54US
Ya7yYFdtmav53uKdTb04YzNP3prKv3dsdwdICFyKUHqiOpOF7sTcwTu4WX6kPxnsv2mUcRgNcf0r
Z7DOCisdY0GtRp8xmJtqqmv0YZlrRacXR8dT6NTCKxfvRJqaWLHfxg077l5EFL6knpSukQ2ooIHy
ZcyY/zYw1/HvkneRlLCwiRYQ2XRv2fBi/LhvW2YfxcDUalwjlHJOSYTATt0oeE2sCKGoqnm/6XYL
7rB6LI3RkFn6BwLDGywztpQiIvW/+7h6v5+ys++Qynd4ZILhAHCb9fzSXJOuzYD+A5T4p8YP9g0B
ufj0TSo5oBsyYCawLxxuzHgM+FzjRwrl4LWawzKYfEiVZM/3nakEVczT0iyQRYXaWgOxKhFGTZh7
FZf3iMMugKSvGeYjAXXLXAey64TxTqgGVf1HkesP3+FWgHP+oLMpHB+Z+70zSAre05dMh6AQ92pn
IJgsU0Lb6jGXr+e1bWpdrn15cm6x3DsusMXpeL1SM7/ppzrkmuU/mcCSYJLJCwILF8fDQq6s36/6
ebTAHpCi1t0rZI74Roi/Py/ImA1vDqiqgtqSewMIixaH2gUH2orl9i8u71ePYUV/OcOsmxf9CnqZ
rRB88YVdPNIs+JfxFq5y7kOUd53E4JVtlhCLKq+UmU1AszpJwqbEJdE2jMATKNo5VHHwAzuZkmlz
4px0HIyd+yS2/H7YpYFzJYXsv0X/decvzu/nJee8kKwSMP7HcEsHIwFEyItOimSNot+2Wb67alYm
llo0XtuS1gEUNkQm5AYwFqSpW5U9C+dI9P6AbGwhUTC7KDDim1q+FDnnpdeu1I6TQbAXJdbd0UBc
b97ae8+Jd9kW/kNymIfY+7GfmNriKo+5CylD7pmWiqJukDBIFRZEgkPp2M3D8+SB14EDAe+t8uKf
IxBDxDFk77IkETE7cCPbV6pMy3SyAXsbz6iDc2rG1fmAEtpxMtYEFE7GVSCYmh4tPwjlwHaRhVU5
0OdKwOJQ9MHzEFsHO+QHEpFmZdBH4JZ1corMCmDb94Q9Rjysl9UN26IFXf0ExDEJD0px0OBqivJ1
P3OJ+HCh55dJm/WS2ug49DsdtBzuswyDEoyVM+Ge7tiAoi29FDupFL8SIkO34O1InVu0abP345+c
S9/D9oDXSn47az/TxCekQPD026LZVFcvVUiZZMAut5CrjS+EcWtLFoIYkvfeBiKyGETvtzsd8dfh
Ki7+tO8jL6t7NHX1sCe4TNteWzcjkyFKds/JdcBkYsWipAMGGdGOw6R+ax4kh0egglzdJ62OgZD9
vrrs4dW77bv35hv0Cnc5PMd8/jq82pUobgMStEV/dQviizEnFU17KJCK+/IkAreIncE0w7jiSqUM
xz/ddIW4bImr44L+G61QCx45uGfvD1hzAsy189Y+JFU/1+z8HADGF7p98faDsaWTSlxJdAthXEuG
rYrFH4gart+JpYjYsdZpuWGyrXBTyvfPBgPh1oMPp1s/9okDiOc/6gqwgw9kUUCiIm2Cgm+wXX+V
Fna94WsSjZ3GbIPbi98q29kE8HiuFKPSNu+7AEXv8mTeygKAOqYWlX6vBojnEZzf8ZohrnIrwBbD
zDXa7+RO2m/v7nsRE475JIQCUDPjNKL9r8VwMnQXJoM6SQNg4LbYC4NNBTZuGTqNtMyeSkHys4Qi
rMMihUZR9vw7k9XQJdvDgSWD5E3EoVB+0b5o9Vm2DKvCCU8a6NLvytzlvQr1RsLzO6TbTvYaCfsC
VzCEWxPTJJQsMnGTGfUe5WEw+DtK40r+iiTpRyMAAfuh8lESk2aqaU+AoF4JANIZfPP5N7y0WkZq
eIJJEZBoAF+KMga8frEvx6bEUGFENdCZNEi3djp5DAPHVWFLucyvtOl7E08T2B4wYrb2RvXrmg3g
Bb3CBBheOQ7KpWV78KxenYNSK/hIW17QkR751JFbs6pRAGzaNADc5++2Roo/CP6dgpxYXEKcauWR
rxy53VY8L3e1PeF5qgbmcVoUPFJTRdOGhGlo7Y1dFk2Hk26T+Q6MJ1aww6VncfQDesWrqsw6xuh9
rDrNWEO1GWoXMBldv4uMQT7U3kRCcYg4K9Ou39zP6YiltOn/BejAWnak+4YyxNTGeUQECiFT4E31
CK72O+sWaMzALBtXv9/QyOc6xdUVnK7ufixquTbVNHAaQSKOv2YsmT75fQZnAIg3Lr/TISs+Q3ew
ctVMX3kXcDGHxywb/yDkPcy0WhvBvToerSpzDrHdcGKlhZtElK7CUlNMkuk0tyLQ8FX04lThnOKZ
Mxh7hCScOh+e81R1yoFmFeeCe5mmpWjsklcYSkd8lAwzNfwCccKhch8ydT9hmGa05BpMIiqNOTX+
UUtQr7uyRouCL6kIcPdYQqjh1pIWL/W6GUj4fotLQRHyG3R3I7Y/8a6XyD/qOkKkA62ZtX3olSWN
SBdPtEbEYo643jJ7l9SUodfNZLV+31+dDHp2/c4gXWlDq7blEHmn1gW8j+JOST18pDfxB67TXNbg
DqkOjcPzayAxu47fj6ReQLhtDNfe0nJXM8jTdOpU+X6YDeWA+SDCM6ZLeok3xTfodJfAwgvSzo8I
8OYHKa01qlORh1Ci1i6TRaQ2Tpfo8jk9GZImegRhq6oO0fCwNi4BeWRZytxj8V05Q6yIjFbunAFF
raGarT27B/q/8N5ahcg72kLoemY9cArGzLIdrAkbkG76wCvVQeXGrqx5YK4hNYKfa6KRUgnkYwMn
00VJUcoXJGNVeZKI3sVjvBDRwxMG6sXZC6v/k4Hi1le63bQABiOOkQl9z+WbqMRRpwJezvopnbRk
jtPhudzBY//M9+ohxpTOjsIT0znwWw+EOcun2w9d7KPYt8nGIjvAKOjnhhNUKO0W3mp8Ol62hPcV
2ILujadVCPD21Gke62jbA5DWYxMBhkxvnyDRvO3R5PKEejD4cQNmKHQpNY/qbOybevodFj854mDD
KuR+Z6r8P/fzFQaPsshHQPyxklGp6nDOQUx00Ht5ohM0agfforkO9zFmZQGt8LxAerUSviky+Rrl
got5DQFdI+qPhYO9wRL6L2/2zsNceDGVabkv8mPnoy2p2xbRiE3I4sq9C7e5l94S9B4tt/WT0K3d
l3zWL5CdtNoXnh2M2ZjT95XpCXogpZqkAa9y80sYtAghD+6urxaYWHljavDDn8OmLod+nE++B+wp
hDS/bbU2Cps+FwaAv/EH8KISkRSudkbEYLa6kDp4TNuYkH/hc29FwZ+u7x3GIdUjqJ+gozKZDK3H
ozVEh0W5G2A0lmjePRwgMFnRdqOSWoCz4fdIPnurtnAs1wz3aIjJ1LixCy5/aX9gQ1shWZbL0lR+
mdnPad1oj0J26Sukpv4i/g3qDhMSS7w78T3qobrzLVk3Hgg7izjc76TaTZoH3odkI2AVAtgYnfKZ
2k7UuzzGBvd5ySmkVYU4HD2H6oml+JEK0qgaQseaj/aX2jtJ+PjbOubEg4nFwISfL69H4tRyBfhP
huLg7sq5QCqJGKWl6yEqWZ3W5WHXAe+Isw5rM7gPqLf0wkR6oG1QA6E/cDXojfISFCO4sXkE2mRb
u4l74bAfCkkNryJYi/dCa1r/hn+OoZhoJjEuFX4bobWNp0a9AZMte8lfCR+EgRVjMevWN95PreR6
+hbfCcW+PUmkDFsb+Cnai1SL55gc+Yoxli/0aUWEUBYKjxcEbpoWqtSFXEC7XZ+5hN4pUxgbD3X0
D1jzMLbxZCFDXjxAk1oqQbpuUWLEOiqKaO3r6AuFEhQAMGEh+7v2+EJP315rGU9W6VV0mJWhkRxj
GJKMbF7pHLGPKcOT5m90qoKdZarxISQikbQzkTc8EwIRIS1iUrq9Dem3el+cWTaV167/4hOeotB+
+h1dSCwwlV37TNiTjukDJ/wt0iaN5hjuQuGfr7kxRn6Gk6LBaJrlomTdsydGTchFpmfjRMWg8TkA
0LEgBb44IRnITgRXWoCfKVpE3w5QsSl72yY/ZpKgoUMrIdRQZdEYLf/clKG9yzyUQi2x7lhBm3E1
+fy83GdyJCLdsdGtyod0DBhBApV/27F4BDEYNbNMYO1Pwkqy0El5KGmhfQolDKkI5F2p9Rbd1Koi
JKg+IURyS5hHPdyzsH2HzvYcQK8w2+wKvDpsXamEQq9JmaIGDX0Uli8oqsHhA4H/yHRVpJUUyvIE
t6P+8JNBtQiysLO07+DchPv+LaT+pCJvYfGCEd2h3w0Zpq9wAjUP5NdRkBxuHmgvVzyOE7h4uymV
JukFfO2rY2rAwHkEyqFZu9Hu/lbdz18HTr6Qw6RhYsblek7JAlT/D8fR67Si1PYLEL4ijQD7L2h+
vrO6+jHPtaIuGAuNL+b4zvIQ8+97Y8dffWH97tT1tsUCVkRLTP/QE1JI7oXmd7lArVQAMXaAgkt9
ux1Uw39DJufDVZIH+nTyeusszIHRFXcg5XlYDgOcAB58xR9ooT8VZb6TNSF8pbU9miplldo7ak6l
oL9mxvdrRmIuwPWTXCDCgxihdPVqfAqJY1e+fWP1XraczUituiTFW9t9q/nz7SugApVI/392JlxY
fnaoKg0y4iDTDFgbo+ueYCEVItrEX2n7/jfJMt3ckWlr2X9z77wmU1a4omV9z2emceBJtIYu1n0E
A25gRCJaaWcRrBDp8T78Tmpqx3FsWB22JaGmkuFHHvA0+5y+j5Fyz5EUfqr5zZzlAujCDWvEmG8K
cy+gZvdoGJ458WSGZaBSA4f7MW+BdcSv+UMc2yy++NtP1ykuXZdfFwflcR5k/GczLluSTbJWVawL
CqyM7j7WSLQIpeR5t5UZ+gPZdUGARAgFhZC9RqjS1+Ru+SpzjNQdyhmHOiW6BM8fFqkqsKKZsK1h
XapHiE7/XY0EPmCHh7bZti983zNuYNuDi4LKB9lIzF6Xlugagb+JQgDHRu6w25jIQuGDHDNeTqf+
4TJxzjTpo/ye+jIHjCiBMaYfuc643ZocMdf74yJzqD1/fZVmX9TiYN8y4ROuy/9baIhOK37LfGBb
rB+678Yigm7ZML4zweD+Q3y0C4Wq6xD0KCuYzlJkiU/cF2K0UKBjVeUoMZJ0yKmOrt702idmUwHQ
T7FGswBVWmuGW89ChqyOJUZTTRU4wFKsIRaxuPb3a0XC5PpdnY7TQX0zV3xmQV41IYZbGdaKmfYj
JPykhzHamtTqtfh9BvTJnMutGdBEXIWxM21kYIX5Y/zAAYdsAJLjocY3OXYgsE11/1KiCPYaveID
Qd3TIHxM7OIthNdahbuuUU21N6hf7pnvYSdD9ZlMOaeBAu9ZLQegdlDfl3s8dBXSQgR3JReyBJRW
ySedoBG6Qt0p7AeT7czYVACnm0Ti8V9QgSWQIAOb3oMCg+BrgqCXvldsyV+DtGHLiGY3uWw+uhcj
vAbNldzSE6j7ZPXvJyj6Dtx/QXbH2aVDRcUNyorgIuXzJ/PdgFZSMo+j+W2HP/QAeCc8JlsYHU00
DKxocu39n1UDXAJS9GVCdGH/Ui4q26b4Y1Q+q4b63sifx8nC6BvWP5TwpffI69sjvxCWLMwX2FQi
kK+LUXzxq1Oikylw7DsU1yJQmQrUDhj+bC1muFvzRda4brKJ5SX6VCVtXlFKCBZVjIospRZ2eeTv
v67WKyZKGCfJ8SKoCRKmrzYZzbBFWh+dhJIVKIRYoL5003A26f65RgT1nx5HNQDE/9H4hxX07DgQ
mSRhatQhguXMs24YVmso3pKXjTyK4TIhp6HxL1qQIY/O1RgWfwKrwA3j40jjK7/TzIqNqo5GhZuR
nHOE1hmxewI3/vMoU3rJSqW2tCq+D9Oc/6shpOhlnNl7liOflx9eZ3DIQT6RJVzCpNmBtF/kvOl9
8mNd68KVOod33kl6VMsF8sJ7Ny7DH7pYaolezPtKOv4Rqu0IC3cD/jlH6uSI5C6ynbRHJWwwiLFf
+6xC08zZrCHjoIFkoDlA1uv1yg9Q1SsjblQL3XonCkSsFAmqnK7wmsWyNWvpRKF4WSz/2doDfBTk
PU54Lq30HodWaCH6fzqFeREUo8kutmqYjBFwA6OlY4CrHaf/U3xsM88xrnpu+DMic66HjEsm+BKx
eGsbDTYPrMF92DcUngCNRbEQuNJccwNKp0vkCqrEL5KCgreETCkx9tML7n+ZildNBoiSqEVVxsN4
Yw2ckNK+NKHB5UmIQcTH/x/wgsbIDiPyIM/aZ9MOAEIi7cT2RaWMLndRT8k+84KPymzfdt9A3Mn+
4BptLuXqVt9cp7cHTjs4bTFMidmY1XXuZtATnIxkgAkBV4JYxYXap9fpP5J7JGAl0dWQCSuzBg/z
srpJH4sji0FrbRN+vsaHWaWkUL6WkTqizQF98L7cAhFPH7DbjMUdojJRcLhfozmSvdykKRVrauyN
vPFZieNE5gOgO2NiTd/Y5LQLecLw7iJfMJFF0w1nhm4pGLCzhsmFZRfn4nRroDDfi/DzkRfV9FCs
vUuHMf5OChs7+EK83UyyfFvpv7M4KJe64pSAgDsUV66PvuoaBck51c0bd/vhs/rT2XZxm8hI2NNV
LbgQznl3Hltb3hmzDE+dz2TTWisjPIHPxDrTBV4xckbaEVfnzssMgbYISZmO2c4qiwInIfOTO7xH
0sU8J3QmClDzKZftlKSWUXADPlS1JoZskKSwuBS3zseA55Fs6gYZvZNGsWX6ARlNPw8YgMoYJhgZ
Y+amoulWElpJXkTBeOvIhr3rbV9V3tb7LWB/6ywrrXMVAAQBeNraGKZiRTNFtAOOYzaFbqLnCK7z
PpEwOT9hHYGXXuOnB4LDHvkQUDByw3R+If0G4m0glh6muqJe285tkunKDU0VKYOMOxD9av85zG7e
pWQ7sZ1LOR0zx3P05r0Fh69i/kc1JuEeXAfW18CqS50rpdjTH8pfii/omVv7fiTi01sdP8M6PkcD
x7Eo1Srw6guQckCPidD3kdqMf9rlRAlvd+FeMGCfRxLktBxtXsm61urFk/W99BmQqd/bEBXOCCdq
OOUv8eH9DU0xwBHLvsWsSXuOuncdQynyuzsulLL0yRsDmKukh5+fcAz+GNukdkRmWQlIDNa+QfX8
AACIqfeyszCs/GkepvvMh/HmP8Hi0pdiTEEXs+dc+kT+J0XgRaRx1moSHiZ2cgdS6VY0PklsAE+V
4Z9Rn2rvYZcbnQdhKZgIYcJDkKWtwx48k4GCzneY26xx9YZ/k47UqukkQvm6CYwNxS4qSNhVvkR1
QDZophpqYvPlZqvDpO4cBVqvbOccLfkEcJwJxfzGr6k0z9s3vq8P49T1ju725Z6RMsOQuc5UK7GM
b9s9jCO0wpMDAp1rSiGvaHE8DCghabqaiKPV2/tTbC6/Zlaf1PssyNY5wAl6+DBkMzKxlqrbt5Fn
kFxI0P2x4j5inGEnqfAz7avMsr8NOSLUMihE9bcywmk6goyUwFzamOMX5gwGZPyeRCJJlAHuB7FX
tpEij5fQZsipZa0c338JMdkSfHVTMJt0pGRUPcxXpAFkwQYDeGNIDmMhVdf0Nf+4weztbdG6GgEj
0iAQuGMGLTYqrGv3Cxfl2pgy4U0oJh8HVb7CRO5i8agE7qejOAU7L42f3bnF/YnEwDidd+2lBOw2
jvS0biygfoYEEtsFJDedPhxRY1MjhcuToR6DOtlYm6iAjpaQTsLZKGkZDsP5kSuwJfXyOP3owZsZ
42iNZE9pCXd3LOP3Iawj8RGpXouhF2Z+Alur8CAk9ESqpFCqaCqlKNbriiR7eNP4xfc+IZxrPpLy
Mn3fQdiLwFfIA8HdofL6z941W5uT38pEEC41pMxTN8Que82jjtk4La1wXviJYMqFMGWfB3CtWYsN
HEXb9qQbgRcw69BJYllv6u777JT5mLWWL+Q+9qoIgRyKpcbE2P4su+zh7AAuMd8OL5T47xjXaLgo
3RY5WTi/bMzDdkuE1A+clRFWnp20cSjNUaZhnOuh72M6J05sqbpuSr5ZvFlGVLma2ZCfRv3t63iE
N5rxZAp10wy3ppgP7AQygHdMkPTSDuWLKfeHWWZx0mXmwzeEtkhD2tAyEK6wofuK4P4Nd1lTY+8q
2EhQk5HGKUK7BOLjnVAZoryYNpVTnAMH6P9wZiTmhkZJ1D0Lmi7vY0C2S+pLTowrrsfOnuMZjJsD
5tCcm4L5QpTxEVsPeYY3SQFqBl6z6TR4+pTy5A6b52EdiIfFJcD2eAn6fRblxS4hyqmQrNis8XUT
pJX6sJEbOJKuMRHeqplyrgMu201hfC11VzUNIYI3azsk5Kigrz2823JSeFx+8iDtlB7em08h4I/J
lRpMcifHzEfL0az3XRKU1YIcWD9kywEet7n9v4eBmSnkHkbHrRhKeQ5Z2cxmK673Qxixg/kBv5IW
pDFsYsv90R37bs+KYQfiMNBJrKMg9rbNx0dY8Ac2UYGspb0CXb94IsOOdfdHuDKG1bf4WGQGyxtR
Avcxusac1ohGppiAuhyV1Sq7zmiLDytqNl3Ggr2XtZ9E83M5kR6RmI6fJLhpb8X97OxjR8nrrhVJ
Ock2PRxVsYcLGJaUUTG8590N1acIotYSZL4MOK9hZrCnNcpoBnZbuUWDjlQLr01HS83Tc2kyOdlZ
vUPdc55gWwL82+L/y0CJHhcZCqIrleSwPPmEFBWcxd7Egm/t79DYvhzNQejQhKTYRzWBTQuAeWin
V8zCmAhJ/cNlQhTp2DSzYATKFPN5B/aC7HEbx0Zv9Z8vz6Y9Xzh31vZk2TeXkF5d45AXKxwFrkJa
M0Rw5DUURaSIiJ/HzAkGv9tgUcLIUTex9gpFUKqQ4C2RhLgo+n94+czBy4GaFPnaY0fXo0ij3deT
23Q7g/VCfi+auO1yoI+ny9d414zTND45ByfAfXxrkSvWLJlUMGA/2/SGyZ5VPGzW6+Wa2S43j/AA
UYigEUDKuQUGWDPUkXuv1Y/CGRytkA79DgUt/EkPzo3liXRyx/F0pPHDQsckbA9mKYzpP9OhYe5E
5y2GZDxpjvy1MtubsPmcFQcNOSHS/DfBbu0R7VSXgmotJp82nGC/Rya0aUK8T0wHXatpFWGK+NcQ
8nghiOsyroZhD9cBl3UiFBRkkVl+R8zPSb98pI8URbe8H4Tb07hS9GTi05PVoqV1kwREROqGFWCK
RDhYbx4xo+cXHe54XdgiNygAali67Dlk2UDP6+/UEWldHu18sUsPQecF9AVwZijy6FvSsOIAmjRD
9o13/oN+2gA5lMPkx9Ye74uz01by1i3NLme7NdcjN77I6qIx6Plc6mxyiz9Enw4squIIqktcFY6V
6kzfdQinp7cezljKYIo9IxA4jtL8mEuFPpkX5UPNcHrem4OylvCOlCV8P/awrULrcE3o3tW9hDdM
GVpWNuU7aNqkDjp4lQmqptwJX43FV+51DpnoRRu/IGjDfQfiHMX83Jl0Y9O3VJKel+olGq2L2j2m
i0PV48j/G8YQoyJfQNG2Ri8EQxMrLzf9J6rALJWqNaJYilhyxdsgnRWTBxOjZgQE05pDNfgBChjz
X+j6V6XuJGNrTesyg5ONR+FldW1Zr4/8AZAe2R2eUNoh9sYDIYIcButcO4XW6QJXbjYQcWXu1WGY
B3pXNr3Vxbma9x9h5zUqg7SeV1TruXbh6eyn1NheO40+FhW7gMiSlxNpLn0tWiiaRX3GbER4txgK
bMPyqAoK/e4RID3nTjV3eqEfyLpwQM7RuN6ifrnn7cz39OE/O910c1QMumdlI+QEyQUlz0WZAxEd
o6YdFilvcOt/2t6LmrDzcnFF7cDvLf/H6itHCPdVbGj6HH41QVyb/GdhK7lW+9N/7s8zBk9FcW0p
8sBcGGU2mhIRdmFMx06PhyGuHJjY9WTUM8xN1kjtfOHjjbuYXMY+OAyOrbS7dYwoj/954v7981e+
ssE8BYW+GWVpaoVqTfjoX6vaNZeeb+EftImF7deFTPYxQ/QwfSvJrLxhmdSMWFDRtr8ZHPxRm/tK
NoPIT4HfvB/dpzuFWfYXGnGoSVzJRTb3dWt1cWwVQ2YiEa/NPgMOqOb/0Fqz67Zk9kvo1z92C37E
2sZhzCMndSFvE8xCBD6dfCr4TNR5XBpqSaVBt1fKRcuuMsM0/t/UrIoM4vr2Cl5PtmMl8eLlqh/B
5k5+fQQHWvk9t6IcCq38EwtlL1GQBZfRMPIXwjipY66zpz2/Q2Cv6tWOxhuCc0d4izj9Qkg5/U/L
NK0kbAGwo2jJNm1WXL9mOgU/inhhn+PmEaFh2HZw2BIUrpWIF5I6Pju3ZYyPNBTgd2aGWG+ZteQE
Oa5JLSEf+XB5aUYymHplIvGmGHd+zX4sRp4zbjBahwLR9dlmiPHjSCpRpzbyIVCDonQlgiu/kV3U
wFstgwF/Zd6gOQy9QuarrdF7Efkt8hwcs59DvwN0NIQIshmexRikwnNGaniyk+93eg1dZ8ZDgi9j
hLfipT2LcN0pJl1XwVu/Ly4QYrCvtE49GTwsAKYT4EwLpcerjzQaFeUmVHjFle662JZsZlaZimBX
UD/D+gvN/aVa2K4jzs+ycnHYf2lePXbE8NeoOYG7Iuh2phgFSlaeNX2Vppp1nILEoxi+ILywx/zg
L0Xe9Shglfdq4dxrVyutTyPLiWOI1J3tm+7LDRKdIY31mQn/k3G5jrAaKJW7fU++9kckMlGT+TOq
ucgAn3NIXVESQobM7yCWg4hFC5LchviONAamHN/QTTVLsfrTKyzmsLheHbpHk6eUlSXjBvGYb6B9
3ftUKXNZtNDFX2134YuicOohNPRK3BeU4ooBQEI6W/lRfA8za+KiNOJP18KgplrKggpaWLtHu+F/
A6XtYoa8Tf07+nbQbwcTNtSlXr5zEqjpApgooSKHwhrgqCwwr0QOL/xnUiZRbSBUV0b8LkoiR+ES
wHJ35Z2HWIcouh1EaNJrvvv8Gjj8VaPgnXgrcHoTBJb5nWtpU10zdmk3IUUuMWRhhgW/cLEZQo7B
orY+5HFlIRpiIC83jWPyKs/dbTrFqxEEbIUMn/VBmGANpQlvrDn6HKTz2X0IiTZK0QGphxrMZ5gA
PGQClg62l+Cg5QK6hI5I2fAvOawS3U0myJUD2K7nji5nzsikqmYH/UDMo314WOUEmfBRwfDy006A
RSQhUH9GWztgAEFknRlTJrNkOtCnrhIbQaDWro8fjZvc2F2aSBdt63lBZe6tllwXdNci02cJaQ1V
OVw+Sei1x5KaIrJrEdKh9ydRbxz99UmC2XEdaSdIIo3IqDtpbm5UGKXkjo9z/p4v0wXAHMJAFbrZ
vR6pR79Rtzg/H0EqY8fGXNe59cP9q6r5e5faf3f5Ky9jVLlU726s3pQTzECmJ3PDXdTDf32/oYK1
6m8BwJSznnzXLpn9SnC/Bn0vIUuKtdwYuVL3tec+Yq23wvWOojsnNDfPVdUKEcOLCQIx8gA7bawt
rqfZ2D3YH6YsNsOEpgO0DarcWk8eMYvIb0d8562/waKfVk/qi16rXx2pWdWfhEG2Eb3aIxvyDChD
u0LiaU+TQl+Wdl6GuiUsPoAjPGfYCesWxWWsDIT1dII4fKErhvAVX/cyGJo4qFkxCLB1mACBse0c
vpQctXP4QRAGs1UkXae14HfqHJFxrrNWO2y/lRP6dpPOpfJja0mE/E3tM0fWlKzb9yIFqK8rVstI
tAqRoRrlbm94g/Je6zRjMpYj43qDrhHwRD31jXokIuTJEJezm2jehqztdm0XOEArFOFUfejjFy3K
hIR5NJIKs5qBTfrMypsYYNVjelyB5yCL14VKZkHSct4sAlAcKcDUZVDojQT19bqHuO1ycwC27vbS
pXf3Tz5Zv78i7bYKdFooRrc7p7yf+7Kdy/r0Q1LgaoDzjgJDVo0Ifhcnmom8+aJeBqAIEXY5zFry
UvZIKz+ApC9JU3VMFzz22Kp2lmOcNLhfgmrbRQGBWqLh0WVszceroVdTGV5xn9udIaW2dNkMAmnc
Nb5Tz7yuaaytkLsPxr3Wpnbo1KUI9RqCVk7N3GoDR1f1KVrihRc5+VdpARDdUUaiRx/1FZvIzPgr
IjYGh6+Af/EudJQ7FgOfZrR/dyS6O1zAHJ8VmhYuuYa414E4+aPKMqQhJLeDGgK0Mb151wbcLaPg
Na0m6XvbCT28iw9+dF85/+mqi3dbzWsuumxDiby5Q1kJ0WZX3tT8tLoulu6LrjZmX/aLflF95Ml3
Zz4viwCah5zeyIOPIaq00YbKIilWQZ1a+gSHn57+MVa7484ehAdCHKU88gf8+KQGQnb29wQG0INi
Q6LW7vFleVoUUxIv8EA+D0rP8nQzubtH17qCa5H77zah3JjJr45CB9p5NjaAoZJjUae5PY1uXCu+
w3GRbPpy5jkhr6czKhTmMNzMzm0viP1s60zC9Y6Zv4ji1rxw8tl8W8CaK3N55BOognGEtE8gDZiB
vVdT8OKP1e0rJUjHYVm+WvjNgj1QEnF+PecTN9RysHujd/0QpmyB5Zcug2nIBQyW1/x+SuQ+w3WV
67vjb48nA9skAL89cSjGwlkLGNq5zoS+rksUCsAWu9qaheCiQ8iAm2hvu0lIDkw85jkoIIA0CHsZ
j4BxQKcGb1hmQnYYO+P/MSTzEBYzf8CSjA2/oNsmdWK5JN53b7aN/PE0hmubN9qgHtX4+zYcxLud
zLcXIJjIbSxfuOuj63oztEb5iBJ0W11/iAghQMfQy2RmaOYyegCNx80Ra0+JjcwW++wR6CS9zPCU
yqA0i6sGR79X5qzTh/1FD3i8bkh5HtAGQUrEx5E4402xOtn/edXwe76d5UgoIiQPx2sdfJvBSCDF
flSr3wcKlVkaweW3WRUKFAuOiIMU2CBgAMN6FoaaNbUFIyJCx4+cQXmFhyxnV/7H1AI7b23f5ZZb
vjkskca/GZaQzOZsRQC4X6UXTJaHGDpV3/19phZ470IgdVivC6oLHKSW2Nm4KZtLF854US0SHpn9
ndyOJCEF1i2+ixJroKUtD9swSuf+eg4rCn2K4yRi2XGr/6lNrQwqkR3x4T2U7rSkdNDDcrRryPHo
HjvMyVsYNV9OHDh0c3lVVkdFMwx5Z6qnIhMf8aRG4QJfn4csisFN8r0DUzGrSz5kLvO4TegqmglF
A2TuHk3AHrN0U7tELzfVwOhLZv6rJcrckhkzYqwxlTg+TjyWcEZzxAXCdM8FcsliiStwtWJFJMyl
5/EbPlP8DH1JMLdoT/Ni3NPpUIBgR13LQ0mecUVSQmqp0tKgIfA1+sXP4COMjJVCA/eKkF8WhgF8
ObdFHtcV0l+CerarE9N9b44rMIkHggKkT8+ir9YLuLqyamUgdcX9ep4ZiY76W/p7vFSKhTOvTEon
Hv5JjQVv3y/IHii7WIpivUC83RW11aPgstbcRF3AfkTq8NRuYhO5xgvI7m8dqK5+ySR9MbxLXHhW
+YSvLcU8SRuG5+uIhpGuxf30Jav1EbfcJgmb2qgbS4dyLxXZi23Bm8mtcxlnMcSt32/35DqBHo4y
lnBvIaRp//N3Z/kH3mGTzHD1qh5lMWEQcAnqBdLHA6BM3BDu9S0cFvsUTUjJgvxrt8csZmR8+OdR
MaxKSYsoTq/NOlqc+RcAbw7J/XXPZ6TYb0acizLml/JiovTlFDds8b+7gegpjqaLt9lMkFcK5k1C
y08kzX8iUd9lbVyerniW3QLAIN5jGZRhQb7ZM8QhDYTamxnBXUiAQfrOCuuFPStn6VZMXzJ+D8MQ
qAbi71IGjK4+4WhKx61mTSdOtIZnUI3gDSt78uVWccxRdNXrvS78pXzyAnS7rsK/8CL3N1sutN/Z
ub/IiFqE6HfIb4hntY4cXec/w3Cn4/tmFnqK+HzwcURAbNH1tswnX7hC9tMG3VGDg+M/MW5+i42g
bRoCntRnZN3e9JgDq5umkKw7xudqxZcdNIDutL1ZFAFJmqoXty4NDHXYoMuyA9/q3T78CiSekw3J
B9HtFyErfCyOjWPmUVNDWqTphfPLyjNTqC2lDaBzMAlJZ/vvmZ4n9J2d7atMvDlgHYK39IEHkwiO
WWokJEVCRrX+LYipuaxk1zmmn8Fx3846vVpH3DprBxNc5XLcBA7dByYdMfIXLGAQUhbRp0pao0WS
i2li9TMxfWfVPTpsqrcjc/FzTDzMpYkERP6Ew53ktkuj0XJYHZedLKAsmGC69tVUFdD83gjqSpi7
ZxkAOmq6rvl5M3tODWWxPI8grN0t/SbjDykABfnVrNDkntBuMIeNDbaGT2U9azTk0pMgYSLpu+7V
PmxzYA0pL/zc08Wob+g6HTR1QmLpI62BUUv00nguh0yPIbrGcGpSKCz+tNE7OlgCa8lGlmODnHND
TDJKStGXATff7H8WezP2IkTSuLjnTDAeVLqYqlsEginkUU8bja71MBMWazEUlrlGUGxgm0oknjD5
SQ0xcCNB3tD1Bbpaa8/Upos56zu7qMhnLFkL1D5mFypQgQdB0JHn5reu38cJBup3Chw07T70hsaP
m3X39osio1uojCYiGqaGF2giNZHToOSXVzOzYalCDZuZXmjQipI+uCcpDOWnyRG9Zq6PSYT2PiJF
bewBY/9P7VJAYVS3LTxwsv2EU36bAQ+NtfwdxygxSE0m/fzqK7t04xdne74duJMTP23uyMt6TMbb
uIpg6hmG5I/17R3VV2ZC0+TOHhJIES1i6PHF8katf1rmydsHF9cDA0WWJou68mcVztpP4fItx6CX
O+DoU37rYW1KYStVRjb7I85XvFNV2Riv3g+dvQDNB+uLVzqHdL2VgZfF9/7J7ih7TSe933xuPzB4
h33iU18t+yBffqNPmxnqyCEh2MK95k9qG/qskbTZM/vz9uBrYv01WuTHRc5mQMR1HKatYL7+JImC
ansGhqQ5ZKSkXYnFiIZnZwr+jFTaxu0j/2ya2wbVmORVyovMIFk/mLlaW8WGWXpy+nYwUAI4xQ9O
6hYO2jmwXU9XlrxP0xrU+r4s+S2YwJLH52ZoZfWUmBDriRs0sXsIb0dgaKKNYhjmh22EeUbHhZY9
Zclj1wg57YirmSJVGxfQRtG2LNU5YkP9klRKuPZRnLMRXAv+7VITM94KUCo4lm6TKm/fcbElgc/y
vsn27KXMNXGgJv03vYmQ0qOHHzrjEHljzelAb0fPGbUR1xe0wylp1SFvilO1HGZ9WITykI9YPLdS
OSTDdQmu0L3xOzP2Ft9STkM+pfTrUJ7FSM6cc0t4icMarVSKhmiBxQIjpqlx9eAXhy62AqUek0H9
IdZOddkvlTddpHboZDP7xaXPnAZilxy8Xq62iTS1dMQQGukrxoiex5J9hnHmZ1XsYjv/e+gdd7f+
dTzJDQZD1Bp9xwGNNILKzquHxu11oJiIEt++nVb/g/4xTIgyHMpmYuolaQikMCBFWyGJol6VXZrC
zloPeVEyWUxaQ2sTG9l1M/GgPN1+N/aibodu1ViR+lWgaXr+5ukO9srh/9dfh95sY/NOWbz0DsKr
t/HtmwN5DqvsbzGgeukrV390L9flULfItwKXUs+4y9TDKmTKtW1OCm/Zn5pNZSlxYWw8aKNNYZVd
wmd7ll8bcFJrhiG4tb5gKgbBQNSWwnq0PguKoEy83JsK0ipFZ5G/O/MKORuYicZZLAGr+Y+VW5BZ
4brBCA/3tHxWj6vlFVgsKRp9X+YG5M8Eyi3nmSo+xTfbf1mSZiGvQPpvvV0VkdV2yko0CJsU1ljj
6tHGyt6mDVgMJlcwq24v1D9l9+L/TzNiMD1yIkzHxdhnXzNzgK7q+NP7SrCjoPlgrC+dcg7btr3p
XSBfmHk+uayiwaJ3bcapGpeDPtp+xDdcVW0BP8cT/o/8lZPDtb7LZtGr0lBS50KQMmU2qAoANvG7
DP9xCC6pvD2msHgu0TOP8zeejX3BNRkVaPKjIjLOgfzbSItrW2DSXhMRJgbvG33u+PsaZSQK2q2A
q9HBX8rDGWR/ipjtvr2gCj6wu/k6YDFmhBVYBWNxM2tVEX2BMUQI1k2i++84KCAeGM0g7qvCZ3jr
hA+1uLcW7RfXv7tmy9zJEC4x0nw0i7JthKcCSjCfXRzxkjUDUKYmWrCeROR4u8IxGDXtfoXHn6vU
gElwX5RraDbV4qV2OvSIQsiGtYZnPksEMzhgmEwL/N35c7vYHq+EcXje/mdUrr4LtwQWfmvgceZM
LntfZ+SV191V4yic0a0PIzbU0YjvYstpjpvDCocHG9ddATk+sI2kwMbiURSqdx9Xke2Uz0bJRafV
hvepp7T1c4g+bsEXySOWhV508RTfcyT+GObFVtThQs/9TksuGqbpCdzI1pKfnje/q9sZHepHbqSN
1JeWwhXS6IG5t9Ic/oDoepp4DttMtWZwePZ/Hreng/a/YHx2bq7L+wV1iaLYF27UMIp/eYBV6UWj
fnDBwdO12rMZyZz+GrbV7hFps/WdVWYzM4MSylQ8OmgBkigYfgUIEHcOMuz0XNIHlOBSPh7aleSI
s/bJIbtVkQtMkNpvpPvNB0FGa3rpa3JpLH4neDDpORIaJu8PTSmQO6weVdaL5vrXVltKCW0hmlhh
X6bvO2gyn+0oZm4GCrg54MzK5sBrT8KpdngKRjFOAvCzK0rqR32VI0BEW1MCaINhI6XxnBlD0/aB
zI5dp4Azputw7dWNfLxlWDwvwZlgyESBw0okaclhx47777E0Z6bdCuT6plCcNw54XWjOHHrnPA8f
nwa1O1DGGZ2sHKELrZX/JoNd30B7u4oYmSmVRJktZ7llrBHbqGg/qhzVjF/W2i05IaINU2Q8E/RM
LSzeWmCUI9AC8GksBOHBbt24X21dCqCpldLT7uvJwvASZocnHyuMx9ceQaEHwjBU4ZbIThvOgFuM
JzoO3wiSkYYrlc9qZsbZ3++euYhvM8g7luSXLRFt3xAd2IdiRPyACiCTBQY8f4tZ9Kg7Y42t0u6s
PVq9Vx0K2XJT9WkdjqWhtkikGDbfALmQZIW+TDEtLk8j/qaShBrEWVlD/J+y8VJkpt0WT1jwZwNi
BIA+MuKrEbeGhv+S49/n1jBwUc+7MXaVG6PvtFQdWJ/8fKH7ksBF6x2h0EN3BSC3T00wQ7Jy8bXg
zeVcMWQ0LybYYcKDr4Xtm+9uK/SAvT7lBVJgkYfzSW93q8zcIdScap7WAq8i8nXkMc9YaGnKKVgG
rOsKuUvuxgJMjdrKvx8w2liZOsj1C00mmFQmOFlawjYfcDrE0xuGGOMOmhGAWBCH2ChUt8J/72LG
oerZhA6bIR644srKLwrrn6zhUtV9dr5KU37ETvnbN1qOFXyZvKSmDlJGG+MYZ02uxJdmMMmXHCQU
Jrk4ELQgH+oy4b/hbMSzH7uO+64H1/fuY1xGkLOLnybhF1HQHjEqPbtxAU5kGvHRVcQt828O7B8g
sGtIz/S4bfPnGQN3I9A9CY41AoHvcFLGK5nWWYD4BZrK5KXemvm5ERjtmsL6pstJK1qunMzKAXfo
DfCGtR/3BLwryIIc425OPpGm/BOOHnJogrh2gGqN+Cv3ChT31SRFxfsSC0xJfbY8mXyIuCgr/WFK
e7ljhcJVMzc086ldHZ6yfus2o1nbl8x/l8jJpHh/Dtu4RYYmFgXFk//9WfaP2PproDhX0tMSsytC
IhoH89w161FYkhJHKl81Q9vs1kjfevbmP4V6HZFeLyETZoVzjRiq1ojhJqetUkILhKAUmjNTjLaP
jWionVjsGS4yCn6tq+rdvzDK+UkRTqAdFob9sPs7QbF0zj9ipM6dfrIsPp92kHjiofpWNLnkinjA
uFnV3Ts7itWIPOcXcw72w7+v020r0vJU4tphrWYVIy/K4T+o6Nnkf/LGf6drzx483iw+m5AQlq8G
PPxBeewAsa0NCmzn4lZBtHWm46hqrMNSPQX7zXiox+fkdysRrnOcQRHvXYnJZUM3e9L8emGEsvcW
8RdnBh4tAJBzbFlqzqrGNlFC1AlgW8SW5EcGvYp6j+rHlolhjVWnA6R3h5hCNBDd49QdRK4aPveQ
PxAcODukApkE2bMIGGYmYKHeFxlXQET8RYP6+COP+3yHWcYNpa3Z3xEYtOY8j6ZDXUoR45J0j/l+
GoFPjrtA0ILW2dI1DCV+oMg1xzdH+3smcU8iREJU22svQj4EYg4WExNUYVzZjVRjy/DaO+3Rl9ZD
YxyrmWdh5cRlbg3LgouGEc4F2ioFAYzS1zA3SJKyjHv5FtI/ebhKMUFXrV0a4lhNmnCRltH/5F2Q
HeDUMaEYZu+ls67p4AJOWbEQwC6bK5x88scpKlPdeWecHwZtH5PMEJi+8Owczu5noD8bSCLmT10U
Ee1rLKohkSYOImPyhc9jP68j2KDdMy1kZFIpiOkF0fWgjPE/ogOuXD2saTE3SafABGxXSliwZKjH
GRe4+SdIlcaQZa+D4Q2tPtRERZGZLBItfy8qyBIMRcbgJH11I8rEOa8Snb0AVnk4fb4uVSR3THkV
V4ZI6SOmzCiZ+/1voYLGAejtHAfii+GVt41/6GojwGoisv1WIuQwLSsYfCsevhqLZka/JBd92Mod
pTK4mfn6zX4tVIKN2t1FrMjVHv1gP3k4/6lGW5hKXGh6rfHPvnY/MpmlTJd0bWYy6mxQFl9uutes
QmvNWC4+CiT/LDsPVN1rm2rbtJtx621TbDT1FpyMawxjh4xXQELjEXGB6SkUV6nizPmGBvlITeVU
4fB/oKSM5TVCUSVCUf6FIXFrY6lGVP6BqeyMIigefOwVEiNzMF46u/Dd5Ycd4NtUrcDMkwKHZjh4
R6lmsqNNutLLeDbwus4JFvA47wzhpd6XMbHcR0e9KF2TuDlpbgRE7CbMmBrsHSsGVjetgMX6p2XR
KUU2IGTGe3sVIN2J6S+rvQo5918cbkH0dFbciZWKF2nf04GTLulDSpKmz/SzNwCq4bg0VpxmjCPV
/jXgo3Mlum6SXAF0gZuv8tQKa5AS9S8waZjLYhMRK+TC2tnKpxqMgQ/FXGSi5s32xRWla06jU6BL
Tb+GAhjx0wm5DljguogbShr2N5fz+bS7GjuWzezZZF5jol+h9zt22wpNibT6Y7eO4sTPQZr0oN7p
7m+IU0e6+HfYr4zYDI3L+XaSIiEK190tHwI60E2hsQBRiw280dfYzMhbPTkDTvw1uLzQR950ezLs
UZQ4GZ9aOT58y9vHvZ+Fnt5gtB30chnNDOQyrDHaWJ6fUCX7xYwYDjBc8Nh0n2+IxBFXCLgPwXS2
lphsqN+o2kGdX1Gq8QQSvN8cEYiv1kSUooNUfLrs8OK2v6d9y0cayDA/T9S9ydkCifoq+qf/NArE
xF/SsetL57IuP1849d7H6T521pxM9heH/W116NQxUCduan+5LXTNo8GAvDfUlcQtWY4fF3zpqCFn
m9wKH0oaxursyzgpcsepZsjPOF/vKMDLN4scVdHqQL3KcV1E/NH/30PGovTr/sfIONBZbFRnAMSs
Dzfho118ncTkWXiW0Bv3j6omXo0XS0K/8nnU5vAChYAInQhdjTT4IEIS55SK9DYeOgU5Ur/iQclI
HeejSrilzjUgzGedVcZhkEutNXN/AtfiJyZVBTbwF3la4c4oDqZ4WBSVqlyvSvhurJ4uV03BP4W6
FNHNraL+92A8jl1p2XWTvgvXeHPHh6zwHtej9gCkVdQAZ3NRs0LwzZ0hnLjIUpMuLgWxJPCQbtKD
xMtT2dKTk+Hzv8K37XV0sqQtzsffG2QfCGrSjAd6S4eeHOGzNOg1FSE4URG+sqMSE7bwRU/jFjh8
W6juASAlZAbW//wXJhbHz3fJ89J/XRGTVsfvZM1H/jfyuKjcHkjr9z3xNUJGGajeWYPwvpq257A+
QT5Fl776TWT5DzVQEbXLvVtyNsI0l3Vff3PnSM6L48rxC1JmTyA334+QGt2hpXbgegLtCQgFfvRQ
wKkYB/zUStxkO4rD5goTnIfWAAodt1zVRetlEb1LzbZkAxplg68xIt5AXfXVVyzkLlHEAAvkat91
V6ljHSrx84MDirgB3wUTLpyn25PrzyZnVWLAPeDAPSFwtPv3ebLueFdRJ+TZomwvf5G1jZnxbAOR
Jrue3wS0vw/UuroaP+r0pycSsKxXW9g4QZ1W9lmVrVgULtTvCB8NrbX+hC9APayWQ/tFMw7EZuI3
wnJ9iJ4ctFWuUwHsQb/MbCrJ0k0WuyOlGCMH+2Yio5sdVAys1eG08TEDeC9GjPbLpbe7zGa8Dssz
t2MKMEwa4g5yb04/VPu4F6YPTP0K8/6HoWvVu33dUgYlk1UUd7wnaSPSy6rIsDoavGaHkDhRiAGE
ytgDCZbP0C5qyUYshlP643uEuwOMrP1bZ47gNJmsVqBdUiX76DANvC5Uk6AedJQ4WxTPyBctMlbP
aqeQ04pue2TtYuqQH2wqOUmrSC9LwjkwjQJ1vN00HfTlCThyrE8dkevPALnRUnj9l2ynfoLaQ1h8
m6GqeCQd4tRa3H/X87Z3HzdRJekNBC4FUdD36R80QFchKo72l8m3oj+ebaASQnwhBZ2gyK1eft4m
COqZWopHZD7ONU4w/uqnWSn60IeoDNUCnNvBtWehYNeC7PeaQRwbi1xgYwJKphcv74DOeSEYRA+z
TY86JAueY1/1BqkBa5SVEUg64y+tX2QTcokGerz8ZR2//zE6BjsKvJy6Fe82MahAztlpbY2Gf9Uv
/m60IkFaPqg3axhcG3n6TNBruKDo5YBgP1thIWTSj/pkMSVfmJ14csjOQwxUoiU7FRIojMvvczpd
GdmwfN9zlTXew5a7cIVXsO/LSgJB7G0t6z5i/z4oOAEYXROTM6ypgVQdMcIjUB1MKjATdtxkq0SS
NHR6zQnbsqdjPDOwrnpwZj7xzVL3tg7ouew1EZkaksKWhbE7Og6sGyXmu/dhELSCWpbl7nulasvI
ewcqW8tKs2zkO/HcG03O5j0sqytkcpI7kW0/7c/Uny+5eicLfo0DwyTxUUeo1cukM1p1UTwTdCQX
Qlkiln+/R8hQk57r5k8xWh6vOZbV4omHywBSRYYsgrq/vQgStUX547cDlAK7RNpiXEFr1ecTH5VT
bokhhxpSVa31QhZ+bSSjUt+MfRHEqlZgQrufnHT22fo9wil9NuN9GllXv6DShQ6+z1XSWebJ2iNK
lSezVBtQXrIBi0E46Kd+BaNCzq1885IUIQLpPCakcreRNclBsSif73iMsMWekHcmKfq4AzmvX32J
67h5yyTE9fAF3MDbBTnVO91X4Hpoa+E+e1GbSX7kCZBYvmcLaVpYYLguZtlM/2vssyHkH5vIyK33
AjD2+ANx5juDald+Bnb/O8aUqlCJ55yA16smWTWr3L3p4jLOn3ehBkeba2c6kAQ2V8NCa1+WpnAp
Q9u/bpii2a0DZN07EaJ9w8Dr8TxhFQ1nQBe/nlL2NoL7pC3PCKVX9wKd37hwZQh2XJ74UElyx1zU
P86IZ73OjuFkqt+mDwZWefN9MPOOq1fVMhQtAGrcXZ4+UMyBCHRst7KB0KloVj2AgTj2NaE+hBf4
BZH2I6N3IgcmlVNRO3oi5w/+Vew89FOFSlo+4Ed4nbN3TpnWuzvpaTqE/y3MBJoVWynaVbyIDY1q
2JqRHyW7e7QGWrCfuabxSPsS46JdMiOw0lGJY35Z0EvGxZBG0vsTs1v6uQNshWlbtfFzm/tJosIZ
oYDvIhS1NOnUtKgu7RUShcSOkEWQAc7hMo8Resd1smD6QjwoUflPP/nU6O7yYOlI85EYalcyoEjy
2KrmheiQ+hK3hCo2QKrW1A8+D2nxl5/kIAfbRpecRrD9rA+/bly/lrUZnBtEHWXHbxOEBuq1tE/O
LPzaykdbSoNt0yhoY0TJHnafOQCe7BD6ZwbplCnJ4/WFd8voborKhArHzy3OIzomTxOqsM7CBTMR
uM76KHLGflN94YrENaSD7XWmfIG3dB7uHVeWcR2kbnM2miTjIG3TsHH3z9sy3067LWpq+3GoTEJx
skOVbIT4REPrpI6uMqll+kZRdV+ZM0b6G4zjmp2H8/lh328RQt5Z9n1w5kr+EcONPkJXJ9hSFCqn
2LYtcrt6/VZFWHyoIsXJa5EuEBQFY3K7WJI/1W7PfUTUT54IC8Wsfk3rKmH/bDzJshZRF3KZchjL
RPbZcvy3K9VE8wAxc7AuyW8tfX6gz/poggssTr0nkkfuy/413Mm3gjQ0CEZZrdHHRa9/TtpZuMKU
uMgJ3mr8J+gsK1ThH3FG5fgg61XbcmjuPzU5CSZms0q7vYdu88YLP+Th33wVU/eH7J9mYg/CTw9e
4lfhvnWZYiPgpR5UyM4Ix9kFgFmvAV8D1+08u6ZUNQEta5IXXWYUaDGzVtuiacYtq6fyHNe6c2/u
Dd4fDGM1SarzpzQT8bXHTQiiexE4aamw0dW1sVLkNGnppAfDMaiZuwOX5rywMBC0afNtOXz488im
iLWtyV82ZGpZU/RA6PMNN04z02T7bMez8NLcM96/2U5gv7DOmE3Q5+cvKxrk1W1tB35Q2jV40AEH
+JH47F2Trvgd6AiynOyoHqd4JgfqTZ49PyrFhy3u21FjPOf0VG2zYCCrDLO5f74gBC/wv+8KAgl7
dMQ9MqB9Y4/Y+I3G0q96RD80zOALbSRiXk21fedKKcDAOJ7pbNdM4+ll7lGo42AOuW3KTkvYys5E
eTu6QrSDdT+Q7xP6L2C3WDUUn+Tx3wqEpHec5VdIiaMhtoPa3R1kXVEYxQzGokT5Z88BWYqCyfBX
SaElEbGj4ZxIy1j4sGTmCi/UXxTwn4skEcBmfSnSB2QbpSh6z5TY+cainqhPFrMxBOkE4YkPclY+
oKY9c7RHaRDi5xDszDbxFjzgB/yk3K81A+BNG6kWDFy6Qidm7eukgjwU8ZrYj8ZAcWS0dHX2slZG
zP1guiDl+PkjFe0sflu0a3qNDF/OpSMm7kyMofP58BcOhpx7eoYyXBnjRlGeWy6gBgW+iR3GThyV
MmnV6N70uCrBLX3fJR4kv581uyTe8s+6cHCCl1vTzAgKyLV02CcMelcohdaPBNCXzo8GYHjQQ8+l
RHV/gWfg5VV9fBJ2q64SKTULSnWS46U72R73uHNNsrFvx4wd44nDqP5sN6q+IYhm6olZyNgvyEKa
hQ2uXedzSctgZZvNgLTbZ9sZwjQgq2yn0t0johsZJLJr50Lr7NOd1Yu8JjM0q7aeSAjuYl+M9ZIY
wYCb1wv3qTX144wtemLfKEpLJUYRzCNRoIOromC8U9HvrIkOdr3cIZed+iB+Oz4jQeCROX10nCik
LGfOQwsuZDqVVMTO0AQ3CWrtmjKHGhpDy8TNNODyHS5r/DGkCwjKw3ycREVsYokEkAeVnCK0+VKm
PrmdJkP2YeOZiBtrg3O85vzYSLtSbX6saKvxbdKge4TpQhWEPkRaJ0TPsKfSzhIKqLf1jNAT14Bl
G8ueIexTJZtcqMivqITSys6J8M3IhaC7hJi21XqgJxeQNHf+HyKtawGa4aI+ygB43dw0BnqFUBt3
A7pH6PzQph3MQ9WjdMjaPpWIBS1qTns86fZq82p8NU1J9fcAhjcI85bNCGWIw46xKD7FwDjEdVT1
Fm8yUjHjvGkm0pe8StPO0Ed3NVn7ZH0C+RLy1MjCjp+mKwqjGfT6BcF5CKm7hRchPDuEs3CNmKI3
yOaXClWB+mVIn/bbwpNrUzEkakOxh7yrJ00oHubYIm3ojYUUEa8sa4AAHSuj8dtDA07mC1N1gIBd
whramjibRWm3tGDwgF+RrCz9W6CZke/IpUJ6DS37Uvy5qALLjhmiB/Tgjvn3DnNT0L7kUGBFxllw
WTFlNsQlCVGxg6+q3zlVoM8Z7ZdiAbEhW44EmMY4Kw75812vZxu4MnPLie48jAEsNE00P9azdOtN
Jj6JzGuV2510K0U25k9Yp35M7VXhB12NRN9dg0ydDZkn2rhwVKJnNHOrrE4iX9Y7rYoenn2ZXAfJ
lwe3i0R67+l6IC8lLNdejb8StfLoKAR/SXKn1fLnlzeFWsGnUck4H3tFcso4ca2klh7IskpUg3nx
w1lBOpmlcIEHiCyCAd1xGGTcnO6+tdXW59sLy2/eCYyXW3Izc7coF16w7Ho9BXHKBDfnqHvZU6JT
Bi7iChxDYSUA0f1b4b0W21FzvlfhAzlRWM09G8zJ8s3teRmIzubk9yU2s8bNfdYiq3nl/YEGkkBf
W2Ycx8QF1y9Enta+gGza4hmDYbP8e2da18wcrj+3YDjvbblGT8smnCF6G/Z+/5AlMoVJg4wSks9D
gtGqamfUEbJ+vAnLPviccwzNGDFDuBhXY0XFq+QF5I3J+l2QaMjqHa/Ov8l55knhzFl6W8mSMy5D
D7r504TL/+9md6H+7WxgBkgmpw5QLOqZ8vV3FVRfOUkq9+UpU6xyMQJ0AbmuGO9eQ+usfNOAMaho
/cMNkHpUS8KzO5EdLoY5x0ODrCqoi8jvYHaBtWEIbfpNq/NlEmK45E2GDDizgD2oC6+kDXAd6cN2
1Ni8A1gGNK1LI01TZYmqrY2FsuJgg/qmzQctSlecG9T6K33HI9yzO9FM5LCJKfGOnqYp02LBwqZ3
e1B7RaiksHLrydhtrtFRXvscp3tYn1RI2d4VLpXnlYRMrVgHYE6/R5i5E0l5CBwwmOUtlfBInQN0
+WSIMqyrGW2JmB31Ehbc0RyMi0Vw6GxGISROM308k8F5ohmzmU8kMGdZNj/0MYQ4kEIFun+AH5pU
6aubyH/c8UwzE8ufR7clKscE59mmKr3m8CSq9FzC8NujgDKEeUKi7WORS8DZjU6Hn9Hxqy2aqApo
oYdyHKm6dl4H8RhPCzlco1y31y/sqmy6pfDzStPPDW7qBL82U+oVlPL0MCJ0X7dI5ZOExCcImRW3
3/UyEdszasYMP+FvFescfe8WwzqQQoGrMlehr73oiEunFdFN2gtG4Q7nNrPOOyqETUktTJ5YYtrI
U9ftD14pb0a8WYYhRONLCQa99VEgCP+vPipk+KeWlduEIEqpAKIdLMxo/ahnCwm/H+Xj0EMYyDxd
UiwfGgMURCj7BzyrL+IHs2VE9Gx6ajxa9DfRVPY/5D7ZqyHmfqlyr9TpHCaKrLq25EXrPh2PG6V0
z7YNiJSqdEFPINtbDaCjVY8ZxekPEtkMYDbYK75rnB+k8mT0a/lQDr43KvtQM68Qvjj9Mkl2kBTR
czEwbyKqzBu5LxEDfBqd7Vu6uwEbm/lfRbJVYjgZjq0A/othhp57WzavQlOV9H3QH9OPnmrFZcx6
EWZbbOl6NX1DwO33St2529ChiNnV+rhf05zzDase6vC1aEWknV/K5xJcXLcdS+dPx4aMuvp4n3F0
G5GvzyG0W4Mixni+3zEZj+ssOdJ3aalzEH67HYGun3PqXmRnlF8MN7YTUDUFYMQbolI7+g37oudd
EhNVJdEdiHniLZl20x3qk1xe5cRvUl+a9k/kkQAV3DQ+sXPTEeoBAXO6FNRd/tLcy/aZzcthTbP4
qR5uIZnftAk9FmcJF6UjefnsJAcmTHw2DYn1vw8RkVJrs/57f0nWcIaWykLCpxUwlD0826usMBN4
lyGuct5GuyKRu/GgAL/srPHUbkUUyaNqeiyydHB7PxDHXknjscz31l+/JMKMKEVv9wGr3lf0ojZQ
Snp8ZiPWK9nsuNcPhmwRF5SgfKNy8J33eCKTlEJS8HqBerAke9gY88esE6GKTMOkbxdtKXyO6de9
LRw0ZlMupU493Q78VrtsF+OUOtlka2AzaLfvgbRXggV7zeyjdo/onavTsXOycimyXVBnLw9c6hEq
aMi1MwOZrHZkSO+0HfCSC3ghz5ODK0tuqnheXryY8VtYck5bcIJFt7+46TxXstdG4IphhPEKWSOP
BWqQdVi7DWhs3fifqKPM07rxcJFZX8mboM/Vlo7wHf5Pn/c54GDlUxWj4P+hPY06M60dzrSECU9D
+aQlv43oIQ8CU2R/qQJP6FlvijAcvCXteUleU5sEOUDjuQSafl9wJstsiMLE0hDaMFqQq9Y9uAbX
ZvyGXznsUb0MrsmxB1hS4cVNi4zFuovb1pKQJI4/4EwTrSgUYigU3hXXs/tjgA9XMee/iHiADenZ
mQlDkpKZBvGi1JvHN8JgcXxVRhGSk8A9N5reSBPT3g2X19KkbpR39dd+4+sdVcOfrfqWqZcNt1qn
MGLKo8hRsmnFmkfTtcSgTzFC1R5byiaMB5o5qYXfnAHiAbm6yPTv/Fnv0GHztCXNFrzIoNNMQjh6
twA9uvUF29hqafyXMcyDsjT9aoPC2E9hh4+9vm1/3QTVAKwJ++kBnokJDvwKwm9sblJDiyK6lbUP
z6KWtYeZ3DRWZfS/31xFItQG8V3NomuNAOKXTjtIfgiGMITh4S5+Bfb5NSHdJ2qPmxTi9Jgy4X3E
JDNSivxdi8tTMX/LpX3PFmTUICxX2pp2H7OokBipvBUcGO79s8uUZD5cOarC40uRvkiCd0NLR+1J
hFbJvGMImtFNGlAkMhMPFiRg+vFi7hg1Xsx8Y0FISV4oqNVqP9DQxwxwusF9uXJKxGPGZe/WyZDc
StulU+yPkIUNDv7zPF1jDlKbjoiTQPH2L01DwQchXEvvusO75WsmVf22Asv7Ia2pTzFF/crGtkb2
JltDM1d3u19kCE6mDPoO93qp3hPSG2rapmrFJEivz/HuFoKiA9EAQG6/BrEdiP+5LKVxdrxg8SXV
vIEOVqe6Z6JcygOqrrTXfuenLVvCiSMuNB9sMjJEXugqgsilb9gpsJ/2iZPTehXzCwqaqeoy7Esz
kzRgmHTt1p+Z+88qpyTuZpUTGt48W5G21+AEUMPQtyB2v94j9YBLYBBa0pbfQGqdwCRsIQvR1hUf
bBU6i1n2iklpNto40hOX+ConrBEs+Z4JYI1zz0hcsiPDO+lcvd/iHbB/V8Peh1Ho/LG/Yv+bJOxB
M1kh2RnKySWdpR1EIiDJTcEMyIpBLYQcCMbBHH6qM3WQgiHK1m51aITqq+HdM10DJJ3FD/hLc7Z/
k48yQSQ4pr0tihNQTdVChqYkENt2ZF2bXG1gvf2yP8YmnWPQP8QiH4wflnYM/6s/aeZOpWbEhu64
MKjN2FQIqptWBrCCjL41353V3/VOPCKeaIL0KV3oNO78COQsNIpOAHOs7iN6EPoAj9Xu+uW0HDPV
d+wvZcAwbAGzKjk+bZ1PwSN91Az1EE6yfLvRJP5fXmC95dTmCQy2wOWGuWrtsrz/nN3XfOjAwwvZ
Rn0N1qJoBf1ZTQz95I5y8KNCsaGcZO7cg7/Ethl5xUGDh4C98unGkfJuwnOg2CEA4ILKlwuGk9YS
Pq+UTrA1yR5HeYW8p+DdVkGGfDSlGtc2lJM20VP5dUUqCiWlAF9QoZRgTDyJRxuu8e+auxV/gfnh
YKLvrGOe7Xe8YUD8lE/beqgzSAa+5tF6ztvOpCRKqZczzku/ANCrQ13k8zn3cXPKUnVTrxDcgFpN
NREkwiWPvrnU9erEJQxLf4oer9wGRTUJ3TSXr9PZvsoU9P3PHSVRTwEbX3Z4rvBd4J6aiuGy5hSz
pqmFpsikEGE4hqYCDQuY1OzDxCuV8tpP11BotegKhRNfdqJqGRd7w7Iy/DAqstU0VnGEQQgUtIhP
PlZ9r4kLla5iroSfzcXEdjW3LMUfB0tarY5UXib7hTYuaGjFR4xBT+vluzSjNP+IVtrKvDx0PTUL
ECt9g6fqkscXHAkAJUO+92nj5GHonI9S/W+RLMj+b9Om6j3qrW6H08r4UZBLAF78H0COqjzpDEtp
scMpwF73qeP5L+UJNUZfCvNdMxwqYnMgcEp1Pn/s8pL94zlS8Tvp8Ko4WiRGagtNgShlBZKFkCF/
3CAZDQPEk4OirHXdIB7wKLWEvRp4nfNYCNWBjMa6rPC5EaqLmsgGwUvE7SDrJ8pDIiXPFidmXr1V
Wh281YKZLXJmpqFJb/IMJbBvstNKEwswf5OlMkAV6KLMpS7/es/iTfRR3HnVlIRu0ZZzJ8QjmFbh
ANw+6+DTZbNj68w2BOjUUStRNgiUZ+QE6cCv274BZaACakvCMpWY8OjNFtT1wl8fThkd40R9UnRd
CsrSpCMoRaRvj6jTWbxIOyTGPytd6d8bwLNVfBJUuzZ5yKZqRC4SF27LzQ3UPmBSXQjupMPEbDIB
Q747ZVSsxK06/XB/4ZOnRd1PlvMqmw2/aX21pzyOcgMsUHAcBtda65Q4Qk6XwHSxA4C4p0fb5uPQ
AkPcTn6jfNVXjeNPup86FPVfNchRH/aW2g3DdFKDRrXDkMbbGys9oExMeMAT99Rjsyhu+FjxHyzl
lV+65cyuZgJhsQfEX6IY/cDBAawCY6sCIXHoWczp8XlSYtUBjmGyO83KVXn8rRmFOF8fdAO90jm4
RnIFDfq6AKvOExyHrIo99mOHIWJjsBu9Iop8W3B/Z3VVAOJHAXRY6zQlpmbqIDsbQTMqKgfJG3L5
QsAqngZhvzYJBRYwwslnUjkpE9hNsVlzSzFBlW+Ik7JvFt9Ffg5mS9Z9rGA3aWlDyJE0DvVOyKe5
1cimreGvzZvies2mFjtH2YgAnKPPqCFMHSQUsQylt5wqP20eUUzzs9ac9RHEmGDah2EizpQ2addF
9FmDDlEpyXlDbNtlOXGCSIp56/8xCQ6hjJTQFoYYCe0VtXZYz8usjrfZXld0DmCvoGccXbPlcLB0
v/LaxYgzy+JH0ZRdmcEJxe+jsWXpzzO9I9/z/W4r+YjmfalzsEr9Vxm0Jl5HcfrAxoS4aJS7i5m1
vHtJVahIe3xsRRtW/aP1Dt2YRJ7qPysgFNR3mUbT+XJLGO8+wCfqXX9yN0mtVek5CmCFA0Bf71m5
L+tR+Qtje6jcR9oSiKpWCzxXyG6G6gfiYCMWs31S6/V8POaB+FOt7T1NJhsP2RbSsdc1Ajbu6tsK
nLbl/wuOrjYL/JvMfTcAm2dxhIM/r+3ZY2psNWurNq1JHdSHkdfr8rVUsGGCBEjwPiXD1bMyHBfh
AQk7N3aI8+2WbrxMDY40q3OKoA5RPrpTJRYk2LBwgMq9i4YIuQmjtz7iXmweYq/KAkYNdbCUepmL
cMEDD+SbmN3otd1vtHzwidB+5fpXzDdZHsOIaKoKofsRFgQSDAh3SE42RNOXHZpenPCPuSFv4Ivh
Te2rFTr1cAIN5hO03DgcTXn5K2RmhZB9RKkyR3AijCKnwfQzOc5kEbd+IeYmc+D1/z6N7UuGrvG3
GGkZH6DmtF8XgVyETryXvMKU9kwwNAwRrATfy9ZGoXbLz4pnFeU2sXrOufAGHLhMAbJd/MWRv+2g
WiQgKFrzboBpkv4p7qrI8/q+6lK4oIlnpaPyvcv1d8bhF2GK076YcU9Ee9aSrMv3khfrHEjvH4R1
5ShhoO/9DILemAFERWwRVoPasMEzYh6ojd2v0fLrxcsIy8nIr44OEOs7qMWH54YVQgos95JLBUym
EY5gzXbE0tifWBpnJ5AZgO4JGdHNfJzR4AdmWIITeXCeJUW+N9s0jn5oVc0PLRp1JR4x4Lf6Vf+p
kMQEKxRbB6QV0FA1n+p3cRontncHtgzVIQcXWKqHw7gvpeBUkbpISHEEGJdHvtCO6eExR6wd+bpT
9VB7rJn1afFitDtsLTlIET3FURYHoNQ/R4YWnvUO1wUEKR+5bHnODtizDA6vPzzKcL+QemMnVYLT
akncNhFEg0pZsJy+KIeQuF3nAcV23JeCEx7dKAMNV5/Ct4FF+DLo6a01Z/W+62SfRTgiaOGXdmUs
DqZ8b6WpxF2aewuwxK0zd2MQHdNlgvav8v5TXoGFygNO6Z12S6dAF5DBAmgk23gvdBuqrMK4GcFs
bVPYi67HcA/i2WIFzIGuhuGAwpP51oBbpWEUziYuh4ZmNjYiGaFP1Zuy7N8cG/ssfsUB/rq3KFAm
PZpBwpMbCoZDLYUeibJSTqHR+4xUPzuz1T7BW4DilI2tdwqDHy6ER/HFuGH83TOQqeK+jXD4hHvi
7+t14FPwlb+h/TnUx0qNrgW3XTOj1ItHLUucUyhHr+xJjeQY+47LqpiSyY8rke8JosytvYjEG7zJ
m7mwkGhZTFN9roJBgirTQjgLIBdDJOzqhvpRTBuuOukCKcpb+nk7Jn/dakrfpllT2kTzumicC27A
dcLm/AaqiJMHjRYs6QzbHmXOyO+/ZKyC9gqgkroNd7AbeieuIChqS0zvBsGy7cbLCEo5MJGuwKgo
CuVzmaxSGQg9O7Et8ZK/Daspa3k6t4jNFKgxwYGQUvcpueATEJY1ytuxH/WoiVcO0gQ6VvUtPfn6
44CLuDim0O7CeEdAvJ5omz/2NSqy5RESroiyc1gIb9Xf+Yx1vKNRnSu0cJxBGANvpdxlchxGkKz2
jdRguUZjmrH8V6g8f3LLaXUN+kl4k0c3udoiYysBdVecL2z0lFfUHI9HTunrqA+mVH/y8NYDODtr
EAXLqIN8ra6gNjQ6zPvImW0HPIN/q5w9hfcIkrfLedTXtn1OJUD3m0+CbFUMsv2kT9Na+WD+y2yp
Vb5KrEvh8AwdYzJqe+epTDyF/56MBg1JwawHCHRI8D2i2u6hnSWChZk2O5GmIz5RvnaiiQnWA5P8
K2Y/EgX6wRzbVxZqnoA89RYfQt4SFVpUl5k2VEFqGh7AYtUJ1BfJkeZoDDaxYmtVNQxJizUL+qkZ
MGf80Q1Cwb5HVLJCgB9fGJ9O99vzg7aYbcRnBtZ9FPSmqFPW4TzAAXdOKooRuzX0493QECw91a73
Wg1qqrjC7N78ZMS4UF0y20NUhGIO12EWZvXY1oHDo71i+Y9vRpdZN3Nt59j+9Nysog92j/RU/dIZ
lITElcV4CWs/vlSheqO2la5u1RMVPOKf63y/LwcSexCvFd4becuvxXuIVHF2bwUDFFjVWANiPgon
Psuxl4qkuVUkUJLt3TwoydIGlQdTvwF0mVlmiFNq22omf1r8lVdf4cOm/2PtREeKAErSu+lwMCuW
CSLWWvoIjig4n9y5gvyVrVHyhXdenAWnj9koto84Iv8sf1wFOzS61A/ppmcep9XbFYWs8kzhuFds
PO38P58gKlzSf1QhsZWJm+oO9HdEgzso/JFeGWCXtF8m+4Qkp+8uQR6Gpi3oop2Mh8mLRnDfcTP4
WnVLGpC9AIOaVoHt4uihzXt+Q5emtI0AuG+9jtCjRt5XdxyeCJ2SZYo9gfrWBXXSTwX/Q147Y89w
xy5zAD3H8XmOypnpqFHkbciCLcK/bmm+2AwF2Ngv019dbnMrb9k7l1jhGqzSojLRA2mAqOce60BU
A25LKh3ODYYCTy0cP+MrsHwJBrr4r1pY4lA1gtM3uQfmDorFYRdCK56vkwSYt1qfFd+Vk2egG93C
4lDHOMDwfvQuQqjQanBgy9oTnZQNDQ52mf+8pu9cboxMORiPCn9NneW+5VcEKZMwGvOQwmuWW5Jj
Fok3f7OZE/cdxkp7bMJ38vElbAeDtXlgqxR0An1SeOz9yW1ycBK2wGPLd/xU+Q51TxsaAuEbnNhs
YCjkbmJ6baDnh2MxFp1syFhkfoY6o/6zsk6ek1/UGu7G98hiUUuTA7jldeOJOQaADjpwjm3kVoWC
SgJe+MecC7m4bXLgveRQO36+RTugFtbwmK2144JuUMQv28UFNHOm66wTE1xucIxCGhlb7clw62c9
RkM97e0Wm4lxKOJhWfmKDrKnbIzIzikCiYtFK2o3AuHr6csHNETYuQ+A80STHkZrhTbLKtQJKbjM
NDVMZwk8fSO5TvEojL0Bm7RwJXsiiFT5+T4ZeFAj/ScHUxSr5SM+mTOOST7aCYLkNrJBP2hV5urk
vrMZItb7AHr52uHG+3kEhXnPStrALeMLJpgGFnVlN5bvOGcN17nsELAAUmT+2D/Zgg/Q7rG5FgxY
zJkvvGORLwWLJPmN9KtUqzRdklM2qNZWJAGOInROtGhT7uVBVm+kUnV5Xqlc/Ye7/UoB2EFptjl0
yd7Uke+raWWszrgXaGEgTqfd4uBMzgG2Qe1q3MmVb4vzKsCpN3qIzb6GQWZcSLcS14XVpWyj/bEn
vUkgaxnq80cyRTc2wtLteRG5itkfiZb5CO83D/6fmdAWhV90CeR4VdIa8VM7mu1LiFbB6Z/mNmCg
DayT7xVSVoaGv0F7xBgnejVmvmJYBoeKZzYK+XNQXZSv2wC+/hezU+mp3895xEug7CIi9f4kRdpk
LK4+8ikLKmOh7hXRmhM/LNpRz6AwPzLNJ/r8hDBLs7pa8u0aLPuNqU+wz0HAiA40zJHoSGePFsW3
S7XI2rqShe3IAt+YjV/gv5XVvDAUtohIasWfeBgvrXvHxjw4PGb+bwAtrV5y+VJUjepwcJFxspJF
7wZ5dw5ouf3bw5riMt/l/UyaGVJpzXGYVOh9OxgKHC4vICbjuPpVfn/dAidE4RbVsTp/Q1RUL4WI
Z2A3UA90uZLpB9Lc5v1Yfkokxcj/iZF22WlRkZDjlJ2YyobQl2YUiYWrnPQ9nEIpeV9cIIBRDeri
5hbG7AiL9RPcRiYDXJrS3dwsI3Kq1U1/l4bZ4fg/YPpi8MVWNLcSBRnHR8iAPZOY8Ow7pAIzwvf8
HvZqkd2WUiQSiAME2iyrpRyl7ti7D89WXSeghjGmqjiw2bP74s/LDeZmUGM354Woj/Zl+cm3HBKr
qR7TJOzqOVc7eugYHybECH9hh7T0APrDYOnjw+U3/kPK5fCVrGYRWGBsBd6haoFFsIZt04lCyPVz
KBWSIl/7yitaZqvAHNem/f9VCjhFP1FiZm3DhL1QiV02KCXujK69nas+v4peerVtOBP2jchNsfdJ
GaSG7zP1CPfIONntB/S7I7iQXweMGKOXBv6lGun6mGUrUzajp8lLSmDvSIuIJPo4YMUUkbKr43gL
F76QyOEkuBjN2ha8Yv+BP0ahiyx8edz5ZEIhEYj3OruhtJybYB/knYhQcmelaIMsFSRc00/QtMbQ
g9aS7+fute4DukdGngQZV17Rqyvp6LDG8GqFWalARWj/2Mtv7+9Ob9CGT1QliGWPqvkz9kwSwPTH
XuQohu6pI0TumNZD/W3hqnRq7J0IJDhqRVLafTKRFrj8wPWE15Bl/X9q9MAIAoJP6w+l819TPsyT
2eeDmDqzqs56lef25eJvLNJDY/oaYCFhphfIk8ijBaAgoHu5YwlZgv3R2/Hwm7ObuvhNNBC9cN8R
pR9vQpypwcz6VPClnntqSdFO126keNsnTu0K9sD1UmTbnAmH3glmBUGHsN5Po05BpWJTMYr8xXcJ
DfHqstAx3G/NlFbpC+ZOI5xpOnGKlTVoRx9FwyOGqH90SyL+fMhlHTowG1IDmVaVnOdbTaUrb4l+
moG6wcGHqu3ZsePpAqbYuWjY3we7YgqVTlcZj2pDUHKnzUcDWiwgKApw0Bi1ZFWOJ1FwG26prVhS
21TOwCed6//42mE7/bVQo2obwf3RNIlyVxmtjTvgnF7X7efXsVGo0F7eIW1PNeuxs7QF4ESqdRf0
ow54UB62xJkUOhEalSphZE3x1GTE4U/9RYlAeq8eH1faFiYibo3VrqQ3uPUJfYEjPK4ivjI0lVMV
yOE84zUnFj8tUdiMoMg7/AVdfcmS1RwA2D/7Tjp7gn/nqAjTYuu3B0fILTFIITsLPLsHXeCGIoBS
Yj5oipV0mx6IkbdcJLAgLoUQCHySMRGiaEyaEtqjHqoLZ048m4g4GSmCgkEbriaOq/YbPxcIuFMI
F1FqKNPXNpToEIsu/kBA/COI1L1YhemDwgVgVilz+WfxSy1YUd1sY6ssv1+cL628mepAow08lsVt
FVSXGOj93bTBHZXQVBj2z+LVkVVRfQyHRgikuyvDFqRuiPymq+4Xp5+iqgoV29gHQK9dy4b89909
pfQ7DHbrziPynp+t+zVvMKQEx0ke/4Paz6GINz+ca6bsZTOxiOv+7vBUhHli/Vw0ydbqeGEdeeV2
m4lrMQsj6RkhuCb8oVvPdh8NCp5lpu72oPNSi0gZa32dW+HafDzeg2BfTAAKSe7ALqHbAwYUh0fM
apd4yTThNipIJWOAVY16kpAJ83JudnfuJJNkTST3QKLBWSAnDF2dITY3tn8N0KS0HUIJ99me5K4u
m4mqBdHahz522NJHZKB2dohXWocxNld5EzNmHZLF2X4H5AzW3wN297+Bov103LVOX+SnoMOh8/+C
PM+f2ei9gK9UvAKe3mEejnBKXnpqZzFeLc1AFg6PWkPwWW7yhpDEUOVjtM2DRuwi1idESIuFQzVP
xRRo5frQkHKr2whj0bPdmhsFE8dzaKOQNhz9OOnnh/8uyvUFcKWvJt928vJuxzkpMqhfbligcywa
kFteJyFSEBvS6Fxu896MNedZMYXmxHdfdM+ovaJR6Ar8w9nfqIEHnSc5aiV+hP4p5Q536pvYNy9l
nX5oXazmM+EwBzb15aBSd8iwu/wsS5gujoeIs7smfyYkXDce1KzIvaRtwooyIxn6pPLKqFdETG1m
8QLPqb2kdh9dcMdczr6w+hPPe3EihlN1UXPLIB/u0PSar+KMNdf2XdgKuWIdw773oMvEJ0exyPAO
si47kbTmZabcWsuTd8KgEyElYGcGSBwntq4M37TnmPGFufhwfOWwaQcgsiC2ygVRgC73H86vM3MB
7iHggIxVkBS2qVZ1wKWyw/rGT6pAA8jgWwV8fkbW1iVlzr2BthD5dStXoNXdGulMZDhXWxZmb7wg
8rm3vqiG1ZbID9N1QdTsA9U/PLq4QafgI0YzSWlCkt1kRO0zigM4hwETh+a2y7LR42UR9I34YYHS
Drdij4OeFwPsBhUGSWIA9mXgnzXCuOmjHe6NutN7LSHxl+6uZXIkC0cb+h7P59khC7AePzNhD0NE
orKL9CYjaHfyBBqgsSYQpoxkFGuouoeaJKbkmQMmUxXC/LU229NwydG9G0NdHdQiirauHwq5QQEN
JFl8SgHbMWo0msyzxJNwLY3BPqek65ujgZwI12+okiaLrFKixWCulp3V0IjMjzxNm2MSJXBDA1PC
w/LED46kL6hBWZL1dw2ecf/WRjXV2hUQyHK3YcG1dQU0/uNqHa1f/gfH4gUD+z3uPUqXl6qYw0ZI
ua+eEQVZP+AgkLlshsUFKDURGaa8FZ0PMY7y5nQannvmwlr7krTDX571cYatXqOYxW9Wi/LeWMDz
I8sGxmitxGHc0qVYUAq4IGuhj132cbtO48e5aX331Vg3nx/IH1W/Bpd9mXJ6EbkeyBYJ2gNR6VBJ
l0QAn+VxqoA6pSMGmgGrv6O3unIWVftTXksHanTlfeBakzTo6vabQg/RyATdEGMpkzoylSa8ceSV
3UY+/1BMNQ7/F8qkN7mTqLsvSEXjj1Vb9KIa4OYVEcZu18Ll3YEl+v1pKyMTfZMXafAxHxRg5dLF
nI0/29PpQtu37wArEIix/vryGmzTiF8ETdnPpqr1smBbjAnLj1K5/ECnJau36zfJ4hga+oRp2vJD
/WWPAEx1YFGNgti3M/l7R/XwV/vP6/FZJC2VRakpQGHxw+dbcOv2ISguF2SB85e8/tjJ+Lb7A6rB
pVKrBn/HCl3Gk+fOiggGax1p1OwsD39mvn7jcJN87e+6nq+uaJKftHmCtRvYJBEOeJ4rfBtX36Gm
akESsr2+ZoYsHxOvR4mX51iGC5eJq1BNDotY4L/wOeW1hSlBw8I5Sik9TRtgW51GqAxS8j0f40e6
Aq5C6BMlIM+bKt6Th8ISWiqlTwUDefj/C9HGErr4miw46gw1BnrCkX7WFApna/U0Hjqfvoo9Mp97
fSmbHlSP56deW86KsLImqVeDGZt0ew7FwJl4DYYPb/FQZKqgvFyw+e9KnMuMiNHwN7xSgghqryls
BIYlzY2uvSogHuUQOGBukh4MBOa6gco4uDZ7KnCpB3ZGdjOHmFIp5/JjkYDE0mW23ndv0ohlMRjV
dUD1CbmwSPl27nUcZM/lo0QPGCQdFkcyWsPq2R7ZfHzd9SqVqNFbCkni5noANSElOzNSa7SnfMf5
ziTC/oi8XbWeXjhXKO0IU9OwwJMaG/LiBUlHCH3x1VRcpRKMTO6EWTIr3YTzmKTWV67Ht1PG6vO6
2MYMnHTrVowktF/60vAFbeOZpyPHh/VIa+xkybtyu8lEfA+yN1Ok44f8ZIU4Eome47XS6gsu+xgV
Fuze0/GsQdgJwuZOfmJM3Albrp+r2cHPA/jv6zneAFCPrx1+nWfqV2UZxSPpYJVzyveEUCw9yFyy
K9yZdtHOpCQYOZrxBUOAjsxv/fYvRXs8MJYGRVjdO6KW+ITpHr965BCf+mBCBVNzPsh2Luf4UD9O
ePXPPiUtzo3BOex7Gzj0i8a951a2/lJx5o9gTUiYYwchNJnxyEDIHDAw0MlVkbr0b0+1vwWdEi1U
4kWOfavlIADvt+vW6EkpWM2JOaDieEeSFWAE0h4bLsw8mEPwVTHQX3edCFw5HAio9WTlSl0caoo4
EUSTb1IYNnKbf0oIL9AI2MTxRwpyqHQ96Pa3GUSch+MVgL3jLzA/ZI0FgGuzSARN0vPth/Anghze
sp3j9nMQoB6wIbN7d8KPou8d4iYED75BCL9OTY+o97U+QxTb9yy5OWyzOvHW313TATkGMGzCbavn
wUu9EhFf3x+pgJmXGeDNMsOLvutJu/IqyvVW4owVE1m1ool2RZzqPktNErUVINQ2gqzCKJ2uUq6W
gXO2+anm/WNyU/zchoP2QAyvzJ5Idn20bJNy+2T/rQu7DOB3IpE9IMvhQkGtbk2Bc2R9qsDwn9mq
Pk/074yv5Pn/CBfTya8VgUOnHe2Zad9+WGqFkPBcVB0F42XavWxD6+16rGWyel3fL2SjPTy2vyFG
NAyQcOuJLdypTWhNfn5tf7IYJZSesnn4D2/TrTbS6YXGA6dsGXdleWc11g1fOEMYIc5MlY0s+ly1
vkvqHtugMx8cZEeky27aqs3GXkGs+4aN4HV+zGqC/0+VukvLAwbN1I/tnJQDR4P3sVl0ol/HE5L9
b5TbkoGsi6o2qeLwfeTt/ZbjO3pjXCseWYEfNRc5CrlRjtqMH0Gplf9O3gxqw0AmKreU8L3Bdbje
IgJwDbS3WBlnEnqChk7XlBwE6AHRXZKZTFUw/Eo8RSKeaPc+4tLsIo+oh6SwcsmyyN/C87RAOs8a
LONfqBsJuh01n0HW5zLi8LPIv72i3IOIhigBj0Rs8s4dFB/QVlSvHFk6OH8xEmJeNEgqzguwvkVQ
pnyeqdyXo5ECvzB4T0fu+GkFCne6vHabCdlhRGkPn6qy8h+dQ8y3/i9tF1OuhAjwApoPtVDUt16U
Hb5eZlzYgzhNTf0XtHHhU6rC1SYTUAmYNJR7OKTBaDFRcKLWBK5p76dy5utT3o2Kz7La3cDWY/xq
XKIk3kHS/crFoM9qSXIYIjQDXlTLrO45C35aUbmNw03n3te9QRehk3upObO1khae0cZnSYDYo1kI
xedPJEkXmBcZzLQeLBZrspnRj7RIaGaV0rBWLDN7akz+39PUK7YdbkbqRx5LpjBwFZki/JG5BEv1
4FT+mfBetdNguMdyPNhBYM/2ObB4/XcbrslPPTxHOD9YpPm/P19kWY0ZGs4iyl9S3rY/0WkSr6fY
OhDCY7yfhJYtzZ0PaHGQ5MWypsLVcxjM/7PAIZP8SZ85A9dfteH7XSArxNR2L/9vaoTaGnN2RAd5
dmXNBuFPCkS+5Hc23EgR8Yce3dfH/8A2LbHTpYdv1hSJjd5mB7rsu6RFm3UiYvHt5jcUSGmX/ogf
pOBa5yu65q5uBFQpKn3YGI/eaqEAhqf1u4lrnKYNvn9hU2ii3rYx+UxwiaKzrnsCtdcGLyKUgg6e
0okNslBlvbnruZ0Fvi8vJnUBKwekOzUPRfQOr1GQJnZTeigrDkYs63Q0Xz4M4b9i3KTuatih0KHS
drsuWBXm30Cx8edjhXSlU4eu26H+m7lghzTpzVQNv8PlMfKfRqzZvTsiUCaKTwGGF/ihMou1zZl6
1lMWT13V17aZ/gPx3vHR76TsJ1XribZz3vaXE8jvGoJqqgC1jJQG8rxiC8/5gK1NZeH6vY1CcOln
5AoAyGcXyTLyxgfJ1ZsD1sG1+6pSF6+D8E5tMVXjHt+Ds7JBKW8hhtn4JVTZv9SrY3Kp40Gs2kVt
mPX1XozbPwEmyH77Yx+NLtNgPyVtqjISQDz93Zaxoz6W3zuX02Eho8+QmDX9sRr1JckXB5dVWKlI
xE9Nq2GNVT/lLZX3TEP8Re+OgxjWLYwPY7Di1z24Q2rZ9D05FPE8KP26lpXwT6olLhsalp4xXWhV
dI9fvY9BrRMKFrO3jYTUhoL7kaw0/vDaGqmMGyuVk2o49C+o5xYEiD8kpLlVrZykd7gVUbpoHGdz
EG5U1bK8mIcFs/SW6Dgai6ue7ggiond5vhBt59eJEi1CHfThVe4mH3E4NdEOGoMlMtoOszRuavzr
ZgMR+c/0cQWElk8gy0yuenduC2hFPNEIMs0xR7iODkT7wEVgZ0iivb90axgROR0XlRGLcPSshEBK
YIIMBVKleTdM4wf+DSmxfZ0fnN0uP1w+Ki5TuNE2KW3dUoXX7M1vtgn4T6MY1s2tb1lgDfSXtiEd
hYwlK+9CzYFp4nKOGO3T+aSh/3YV9ni1uSk6Kjy6EdvD0YbHAJiD6c/bvQs4k5nIUvgn4AqXp/By
qQkodXqkYrF5rvvpdnSOll5svt65mRl9ccqPprr2YPujwe9NAyNXR4F7GX2VQiU9O6sM+lZzXT4D
nTaF9Gq5GQdoICjE+t+ViYYr0oHr70yA2V6HyL5Y+/XJZCLBd34gtsMrSKBbQFQixWiUMTvy8PmL
vDzvFbfCoJeEknGNuCtuQqs+twpVp6lJ7MWrQqbXzXpBs8pAGWLNXf42yMXDJrJECKftcYJkoBxU
HeCxQN2rhuzpO5oU7ytx/vYfC08h2uWnVnAg89zZioMhY7P6ZqVsR3E4zwcz2PmqiOasPWAsVVC2
3XSBF4DT/JUGcl7QM7eeEGzf5WkITXmnyXPBxq5ka0/B65DlEVPApY47V67FzLUfCECRuXGHqBrD
I4cxodgcoFyTe+pLTFk7koZNUuteBNkgGNduD18QTJdBnTk/+Br7VaWkl6BSJtRttS19vLtu8pEp
r8/QRGa2TRcsC7aTZk7r/Px3pkKpQ9+OC1WL4pI0WOE/T2Cpve0qmqj4qLIUhkL11zVj7fbJmObS
o4CF/IU1YeE2FAnr3WUjVYzzREAk+DS+o7sGUxupEdQuyN1TMDY+W30y/eEg5hMnuMdcSUiHtCZv
qihJxnRHXITbHX2Uhg8/2XLcpDY6+WhHuDsnjcFInUjeTdP34oJ48UXP+KiaHT8yW/6QQ6MnYFFv
7A0FwsAjwIDlcfMrIPyrzpawo/x+WXrD1SsFlM0qm41kfTxDaxNMqfh76+ptt8Xhic9vTHjFGGJQ
ujtLijfKnt4gRp4WHSIKCmjJejxfAbJxsh2V0JurQJETf2YujIitkc4QFJKNdY1ATSZ9z7ae3whr
Vy2NU53xmwtz80siJQ7DsLXfR5STolcKgd1ega8j8G0oYBnBtQchoihF5g3ongpyjGinpmE1pLUV
WJZAXsMioxtABF6v6nmLSqZSNi5RvF+YyBqQxRYH3B5yPLKiM62hlTreX2w+yYCSwZTnTSEncGIs
COitUaHC3Mf/rzHWteaUDkDtl5AZ8bggNGNjl1JydyqVEcw004RtA7l0SkPwOs41NwOU4lyohWLd
YIKQjAnQEElGk67cC0rzUkx2Vwjv9wYsUs7l2IjFBZT25w3jvCZQcgVZDfBbp/O6qSfZHqURASPE
ihsdEQd1CLGAndchWUEjsbCg+x6mmucXS0UdYr/RhfIEOv9RQdX6rfHiENcQ7izBngHJTR3/c2MD
03R18SV8Iohb0eBFPqoPYhWjra1cxVU0jzJOHkIb7b5A+3HZ38JdLaMBJxM9vFQ6id2gJTEfxmQJ
bJ9J5hoXfkzKkKDt3NQ21ipow9iSd6ZsSScB4n53kGNEg/oZNySjZxWPcabGsNIWYSs4se7mR01X
gFO/H+yLstOJ/suYLjtPCO7m+Ks/NPPQiMQMR+N4CQqeWcg5VS2C1F1o/tWFaWruWcczik3yOVK4
P3+4MgnuE53k83rdw1g48YGS4tuHGTz3RRT+G9e8xC4NAO55KKhYRL63D/FnhCrrL4RIOKiz2NYV
qUN6TUjOVvEoumBKat+W2sAEGcuPpxADJeVmLMnQ+LEw+SqeMpz9tRD/LW82rt+MZqQKo54k3l3m
CgCQMzjLUeYF2TCD0LmR+wiB3LDiI9YEjw7zhQ7xxgqL++MoqWIemPSt9sUSXljh4MK0kcR/4kZL
MHu7/OH8Im86IE8Rs2qSlR1k5+Rwt/ee/Sble96L0IEVBnW4JkytsjRcL8qTdK3kWGKVbHGtmzHX
34phRNuERtcPktz4TKkrveE0E0gNOtPlr7YASvyFfnPhv+FMfo6lAjJfq5GqsiB1W7IC0ZCftYWB
KljM24COjI52SgBvo0Sp+12KdDxAekU+i8Yz8VitUyVdkIzmjEQIg6cvD5hT7ZYSUe8VeznqQnxT
Bwh+0OwGa6PeWvJAIdG70pQJr5eMPN2cTLA51+5WYlPQBjVFkAd8KvA2vGDF8+vmd61Iy9JBW+Pb
H9v8UEVNxmD8dm7qNFOxAe49RwGAQQPmC0I36KVPjk5NXFabhgSY41GYxT6E5wnTnYneW7kf/mc7
Y8ddH2tNtcb9mtzDSFlZRGRGFaS6e40nh3z6AIyraY1TG5MIV8RcuHryRU+7H3RPohlgn0l4CLHi
nLALC46F1ZJpDLdouxJJgw7NHftp1yQsRGvYJuS+RE+/uV88xbxnlyhmyNPPaPIgTEIHSQURjEhw
6QtJTopO7ZKShj7rl7sue5jgF/kwhds8etpj4yMenqeP18/kEk5MDp/25bw2/Kn3r7IMpzZOhwFG
6QqecLd/ChqqrHZLpvFRLvlWt+u/hKqwJEyhHP4/Fhkr+OO3urZjKz+ZiYNVnwz3hcTuDCY1VjII
QG7jDZPDklzPvC3IW2VpoFS65PHNhrulbdvHlOd3BMkL0uYW98SH1G9H0zeLdglOG38IMj9GCdRG
Kt3ZyJENVGZ/zIQLsCesz5ZhNT2Iu+gsdmeTmSnKMrrNUZyrVu4JojX4bJvZ+FEbqiMAbX53BYTl
Oo3fFyIb2+szoIriOlcTze/ROFb5yxfvBFXP//O/E/JBAP1+vJMI1/q+hJvGYr2BnlFkBhmZ1ZAX
pIGcGvGqGOPNGriLo3eV+0glOOK0c2xINDyy7oO7sBNSLm6OZQReKGP36pRL4VlNa3vvnup1TCpq
K1qHAZyp+xkrH3Q3qNKVwEXVX3rSbkQqgduOyiZ9c3K9crpXKyr5kzjyhLcOiHKS53r0sOSvxzm4
sqSeH4MTpD3KCAzJBVMJ3IHTC/8O2mpz/cQ/ai+vM2vwiG25q/JzKymD135ZmfvChbIEltUCNDZK
alCj/kZmybmm9lPNHBm6pLtNDzIZ5dGD6syHIcGhjokdLTjXyh+y3Niqp6tsoAtchP7Kl14Wkxe3
JZsiOtxojWl67EgL/kXGTQTbF3r1kWEbGyVoivyKfr8ZeKJWgCwV3Fq6TbagSb1JhUgnJFUrVaR2
31aBg7O44pJuh8VseEuGfAgL+NN5upm9RBkHEeHbXCBpjG0j7kKvaZ+pdjk+vva2dSeMx3P2fB56
pEh1ZrRhT0F5uJ0SvdN9gbGBpCqAAaWyKIE++VpGKfHHo+yW7+JxBn+zGyL8XgFo05z1K9MwSHnQ
XV2vg7unDKdmMKRVSjjqEJqOMWb4a78chtyco8v4ClMJ4nRiORgsmS7Je8ObU3ABOxtI8eXYDJyG
qKZhL2sGFh2R5lKopn0HpPIn6j3j0VVShykIuA9ZX/dvpfiKOEkp6fbg9QePUCIPMGacWaCKBwQR
ozHozyS4EkdxjUR7tHVk/7DlHkCsvwT6iDcjMsUbnbNzVifkR0xHTHIBVgHvsUwqlPXv2g/mS7bK
nQxOrgtHobT/vdZUhyUIn38/5QnF4WZ3v8gstNaMUKPRoz1SpViuinJr/w5M+poRk4nyIhSxns4d
OPIkp9cIIMBIK+v4IoUYSw9RjbGgfbwMwWRDUaoYag9F1NBBUvHsGce+gbBn8tcgelXwy1YSyUmx
KLzR06/cQvCR5Y6x1VA/RhxXtJIMRtG6kNgP9o5FbpodH6WOXQ3qpScbGXP03LB1w9N2V7r5LA7z
d7NIKN6ZL/WTYkqU9fqRtGgcSwB4/LFqyDns/m6eqwwJRXlzeswvZ0P4C2+lFAdnLO3tgoAJ/TRG
c2nsU76jUvGLMnWo099oeUau4IT06oafBVvd2QtyUV8ixu+QF1JqtfBaCb1utxUzG6swUzK+cfJz
Y3jv866NqDAG7Jh0guvK8eQ9pTFNP1QSah3Rxbuzzp7Uvc5cS8FYCr5+uhWiTETbLMlTgN3U7Xm9
9J6ap9yN4rhM56/SNBkLrLgHtc35cOSs+9SErFTkrg2AkjQnkhSOeCeZYBazKQQjEfiXA3/SIx5s
UHWiYJmO6W9W8cH3Q3Fy5JnskgT938GuEy6J1gsDnp2qhqgdLFKb9hzvNRiegPN9ketdigtYaCry
j7qexdRE4gCoPgOkKI0UvysP9t2ao6KnCoFKOmQkXJEtxNiGB99RN5A88OAjHGhEJh33s4wSqHEA
iBhdeECO5I5b6lZUJLF4vWsE6fsEU7PqHDBSxKqA11QW8t4raxNO0OVGA35wyxKQiXlrg+WaCJaE
XahINJ5h9J6AJZQnuKI7JkKRDUTfuqaHNMGebZrNMDJtrIM7GJF2YFDgqJAn4HQ/Mmsytml/ra01
RX9NjZK59ABSiJdrCw3X5M5VJwvVlCcc8LOSd+KmQPag7IMbD5TUQPGSz7UGytUDR1V3ImoFILTo
jx9blk+ZYO5/neGOAkGWptMccGsn/gaKzDwjkDP1I5siXvGvlIXenijC5s8KxGS7v/bdV6nTTi0P
K7C/Ou8STJYsBh5jUftSTYDBnvq4bHYzBTvAiuWoKfhqfY0uyfEFUaz9vMuACv024oa3EhlWMrgH
+YAumVrm8Kd2P6bmlGT4rjCAitYsiyY1X8TlHisoiWlYpFmyLmK/quWmPzB1hPhtykzqIe8Y+QVy
WzUsM+tnJlxvPi5KXCibCbkO7XQrnf7O8P3mN/pOCGNco3mZ39T1B+2YH+fxtV6lsuhCrWH+cVa3
gAo+r/2Q8+psFHcOKSEukurabRd7BNr+OkbMX7cmGjTSIDdrx3NxrEJs9YbeoWr6xEXVUemYZ4tv
Bte9sI5t2hF05isiqhvsnfRQV4QJNY6Ca/taFxxOCh0wnlcP0N+e0OqOTbli+KW/CpRz58bKjuj8
Ik+efamBiBd7FSiGOyiyeRXwN0x6R9PEsaomPJeA2oOVXHqPFX2CdrPubwL3ie7wNz8woRK53h24
ccUFbftRIKJgyowt+4boN7h40calopnEM57Xn4XQuCyRNGKDHiy3Y+RaxrWyH5fXlBKvcOqC2b5s
RPZQA+FsPfHw1Ez6sxNSVcTD/eYFAzsVJjdSrl7fyv7xU/kTau+96jjZVtcleZQ4FD5t7xgMSmY+
K3a3Tz5+kb62+u/mjNS6nJ5ilW7YmGPDO4mpGio8JFEJa8urcXDSCBbPiyfEX+nt1KYgfhBf0Utb
olkRUJXgACwvnZuMWyJnvJPMBxJAe297kjkuHhwNWLbLujlPCj0ZDQMOAEKBUY0XSAxoFETVHpFV
MLeFzJYB9rH0NrP6mYEN9y7S1qoPScVIitGu8phwA5FH5561jcjddKBe5O+h7kbeTWXB3V8qPzEe
fq53Tpg72IX7/fg/H/l9SYwhv4z7ce0QvkNQrfbtgno88LhTZRAjgJ1Ww8bM0ZPTUGcnDZkxnd1L
Y00r1kw1pQGEnOKcmixlhFwDzrESltCmspn+L/WakJ3hrX3zVMCGLzRsW+3Ti4TxeenAytLuGyu5
9B02YnXm/jYnKtqsOd+qk4HRogWfl7/TA/IOw5ZCyXBLfjSzHzKheMS1e6yFqvzSTTvo3KZie4jJ
O/mqfTKEDQ4EoeAkWJmaFpelaUxYBb0Ei10o/N+V2QnTBSrkaOxV5/EF2y1czNfMlh7xZAdDcRPg
rLHSfb2jTZlyTUzBFFb+Lio3MFBq9BlHb0DWFfKZNIK9eVbbYIdCDjRBkTd6QTfg7t+XwTNH7vTJ
xiWz2kB7CqO1oScEJ2j35tHybQRSEJ1/7N7IutDbrhv5bWHCXb+MFuDACA7qQ7LU6kcltHUWR1zm
Q/7oH76o1GKa5N2g4iXrYoejjhmD3Gu0lkYhJyLLvJ/PZ+ZnhNe8NX/QaHj3mLt29m9wZTvUYgC7
49iHz74O4B54bYRaA1rWadwWFxnTjYQDr14qiCiDvdqGxQGZKRPRWr2nzCgl3wstu77un1Rjf4IL
nd/U8tI/rGugTH2rVSzZD/APNOagdfE/jUzFbytS1WmeLrkgNMRievH7u3tXBqjmrsGu0+Eo5fwf
nEuYXfoFO+vx9sXMVCPivPkrBVd8WBS1ghny6L5iSWeRkDxQDfpJ6165WWeLyK+0OqCp4uoRWJcl
TDEvdyG//DyI0l2sNw8UOmND2s2Kbxj17XftGLceyE0tbM70O0OPU/mVhHwX5mpPEXF+Y/A2N/Re
3gybloXNDMFCEJSswSChIL13SbnclaQrUVSYUjtcBhyiuutKbJVoLnHpGPA5O4+kU+YRcthK2nF4
NpseO3FNw1AkzZ96KJFMKK/Pd8oMfOweFjfcOvwKO4OIjlE/FuI5lsYZMb5XGgT2dnutO8h7U9US
hhaeffzWQsiP99nzj/R4yq3n78CdiPnDlIWK8npMo7ghBFrL6T9QfIrONl1ud1iGfzoZgA9EXqQ7
EkZIUaAku8apPzIrac69XlS0OyvGWEJo9l0nVQz6oIYGZ/VLlQ0uHPG7fbU7MaYk2Bk2h0QCyRJt
hxKkoaqMoWWNimwy40a/Nog1Rq6jdzr2QS6QYw8eLZnGS98CLeadtK05PEb9qi/hU5IYaFsAPpF/
KII2FJ/ZkEqhCdEOljrucRmLp9SS4Wd+TF6T/Qp1mTcci+NaNS0BEVh0hLWAzrwrLyZ3tnLkZaD0
KxfUof0CNfn3tSlSUECADfz3QCtJEvnfHkKu7VhMDhpUMOrvJmSCDpfg8YD+T6dW6a1OKrDHZl9j
u2PAlkcjES9C7eHfBj8PqABAaOGn0GmDXXnVeR/GRmo+lRhRaxZGxDSjy1LWAsHkN9rZMMm8aW/2
TAX/cw6Dbx+KL2d2F/Pfcooc5eubavwLvTaN4XRyAGVatlfLzCdZUtH4tyNFc9z3UrNNIAvyx8jZ
ThyUnI1zhlNoguqBjw8DdvUhnDlfDjd+TCiWhWFKTTW/EbVOUdfbQh6PSga1m3XCnnHsQ/mgSAR+
YKkDaIjc3GH1Bpilfm2mokjUc30O30x4tP6GidLTLuLyWFiqpOtX7iK2QM4N8NKdj1164E8iVVXd
vdAtNgLRa9X6UBc7nXWps3veUOZuN1+uuufark5Gvn5kdqAEkwNu2SCV+GOfGfbmSJl/Np5ctFhk
ioVapQtc00LRNVork8KusXpraYcgXE4Y3+trLPcSUHjClkAwfhCS9e9Yr6wm37x4496X+kjolVOV
Ig57U6cpRVvV75umFHdIgss2qiCMUeZD5IzDeXwhae6mn8yTZFhAXwlVb187nnoNCxfDkZvb00qI
t6CjFZPONswlgJzWOVLlzmxZZV+1OhpT5KMxIufuq8QhTXXT3Qrftp2/k2IE+sNpJLlmoB58OAM/
YE8WsXyZ51Dv4GfNp3Fp0eccwD7BULlgXhL7AHEQseQB/1C6KIZFdRgTgcaWHDFIgGL8JF8yLZEB
8A0AI2pU/HzwLj0XU3wnDZLEcFMWkDsDU2qwVBYzNONi67qHv1VQfcRn2qlx+T9cqaj5cMxJEpo5
MZSCUgGR4WY/a+tBTNnZVUmceZs5Me7l+pw1jiqUBFxKPKzfunyJykE1X5adV7Xkdq87afQnmRPA
5XjaQkZUjhOGxyE5Q3YsEZzV+xIPdpG3hf7ts/YbF9PHIGOuSBVvgCzVci9g3Mv7tqztqERMdJ+8
hmPLDVqbwNULNsvel/f9fJ6fv7NWpwzGmxdCyN3a85QCMAPHDWVFJhEgMEjhYr5ASfyrfB4snGM2
OHMNvRJQd9DGLN2CyiMlPOEyAUKVUWY3MYFhvNn/aTyakFio/Pr3GDQ9iwEKk+zxU3L4Jwmc5Iq2
Cs1yjRyor+8rMA9Cbs6FuzsZpcO/pgoj/k0Q/vBu1fmuwrexNHGL3GZSqjPhv1BZoAqdVB+x0sVr
99l9rPi6hzzqwHUoX+4VtMmQpbygSwPOb8+0bnpWj+YKjlx4s3uyzE/YmkJ/ZiNOV21Aq6WLknSI
G+3WZAbxjfUf7N7x2ON+L1VX64EEMA6VoMSTZfyXol7I3RP7Jg4O1Jn69To3lgXXCBPHLeI3xD26
xtHb8EC1ATKJ1IY6iilGl6TnObLtW3I/LYk/lutrUKHNHEr1hfzEHHDey1kDT++jaLpiEW1jhxpo
nuzTRDfs7q9qwM8UV2ujTgbAWx9Qtgrb9WQRPzPl13Z9zKu2mmSzlPk0mLEtk6Ro0ilbrP29y8Fm
FtGmBtidV259yMckFTG1xv4Jnsh/cqnGYhtLzozIe77HdOxfOCWIzFj3HmyeIopIzqwrJXznbb/R
8s1cOZqKtcSLwdEYDB7WwB1EoPGxwz9YrLL7PrgoWwZjK02myYwu+sV5mO4zeXupxBiezQ/b7mQ0
C+Hyain+7K28W4YMgkpurSJGkSJktjQKUJzVor3wnCE3dCz+9ms83CC/JbosTH8zDn/HyBeVoTb1
0hJkfcafV27xajWfz7HvA8rN6Mj7JhcDlf5tWrbKd5PFQsF8H4jg2FR2Ngk1/eaNyPXMP8Schsbb
kgwGr7o1+nWsYK5ehQCI2x/LiweyNLCcp3v9k3Nocxba4GHHUftNDzsJj/G3KsrTuEV3SgmLQs7y
mTLX7lufLT676NZCzwA/KOpcyI8vEOlwmJquSqiwTO78x1Ywrshflp5RLctKMl+eZHD3TqgPSZ6U
KeNESkC8rdhvYPTY94BbrAvFsEnuHfeILye8HgVzckzKZUjggeO+QbUzYEnko7gvVKoccnPrGLZB
RN44nEPG5Ysz9mhoJpSN0pRKeRmhK0nRxFbyF3QCHkg26//NIaL6twhx50UT8amdMZp4jZ+TLIYO
pWCgf+1GaoHArYuJVEX+Hg4rL7zAdc/44+jVEW+UAL3eC5QtdWC22vIABNN+nAVs41Go8G1EnxTP
YGphfQGWyT5W2qS1lkEWSgqU0+uOtxR0/i+H04utxh4Z5B32u/kLAULsKBWdNAerWORXu0mpnkK6
m4GwPsprsspTDtpTSGeQ4irtQqXN9LkhbfDSAfkjB/v3BtwBBd3ZlkerGEucAH+xRWQUvhjnzXV1
JgArwSqDX+AuCWlcdd5q5+aRkNHKvJFcZX0+IOHLHTKdfGZjKzetg+KuYK6MgX08bSNlgGFSodSY
eDHMPvXqSCicQtgFmwtMfTjWKTpPBGpT3VWv6fl34H4Dpel7xEwsJj34OLpghvrzRfY/hWL+i1ur
dpv8yF6WuAyVWZh2AB6TKoMgd8Fu4bwOOpnAmV8K/plSMjZv8roGwAVxGbFRlsPOHb+xoW6G5BBO
u/IQJ6eLF98zSHJshkl/b7J9rwXNRhMb7sSrRXXZ/7jDTMFdxL+SL5NwfRmTSYtnOTsitX/x7KR/
t345NMrggaz7lKKmtYXstV58Jilitj00HnrAjcceg/qnw4A6YTM5F0AYYHuT+bc/7xdGdCEL5zcd
0YVFUaSrr22lQ6dJ1SFTsQa3J2xa1hr9lS0XRAENHNCp0uWX9jUm1P2BvvLaW4z803TCn9GGpHwT
bzOJhYBQP+ZTfQonGdUgvvS5QmcCEMQ65K9fuDcEeHEUJI0nfkAUqeR/NtKVZCmNOASZEm6SUfD0
lRNBholUA8Sfiu/cumN0TvK2vd8tJnNBiyHa9hMMFToJR2fgsA+xatopshMd+29kjhF2KNXLf4Xe
Bu8ccvot+dVKHXoUDGvOCzo3K1wf3cTphqk9BB8MkpDS+s2SV3jh8bmR/CJQUQjdjIwPBcbPKk7T
BwviFaf8DJJr64bttBatNdIoVkwVfC2YJKWY8XTNK8pJe2sCtHz8rebkV4oVMAk9tGfNz4g8KcOX
Vj5cPCkFbpNw+dztitzoAiU3vC3dF5JOnEWtDp4r8xL+4BlLBXZW6yCzl26GPPj327WL2kdHtNHU
2lhYqTq7u2aR/9C0SK3v3F5mkOw+1TOfLZMDyX7GkXncqv4Qe8NEEmeLQDnj6YVBFdZOSYjI9SOo
KjMhhJo31zbU1+NAwuH2HIacWnK5ZRxdyTgTGn92nUF+d2rbvZN1hkwHGUMKNQ671IzeCa4y9KHG
IokxnrGhW8LYEt38NLVA00MPOhnmuUBsrKYevDtyMOtkIvMsUpp1LWcT6daTmmZI34t+hSKZDQ4L
sggqbtpT4p7lL2U+mG5iH1HW/U2ZYShfqpPIZ+jxCv0hBKoUwzIQshxRow0C0O5ON0fVZYafEN7W
PC+8bznwIOcP6rxfFq06NRou1hd+Xskm5rAOFYUFb2ptL7nR9QeekzhkOUM1SN75+y4pVid9Cv7B
eKq9jpCbJ9jh6+IcKUYUmwvlBNO8GVQTJdqWlEM18Ip8ashE8lnfBKJ4HCzCC7QihjcZS0cKc4l4
igLDyzNDcGXu6smjKsesCJb9LmUrcX27dwoWqhNvIqxobt0LyVb5JoHBGrigmOfnetbhGgx/hgIs
Y69isd+Eo+++VWX2fzcsKCZ1B6M+A3BUSUoPsS7Dbadz+a+nHET600pgR49jMfW8qbf5wGQzkoYC
ZHWETsdozNfIt/S9/xonr4vP2KS3DMbPcZTc+sh89otHyXLWbYneSxESdBkev4ik1EOPtWA6ascv
0VpiR/e01QDuNxkkG/f33vf9xrBRpEGLILmzf+HmX+G0ufCw5HwfrK8mJEYz/5aFCG1K9IXC8af0
cQ3vinA8Z6EfzEGd05XC6o2jN/HS7PaGQdNARW32144koxRLcx8m5xDrP80lnLNTCN1EcztbApjn
v4btvNe+EgFvCOvpqXJzWFXMn7J862VV4+fcly2viItF8+ebNyKdW6zj+who6rP6GzkaSZMHoQYK
ngq2DWBrL/NnUglc5wW7Jr4BFABLF4tKsQYW00i8FAfEljFVGl6osIAe8Ur40aJ+rT1oQeKy4kih
avgehyU4tlwZjOkYCoqUrqiLbMg0E8PfkVu25TpeHOVKNzApwUuA8R4Ho/lDPHAasr439vjV9Ff0
ZpcC8FG5gmQk0TPKSz/WHt5axW4wZvgfcu7j4mC/TiJpauZ6/dm8tj9Ui62bIHdprp0gUrz8c4nw
1FPmZFWif3lDmAwlysXJ02gSS7N2jmCi65XJXh/YbHGa+PG6llgqS70cBK8E7Xs8OqC4W4w/YTaM
Fy/S0hPlgRM8QDsIDt1iQmqKXxU0VuWzkXx9MiBVoyl6wV4g2b5reT1OBCJIiRndlk47Pn7UAez0
AwPQUAhpHI312Jf07DHeHWYLSJrZlsJ5nv8UrBgdojFHv0Di+5FG976HmBlVPupMzc7w9n2GOeKR
sA4/T5QYzQFKlGnQ3Chyge6K0jO7bswfSBZ3lu7SZjUDV4nGZilUUYg3fld5JtWcCJ2iepVzPN+1
MAsgxvBBZZccNk0gBGV+SgpHJrguWTke73TEknKysLy47tdFBERxzy/tXBLsdcyz2MKIZChF3cJe
6m6y9VImf5xNT67jPu9aN7LwztijQ5YwfsPY/HA3yr0YR3/MKRHLeHGYga3KZaQdP/wx0uXi2S7j
xBm2WV/U7ltByRTgoJsuChO1nBI+BZ2qW5g5vY65wtcQOuBXh6uI73MFHVnjFUDi9bWOqqHW944l
zZocHU2giuYpkRCpJTmcTPCVmTs22NDcgJNumhZUFTiVBIjpJlN+fPbukhsil/K8u03uVFovQ+nw
uc0bH2axr+d7G6N+HAdSMRsf9MHTO+bkmbdg7VfnLg1SEONFFBz84AExYsRVPGGx6bVSw8T00W4l
WIDK0a8to/EAa0tciD5TQzG/oAF7H3JWf7tJn6eAtH2ebp7qzzPd9kmSa2NdhJU/toYG900bPhKq
2Fvzxvd7ZgChLHYcxzs0r3wO2NFRgwrH1B3diwWHTMpBAvmYiN5/JsXt1LY/vGNW0dCh3yE9y3kT
hwDqKQ9jMjvNjDCDqrCS2jBKufAmO+wzpmIWxyL8iPW2ar4Z1W9ZkdmazN60JlngnxYF/7xzFuRt
0W2FVaoBG41WeeS17E04aiVw1sFVwJR8V6Gj05SmruanIqcMq3jJSdL0OWdpfyLDm46FQt6q8G78
Ud90vBW7643+wkS0ZcaNS2jr/5EoDQytVJdtknR9PIRGV+mLZ6UfX8l6Aaf+sBtlMGdpup8PSHM9
32/uo3ZZ202P3ak4qVBnpQk1I0lSm3QTmnonUkaKZ5NWFqgbXd3EsFQldL3P78Ad6EMocYEagDku
4ZwrNBrzQSSwr467b7Uq3qDNwfZ+t1jW4NM3WtgbU3zyy0jzXp0RwAv7qxD4awpHfXM4qG3Zyz+N
fFd08j4qXbhL4OLL9ozFZQlDZUrw1GYja/AD2Zs8ldoqtJrzNDCmTVjaQuDdwrr4Ivt90LzJOIpT
n55VRb/+nUwGo21PhacKysBj5La9o9KXzWMmMnw3F+rKeDCfiCnDn9Fo2/thuCSCl27lucxWTF5w
vcCkCFvCU0G8ajjNmPtbKyc029837dpM17vHJtTDApc2oc5lIS2emWHkhhTRj2SYEhHg8dB/u86M
f/XXQNIyu6mOBm/x6G8bFa80oOzHdBwssFFKnCV8zqyR9Y0+FrNCvT562be7Xa3Fy28i7HYZUX4e
7dMwXhQmmxPWUBkYAQNHpZGWj1JEI6oepuymydwb5PrF44jrhsE7K8ft4Mwp11GQnVQVcEg6FmQc
e4xiYtVYXIS0DSqUWfM8nnVedBl+PTjCymjBO5D+vRuE+vcDlip/G3hcuGF4hWBaAAL+I/u4WkBo
RslOcSw3ts40yGlbTsGSKfiPCK2rEjrRv5BM5mRLB0oi8dDoEGxS/15BmybqBRKRpllu9YFshU98
8YMVC5E840hfAsebuqc4cGSTLulYZ8KXEkFwH2SDx5/2cQ0kT35JMKXUrtjxpWw/nc6S/QT6WksN
Eyqrq1v3RmAhTBSMs5OUvKoBQbIjWO25s6AwhAmj3tnvA0MkgWO0gFk+ONrDY2a6KRKt1UxqQ06E
hZ7YQVRNNfBnpgZQHX4RVqjCXh6y1LTzjX690VDYXZGXe+2je53kjlmqQsD0328wNZHF2wT7/AZd
bGZFmXpCAE+RtCkiKduaYQkI949scNKJqkepUHHIKDdTQZWD2uWUmEIef+1JYWWNV/hJ997cxAiM
4Kw+yLn8r3YEwUbS+D9/ucIgYYFi21pIvtxfiDYlug4TMqHLOhn8dj2EJ7qb9OhQ+efr3JyqTAIZ
VlpnsXa3ID6PRZoE+bifUEUO5XCMVm8GmSqqrv7Q84KIS7/4CoJwzSyEygWN6lt+D/GdEKD24svt
Fe4mNWX95O4D4UdMEsNqJNXJ32g8Z3wcfs1EzArBgWaxS8J185jHMdu+Ah7ieDEpNkXBGAuKvpda
KLJRI53jRGYEmUQAESvPKChP20GQXA2J+J23ygkHcTFysBSWmnyLo5bzpxNTYgV/gEeVSCINCVO8
BhdTC6OER3cwTpWex4fTgyrTFoHtxN8bC7/GDtqYps9c6G0OuV/si9haQ/yBQ47Nmp0awe5sTW2I
E2ZsAu/+ISCAGOp3hd5nC2DIiAoxXlQ5M/QUOALBq5YuZVogTDh9RUL4Voa+1/hgt19tVi/wYZI6
eyf7y80CAC8t1pVFUerqKrMxdZwaJCxEZdm8keOiHs4HiP8f0b9d3IHlmjBq5zmEFDN9SGCZUTQp
tjwOVL0tEBAteBHp1uQ40q1ZaSa5jZQ2dN2i4+7pub8bWouqXtL5250PEKJxi9hE+21whcFWEC4P
r8d5o2zraifq6D37sXXzKdakvZBwkdewz8Xi0kp7T1M2RjSJQiNav02T4omxVDydPGKcYMiJnqut
kPA/2za0TvNWLhsawpZdUyX+rKuqyxiLPKx4GxVZpOJcWlAtoBToMOe0f0/HRtfTmK0S4PdWPqjn
fqSLUmFJ0QE5Hta6MZni197wcg1P+CNY3I8bgbYMM4NrECjCuw6mRFqC7d5656btunHPWSHEl9CF
iX+sW42mmeTth7OGx0FPM7R7fe11gR2CUHUzbjPLIwc10gDsxjv6UgKk1tEwgp3lR6qjeVvZlxdY
7c0nFEN5ZDOv3OBFiJddm0zsQyYT5Vvc3Dfb+iMALd8IfARUOWrcGy35b0I9PZV8IiwvInneHBjG
TN1nKraqFiXfDVIPPKf/jcLGNIMjXqo0Oq7EVohpf8+LrWvZIyKKlmyWUA1zF0fgfcW+KIITjQW7
cJ0mt6P/kIB50Rr4GSJC3XUamevNFNnsRW6P64ZoNu/AIS1wUwWt2R2BOFJUXJAGDikFfItW6+Rn
95n67LJbvM7PL95BRjBdT3/2OGVuo/DqIpgTxSxhVPeuQUpM2O2MJ4o+8sLY0ldVmnlt0px9E6fY
OGPu41e91hDzU/43esOA6a90QvX9Q93LrtD2ZmskvpEJ7MQz3SPLgyvTW5HFgAJIzUJh35Rh1aGD
43CtCPKL5iLi0J36IIhOIIdxO7pgdmcOh0V4yBIDjyKqemwj1suZTNEsx7sY4o+Bmgcp4V8mT4F2
LcpQQyX7d1SmUiGowGTRekEsdsCNgo9Ls0Fs/PSAGVIQGnAlLcEFAbNsNQk7lJhohOgGVk6benTK
Jyx2ZVbaDh2vgQkwLAqN36k+YmzjyuIYHVhptVW4LHqfl+LmgU9Jv0vzl7Om5VgseH43dvO2Jk8L
bT4YHpLbHZxJ2gbR376ObQnb0tmb6HNHqjg6rqOYkGwXCbJK5d3HxOWAhbQcGSrFxQ0QJrsjRpFs
StgqPJygZ1cLruDpHseX9D2WPL1m3UCNha8IAM2ejZerfuUj4FluoRvedP1duU3OLBShw6BG8juP
7nGg9oPMzqNwVY4pS4Xlf5IKsL1eSJCDQmHJuZIhMvBAZ9TkKh3XGjte2dySvaGtHFqgW0cJdyQM
xNDM0X9ydERRgKxGQCXwRcJ4maD9xFaR0i00WGg0pTsSIOydyQSFXRaSS7/QvJodWZ0xQBd7+VuM
aF+FNHsHa3zc+btaVhVQB1WiEeGbpZTUjRDZ9jtA9U2sUq3I76YIwX7VlO/CmnEfR4iGVCQoaTF3
4Zv3x+w1dXL0aGPtPeQvhWRXpClbeHV/U72SJMzHUh+bSKyupzfdLA9gkNefL6bBIZpmzeHsoDZv
0ldBdNJt94QGAdYM11sDZrpbkpEYM3Zp4EzQn/6VOVbQsEikEUU+jBGf500rNJ1qjcrdkES93ZDQ
F97xdu7aSoJe1r1X9Rj2tJRx2ngcd/Eccu3wBlUSkUNFDlte/JSYZ+dIbxCICagXqQbZF8epx9Eo
gNmHRczBQDUcFVX2KSxd+wcMcj/4Qw0gGc8fczjOtqm36plPIbe/j0SEDh2okz3ldzCIhr+8RRt4
hqax9BoVN92reQWk3MP2KGHbkctRSjNX6KfC2xxqhMenDhc979KSJkiAxO329aQYxqzlhIGVJQA/
STbf0gSDhRp1m2OG0M7xpYXeIGEpGAWbbOJKBdLApv2QwYaqPSNjIar7sR1Q8RZWiPmOwoWS4ipG
byvXHdzgv3n/w9O41+M4nka9MXZ4p562lXIvkkI8yWNmRKGF41PDWbhj+LK7QN4yBXl+kx+0exr2
RRl/uPYZDQmvPRGumlF2QPvIUPmyifXSJy3Eybvmjffcgi6VNZsc/TYI2lGX/UREacOnvb01kbbf
nQ0Ut50wp3BSxg8vlx7ORhRfC1N6MnX9+Z2LqRz1eZqqY+RynajoXwCl/4X001WdsH9XxiZEvYga
2cqHxnYXyep559y5sbtemmGBi24j+GaMlMaQSHvFwDb4vzvqRhVKL0kQ6uDucBmtiOQEdgR2g9po
rMbRp5q4jluff6rX4ivMFpG9Iqpmjqd6MGQorU9CrxzCAWRwlMx7ahXhMEvBgVAWQzyEWYoTUAnX
Vk8dyu/+XeAECsqoLwhSAe40rb9skkfkMrVyVoPb25CBDco6oNzzvjraC5dCZhmZD9KHZbuncCd/
aare26Ms/y5Esk0RF4n7x4Nnc5Z/SJcnRbEtBlsl6wYhFvZPdkxms3msr2rUKF6RmL98PnMdu8AZ
DVHWS+rc5ULAqDPKL4fpmN1u4REymdxQj1BZK8PhM01/tIp5tbupsWcbBW0AStP0JPJmoZzHMjzt
QIe6ncx6+CzrAh427e8jz/jwWnSSd9TiK9Ezb+SdWLMwZOw3YCPlNxmkXj6xkG1zfPnYiXKstdBo
4jvpR1oMRImGupL/egrHL2H8H6fjrK/wpL8dJOkqmCR69TE8o2yyGWfKSrsjQNpBLJHoiz4/ecUm
XVzCYmndnUNGDmqd9dC1u7fbEbEIh8XFqzmYbUnM8bf+SpOqrvfHbUmN+ffoag6YKIrFWIRzO6G9
45lzlXLQ1byt8uL6mbrGbbS1Q5FQj6dRKtmqgx6tsGoa14c6VzoPlBrrAOQzAL236575Hfr+1Yhw
BquFJ/Vb7wMeEejeGVzFBy4dk1rBTTjORsdKVzA9iNDqsDVfkTurKw+tr4PqEJN2fQJe3FMBf8AS
EZLlVOIGWf4GretZlbeDRKuPFEgMZ8gW2SUePT2QjGE7ajyCxqzXg5RVlHopT4mwVTme/Zwna+z0
DdelE/3A8lrfhrg/tIbKnQzCuy0Q9OS+OeRnQ3Aci45LgLXVC5B00eOIeYutG1Q99DoIHy7do6Re
7vJBpSeMbzg/kIjbSEaHcUYD0uIMC9aHkFsr6PUVhJibeNmPmbSbVQ/meMhZcEqOeQLPX13ocD2h
QOnwh5tPgEhnNUAIMO0G607Zv1NCAuKoa7sWfwKV1is3yGkhogdBoqYFeTr6xqlWpoRccfaqV0DV
r1GjatxJMASsS19cBIKJ5VnTxoJZceHzMSIudao6NjYQ6S4MGCyECk96BMnWhtvPlgO5362hvE1S
sI2ZKxF2dxvFY1X9BGX0rl2i0SK4UFuZjxywBq+ChNRmaI56ENxgp4N8ghuW5HYZ11ATRy3/Vu1H
8eBfYK0VolBYVZmiH96QAIJfLPHC5lB1n3un5QUzEGAWPqeykWiZ+1jcX+4IpAJU+axPgxChGUik
t+82tbAePLOcemayA2dW/S2xAlPpMIullDZsqde8tZsz8qymCIJeuNxOU52E//zaCm88TX8qHq0p
muV6T/9Nmy3QRXSugdFKUIKNNqgP9SMGT+B3BhdewNMpxeG8o0VtnO0iqRR5zHLduM9ovnkNIft9
J4sbMW+ag8qZ1FjYe7Ulcb3FRM5AG+QACkuCySk48ft1RST3QGgjwI+ePvR6WFn0fNNRKiQJLXOz
FDzLvQg3mDJPtRNQ/RHCua0Q9GkODXhrtQ9hdvWMTSklk4sknYqNqAK7SFAlL4wapCd66knn/Lpu
p1oSKvJCYYbiVuHsj9shKFcE7GsdJICMVJSVHtsgJj6MpJVR3IS/Q8Xlr9mKnxzeq7+x6GueSNLM
WUYUHYAXBr+utMcXu1D/15GOA0DXD1vpH0YtvxALT4UfYK3FTivIkdrc/ckcFrAw2zlsyK0DA/X+
MA7BziTYiNIB/higgQT/fQGphH1/QkYrVuKh2XHrFDrSk/q4qu1psWOjiV662vCG1ggfj09AFlrw
6T4AHToqzLHRJUsr7nfaI2qsf6uNE0ZvT58u78QvO4eRBgZqlP8i7cOgEOPiDkYNCiqTHa9gW4OA
qjvmy8ELSA5u8Uph4pjYPE3fb9qgfXqiIUajT6lIO4p4xXiX0oDcQUVqnY/sWudAjV+UhVR4WV5O
bGzJEioLUN4VRhYNbQWcdjoCBKA7aIDtfMvwnD8hlahmZgaIDOVA04E4XV5TioU/I3ejiF9AZF+s
EfkIcNZw/ul2pZQAz1B+HojEB5H5F9bSJRujLT/rGMH8QJv3Vh0SH3lOT1jJfRF6+5SOMMiqSuxz
F0B2M3HOK8g5qz5p+TiPVbWOYPFUD9+pMIT6GydY4llhb0ZsAx0DXh4zabQVVEPf0YDmcEq4i+XX
gkfsw3gHqy95157/1Mh2DUrUnTK6W9Y0NfmIbhcIwx8KsZupSpVLqt+0n1tHqfnQCvZADF8l1HpN
dctKUxLB5T/G9QNsLGazfdjqY+oFLcyvq3Psff+D6U+wJKSjnEnIOKBTz+TW3b0FcffuQmNInyJQ
yF04mcp1+KC1EoyDCtKbjutkkraLVVBF0MtbFNfxrJzdFxqG80NyyAus4NWqty5jJKIzlwb/W5c/
YpsxFIJhl+x6htGhSkACNy/clXexgbhxcmsurTmaMRyWevYDBC1MhsjmROegFWHJTxzsHcux6SaB
Smza7ONMs4g278kVSbtV8EK7npWRzpmqX4XDs2zK490MK7eNw2lkJ9/YszbL65KsBKa0UxsdtM+G
K9bvQ9RXV/BYV7puEKKpcbEJwSYHkL9aK/17EIGmWkpA2t67ZnTL2Mm+fAuPHSMnz+YKQSVkT3Bb
XjMs1GDu64g6gYxdpSY0z+siU99sWIW/bdBbkHmZJfrIw+N3EI1QO/nHku7GooBfaXpIIcZna3zM
Ano6XSCCGo/tx1HpUYqN5gILnPlML55TRj0NXG/P0XcUcpfXDcbKwfYIIW3wDk3yDZZ3S0YcSUub
t9/KQ3HusRM/nwvf6lOeTNUHaBGGc8NWBX/zHxdDO2Ey1Bxik+j6M8b5C8EZN4y5Ct3Ui8Xh6Znf
7r9BbenUJCHiY7Nf5B5uqFSL++VYRjPrPwsOxeAu/r6zwcW05Lzs1T6GtEWgrpPAsLX6ZzH3N1k6
MO7zXgtUG6VEBSxvO6yH65GGW1js0LZn3ffeX9rRxjd7Hb73vLC0R5z5QlCDBUaRF+qlCsTxYUNi
0cloTlWrFfG8Utm8xCs+06L3hACYRsZ4VY4lly4FbwaulI5Fviz6qYaa5007pp+5di8Lo6sE5AEp
vbVzDgNfXZwpd7qWjcaVwdg+Ynk5ILN8fZXT9YX8snl4uGO4075TZr5jVlYiiIyr0PAsA4yYX03o
ItqDpMxcalOJdWiqnNa8bSSfJKgSg6NaX2ncxMJLyp399QYjKK4oSHu0vUwD5lv8r+o7DVxuIC+g
MjI+D4HfZFtzXvQZ7BN3tTQcDNGsEf1qQauBU4HIfCxpClDuXWVFRPJTSNN8MJCg7S2DVDqPB6yW
X80jSeVChHNxaSpemTz4u+L2D/McX46NsqlStcIjV2QlmSqtGFgTTBQ6qv3M7hsr5eYUXXl6mCrN
iW+aAN0ELyhieqmAF/qRqs0wKb2mIzWHCA/IestuL+/6TBppOTwYOMrpRs7X8stUzsmNS/Si2Dxa
/pEMn+Xw8R1AH+oshrwKz6Z52KlTabgdNdxFNkThihAN26XV/7p2RiGo9Mptdyi7PTYLH/7jfMMk
CpI2Gbw2iIMO4ixFKPJ16J0M04HI2kwa7Pk/0ZLDllY5n0slGucX4xAphIT4urb3MzWmTCi6adQ/
Tb5vudeHgNOf8+BDhGpPWJDPeBdmL44wYSJQ8OIDaFVDaqwp9N7S6izA1Gcs051gYbQAtLKa7Tcp
7aIlxxaZTv5WeLUTklJpt0gmgVk/Yg42bopOpjf8A6aRI+90esue91o/opoM9vGQSsbIs9jdCErf
xnR+Pr7Px0aiSRSZNa2Krm6gILy1smdY1Y/5g0qaGg6BqI/030cQPDPHWJTZvHpProsOttXJL4iq
oE+NswBi47d5D61cwqhOFT02uHgOk/iHyM93pWnfNowPCt7eeMcz0W0SREoTIbJLN+ZE3SSjXF1b
7WeHKp6iQeIGltoSDCWJ/RIWrJMha0oPjHSeDy+TwrSeW/9jGoi/tAld8UWcE8P4Ibt+BvVi3c/Q
c4GMMChtlLznn/UOnTLOvBfpKDYewmxtGqj0TGdFqsvy7uNTMKNOCHR9axWJ/TvcAL7VG7eGCf/v
0jOuYrvt5DiaSKWHmgZvJwtWtiYQjluDX9EMvgR6V7QI5ha5/hEZzLdw82wi9P0g1ZLbXkTHJCDm
9asvEw7nhw9vY/yvHDqGDiSlED5LRFyhH4KPrJn6RAOPP0S88urGHSeoINc/0ocFtHw1Tnj4P4qX
JCcGXw4ssjyNM0f6egT/sx26LEfaoyBQYaqtPtypqsn8ypj6p0rYD49eIGZyoCIFsAcvJVdEDWih
SZxqbVZnaUboTqX/t85KXxpLAsE4SBi/R6wTw8imx1SVMiZQkdOf4C3qkllZs2usq4FCoILVnnoO
P1yv9tDJ3vJYP5BvIdX9tBq02WsYZaLRIwnnR4+PPbjrlzttfTeMIHAHFTPspLi7cRetw8aYTgU1
oUGLte3pf6V/9WZnPCnObpof5MuFyqGVRIwIAJAYYfUBX4Pm4apGSOROGVdBt7+MqHt+aLr/SEcw
ZFxsVJar4gFc3RpE8XRAZ+gGGt9o89cc76fIcTR22+GnBZ1R1t6wUK+7l9yKthjv0savqPZWQABb
PMiMt9IvnISuOhBvTL+SwyJ1zYHYNHQKVBJI+RT8DueHAYXFwXrUjBQmBdkGWzFCHa1liod/Cnyu
Ci4k8U9wQ7hib4DFPKCPJbQbL66Y7EpBoLpqpJ0Bdzes2OSEE2eOeBNoBY7whZkoWJFp3Bzl1f/F
nJd8lKBnBWVjRwKfWwDMEcmPhZ3+QBEiyrWq38F6/RPbuG+qva0qeaOhBLYgImGsf7TuSwLwwD4t
szd9F0q9biazwUHIMAYfhL6ueWYwFQ5oX7HXPTgbkjv91YPfVxneaegc1Zy1LaTGlCETG90p1Np7
OOQrWSD0hXeRCTok4W7jfj8vUraX5ZR8VsXLy+1MxR49hcZuoklgNSHH7kEGED4lMkLE+KywTmkI
r4sWJ3Wf3hG+qyZ4bpG8qHfC7tIvQNeyAprkS7MjUksQCe+il9iO3XpCKpYOglr9ILstpxE+D+jH
SmcIuoBtaPQ1/uDNsu+Enjs/uCERuJ6xtGNRZh6mCXdd1OFFC1ajAch3C5oniQe+vejuhuFbtzRS
kSyDOWcp7Cb0ZHGO/93S7CaFE1z6Pnh47oeAUDiMhx9pC/WTwUksFFeM3Xz7QD/HF5Ok5nQEkI1/
p+TAEXGOIwJrONBIPbOFNJxH86MHcaN5PE6aCjwVrA/vqRk2YUlwx6RV/2NJ15V+ChkSPvxBiAon
rgdNlU12kLSWigBb9b5p19R5DDv9pk6PGZOUwzWw0pZA4lfJjiQcuzzIYcvhwpiIejgEihR9IRod
FZabi0WnJj3yZU8FZwJYGa8EdkXDFVHhJ6XdIYIE/UNJAKPzWFIvLPNq+p6QROchtfzS+07IFtzs
FaJuW3Awch3cgPBt/gkC1K+7FEl4IvqM+Cmo2k7/42aOsV79kPZOx6cdVVnt6iOF4tV8CMcPjC7e
Jwpt0AAufRt084y880qzXzhR5glS4yiK91FtkMOSIimCqE7fmPe1NuxE4/lint4lG/DD4PlVUAsT
ElcTTkjrMN+M2Xu2MhiETzNtr0luyZBlTZzeBb/vJXQbnawjaYhF5FDJKaLBAtMZ3OQqF0eeer+U
BFkwgwm1IB0qWyhl/E3CBWlE/BNJ8LytSSvHqQKLPdW8P7K5DBc7D+Q5b0SZ4axx8XxMlNrp8f06
KYHdFvcnidzJyGyMZhjyaGvkLnrJ9cNBbzTCLW8FSWIu1XVKiFQXW8lWXuggCTWHkzagcLl1Ne2B
WBz49vrWyBOrxHFbMaBRBxt/FWSiTMle2xYuwoTKlHi3ifbeJ57hS1SkGQm4hJOUWwbM99ifDYkA
OH9fpoCDVFhrt/X9mzZ8EHOgimaIUMbg6n5Vi11fH5yzkTO5+QsXaQt8AAbrw8Uz/6K5iduN4/8h
BUW+K+PA04Nr72HP/ElXA7yQ0pWHNUT/Mt36qY7mSy15RNCgKuq5L0lEu7dX4k3L3SSHRs6FxN72
xGKLIrV/kFhL26mlJtoTa724GriuQs+J1f++aQawj/+5fIcLoigcy7LlpcJb5yubDMWSjIyinZvN
RVmHz4Rvd95xiZzxXbWNyVFeqcTqr55LCoFigXjwS6vod0AG2Sqi835z64CWdtTSswaME01pgTei
7XMRUr54TP2I0tb/neQ7r7gFcd/nr4GGn6myuwlBFtSb4GmYreoJIjmRsrRNRwRmI+8GfFEkAyUY
BOSyIqdy6i1gPOMqIAfdenbGsHuT5iLKKucuJwX79Iy3R0PFjW59DmiIHGmN6B444l5Qa77qYkN4
hFSSxZsFeeihkmml7IZRej3gn0qGe5yC62CK5W7veHoANxnt+ByUBsPscVCMFwAKmz9QgSBvRiYA
mxOxrb254L5G5WSciAx5SlUz0B42JYhWxnvu5zQffhKktkO2K+uxWmve0KzI5VwmV5WQaeRSZk5k
aGXhYwDLY6XN3boUasb6h5GBnzYKmUierVP7TwriTKPDFA/Jc9lNwHRtW9mSHjxwerw9NR3vlBng
eV2WfenGng/dtYuYEceoSpsTp0WRsnAv9+dDV7gcMKDuHrmvnPCmSb2Kr20CvF7h1nNiiq6hQFd1
n3SwfE5N9VGT0EWxnPvgDlkVCPhB54selSnThMdfy+ZWnc9kGGPkiMUlIE3RnJtBorkptzM19Bpq
/qW5AsiNQn8XFc44SeIbXxqTAJLPav2w8z3IDR06ohsZiPQ1Rqa8gDsLhc/arhynH5tFRfsAkQ6I
YVqMhFDwZaQKPB+SzBjtQZqYCRNfJfS0hECoaEZVu8BF848eNf46J3xk0AA2pmg2YY8EHvD8jKyZ
fEsULUe1wsp4pUKyGOppvIqEbcvnPqG+Z/ohV7iz2N8PgkX1jKWPrgEJpHWNyRSeykYJNjyh+HNw
eor3tohO1GTU2tS1ygKF8HeD0XXb24o8Yza2q9dA1lvy7mr+Wh+Q5ZL0/r8wXNNy87FhJrDnPC2I
Dh6YrvdofbcFhJXR40+3HUSEY+MP+nlMhVLZwj+lMWIIMCpInDdTy2fGHhYhLQLE/zetpafhLMqp
orqjhJp9psps0aeAMgCrsiQPZIyNx7AwGTfEYwCZO90lbvMqu5I0ZFWc7/Fmm+e2zvMjmJsoGF/K
5NBckKZ2HckESMrkQaxmrePQ2NNeC5hFQSGfGHBb0VloC9FeHmSoiqtDrM6zKtoNI+PFg8d6z3nR
iZVTMEMTRXooRMVb4JFfhoLmRU2Z81szpbhmr/9umqqZ58K8eZe3LFMVd4ZlIA0hAGtTI/rbMt6v
Ny3soRRt7PAm6sTgCqOsauVmTNmQx7EX0D+og6Ak3qE6gY5jNPYNILzv6Im9VGdciwB/Yi6CxhGc
EPFHZSxFC69M5Kw+WKMjC4PIpWxjzbVy/XHg3Dffx1en6woCuJeVqgzhD/Y09WIDpUZ1SMH/dDTg
/DMjj9ARU4ey34Vw7bvxWzXfvWdO2uUBpoJrxo3ljnu3GcE91ykuJQcKtuwSIf+E4Zo8PWUh/mHd
tjfZ06ANwByEJze5pcAFR62M84shgrvqUMaCFnuY5Usq/Lo0Q2T4wkVXfmroXMRZPRkVcy2H0BGA
ApOTTxMoNPGzv9ndEJt5/N8bzO1L1gyCuZS155ko4IxiEem+ZF4+/O1UEbXRtk5zBoVULCkH+VS/
7icehBmuYGjRcAJmDBQIPT6ERRlhZnYZNh3wc3IHmsVzxfAQMakWV2cOTwcW3tqTncztALl4OspH
3hJOP8+u8MWpeVUiAv9zrte0ON3Lwgd66g0SoTKTYu5iA0CQSTsCre2YDZVkTgEi1izeRi+yBZk4
8ZabPllQft0NstH1VHmhyzs1NmFprI6ZjUvgSJJjUmzMQLP/Bc3/J6cYEdJ5qJHhWV3JTFkqnND2
dR6eh5AK7V/rYcMquVvhecZ1sqDxbxmExp0ELjBfjdET5zp3PZZBLzV0ONjkQnYQi0lhHZf3ZWDX
++gOmOJa2EkSB57ULy8Gu6URae2tgC9CcyNOjk2yX3/a69ZZ4uGKh29PVNfRUgjHALP/cPB+w6xM
b9jrpJvrn4ef4wMTZm20t3WEPAzuMfDuvLgGoMvb62DpliWUw9ewimaexA5e6t/TI5sz5tiGK1a8
b38u5sT2Z3+Jbv6hUzO3RkRFEPtkGkqM0deutWHt0ScbZ28Nb/QN+h1OuJSy0eSDKYSGfMHCLvbv
D3zxDgTjb345K1Hc7p/lwm7bOUBpzf/Epd+rOfP9T+2uVC5+EXbvgBQ6KsOqgPJDHhbIGo4FmM9D
wnLDgBMnVD6tla+nkLg1Wpb9oU9SyHa1LEcZ5HkImbbI+qVJjoVTbjXn8Aez3VT/b7BYJ0LIUjka
WlYtoSJx8K1oLWSnf7bt8XM4yn0LXAtJJY0Ih07CPGWEAERDkTRmCz65Cbm0D3iY6+VDHZe0h1J8
Kk5B12OmmWmHeWgi3hr/zqgK9Mszx0/694W0BUSnFTn5LvyEsYlcAojYboKBr5qua7XuoYzjyyna
9vwImXOSawjWAYRHOVsjYD/ofU+GcJvcj4BarOdYllgGcexRT74Ue1GnscAHkjGg7v3aLOIlnKyG
665A0HpEda6Km5Nq9nRfnPQFpUKT94QfZlotilq+fWxdsC/K22ccMz9bSzQCcOaYDaAEh6OQpCM/
gpJ4K6kYDaeZ5qb8ccDtcEeR+88ipE+U3EZKYl/SNXOz3etjbpRrSccCk0jk6Xo4EeIsf/hO5j/o
BNM76oLyOcUr7v+K+6IJz4v8jdbcyrAQ/6nSFTzdboZAFZc1AvFdP2xZJ0ppWHTzMdwDyitaiWXY
aZPNCgOSd60usM1uUFoXdHWgJox4+wPEgVOkWGk/AInnr0LRrCcnj6GW71WsbVCrjfIYrqVI+4WW
CQh1sgSPLrxnjxykXKZ9uPlOHG/NBe5QWzlYcBzjWq4Fq9ADU1Fta3vP9VRz2LLj+nd1fT3zFAdR
SSbRZBlv5R5W55BPTvAC4O0kSx39AGC86QQ8Q7ETXhLivyOdbuc71FQxdhVCAHYCXRW8XOG+gfFj
1d0Sbze/fLvGC4H8Zak1vW2s/kMLY5AOOg6JEsUSVSZcfP1apSbv+VzoG/6a4pxqhNRfUhOT4INt
E+buItLmoUWTqOmSVXnyZ4ehGfl9A/AAuFc4kfnqTNeDXtGeBinz/gQC8v4CKRchaYOeqtVeq3aG
SI7zcOll727hiMg6vQb0d+TL8UfmE8NB/yMa79Q94rV6BEPsYZvOTt+ZGDAMQWwQ36HT7KbuZigU
BuQJZH6imxtTYa4/lU6h6F7V7G9y3gnQDzcKIqihau3P6BBC2niRFewNTBWcpQ7e6W5KQnv74S1x
3th27Ggg9WBYB1Ml7VvL7Q9w5csMpjUP/JcPmynwm8MdRnFOSWO2cisGk1/A7otA5wKX3SlyzLti
efSxg8+YBgR+Ig5xWX9sCdtI7uq8AFw84+CAVH9S+6AMEj32P7hWbyNqv4dDTLCzxMPvJwFFLOgm
2kceNNpW4GMj4bkAO/kx2NE7YyIsLXTf/U2yE9SNhe4WYQklwOrx95fElehmWNdS6NNnxzgnOb7o
GuHGUfyliHc7ocLdl/0bg5jAAX7idjeXQMf4h0EscQh0TQeX0lz7lz4bSga5sHkeXF7M1oSmzW+S
fF1k+LUVZtzqGSzT+9cel6bffLTBOzfxJySJpdVt7R2Srv0+jGFchSV7TndKQbqMM90U8oVz+A4S
0q4Zd43LP+OegUK97etycWfv5aWFWpy1NOuRyCouKtaHVdIKZ9je7yYb5XwfTAljPJixbM9uqjl6
imtYuQpCLD4IigIk7QYxzoNtOrXrJ1W5iz38o6EsN74aD/Fwbw4S6Vf6bDjQQj+qXsIKQmY7enXQ
xHnFqH/ocI2HYCPdZ6XJ0SmFtDRhGUnSHm64Hl6cp7+YhIORwzKsLmu/Igpio7gK6CUYe6URMKnG
F5f1NmiESQQBvQyhy8LPzqosyJ1NHAmOks/rczFhVSePUMM+MrMB9+Am1hyV1d0tnJibXd0TfaGM
n74ZVisVacV7qjZoAkaQ+nZoEMkibA0NHz7dMC4u2SFa65YZxcxIQSW+O/K6fRFquCuJxJfkp+yL
uBtFT0KXFxXqFzhYqsYAWr4XEnGl4D+IlJNKJ2LrFF3/uDzNAYp67gNJ2VBO+506byPsWqVG4qYT
zrW/x2H5c5vwfX/OrZNNa7pecgmuK3MHE55hmQuwN8UeQ75hRVyNL7wRFM9X1tBkzS792+tSYonN
MZx9om/bjnNFbJJHOwmenghLyG4sJzEhAD1yRtB7VDzz7p65/VEgI3pEk7NydhmsRg9qH8fFl/a2
D2wChLsgK3KC0yji205pQUsNn4/dI6RqVxnxmHqdOPQiAni2aH5D7GbdyApbDPR/0779pRbCxns4
eiIKG+m4hO4GxluNrup7rJta2oSifIJ2NwVRYiBbjof6ubE0vPMaJy9XWVVg7jTifrRJjz8M6Cxy
wstzYrInMBrGWczhb5Ty/o/3CqTvSXfqFMTB5poU04B5vUSs/ao+3KBvrpTUHqOGepHD6RJPzuJm
FfUKhh+sTJyZ8vJ6pnQl8y07Lma2k8XEyE94mP/MiIsy6f48qS/m4DP5DNb5PI+Pve3J672ieful
R0A1MsURUFfIGPEgtk4CE7srrobyoRD3lg459d4uM2biNmoD1MhSRY4fkt8DLVlfSVuZfupDjU5h
eQm8lXDN7b4yDe/KFjGExzNW0tsemXEXrPLkr2GZezmNYDd31xuCb50lYh9fbwhELSOVLzxfnbzH
a96izxDLYdrXHXcgt3C5ZfzA8c8BslxEoYeGDoE/utwCRuuTW+L/DK0hRlaV6T7/W0OeluUNL2CB
43yiDC54qrAcOE6TXOtHF5rP/KKkSJVZ5oYFONX1D0daFVMdmgKwFu3FN2x09oe6mUKTnnwqTk90
pg0+t7E8/SsDiJoEElZZCLAc0QcB5q7XYUBTRPoNK07+hrKjYUexoVteyhm8DwN1po3E5LunmllE
zNYTrhAqYHBRAFjHMyDNn6juQq6mauZunA2OvZsLX5K2Jb5reUVZk6BnnLdHrQ1pMB49jnI/Yekt
xUlcODFnxtedHzGKgf5/2S6EZlS63ZNc+8patL286sFsyAu2A4UPWPCMMUhTVCaaSlsWA+LQSi3x
ciy7r9JlynJRFXJaCbBFjFtQvLhuB0K8dp94wig/TIVIAXesTLHQ1RIcVJpgLq9bQQOmYv7zgI79
b34rjXVzqdvB0BSmhfMaDbOW8UnsnC/65h4bj3Up2Z5AtxKvzkMlQx/Cb/ggMAodi5JcadcZ8Gh6
AE8DO+xM6AZ716q4zw/vmc5R5hDeJ/2T6/roSLkDyWEbLXQqWh5vemzlVH0zluWT69aCvdeQsZ9S
umhPe+YeWaSXsgmEI2J1pl1ITJNCIaw6ZrDjAsBgZ6fRjE6kIMfxHbN5yguOR9oZ0kMyvNf78INr
ULCCJPgfaZU3FVun4go3WeLCwWJmhqYK2MOtsbn3tpU5eF9QXV9VK+y1SmIcDp25zFqZrheKwiva
bZaltrZFasfvA2yak5tYFAfc9oaJJZJJwdxNXkrpi/U5mfzf+PQ/LVsa9mvo56Yfs+c+q+vQb4M7
65lUjjSoOGf06MHSxo8ZUT/2dMXOJ8XyV+12cCs1nlm0oBErcJGD+F0BZPSs7iGRlz8Wl/J8a+IU
sd45xkX2fkFz4RPRkyH9maTSh5LfGmtbLus7hElfSYaQDJl5DxDYv6Pm8fKO+FM3UJu6dIC8P+5u
bQNwWpkMIU2KXXD3oU0Kw29IBTTfCGpqiHBqZU+BrS5mAMeKYBPPNszezZgTKLxjRBIQeCrrfF1Z
WPsdgHUJxt1e2WlU+yZFZykDt7itLtannr/myVyLp4yCLkIi3sZPJu2ggB45RfHYuVXW3c0BR3GD
8DXx27IvWIKUuSzyWXwLTbGsQ9sG7RMoVpoJi+rKppV21gkMFfhmNYStxhre9FpdR5rJTWO3h0Vz
t+T+Vs85x0123EjxxVByqf16uLRIjZ9sz5CQHppaIQQWs8wdUzdEoh5oO1S7FB9SGUxNRXzgSnFs
JrjOFVmOmDyhZyT+WUeHDB8Irv85oSRpxWjA/MOj1gzntRkn06o/QyC5UBXVO26SffcRujwijgzf
piHCnR3iZ9yV/RI5qZTcp7wbwxM2J8W2sEOyX/85jUJkuL5fAW06l6jwZp29e4GtlKvO4W2JFbsY
+wgwkicv9aQJ/J2lEKY7xICdNp15zEDNwktb5bcy53bvkAJPsadusfc7EKMqb/7nEmkpy7ZXjFqr
1rKHIPxgyn2LWVYYdHA6cvnvtVLrMID2SsQO49LMv0hEoLSNtLKNbRXkigiF7WyZ197zLIO1d6D5
N8dtyQPfPNYEfWMiQ5hFM0uMYxKwGgJ5YVVG+QeCJIjp3JqbEC2p8aGMz+sKJo2eiKcA6vYu2oz2
VUGmmr7G0NKiGMAX0cT4mXVsdfVd2Ewz1UjOO35RsWJG8SGvSxgDrFerPjdAi2fAjuk9ACpzA/wt
A9K7mn3jT9O28iUuSZ1nePSD1X2KENgd6aReesDO7kejaarh08BYVo4d2R8GZl14ugwBv2bIFQv7
LwxMz8POHrM27o7iD2UrXzalyi2/GXt8a7HR5839iA+5zINYXYoJn4A/lukCJtEupXloc4LSlQgB
dN/5zi/XBImH5yVCfR5PUe6LzIdgaNDPYqEBZDRZWeWpOx3HtVZBt/MBvVclzs4/cmqd4VfnFdPk
YIWollT4EvGUBRVFkY9ZYnW1/ACsW+AZ5z9ZVi3EvKIRlKVXPGxaL3mF93FfTP9bTdiyNKkrkDL4
7JD/952jezsD4KjQnAuycIMr3c5Wpi/XIGNlHmX6xan8IUcHw4RTQdP9s2WWz4HQSOarId6B3GLY
vQq4qVDMgU8oOGzjpqSn72bgCMq/vwdKVw2121UVTr31R9ew+TlZCpCipwR0dQCetLLgJubHXIKg
K+d+BvL5cjnkba/1DsgK4+sGtPo6zrszhtLetEVD6HSBVTZcs9I6O0Isy8+OiuKg4S3evYzpfx4a
4Wrq7c5cCEKXcMg6RscVSG03shjNVTZt85NH/ziGnzico8B+3KPNKYW+jtGOwU68MfsjhcS9vZlu
3khQ69GUfuXaFHDBEZfOnfxq2ceXt5j6WWJ/3yLYJKawGVhI+fKz+iEaRNKrTS+STrrWMB0fBYKr
Ngk7Hn+7sMUFN9cgHzIjjYkZfNiMcVTAPjoYW8z5c3Mj2gRTOHFvIMj4AOvSxhYdkDjZ7h+bYqf4
lTrfNQcsjBK6HvOW3f1jF4lkRZs8GElR/nsmVQMlPw30+pdsHcH1LexTCBrdRwGGEFH433TygAGk
0jevNYr05lN9HA1vLRQHcuWQ8cLwjsu4rAbmK7+VwW2QcvPHah0OLp/wPOwYJ/khore4HlBMZMQb
zxM7DO+RmBB4St6/aKpNvBb/dh2a0hS4EZpQFXdV/s9Gtwd8wRkPeglGy36o0Jt4JMdR38UDJAOP
siFH4iaA0c71bWUcnwY7+aiHwHbzKgoN6bZibmobIyzDeQeDxT8tx7JCgO0NMgbVEsVJm95k0aYT
Mqloi/PHv0sRv+5zpQ688zw+tG9c/GDssVhingMc/NxPObKXF4JZFpGIW+bCRq3GD3bW0ONJJcYW
2e+K/8HhQTS78j8FTcUgyDBD7AUvzNDDIy82l4AeXigaE/qlZBzcNhETpapxvIUig9qZETCh9FPZ
n4SXxoLwpQbaX2hrCq4Q2GmFn4k9nofTFM10Ap3BwEo56HLtHPLET+EzUO//2CLEcj0P00cLoiws
0Tf7tlwOMvIQOlcJyI02CSO+zUbufLiy5wiWe60BXkmo0Hmt+6b2p/Anum/OfVXrBWiqgmaNgBlu
8CgN9rIEF+yMeVG3MmzHLM1I1ibcA2hjNVEbgc5G+5AuI6YBt3vOGUR+9xMrbMh9d6dY0X9KesQI
HswsmLW4NiAY0K36IY7y04G5A2tf4AFpnjGHH7dj/bA+knFLEkxcn1em5yPHHpose2f1NNQXcicy
S+cMseyRuKSOKjUMZIEDBvPXKbr2MWyCM66qEty34KRRPFWXZJO+2BtwHLg2TB+L8swifWliK/pP
BlghbyLlJC+oZPTHKPYw/koCn73ijdaHJI4vXJoOe2zQOAOlu0jAPUHWKPsGzeo/mvOyh7YsQAIB
x9SWDsRbaDWI1hDja/rfwcNiW3len1183SzBKYIt5y9Ug7FdWhwmohevSVE434bhQgsI4vzsFwH8
gn3h4LlD25mQgsRg0q3SKH2RdtTcxazclqKkinOxJ6PoITnZ1RT7d+wyXl+NnOiSrgZzTCeaPdzt
36230iljxSl+TVoU0m/mrD5Asmw2imN8Z9+nNTZ+XXaUgRMM9Yq+bpK+LdXpvzqKNQud/JsHPx0n
61u5cN9XOqY3QQsHMY2Qp6sp3uRtu4KUtvjLHgWQJLtWOVyi9u77qhvzR9RPcL0D28YkNPewHsFr
JnBiwDi6CkbPGkB7YD4w0mwmyvCeRuZ2SAk5IhBSpHt6/g0Wam4kxMLiD/4DiHJyHA4031HKcFY+
WsUzn5sA2n1i7YJfrE8aDosAjCEicvwa29LMd7/ONUiB4GKFonwe9Vd08c8eLn5qSzzE7HxpEoWq
tgJyD5MtFZM9hcbUBBD3yIR2FJCoS6F7TYKqAHURRAkGAsFFNiYUaFT90pTcsZG/WskkfJYHeJQA
VwqKDtxSjZumClb5UgDDbx+jO4bqHE2UOaG8Me8gQr4vB583ZujV9H1MbfoVvbnbOsQJXBFEu+jn
jwo8ogGsNCpC8YjN0REO8boW2uOFkHVXy67EhNIXWnpnm7NlmP8UhyVSfwrcYUJ2zrNkoacTBgc+
X10MyG0vSVi4TaiyXLxUPLbv9E5Ko6xHg0KdfB/saohy72pMPZwVljXIxRNg9a6hXp8AaqI3BQ7n
ceqggO1lD/B2BBQwots78ECsQkTQNJXrT0/uGTPGpWwfHE7OSiTi5L/ZFwI+/0TLnMVrp0szBXXi
G9vHEz0jh8JEHMz1+i9j8ZoPuAoRY6TvVCVwwm+5kM/z3pZVTD8PeKFM6UmMskhStQjtZom1wVsj
i+xUPuKfBa9IDRVf8ckr5j+oQCgLFeYYy6Y7Ps0bsfubI/dBKrajMrsbCulc3R+bGbFAozFFob+i
9jSKvAXpESeKO2vNGFT6fCJurOReKQgQRNzsYmdfYyjqmeVGY10rmzOpxFZ4YBAhniiqu2cZPuZl
0iRjhtv5+F7f1TaBfhbFmJJpBdOYT0Rg+jZJlzUDQ4GAYq3t8SoVFUjeX3OqcVOWLcKeD97GHO3Y
1+GqpqOSmsmZv+/6Nz64pmJjjJRSAF1olI+GnovxAW8skE8FLYXCWK+jgyVcj2hSVLUY9z4waDEd
ngVfacmXaQrgsXl5ObuE+yAbEPvue9fMZY5peicxSAKuoPO2jalJ8ArE3mdKFhg9vOogOxzJcCmE
ownVQXL2PWeDOk5ADUcmDhHofjcm8BGLgGrDlIL+vEIcboJYUtnbb0HpJLwuimspDWYFztM6ZYvF
BRIzofBC8f+K5qtLNZ+531Sh89GlDUQLDqxeHKxGNqoFjCCBkxASOJ9dC3e+N0Qnxh55jeFxFWKf
aX9HcCkE2X0Bl4lBFV5Yokj4TGwZ7AbJZqqC1V1vFwnLGfyQW1c5Pct78ivYdU11jsVFvSvmIZ/I
/cjiA650i94ymhRH0ovv+vGl6A7aGB7xedS83o9HEYDGwngEBCI5iAfDRrTnw9DFvh/KJD3Sk5LK
E23iVCdWw8Qvvv6D9zQXqpN/qh4dyCxUbqtC28YCwS149jWLb1vga/Ls1vy6Bgus4pee9ky/imND
n2SM6JSCIRUbmqIb7KIJkpyhrkY4PyFAkOObjafjEgOnED8uepbtZOq49ZhRO3/rd1hq9BCi+oyX
D1t7HC30nYuiRWqe/H3dSftp6u+aaCn8Y3jid8RuM3rD39+/O9Il3q80MruM7CC5kgH/lbuj4BYS
dNAcyNqHtbQ4gYT5Naa8sTYGA2QgAwygSfun0ix6veEOZm5tXqViYlTKvLM/5xSQpzWgtDcxwFva
ZwgXTIOTUmrhIQhZpKfAArCu/CeegEloebVO3Z2DFaV9jjaqBzfycunnCIvvaras9YrVbOcz/rBZ
Ao10xr5GbZ6MZGq4mkfCxUekF2uLGLOi6OwcM/mXD6fxiq4OskLVytkazAzNUdF1qQGHAQ36rdp3
5wMQIjtgtUju7c2f7pdmckESDBR3RLICQ+bT3xFSm/WitPC+bsimi7L/HXjGpDRojWxgdzjyF4M/
YY0Q51hURBcz+3wufDH1oN8kj34IFtqoo3hpkm1oKqA+KnY7rXPsOe9cuu1625YLElkoI848kDPB
ADOnNm20rgbY732ROqBVQBWLYbuXFLCPYZB77hCiplgqXz7mneR4baFwsndjRjRnmzJdGmz+D7JN
ZsqQYp3aQNxbdpXdACufWf5rkKj2xUUOr/m0hqazbBUKxk7f8gPm3VabZrWVwv716k8LEHcHP4FQ
TE1g7NRCGSRlZIiIDQ/geKMIZmN4IuTTceHdxYcQmhJz+YcGvgSnZiv9lxnm54BcGAtd4KQ6Qfn6
uPmU0vUpgxKoNgIFaIr4/tVM7bcn4JEWwUnA/4xnC9FbboDEdaCXOErAvPpI8AcRN/2zn4xUMcCx
wg9lbj+mx9ExMgnRz5HtfPdSlc8kJPYsF9qYcWh1QA/63yWZ8Fn/L+YJffjdwYtUsipkO0XEtxXz
6FQfQiAUwQjyLs3MiH8arvOuOq2ojUUXymSDAVKc+doZFkan6/PBH1lOeS4Uohogmq1n4iFPAQWw
JyutiGlSi5DFE9L9s0RKk0i0bm5T4/Evw7NOEQ1s+OqZsZBRhA7gpOL1QDPnv/D+DR+I1OOGhrVq
xoXUVpvcMNRj4c1f4ClSTiEstapt8n9vU65jozT4Q2patuk/BQSAcEkNZoeE0v+6Wqo4xeetswJM
i+vqbp8GKM6kWJcgJfGyNdJjl8gVqMWyfRTPtAHQH0lt0Q3+yp+boD7Q5MP9fjV5piolIL4ievMd
sqG3FGbWRjOJBWfFFuuX5C5iulkU7kFHXCxVeLh1rpbC7OJyoPq1sG+ZNd0RJ+/ev1X/vekG3Wqs
6mmot9Oqh0ekihKzvq09LTKG30Hq+EeXN7Do2cCSsgY858/kmob35RTTS0YBMV8aqeJLYy5AedVl
pz27qgWB7pY2LDvFiOYTkf7Dau1J1PerIAS+BA9TVPwwEdeyZhY0c/tq/w4SYiOIdxGurm88INYp
x2rc06Xia3LA1nJgiAOOiIYldsGjJW3dKK9oIuYukv39W+fE0HFE/liG2dz8wkkXbBXYQNWaHD49
HnIrib0Cz0FTgUmdjPhMOa5xkIMni+XSBml9YUIbmhelBMcaQWSNQeCwBVbHrQ+IKERg6Xn8/Ai5
b4q+NNCDkVGzvYn9BMFisbKFtfOndyn3pKvu83YXszaWABX0jvhuP/1xgpNoN/ZqN27/ik1eRKyK
ZdemxIUZLFsafOQlNcY2SATnpD9+PN/NIoU76kZ0icc4zFX9ZDDAGy6Sz3BtirkuXXzcnh32wgki
MDIR5ZHlzHXI+ad+0QdN1DZONTK10U9BVC+m/5H0MCx/zq3iyqPQ4xWYBczRVWgQjA9mjRP7EQeA
x5Y0iiIDffCzpwV5Bhe1kpfNxyn20MhHtL4M4lM6MMRoRntseZRPFohReG1xSixqR9Edpe+K55of
q5SllKDEjlOFvmIDTGCcyHimyz3JYGipyCmQHyXKqKAiKX3YC+jlMbZi4a3r4WTZ3l13qwrd/+cp
dXq9GjyskU6wIvPWP01bmXHzr+44A5V1c+sro0FQEVL1nD+Bkcc4bLK4gmRWAj81vVvZj40qq+UQ
rLiy0eTyibccF91eL35CaJqQtvNM+fKsdo8PHy0aQZaeM2cjlvIzoPdA5iRSpzpZsXtIr1sVA4Yn
H9NQCaSY2YKiShbkhGodtglg3L/D7w7u2GXhEWO8A0+Z+jWtC1CVSERXVmR9WCg3fIQTbn0+JKVF
Rt9S9zKM+FQ0kM6OvGlUbbByakA8ePGYR/E//JIbcypr5BFpIIrBauhoOcGoaqmrGdxGKOUZkKSL
bUmzgpZsMlf4Bop7h2FJzvtT4aLuJZfzP31CH7udgMO/sQb6brBWifIIjiMzPeUdhc4afMAeBjyz
Gsa289txGUQWiMHxhMyZVL5k3ikzuhryV2C4ALrkiJgTZu8sEzl7OoSeMYHr5pS1dtbfBYOFFbgi
JcRLfu/Mw7Cxy4lX9r0OToJzP1/8Scrj8zOUiXrNMa2mbHagKfRD04fUYgbbqM4aFo1Z3TqmguhH
np2Rklh8PfgzvgbrX392tSNTYevi4QT4kW6vf74hJYM58ZG82jbWhhx1+lOrYrzmSX6CwxjbMokR
X+mQgHGL+RwqubioZZMF52gr4IuEWrk5bOPuRuAsEE9V0uwssPnwXfoWgV5foxSu55wh5e2MCmhh
yM5a5w3mp6z/mP26q4pS34AnEOLcmAlXH2I2tweXgoM9tn2vYnHpgnqcsOe558u6dv7dJNobLe7G
1RwtIAO+ECvaQCbMyoCBq0Md9AS6n2/mqKp7viZxErl9wY3HcIQa6FQnC3iQguh+jN7JS3lgFZxA
CmI2Ow3eWjH0e03TLlyTFPjheJ99WJjNGUo6/+Orbyb3gAFv7SNHiNNLBj0QrgoqRKQ54jKyJ7Ri
NKxtYKTo9TKW2bN3XcdW6yJzVHW1nDMk5cW1+a+PJlQjRPJ1VxzD+Ez/kpI+B9D9syXkipyJVMXJ
m7OW4XKujO5M5gW7bgCnOKzYAFNRjl/XLrcG1VI/q1GZDF7MZSzAEBmqeNh1fP9z8Sj+8wXDdcmo
jbgRq+JcnIGKSvc3AJvs2n1d0P8eODfATw5La70OtOj/cBWONu0TbUXafxUa5groZl1W8pFD/eIc
zGGtn0sq2qzeR3Rt6IzG3yqeH71ofiekqeG5iqKTOr0JJBf49fMO+XFcpnYQgchMQHO8IKP2yg3R
md0x4m+YV9Ixg+LHsIFjd6fZwtDhRgCRvZwvX38lYd+t/swGDTY482Z2RepaOjukihslygXAhPRQ
+QkBnGUeH43oVFklL14v2RepugJue5DEcLZTlLXzuACj3RZvbye7zbEMtTRQhhFig2UWl41fs6R8
+rPJWGEERqs+IINEr8fy1nzxbVyLaSXY8GXXNxAWQL5/5LuMT3213qch4U8fmhsS/LvSHwI98Vy6
DPqWJSI9LPhVSl/9PNBmTIJ+XUo1yfta2IUhPskwbDeqBxQU82ZstxxIgcaeSjUf0JuM5D10xcb+
X6/Ym5RpALX9/QafaRU0uQt//mE+9JTr/mjXjKd/RKgSxliEEKL4JynCFzkIq00SKS/ZyFyBqYz7
iprKPL/lltUipivDKoR6f66dNoT48qLXQhd41b7Na4RyWahGsO1C8u9rbqy9H3YMNF6o4W40N57V
racsKmbcVuPVzDLXjeKGQUxZOGAbOCHi2MkkhlXJfeqmtUWmvkSCbr8dAqitAkWPCXchz2Y5ygij
st5G+H4Z2YUQGEW01GkeAIUfJZZJ21CJ04yH0FmnEgOBcHtRn1xcJg1L48skKzy2U/MlTv+Wwdak
BCl6Fkg+tBgttn+PQwbSjn0xEUZ0gIyo7Qd3DQq8FWsI10CXm5Mp5p5kJAHwkj6I2NHPkprZiGbu
HFVrB0HL1B49RL5yCBGHmdcuE13n4qDXq9CPQPBl3UmTRiW0RlsZQ5kYvRhLUTv7nud60eDnsWpR
nxpgqLTlr86gJs5XG5Z0D2ERL3KmS/ZehP3+sskghtI9SG1VL1wg+2pwG1h5thiIxwjUhGNrXtmM
+MGYKVB/uICT65v4Y09RTds49GRjL11YgKNjA4vIQUYnO4m7ceK0rkOrlqpdd+2Mi1GEaxGn5I6b
XacV/9fuDbXJ3dqQSdV/2kK308joPf9yYAP8XQufmYUgcrM1i60++zJq9Y99Z/xi6bYH/+kvORm0
9gEEZP5eCGEXyl9ptsxuP9CUy+ormh52Lxg+eZgvXMmrkuSM8vQ3kw9GzSjY67p6uu0/YLMcqBnl
4jWnaTojaSFBj6LqNDhIaVh3/CnUYILU3ib3Ssajqp2cyO18axEKXPx4avEplB+L8BmDhZmW8NWJ
CBns+EqmzcPq9dmzGa2slXe+uu3Ho/VXLIfLIibWwircUuJBDYyNsHxrvMvNtmRW2vIz6YM70sI0
fA+CZ/AAzruJfPVc5jyl3Jct5KcZ5Ac7/QP3o3g0+ru+djWRh0JSYWqo6RIku06rVOm1c+dDo5sr
MCmXu+Eqx8tM/Oi94QMqTUc7gzAm+m0W2ii5dVdQ7//knwj+oG6EA7VGngmJQOGc9gAMih5+OpXx
VDfP0t5i0Riof+ZkNq20iwngoxtpycUUF1kh2BsTQ6Rka/hPO3iJV/SC9Hd/DC6b6BATMAXWWFSB
88b5MaAdWyg4oouC2bHQpDd2Avn+4TJWpQUanq/NXhfhe32Xsg6GM7HFzsJBJX6myEdT8X7LnvgE
Hgye/TMPRkTPWbVwUIEghHcGiq1Nu6J7YJfww3k+xuFTtQZpDKQSU8SCKSdpvvbh4VaPnP+8+Yvv
HIQ3wotMLHKnFL6X7QO+WAsDDpJzjPsRpwZnYziiAzZfOWWjqWgNquTnYSDpLleGzCCoFZwsO5Yg
yZQQFKha+mp0NfK3wt3yWLcFG2EUCY8ocu7+3GSaoUHCOqJAts6hXMC1dbkGTZBDK8HtVQXNGbnj
CmE4MX/DZrdoj07Qr8M5hH42hl+BnoFuEnOiq8Duwx+TnueFZX+7UTIANGRacgjIBeyO9TwobbWj
2HfDEcp+L6LeQlLzct8K7X0YQ6dsl63DzxonxM2jVkSAMM+C6BGPwMKBQxE2QNhm59jn7jmy5rRH
lcEyInjS+sElcOq3SeJbErgPqUwILWSPrF8y64+c7eXb17Qg1QcpfXNUbJb2/m/iC3iIU1KGH5kv
OKeQX4LCH4qvdT9WmNUd/x+xPEq0/uDG1kVZwKoNz7DK6U1mg4cyxhZ0V/PNZEwVJ9x3SbRsrvar
A0ivX/FauQLfrb735n7CAJaB9DpetsPOAS61XWoHwoxgppwlyyVrBxCm6A/bixapIk8mYRQ9SYH+
e7xNHd5h44KJ5z0rDK5Ibvu0ZjNFQlUsZQQGPS/a/YVjrI+CtjqR7hV6ZgHbEhPnQnsLM9fx7npr
a0reR5xTXZWZfTUUXA/MNl1V2v2L9137OTImhx06ILA2Vy7jbirxF5T4EJMfr9YesKXvrdjbDFrm
UVRS/rciHXB8ZxgdDXwj0shZPgliCFE0s9MWImUeOuH72xWedLPBsJLcNK0aBHVOTGG/lS5wcsI3
TC7DX6sNipNMgOYwJtb1ZpevGXak77TIxAMNIkbVmycuu9GBVH6PVknF3Wuxj7x0ZcSWnaL4ksb4
pv2cMZy97S5T4Em0kLHJxTttO78F+HjE7Z6tibZCbxrWUk2H36LndSpwwjbCOIS/5MAq+Z+V1IC2
HUaF99G9+JkCriv/Pvc0dzf4i+SLe1QkNNIYJjYu9J8VELe3UP1HkamXN1NPigozqulC/XS2vhcx
N8sp0o+zSBX62ac+t+gTz/9FyKE9LeWKATfRdV4CtYzIg6QiIFWCjREIiRVmvbFPD5obBUygtjyN
UXLCpbdyBxIHbRx6sJirBoSljK4eQTdtr5DHZZ3tQAsyz66dN8c2ES8WisHrWpDzUINBtoyFe3HN
9QFRn3pBoAiCmKxyIcY7FI/2XJQMozAVPbwVVRQhaBqnbn/VnbQ1mv14YHk2fpNuWwfWxtDeZKUq
KK8Gyh7ry1U3zvq+2IAzn/cMzvef1nnQlGh9E5hfHU/bty8lML2ifsBASUGHyiy1q1t+6tsTf7U6
gw/LicbUsnXyyQdoOO01B8X/kQZA4yi6klqX58NCktyyxaLZvZD9iRYSjk5Wbs0IQJvoOTyIa50y
zmi/Fx0rFW3/wKhdetOJQDbQjOSmjj90Mn6Xrv34dmqosc6dS7yMAvUokGZrg21S1tIxwwT5xLav
+dJcyblg6109ThQpGZe7MjnN+NcfnpMLMcF0gvcCv4dzPyR4E/St32/OL0i5xLNEiqz0T95eLtfc
tJnvhE51XScVie68/pu3tZ88cKhtaqYjyoWVgMVrg+/UbHWXgzTo/cLEgpkr9PnsNlrdIYzjSdHM
9I5Y1AR41gLZdT0ieSPDm5WFz0bi9snWtFGQlHMRcS/pAoNJ1lnSQdaUb7HzUd5/a5dJDATE7OxN
qXIYS27U+6KaIeag/tqI8XQ36tc/q36NYtiVeFb1ogrhXvFgSy4R/Ws4ceXulHImwgdlEXCSqAoG
JGlE6bbMicluOWqvDtz/Wb7yADd1Hk3Uyir+K0So2Jq6jst8xJ/aSWevjTDmABKxoU3sF9/lKIyk
5D+1qWIhR1XbaCVoZY3p9o4CR63i8Jwd4YxwC6BEq6g+sE3zpbCRF0uY6/uTToAHlQxN3wuuUCZQ
u8wp6endc16k1RY9XsyklW45VLAIYHB0e1mDEPVlPh1CzlpH6V62UubbwPSBEeJAoie3Cdx8v3Ni
YNa2SgflU29/JyvXNMKQ2eUIjMLWoiYA3vJ+Rp54iQDHwkzAiME+5tMpy04HVpV4EGfqOzyX2RMt
clC4zP593pGh5C2LSDSGR/eSVg2ZokzW4Hj6luo0QdsqmnysLd6pWlRBBhWUaWkZ0oKWkKDDHRmj
hlDIVxXPiSqaUrRkVrQC6ZSPPaWJ9JdOO67Kwn/vg5n8Mjmn8PS1TFqnKCMqfGIcku0qCzp2iH3d
ktck01yajpG1a5UnU47LahpsdekGuZ9X/Gu7uks8e8KoLBu19Qun93Bylua65h8NqMECie7Ynm+k
ejM/Mfj8VzzEPJa4xGpmRM9ErlZNXxZKKyXCfhmovbw/zWXelv1edEjb1G17wTOAkln49AauJ2CW
lIm/xkR8hgXSiIF4jj1OTX8cUUxme7eQ776kiKcINwLvGqugfpllxfZK+RCZV6PDp3oRO4j5EzXO
OXO17EQrpHuUQiuUAwovSFhxbe09toePBhBbDs7pHYeZecGSlrgPowBsGkvuNbE0KxHhwLgfo6EX
mTqcogejx9wpPb3uWhHNvDqyK7kFiw8QWO7E5MqjsQW6rjMMbEC+ImAbQcTrZcmc+ZaJXQNGdgax
T7ZYhHTDk2gfrShutwunQcJOWjyjvS12EiKfktK0XP4abyQUmk7dukIRhp3/D6DnKF6zVcW6QWV0
uuP3XmbJ4UwoJNCyjKXTNpdkEO9VczLGOnqQhTH6gs17G02DZtcm83Ibg3GjZfGM74mSrSjIJjzU
Ma6h8ZldA6BD0d9vK1oQo7/L0RPsdPoAJaW7XC2oJ2PWs0QkVc4LSmNubne0IyqB6CCtJ8lwdBCi
LFud+LLfGvYwxxPY2B6N91OwgT5DArM7Cy5pMqmG+RBIAUtkadALXst0CIFrIfFf8RB091WD6Ina
7poZPOD5ZnjI/sinGuQxaarBYQCIMkOnUnJFN3TS3KzJeobaar1na7Cppt5WxRVGchPXK7d7qkY6
XDkHyrh1kuM8pZnkgbDft0RWtUF+D7JaGwb/WwWu0Ea2E1hPOzbMZ1nKfapa+SxnTd662TX8TeM2
dLw2jA7I/NT1tth3BYtiX/Sm7JvLz/z0ZKq1kk2Mc2/58Qc2CGB9J0C8100a93rIWUgeDYemTJn2
lghBRvMWPqgtCW825IGhrNKY6QMMdo5nDfv+gMipE7vcXhDNqrqeN+gC0RTF0klChSFcxMGtq9K5
OywbHBiJg6PeDrMwApHpMQGPC+wZarvgwzgNup+cdkCSgOAencen2VPmSQz/q69HEXlP66EvZQCh
XCMlorTcuIPlLpvBwGKTEMW9xrz2TaTbzJJj3ENjtPp85PeWuWdzeHfo362MC8siAuAwNVgDD6y5
HXHaTjn/blgJBBdmbEePFxK/LtjeO/QNnhEg52I7Q08qxjZNfiyyXOyQAeOtBeNWoR/adN1M66g0
+pBC0DFkiYkNlZqXrpY6hgsSIywMsjcaYgkB9SojZSuNLFO9IHTeda5KC8hh0tIKCfX+Wme3Xarl
u/PwFPvwPDJPJzGh4vz8EHn6p0LrodXQoGimaMzxaCoflR9pidlscOVmDO/xzNVXtOZ0+Hhrf20y
4l4vpgJPzPBoyr9eXdYenrdYzm5nURaetUcwOyqTjSO96Xv/w8uFQyyI3G6ozRPhFjS/sy+nIRCs
67iQI6ONpYDYo77ylhz1pFXkeVB7pdP5zWg9sVG1QSnGuTH2FaUxtwxFauProdYQKhqs68iRBeVT
Ai6kPTDuKkKDJjMXxLm2/xyftQ1W/azzge0Z62yChq4YqijqAReZM9lhAoVOFPycll5pROKGPE3O
9zgJoNDI2uBZXhklYWm3R6chHC/inzhKEwtIyO94Qi9n0xozlGr26ovXz/y5J4khuAFnGHEv95jy
J4wMLboEVncTbdxTOgD11pdEULk/6fEQb8kRmX1ijeMUhgUUK2t0reBLwTKJdUd0cclhmpCGb/b5
34YmJXOo9uEq7WOL41rQaI2fOopk57if+w6Merf2yrBTHDJ1Qnd8V0L2wb1W0VoFMIzzgSZWwDYV
tBAcfIIVeIrjcc/qm31grKAOjW/MnfOhq09fQLQ0O1m+bCDCQUXD6/P8WVMmH4ruP+5raAOfy78v
VDgNE82RwR+kIPVuZW3PptLh26dJNlT6M6hvpLUCSAs0VPDlwQ3h0csbVPjopLQXX7ByVKdztwmj
l4XXQBt57NAhfDkQbv4jFf4LD57yDb576yh8lbVWEvXO2GD7OzuI79oK8kwQSup+aSATOooWaw+2
pH7TpgMVGJlYyA47VGdjAUoUCHfY0D8KcKnKgUvlSJs9/EFbKLnr/nozJtgPwBFP52we7L9Bi6Gp
7IzHxafN7mMPQhkc012BXApX2j9feu+3DLyBiGvWtKZ4cKji4XAa8IIgcjoekiXJd1xeBnew4nTw
gd3KfZj9OnMmbHcRChhRewheUTuKV/VET37UrIa5FftyHRoHNL00N0G45w2kxwpIAV6OcfE9lVui
NR1vo8GE3Eeh2P3IpNC3E8qTQ6LvW273MgbkMLDtY2iNr8SXpI0Rs3lRS2qYyPKmM86RRI9yifS2
RVo7B22kj+wtECOUNuHMsXM1K5pQc57VBtXGl+5mKHWyoMIjD+WP4tLoodrtqBlBKZq5wfRG4x8P
kvODQr8a5FhmXolj9m0BktbHZzyxP4WHUTkJDVGOjpn9mBjVomJQ2Fz2iZlUIkygk6D5W9rADYcO
qsq3ploLSjYzWgoyAixbJ60d5ZbNncmofeEnKfp0Bevvq8gI3Fkzg5k5hG9JGnqgBv8XwyOSNcfU
gtKbH8/VbtXGsUVlocSGCXJkCwmI3f7gh6jXHqLxJQsalNuh4ZAw6cMXiRsh8L0txacBt9WFSU8F
Hkfaiu+GXsBGY6S2v+cLwOcpJ+ZAim4woI2s4UK4wBWhaNiFEO5D/WMZ5FrbcRBBN3sSoeP4U8mb
GgZue/uf67Jy/aEJowuGmO6OX0KpazC2naKM2oZlTP88rzP7O1aGGcjtZjMknx4eKQ0aFCJ3ZwG6
ifC9K/CoKwBHkubBxEojw8JwZ+/NTQTu3A6LmA14g8pcX05bMbZs6NReqXmYVNhFM35sIta815Es
rbfVL4WORNQyduYXLnja4BU/0LY/xypTIZf2tnVnV4A9EZYfr7lAfiqXur8XaYRyXtUQYJhbx288
/zmTt+CVu6ohMKj/z8CJXQuiSuvaZv2rKgcvpRe2whTnbqcB+6TLWiBhXQaHpPc3za/n3VLtMPqn
jMupCe9UAp2MNk1HTMRwRyfZTMWiw7qCggo56PV90X2sL1FhknKYpmJDmrLzX4bI8uj0+43sm5OE
6FEINbAE66996f+8kwKHTsCwqUQK8rsmqot202ZIo++iU6Si43fNptQbNWxZf9zodzgBoF7Adr9M
vwNZMMsk85pL9ABaw6eWX5kiTbYZBmFFwwjKgIyZlfxFZAi4/fQDtevUqZIbF0DQlB74yupQm1SE
9DCAyUPVJx2Wr4p5CdurEq+PnZTFtMpRFRDxzNTDXAaEF2XL1K/QUyFjxNIqYM8hSQyvDjCYK7IG
2MBeji9IEGGVPY3a1bHacPhiwO8DVpu6SONAfflFOZl2/FkkHsFoHRmuGD33y9ePaS+j7oJEEo1k
McTDKLd7yP0qMdqrCLElTUMQCCqOWVUerW1ynvAP2afkqKGNKQbxO31PPIfRkhX3r7dCkxCLhMP6
NIJ1vZJB1N+rPnc1JSClWsiFMc/3IiKbmkU+a3qRss5JdRBt8DTVN9whzChhukdPCEAL/oz3XPkT
zcJGsdQ9Q7Gs70QQ8r/nk0U2qSv65PyPA+YTrU9WFGRG2zzYGeJvFi1b9l7tCn6evcGl8G+29ZJa
TYYPrhPgefRWoprAMlWfHop8xgHGnIs7z9tc7V/cnQ5t2Cn85PfUB+4YY59u85KxxPGGUrrY844t
CyfTx2ouZqIA/+gEj1rkTM0sBI2loNbWA3UrOu/tA0OFWAgLI1os1FAbJUuhhDrB3eesk6WegPIk
ph7ZOFSzoYMv33wPZjSCaSacLWKe82aI0iJrxvJkM4nrKHauZd8kXOQPoO4mB+JCItxRT9GGrZ2a
bfk3S5D3oImVWFbzr72XAuWs5KsImS0m7rSSbfEVqba5w4AT9ujAyXEmErV6aDuV+XHwAjNbT5e7
d8I2beZsemmuvHUuJMjjirrf3i12c/kexSYTQ8b6ow6sgWuWXAPCbWIzcwvK12uZ35PZXxQUcYpO
BNI0mIbMfhZQyJXwveMgEnHVVgupjj2LFEaL1AegQLelHibBDQn93QhLoWOibqhVmGk8G6qB/M/5
zL7TyBQcEH0misOh5NtDpI90d1Cs93WyIm5RCHGsPvrj3gSMWtLo6Mrrb3/OJMQd90k9fqzKWyth
0G+YAVXN3qtK9cKPM45TbDv9Qq1CFvhGTlfE9TnxyNx2BnaR7sYYh1pR0YWtkozjls2P8s2Gw4px
Sy+IuWUun6XQFYxZcx/YfONOI4Q+BO6yJ/J+ZPoVJfUivqPJDKqflS+/+wmlT5ehwA16TCj3CzJK
Qa5riGLyzb1R3PkX8FEoLou0PmBpoUlUb7nwp1nEuaxcJKzFHOS3ctCgA2D3AQ68VBrLaqP9pKLj
4fvOm4ylKlJUts3Q0n4ZWdIsaaVt/55u72WhUEDeXdYRXQ4ejcdPR0hijnjvgFPVKOOff+B9eV3O
bbi8e6RGVElzDdFtOEN6RZGvJkPlc8M+5fiKKkNBYNXOHWS54UqfHiQYbmAusF1Cjg+mjg6LgBI0
1PC0kYP5hBvO5vGS/dEoBoIImFfWo2mio1cA9NQ0IXo8vQxUf6rme7ry7iXSyhZGtuOSKkrOKWaC
3FCTxuJ/pRf7zss2LUY4KsWKrAPtjA/J9kg5cyjhjfVlsqVkTaa8fZw9XPdLR4pijtwQlkxq8JH5
yD/N8u8VpuLXKeiQOB4SHRbsaWJ3Y1ibWQYjFbnO59UK72s3feJ1glgjX339wZpUa2dU7M+CVtjA
8RXdJ1xtrxa0Y3HSYWytY/thNAHYKcvmqNrrevwCF/Ez0Lav4Zn6i5SxEkBrDGF5isPI5UPmSxwi
brT/a1Z/nX5p0eUQohf5QxzfnzxnROJuIUUQPZm0P8EXpIcGSEKbvbz4Gx9a9DERglyC3bpgBbN/
8wS354oVSwQpurjMVxSAf9fjwrx7W3ErkgjoCSRD4HI8njGXBgpgUeKXikZPAZDHD9wuqDhZjjMC
TfwZfeL5DJBacKSF+9NguLQI4mMDNPk1Shr9v5jrBa3Ri5qHUIFhPpDBfinlpoBIn9wU48UIdWXQ
aHaUP1K6thATBL0Z/imAJVrGjzl9IZ0V4I0Ghpfr/ad1/yE3L34LUXntGGs3X9BJJAoGCKxFX90Y
dhciT3nXqysiui5dtx+/UYwbpV3vSGbAV/ne+kJ9HOb164Vkm+ojfV18BRtEWpM6XVMB0eNychXf
fH97p+w0D2SxV3KkrtXonrfnSgk2EqmGLWuyjZgLzrXkXBmmezmcFSIXaDRpnL2HI8LoN7kCcd8n
07sVQPr2r28SXVSEZ9QDgz0NkDGQwXPtYLwlZ9gvXd8Bwdo+404zTMq9Rl1U555I5CesCz9Mq9ds
6cIyRRzdNni4U6Cs5J0KNzTkydDEsYLEqVfTky02f7qGhUnb8LVDRZ1yZGUs42/HJy1nqmrKoMI7
rdSDGw2xntudrP0KeUWvfiZAb08jL5YdpKbc2PyFJZT44Dwrx4w9nfnUg2TsBZAt8vxu8DQqDaLE
iop69rNqYx+F5z+VrzepPUYzfm7I3IevLNN4Uu/5isQiPo5MczT4QAhXpZ6zhSUhIaYhc/wfrUO2
T41G5tv3E7DLlwYeM/8R31Ovd5ye3usOuX5fRCRcdYVnPFFHpKaQ2i+Eo6435K0b3miTba582p7M
xnHYGHXPrj2fpbkPvcvi1cpV8ROAGf/fjAvTGdqKKAAZebqs4GnGd7CBV6VrS6AARP3Ym2nvWC5h
AIfVwHQeKuMOdQtXEJJSji4pw2nxrwy/CKhHHkeyGtYcihlBMw+chd+YR7Xf+ry3+fM5vD2A6pQq
yQNEhD99R9ry8aCSBpkN4OZkd2Bry2E71xvG63jpBREEUAFeju9gcFuz2i6lRYNZUakX1Addklt6
j8LjgdqMOh7lZ1VVSg/3VdjeGGHLVXs+mB72++OznLoOdg4tMb0Cn65ubFqF1LFCx4NpDTMsL+Bl
0F2/lTQxv+zSrvtgACet3D/18YcBkVRjkmQzKgBU2oGXVG756PHEizB0pW6B7O1EotUwsoIYyTS5
Cy8vjd8m/6coAisarr0ln481J5XUuvcAPNnc1aJWhBIUX8CItam0nMFFUyPXJ4oP7g6YnLNbI3Nt
pII/8iR8TrJ42RQoS7nky6iWifQHzOVWXHgqzoWGumzLmBRxOQ88hUL64Fx/8Lf/6/iYsDk3g79o
0YKy4TCPkCbF5N0qFXvD8W/CC8QT4kldSM0G2bw2NQgcVLOPt8zWAJnGsamXSqC5dbkiXB9E1CDt
9CF1juhSVG7gILOe3Q8LkKcbcyZZ3lA3B3/z22fUfG3TGaBJ99l8SG2VujAdZ4mH6pnS92mQVPju
1nwSkO33davWqmQf9Tygc7B8u9GOYYmphG6+e61mlaD/tM/AGrbI64vQkcS0oLeoDHnHhRGP5BEY
q0E4SKrtdlHBi/8q+e6t9AV6a4ADQLralHwH0fxXk+vn6XQZs6xkRhTESOC7F1jibzt6wFTCpZZz
BHSb2ur7sQaKlLFcIx0+PBEftjgRlJkaqjayyMuT837rfKyuw45mvICgCtu78oOA1TKgXothbz8V
CYOOB99uRkxuv7ca/fhqPALdB3Lna6NVrVlOr3+g/Y+2gvPGWjDHT6NVebJwCtZgE03wCqHx/7U0
cc6wwQ0ng/gnicRRR/rew02/APRMmtkMSkZs0sSrCQuFwi0vBCXnjoy/fcvNt+RgwdEVb5ns5fx+
jvrSlxzy3yn115MiCYeG8bticHLJ/VSCvHf4SWHseP46eRGWaY1UJGBqj74vTj6FwO/n/SQpdBiJ
cLRovju8Gla/WYPWERYa8uvlmr2o8PGHcZ5lWwpzcURS1eyLUo5M5wlJVITM9MXqo7wo/tMCn6jQ
e3l20+OP8BsVpqEjtBobKcT4JY0AD5jWzLxWAgNmZwwHILlgBH5mTHYUTw8Q96nlTGfNaBSgAOXx
f9o3z6C9IL4SywREvgrJcDgKtUbxvyqaFF0P3CkHRcCPx6eLCRqrtSTzdd6jG1ZFwQwC07EHLcqD
ZJhImyBgsrki9ny2SA8ztb3Nk1uoxNfzSk98xAZGBSdnBTIYscvprXlfl/XHosrrwd4IvNPaqjfF
afeycO6Szp3ORkuGDTXOoD++smEFvIahl/JtvZXOD9RhxILKSh4QE90hV1JTGvmhISz+mKNwg+gR
AEVbqAMtGdsjbeK40KO5lKqdke/nbAzubtWe5JpmzP5Pvly50S/TcuWdVsK631v2nqABV3QZpC/1
OogYvEjhId8+fmkGD9JjHkdRl3j9Jpgwj9P1VbZogC+k/5hKv0xoq3KYqUJqWgYqweRGRXXHlmVZ
c67uua5wI/vF36mFiK8d07QFOweJ8+Ndrxg/CjW2YjqN8GWpICx7UsIOzxmgPAJVeqMdM6s7Uqod
fI+zckXeU5kuMduqbkqx5iAvZ5BmAIDfK38aYVvM1G3XHnr4tpw2mCy6+k4nvB7FywbPh/3yPPoG
NgOmspglIEfmCFc1RfAfAz6+QYqnQ4JA8N4k79xOcb7jhK94mlr/R+Pn65tG2VlWz/Rpz3MQLLmQ
nyYEltv52JFVE4HwBQ2RbCdgvZMbQU9tbTtLlD5hNZDXOj18mbH4EIswz21CL/mgl1AbqxbigFw2
jXQycQNPoB1ewL/5vuBSRIu5iw0EihLETQ17hjAnBTLrVR+1mrxoVFT1QDGX5OxF0YRcgT9Uf3f9
SAy0zm4lAAYOihJ6RYArWECvS3c6tWWbiv9wxYdM96shxoLNwf244YPmdUfiSxMhrt9uw3T7H7Xv
YkZIWM3XF6nGb7LkNaWyEaObZ/eQKY8PMvsX5MoZoOjekMD+AlVK4jjOXt8Z+zEY2+QQdVCsbvaF
EYwsbkUXRT2hk2DhZjvVZco+KKlrvfqYWYNdvnr4Rg7tAN5nFdFohJHWprHv1/89ljna9/bgLr3t
R6pUBcIgPyiNn6b7DZzAfZ5Fr2wTlSlNfHCkhcMStwuM4OZRpz1v8JCfe1Jz+hmx+HqbPFE7tA8H
KlNbdHtMhBPF9TEE1eJ0LV845SZPfRxu6pKZNzxgGptbA1k/xHn7bXnUmAaRpJ1pxhDL3OnK5p/4
NeuYPBLnLIz9DTm9JezSgQfqZ7v5eZPvPBZLXP7xmdKmTvUlaNjtlPG9bmyOTSKpQv0MQ1q628IP
KWe6bOwYdVWyvTwKk34lxdAo2P2Bc5ioik92zcjkguWBoBFkEla/DzrFmoso8u/KJlFCxW4qkWzx
IeSo9bLlq+H6zrm+cGsp2ID6NfK7FhVYtUyvCPJSmIQPsBVYgd69oF5HGM8rvtuXlDQ3ZiwllHUw
vm1DhekOtgrkWuWfCY3SpZDtXp021+Rsdp1v5dbrdS8EvD3bkhtcv3ua5ZaFKDyaO1g9sSqv3eeb
rSdLKvAi3U+HGtr6wd7LSwj7A3BATAQH8ZX9N3jk3H7VjjitYiYC9x66iiIZhvIRo72XnQuFgNrS
EWJodM3i9PknynCmbGofVtydo6qxGUdtqvztU4Z8F5RAn+pzXqPmzflAU7eO2heBLIGEpLslUJ7n
hEP3VwoFyiWF/KdWoHMgHxWnAlKhfMi0liApUN/Fh4WlUfOItb3vG2Ov3zfgb1WONk/l/rZmVwi/
nSRTsxAGMU4NXRpz0bPPcvLLFrzuDb2tM0F2js7k4tJr/khgE0jotd2MKmsnEROgL7k9+JspLDav
xpuPI+DTEO4cPSCwwpjDogq5BCniZVVJ5MUy5chXJXj17KoNCkVPp3SOXu5RQ/xGo0TEGf0B+m5R
lPCcrdvzS/nskohkiathYdwA+B/KJXoRiWZTvefrGnG/zMHfLNTTcOi+8TODPTZKl2fachLpvmde
pMJzmiTT/XZNd9OAxx21M7uXHMpGtRC9KChhBiXJkaz8Y9kLumsYth8sjuXezCTkUaG3VSxbVHmg
hQVJCRozqpt77uFDuAEhpfo9fzKpRebxsfRhocVWIm2Ujfa3Ff0odQ4OqgmIGnIuvFxBP7bBFMpX
mwQuV0CwkNJBZYBZtyOhKfIOxWgk3239pTAyVbsJgALSMWwALPs98nTCz57wUhaq0/hZs6qdrJZh
QX41Xg1c3N01x/AieZKT9WEvqhO9hizgukCrTlUn3TwxkbqENo/t49VbFKNecO5klsSc8objshUM
n0cE5jnIbeMnRk3DBdS1YjpQG5B41mBPL8zKonYbxW0xVucrc0ncwSoWdtR/g0NkGsGkIS3N+eg9
m7g0Y8kAaLRCAim3Y+VIsfDTUZ8XjJ7m5vhu1jQNPtMEq3KT1w/EyOOj09g0A31HlvRgTQBsB2PW
WL7CQaPOze9R3Ye+ei20yb1peiTv2cV72Mldbw/0NZTYm4NCaJCfL4NR5GOmgdIfs45TWixLEMkw
i2BFnJfbZDOCnRzBL51y2cHbfJqbGBggUFxkZ1e7tQAyqmIuSZ6fuFhqFT1NP1GMssGE8qKG9UI6
pzjqzCVoGxdC+kHkQGS3JCeX1gWGmGVvAenKDmSXP5pI43pNdbDD7wnEitoRpLfqp7XL9+zT8742
IICVsjE5o/6CLM/jniyTJQmC4vTm7oXj6+xX8u3g+QrXNI3sW04q9uh2qRmSpadGBpeFgBM8Gbcl
24Paxp1E6mcRV42SM0fGIPBhJRO4NmrPnKvKT5dFy8dCwsb9DBy2kKB3mthiRetoNUmQWndN5j9P
nj3hHPVs53RAyrSJRNam4Kkv+lQ4Kgih2RIp8HTFqCmWbzOE66/ig5b8uuqLRX6PDFpTM9XmGvgz
hj/bA3Asz68merbs9g5WGiuS39sinQ8QhU41gqIm5GlQcV/Gmpl5WEgQ01xcVjft8zWGZCXWRBP9
a9qMgAWzkzbqRljoRXcgbIOnkFSJc1sYo4xgGbO5p+A3z0HszGmH/bpqTrGR6nGLYi+r9i0W3xDZ
XNR3vfe75/MX0i4ykAjwttL6R0V3NXNhghaMgR/Z35vv0f7mpvty4+hY17PDg5Uz+liNTZrqaZac
w594uclIhXXHNhhkH0m8BSn1D0zg/anD061dAZN0iPDHqkeqlU6HXoJbnDtZox2aGE1EJDA2ik12
zd7sOtWGlPYFlqxogeXdZ5IkaENsozK5M8nRkeCTt1pZhnHsx9d//kzBIC1Rira7ETnRNpnDoMko
jdhHnLnRMLcVX7yal5WdfFxCDfIGLpF/0dGvwPgi7QhTwAKVgfA5MlY0NlD3knHiAJJHBtunoKEr
jvZGdxwFGy20OySSxQh6idTmjSKAksRHdOi6PQhONXgLeIZs5+3Kgv+ujbyplTa3HNAuH8GXh8SI
o3qmU5hrX7o8aJO6MlXiHbXr9aYefcHFxIUqkmuY3axHPz8asMXvnxpZoINqAOxnA1xDvmj5U47X
zFmWLuxnuByPJzXYKEne6n/mcm0htGv11uyp/XXy1PDdBNsOTk3vt6yFdc3caDBcOveMgyKOsJH+
9M4h0tK8wbN3kGqtDb2TF/gwW0oFAfkSWQTk3gq9bjttH/HorDwqJ7zV+emCuxELzIJFMIL7aE5m
Z02k6bA8D0ekcQWKq+YV22Jf26MKnPcCpj+mycAkYk7/9M2k488Lim7CLG9PDhzULCLjTJFoFozq
EKyFIgj7Kqw75U2Xte4wDCDq1+okcHtn6E5HjbpfARIsDOP3AttephODyLEA7vGnQyvMTG30SrLp
/cMJI9UkINKaLYSUUJnQGzN52zxA9W3wIu5EX0UVVAZOrWkIR10XS386Mx4pPrSFYuJ8omT3le5t
O8Tp/TevVr2Azj7Mv0cSIi4r683yYZMBPWB7kD0abJUCOpMavToE82fPmj9iRSfd4MnSMfVI5jMI
vr8MopEMeQYduKxMx6IQMo9it3Fj7W+auQ7zJwOV4e1XR4s0wWJO/f8wNZ8KRCgPnhTWJADDfLhi
SkHjow5UNFqC86ufcCmmdu5dYANrdyFn1sfuoCRJ4fRCLWfZzXu9VOZgAIqaalIpmAi40NA25Hc5
s85527u5981euYCS+gM8jvoPSwYUEVJcHrrENGOorY8qHB0Gkmv1sNcqj+toCZDdN1iHSGN8C8Av
D5x3FQXZmU5+HBEYpJLaVYXDicTXbvqVvfXNY6dcg2ErEWsyo/395iSW5ycJa4EFNHwvRblkS3tz
9vpozXuZNZaFWk6cCX3a8xNn57YdsRZUI0+lix93djQ7opva9WAYvDD+3lptPxU2LiCBzoWrFxVH
UrKSimDQqv9OpG427rJ/cUqERlqDEkDekMljW1KymPzZoCRUUIp089/XRb3QQZ5xGnAby7Sc5NEZ
TsqeEaXRXz9Wt6Wspwq28zpnVYIr+yAcwVWn6VVD3rO3piSijBvP8HdaMv70f1Aym845YBZW9uuI
F2zVSNVzb24sLqBzIbNs6ir74KNywTyOIq1sSk4EYsQwbXLsFOF37jAINMwZL/Lygjs7vqBwyeeH
5mL/lxrlTx2Mfph0vJaQPaNsQIX1YAIAUVtAiUtS9N5n2E67RtgHxwJ+/J7kMmHsE/C+z4oMC8z8
jaIfdvca9pbehVtFjEMejJkreTPhDbnGWIyWqu5F2WiHjbRt8qUkKxs7p4SBzN1/xzl2T8bZ5cyf
dVYi6irq+SKNKNIoI6OSlnKPuPWNiE5UAHx+sjY/oEuut1Opa3VCDxGRG9SqdijDj+QlN5+46Xhg
/C/eVC1jOtPVwvTPl+9hDCO9Xy66YB5e0MjalGpVzbH6X3zqR4JM2A9h/qkzCOsfpblr3kFdVCYn
/+PQQj5uNQBbpmH2vvVDFqJFx6DSY0kZigYu7sZ/Q2OOkiYG6wO+pbDV5j4HUv0ZTqA0R7/xEBl0
vLtOp2RFySdP6I3asRenjhk3imus9JWOymhaCPCLCNhptuF71IKBHO8GI7kLtpOfyutzAmDD0yUc
2vm90RtLK3P4AfqDevLXINJiUyM66if/fb8k2IEH1Gc9fKZd1EENctkiNub4sqpPDW41d39YyOPX
o6fzuT9mFm682k4CkcEZavuUt8aFy0TgGKvaCVGpGwfXbkjy6X8ijuEAK/Kk8A3mkbLyYrWAJAwC
fJxheMoqiqQFa1nJzlJcrWk/38zGav1y0vhey6+Ro5b27PpJpANRgw/XTFlMYociy5xBcHoyBnZI
dgWNpIkFD7CQhsUsSkbf2+8vEuZ+EZvJHsPOO6qac9EDIA8slEpSCQ9J5LiMPmA+q1a8iNbV0BXr
S1sxGOAHR6OAWirvDZ0YpxlAofBc9s0JU0gZRm+SOF9NdiePD24CnVWFchEwQ4Hzuyht8gGpGsxr
okwwy3kIYQKyr6rU4wEmqtEBGsy/1mbWtVXvpvpu3t+dxAm2FcSek06Cir7fcae9toN6GLQXiJkK
aMe/iXOkvV8ph/aZlYrPT06OTL5UrjXKvstA5NYO/NWlkMFiZjQ+6/G4gEyYMteq00O61eDvgDn5
tucw36QSh/HFJ3kakrZxMM8ooCMm6NMcRwsXFUPS4j5MxqpEh6SPS/3NnfGggbO6fmzfsJdBTlsD
vzuCJDiTWyCRwhHf8wBzgE/c79VlXMumexxV++2Rc6XabCwAnufWRAhfbLgigMI7I8/Xu2Vpftj0
dEo012zQ+gbpyvU43jv1r7daIllyaXpxwaT6Z026Y+xJoFDZzvIclim5YyHSINTpy7fva/Thw1g+
NZO57vx80GLyvopsEwatbAjgTfqNHwgVrl0GheYlQ7+729h+uKnJ7C6v5+Z587OnUXn93BcmkiBY
wcdmudUmIks+12nIASCAl7GgULFqCerG/eAnd688N85elRdD3hclcxcJfNRTX6We/9K+Dm7sc3IY
1okpts8MSnPRxn+AzRhlbSR3DuRWtA/zV17fxcw0yszNb7zhhExWPuRzf0wWdbNOs+m7+PAwFOYN
NZ/ToVzrOXQiFOJOl/v2YNOftlxTpCLJhehdR/askU4AKVJqB0AiExIlwbnQZe/PYEqrjRj4zEQq
z8/smuJ8vKVja10IR284Qasw600ykaGYJBrsmNd4w6I6owfDUXs3dNI1Yeud/FE7+4TH6UcTEWQ4
gn5kW5g3pwG6AJvXEy+ltsqCe5O65/gvD2+qYPO+opc805B4LLOCWjGlnj//HwDPXcgi8TRL95JA
FGSnXs5mBEsh0OKdO5L1R12UOmXn2MwP2UwSLlZktjrKfn6E2BtN2rIpuEXduzBHpr1+3MGyKrh6
bD+RqZht2TQJz/0h95aBw34S8ZsGG0Km0we4GM8xO0VU3njvkVdt/TFUr9cwevL+l3JnmwuI1xUY
BX17JkK8ZDVLT06WjgyDtFZED1g+khPtTivdbudz9yCbCWobOkD5UtcEYwSjk2m15bPUig4IL6jc
lRhqs+YSdpF+osbJbU3072j+RSrEOyu6ZaWu1jCx0eM6lKISEes4yO6yZN6qv2gFGNNTQyw4lIFd
jbIrB2fMk81+9bnZn/Cu2IPh2UyEfkeYB+HELeBp+n8CZxYBZfsymeIcXSneX05ACtmkax16aP3h
x1gdhtZSMHOlLbU+uifqBEc4jfTsSvjb+5x38Dvjhn1p/Ab4m0a8qdWiO0PUHgyX0o8Jp+qoF/9a
x4aRUibLVDlgSWEEBju6KFOcB7EfxfMqtzRBWS9v0PW7aZyKVTSFn6A3jwxCzhJCGicVBacbjd5f
1JGgtZXZQ9JHpFIH4TO+B9pFZP8dzWwQARSUoX+DZSQObzSy5v6//MIwYb8DSVXkRpgdKiwIYIk8
iK0imr7izyuRCcJRbnIAhr3UWo8V6sMqXFwRWIxlqGkLLew+DVgS2h2AuDlHa+irlopWmMZ0lrFU
SCPJMC+rupDxM+rIHR07pldtzlNAol8A4j6GT7xLH8YhQblu26Wj8BBaYWFws9SRpnHb240oNNt8
HyJttoNWKuJfVXj5RFECYs4jfK0c5ZsyJfhEpASpnHr5l2USMjrff60xbPAbY77W5uPUz+/FPE2q
hcK9O+/fqYyUBgUTH6jF46/DNclMMBQdbWItHJ0W5nY9CNUi/iRL3Rqdtjq5AHJhk7lzOUdtbE8w
rFqUapJ/ftiIWBQVf9YvLqm5v8yQVMU0YN2eqXUjR7sIQ6kT5LDjZu2TnLOpf+8Ds0mnZqXnIXgl
svrUGOKCfwLEH/h2x/mvZOggMcRa7fNa6paHNU3HktweIgyFQ4Xh3y6zESTJF6zr+2hJKypbjkIA
XKZWinBxeCkVkRPCItXCmr94yD9nyxMgsgWz9I0T4TPdaPlr7vPOYDAmwbbjk/M1AVsu5+LTHubM
N1Ykzb8YL7RpUyT+NaMngmKZ7eV6CznsRy0AsJl9tok2vr21fNp1d3E2t0YiaQk8tvM/GIAh+oSO
11EDczzD0dq3Ehoxsi5qbSY4FD+6kaoymNHGUBCwnZqTcWgArJ+3B7Iu/Tq2zuSq7oEUv8ZXlU0W
lMIDxgpurZoEebMR60IIPl0tIsXFcoCz+L3pZvMKfk99VCKAm694t8SRh4KX4we3XZ5o4gK6QRDm
DwQ/LjhcZ8rB71ewWBA9DEbUcEhlAE12eX0OGwh1T0DHenlAovhyIk4/UTNyeN3T9d0gjofnt5G1
Ottykt89Jb88IwHDeZKSuhmUA2tJktFQuPArcmfRL8N4ysdCO/YfHGyXt0cG+ArzvhaBfGtLhxUl
BLRU3Yhxhuy/CwEMTMMpi9XTlwXa8Io7IzyEjuZmeBML4Y+nSQsQ1UcFg+EVJcg6pl5WtNpoFqAh
umt/gOS1DqK+kOnXBmwKw/oCFYZJaNsra0ibGTOYQ7XZ/nVQafLGlqn7ceNsDJGKfcDQdq4g/0l4
ale5QJOqUhTv0BEq6j8R1nNHD2Z1Osr8PqhQjY5iGBWY19vIJ6XtvQpA64sgeBcH1yM8OloFk9Ye
E/k6sYN2UBvsCrd0VuDJtzbOU3wHTgc5jINTpkXZV7H01A/T2y/rXRA/7Mu2cN/aNliyor6kAuHC
t9iAUryUsAf57VQ4TmHJ9UxYDlLEtQ358kZ6WNjKZd8+hersjMikOm2JZlmBLyNMm+DTjJIkKFjA
Sf5ACcfMjGWonnzbkGErc+seMeTQZF1fdv0CaNEQCgSRe04ZYlgb5mrrYyJF7Rs1Hw0pFUTa3Cf2
vf1pLhB2e4el2iLBM8XmUFzctMgSPt9nbgYJDy+dxmC+kln8u0HLXItqRiX8Fjq0ZDUgZ8gRRLQk
gpSrdNxvcc+ib6xe1AHH5BW8cgfKEB7iLzXgQzDSp8nbIH+raNEiLifc2K7WrCVQ1nZGLbC43BW3
IDLTJCL3Ji1rZROEYPGCsKlgwsgugIMarlkBXC2o95FrdLUBKKWBssEuAjhGiVbnOymGe0cyYvYG
Bnx6mZ4rkYN2XX8bBuNrhk1uqmblnvqYin5l5Jtvd7UqoYn9KfQ45Ee5isoY/Kt1pjCohhhFyQ/W
y3JD0D33AXsG7jZsa0tWp3p3qO0hUBQLDeavU6nsSXtFjvdBzQEkMuWVlX55U7NwoPrqjUU98i0m
mFR4mNf31fSI0u4hFoDwubi/BvtQwzcIK4DSDdT0LeL4ReeJt+bS7xGUe6B+TSZ3TdPclxCfr3yQ
EhqKuo1Phvk08d3HXB8pSeY4JcVwx4tRDAqBXv0aC6qRNkhJl5mo/3ujiWfYOzbYuF4DUs8L2DJY
av4hb3+2zZCHz0+lKNjEcHy3txFu6jAxNFL2PsvkOFFX5u9LV+RD7+fOD+xIMGr3gcXiRH8XUpJe
nFVKmhQn730Ep+LArzC8TGkp7hcYb6zBhu1tcEzsJS/jdpzOO9xjqWfAaojRI4PsKyliK5O++3mz
n+o+Cm+Ik3m86ur6epwycONorBIpZKiaomI7RT0jU9pbT4g0NFnP3p7UNrdr/gvGm/yPPstWVEKr
WYN6y26/FP2LWII+LojEn0Sbn2Nmkh6xk7xIjVUs1wsz4/VDdwvmV8+DgsIyW+wvfbhigQHRxUOD
hZ6qW9rZigmXS3rJCaYM2+EpUFJPKfXCMOpFmo+hig8Y+JUKfOWMqYwbEnpGW5H9B1nYFNdwYCYn
Way5LhXpFADKvqw6HQbK7OOAJs+0FfETsqiYnGZCaFFhmMUW1Nd5pK/zfeEHtd8xqrjpT5zRjAAo
A/liF4+Mf4A61Kdv14FJhkRLe+KnDMXOzrurfoeGpEZVWpGWWDkzQP0Vbp5eJrRosnpikkn/TS9t
90R//1SuPL6bWcG9vUXiBZjrodnz+psLjGjASufqZzmhaoZ2iDp2SBbe9Zge3/sxrDz4rpNFYrpj
9qS104YObZycVQ5/FqFANvygqFYA+Dpv9yZY1zu8E1lsCpu0e1cYaF5lIHhNFVLpHbhfWzove+Cv
VeP93J+lRaS9CNit4wFtOkOaBnEqySwy6goEj/d1GxPl573Y+p7q3V1n4Vr/N346m4lSAc0sN1At
RFs4qrWKMVSncgQgeYNDRK6R+CktOB9vTQNCzXiMTHJSw3gKhAlSingDwIad5wVtarbPteVXJ7Se
gFiRyxz9Yi7G2T7mBbwDbI+abPZeuogFP0QjgQYP6oms42L86mWyrm23aUD8wSz2af3hpe1mW//J
KfRXbJhJ0t0nWKp7FDeR2jLC3cwl4InFY3909wkRZNCGAGCa2twwauWXECE0iZwsle7kjaul3Tkd
mNdG8pQQK09CqEM5gZqV8b4GKQ6UEPbBMQCvhAcXFY5/wMXY0GEpRs0xTP8wuk7WK5dl1vhtrmlo
NB0tVI3hNOAnTjSJvsHzLYazaJEBlcdvQNhLEbzkMDLoLgHT4KFAkkuwErN4VNcbWSQnrzGO69fa
+D5YEauf2Fs0/ZdAH4DaCaIXs7JiAjABM0OfCLv2FEbV+eB8qsNitMdUDMndgeyAUEJsAhNu4qHC
ydWwcJFMEj0WngJ3PNxCJL0nggdj4X3QS8gHaPgV4sExvTdUgKvu2OyEA/HaHmgSRduRoVz0qpud
Xn71cF3k6RJhpGdEUPIj4XJEiFN7dxvEpX7xyEf+RZu7tQzwaZbh522b1n5caUdM9g7fOTVYsdcs
cVskzJr7yubmzdPLcexdjGO9xe2sfAODVLYEJb6VeX7LHPnSfJ4+r583jVWKnAueYb4/YIIGZhpB
kL6KSN3G4pRhPd2VlZUACXWd+kfjkol0dM5V4jgkfRkDKiuo2RTZIF0YIu/BpHKwMo02JFpRP6bR
TcMdEdz9Y68qfgE+JplbRWthEt7psrKu1bekKCpeRgw2sKXO8kk00C50Uw+OGgwsEdlednk6HA40
sk7MP7fyNlU6/tkNpog2Ab70lqyC0F47oE2t4TphPicfIaltxecBi06ztuq3dDWMl3VYbIpmG3ks
+jIoqJJVqDSj1opNZIIoUu8f0BITh+LSvtFNR+Q+CXxoFJZoGc1HMEbnxRFm6+O/Y/yMUaqEUElN
BoVwojMGhA/xVkuEGazE9fiBQaq6QuOqMCzsjYZriW8eRLJLj2m9USt00M59eN++NMpFQEQUZHlV
2s2L8DMeBVKl3txXE4bW2PGf9y0oHd6vNfBNf20tq3xE+61NaSv7HW3HJSBdP1sUEyvmm6s4ZdKG
5GdJCYYivczKcxnsd1SDoBseSc6+mKaFDYRT2gLC1HXUOUVyF6+ODyRGlVa15GIdHSHZGVrrJNdV
M7rbzDxKyWCCcb+iXjuSpPgUDzr1Yjz8c0Eyn3IIo8tXJugWnwbwgVNRe5HI9JRXqQQKieuqmOCx
JXNI6sTBPDolhX+H43TbswL07PnFsqerIKs521A7ony4sseMGHi6pJ3wx3Ht3OgtoM2EaQ/XGZyR
XO7GDUdMzL6FaSDeka1KH3MVfwvzXiwdG4k3RZeWQiI4FytEpj63fpH/JHlIo4LEZgMCh1HPMg+s
kBmyUelpTFA8mX5ikxXVhq1uNkxkef86o4shyQRhzj8w/pfnHbhQEmzp6MzZX8Tzz6hpl6UaiXRD
vQ67sRpouqlxOoKy+nP2oFd3zQ94zZZkDND+XZgg8TejIf4RJUtqq2l8wGQTTNi2XoqC49CuJB0J
cDkTuexsPuVB1wUUrkR3HHf0QoJJ5PMXnmptbtU8kW9AxUxgplxUjiO1VJBaKm8b01D30qNofKL4
1zLX/k2CPqR6vEjHVshKT+C9G8auCGO9kuXV3fOriOOMr+9lAuoA6c2HYwm7n64HCOqyVDaeDKHQ
kCBgUJjRMbLeQ21ooIALHqwC9p5LGMX2Q7PRmohu4K6KnQaGAH2NryJGZjBC0Eie1cXKAhvCTdTP
zdr2qPy87l+C9KMiRDbCjscmLcf2fq3jL6LiH1IXNaqXQ+YBNwbHjW+wYpf+utdUqxkmPOYsUvmG
pDS0YfteQONUutBPEFXQtYDyocu5SfYAJy0RYTge+xSo9/VPLlQ0zQvnHDo5Jsgh+ZfADEObnCDC
jDndqqjaWCQ/rD05mtre8xrYHnkICEpFbY6aSHDOobn9wKUgHJ8scArhB2c+PqGVU71H7bFWNz9e
bvM87r0dSqQdjjsXmKIrrk4DS2UOuYA0ZKnifPFeLWEAYn2MEX3YBVMGUD5NEdJWszMR1RZkBQu6
pMEuLkIOupXw/njsiYwlclVBQ1oycIxXqIxQCJvyQBC8itJDpa40sV0gGWMGnR4wILSHh+hm901O
3Uaoq8YW67H2PxoADJ6PuXBWaIpJxPNexJBobxvwGIKqd/uDos25eXVG6IZgKyx+TyF8KFYTTozU
71mso4aQhL7JwH/nnmFo0vMRP/JXMGlQyav2jXIJnF6P8a2KLURSYbCRHVorGeFxCCnlG3hR9iPr
i3Z8vHTpN//XxI5l22nwpK4eyd28MrGxXJZbS6x7/Hut4sbEfad6zODuNzoiXy0+Wy+DbHoOz0rw
AWQGa+ourDwqb7kAb0xRjQosMetQ4lyeNNNjjhb7qK8RZYWYw0Ru25jPu4g4T1x6kehUnE82FyJ3
TBl1RFxVYOKXq4AGw6sQmxj97OfNUKiX8U7wwhe1ze+DynCUCPdcuazjK6srPYbrzPDvx5pxVIxZ
RFo/3SIpAvcIa4emAKBjmBRPosAbhL823LOSJT1IeKqJugxMqistXWqndsMD1jha7o7vv1CjYw6v
Q3fbfuzpxp8cjZlbJW1fWWbU3U8RzAxBKsMinLwnbKBSBeSEf1x4K1cexfyucUFSOih39MBtu7HD
7eZY9QdDyghEPcGX0e8AQnw0DD4P+cq1nvHBnLivjP+SSYAFivUZRidl+KNzHYAwlhvMJMdo3gLN
/RY+Pzbjq6upzncBxNs+dPZJ/PILQj6o0LY1OOenulQaNws2QjG7lrQP6J96ff57UukFRuOMH5Uv
VaIHhaN1uMcRo1IHWlRtQ2rXh0A91UsjdvO8YBpqV/Zg9XG+VLeUSwPDhvjV3/IYbblnkJhf3I67
v4EEKg6ahhy0mvvzPD2nVt/cZC0r+tW7AYzUrKGe4I0XHwbQ7ZzqR1V5U2pnbEpn4r3aTTsMba6W
pbne4axCJSHrv5IWONEJXIev/QaAgTl+Go9UdUNhJ/n4LffLRK50qkus709gJ7vpL87GaQaY5NTq
vvrYOLrDYqEKhuI3Y1LVer3rSJN244EwQ1y95BXMrHJeMA+bawWdKbiLkEKOR3H7VDH2BHPRs3/G
EaasPMTx8doghjnyLdjELpAZAYGDFU9fl0SPwNPoG/63MM+CqiT5qm2TwYKYgSQP1fVyxplpQRds
tpPThN1AYeP5761c71/y9Qq3G2MgVNM++EflbJMmkdWNQlJJGRj8sisjSO4V5dJyAPO+7sPTTtji
D6FC7ouTpvlnDWibJOynV6WrgRbmSt/Ri1bcMRRd+cDrlQIXNYoAlKVRiAg7hsqpwudxzWOzakBI
Jf2CLnuZojfwpyICuW5WAwsYFwKzr9skEyV7kmbssy7DnUm7Ycy67NAwQwTshqH4bvCdts8LbOsc
ZLc+AdGVsXUboXT0psMpsgxSNKQY0/IIYCpxmLveJB7o+8/gKPQwky5mE2UTBrCZSc8+RydSN2w1
8wNHPlu7ycQDUug/AR26JzUX5HRoVPRpDGBO+fegXnroWcO0xtaoD8ICXqX+9eyfWgPskv/cOBNk
YhBlE3Nc9gD1LxrRUDn53GBfb9d3NeqIxIFmHQPaANBAU8Zc5j3qyarda8eJZ1QNcRcktAcgajVT
mQX8kcJxM7TwFkfd0s8pBgEVlj8XSqjkPTZHA2GSV9npWPmFk6uOTMXNIy13mQ8mZnjAfzgW2K/A
ztKpCRFnusBhyu6MHHzC293D9bbOjYTsGILPRTAGV7Bl1sl0J+tecq4HzDfwGY9dP56YI/N3SajF
uZoQlXdkEdNA7MN4wJZ49aNPK1cr9Y2U7OdyRHGqDFnLnHjIDO5K9FwDV1iGfR8X0ajXf/K3W7L1
BkBn59wuqn9cuRpyggrZ8BaZrYHP3/vlr7s4BIi93Wn+GDWIRmNKjPylB4JgWDmRZgwdZ+hVSqT3
+qvY6nXYxWSIETty8RiRNBGfF1W9Gn0JOC4/YRTdGAedVCN2dOyiH8Qy6S9TFFuQ60Bb9TL7UdNy
aa4bLTm5u3fSgpHwDWyG1q4ClFA4GQVwYZep4yZm176rWij4xyaUdL/i2cp1udXkA1TRPtYhdLS7
DEKRrh0poCzVqOUHDt8ToT/zNWfJBQ5Kc4gVUR6fr6tdOwDvxsQjAl+cntyH8XG/D9Hr/d7/Ml97
YbpkLJNksgojIHnmi9W+/qCZkiHEEAvZdEsflK2hhq4s4qjnsLl1DNS7o1NZA8K22Ld5h40NF/qW
ybb4dxuF8zx7SyRvOjDzuabNFryHxsMrGaM7XthHoakBRKWMHq25bnGCWlMfklZ7VfnM/m8R55uX
dXME6UUUupZYMw0BY9eGZLMDMLkN3Srtyl8OIFG3YiLzr7lNGCH0w2Ne4y4tOIAP+F3Vauftmwst
zB4u6ACPklN5f59oAv+MSCa/9kUMamNcNezLZdsob3vXuBun5/Xyih4jh5Ab10DkVbXSKpm+pDMG
5SKO/hZHVQDPe2+OdC7yOhr6iacfA6lkxz2MuILgikzFUMXzaQeSyRm2gpeB/+o98IaUmljmgH80
M2nslO6RHhN+l0bLBZ4kOHX3on9G3sNzQbYLi9S3PrtmfNClNOqvlbc5WEtW8nePJeG1a3AUplaR
cinF0BJwglv0VtbC2HHw9hHSjera5aqaz63Z4nfePMX0w3Y90M4PYWSdORXWL26vb5nESnebDl2D
7JfKkBVrWtWGwTJWF6w4KPU6MT5SSHBnlANT3l/XD26XJ5oMixH16fk+jRoSOmmmGHatoE833Ip8
c1WDgjmLnhwnvRFx6bs+YAoD1nawP5vfIYEFLNos1i9lfUViCLhRn2OHc9GZhc1m+DrzucUZSSNg
HW5m+TfNB42DNKECT8ZB09PTFsBvWYTfN1rlaHACjMcb72nU+SziuNTiX+QKsnKSrpd4LGuEMeEH
0ks3NcnrwigW8m4WygEdDpa/opqrN8fGgx86WgMV7OeiQgHcoqo+4hTrr4Vf2RIhCiSVJgKhFdNo
fEsnxsENgS0vee/mjYFMwR5OHodvB3oTvt9U2om86t89cVS5o5Oq58TOsL4t5/3RPoVga6wxFB4j
Ho3Jom4SpLlKmdmDDDlTaD1tpjTQl1m/FVa/mIgSDwGdvB910KqOBZ2JereudoIhWaQBOuSufwIz
cMsGSNT/7ms/CFFCfnPiCTjhAMSMqerl4Hnhb2OmoW49Tg6ZJCRyr8SrM1sCBc2O00KLgdoM8NTq
XNs/cJ5Xt1xCaXkn0uZFKi1kddz6F9yAkGZMMhVO3IlGgsaZi0cQ0xY2ko1XoY5j7f1zb5G1wOKo
Gqo4nICrMF5lkAeiPaby+/0xk8AZE10LVSJVi2C6PMS9Dxe1Pv+w8ijgUqTfNhYlobUJnD3WYeXK
WpTHzixRcKJ/5ttAxGT5mYUxtgdLX75S1k1tuS+d17J/A9GJ3FD/z+4EYJ8DGoRyHTcJfiOoCOkE
9nPbrVuptRpF0Y8yV6gUQsE4fK+Kq5jiU/i8hL+JCj2lC7OAJ9fS/8hJzcxhbJuMdCd7t40hyVXc
EimltFqNF/rCTL++R01z69yGVtG+1+asUZAtoFXHfVCG+cNIFjIbuxPfz7JJaI54gl4tDoKz5DyP
+68axqDdEWsw9bqlS2kNsLGPRDDJY3nq8JUvastwm3mgeZSjs3uDLCvJqu7KaEUO/Cob0/KGfXkD
9UEv7op2DXFSvgg8ItuYz0MJSkUDKqkCOaj3ZnL6YtKpzOjqh7loKk8sKKPGQQI0leVMug35kVSh
Nq6hxJXtLKB28+7OC7b3KtZ2J/eZP0hhnwCIRD5zcjkOx/z4sbkLO7gtNC7bYhYEmhS6zTSkNOr4
07tqwzBmpv4fB3cpWqMaxDQHV6jMBWY63NO2tXmRlE2OmFdPZAmvj3wJsL5Wi1T8CvcptC9xIjGf
+p14nZl9PJCc/Rh0vRHVZZD0cal1RDuz54BL4mJ+Crj6l8lVBktzlpLiK82btf0pP7/r3QqGBP+i
Go/QztXM/Eqh7206SVqo3EP4fPetTqobE8TH5fGbgwwNiBuPWqi8wwTEn+d1+f3HnSP+OghO3auy
S3e2qViTsUfrSchRsZyBmjwK0lAIbLmxFTIxIU2v5Ii0lLys5mnX2kqB4TN1RnVyalgVTISYhMai
EslXN4G/FFWBWz+AKKRNGS/lAbRB+Rd1kdI+DyEsehONJ91MzlNo2TmAy6sjatVSv/t8sQNZxez+
TgX10FWSLRIxUR8Oa4cPIx1dNUp9pJM9mTaoJDMgl3bOMre3YHAtfY+bFd8cvETJvY42G7+nUPu8
iQTd0jvkBGZioETyLvebdY9/x4R+Ec8QGwSKlezsaGZOu4u6gGjKg4JOISDXTtqY0aTzPM6afhcJ
TVdmbU5EKmAH14yikLtT02Fi0gd+E6OlSgFW3fh7LXkD0JdLySZpnX7mSyI5jIIyUc6jtNoOo6lT
X2/NT07SMJDY6tDa8nYhVO0MIThDGLASSCtgwjzGSG1z/ZGmYL5mZpk8NjWnQ/OaG7QNiwDOvIMB
DhrfD/5KLcjmu3+5+RzGPB5so+moT/Bg4RjjfGes0yPtPagR5ENRo//Y+SYFTf4CtpOQ679Qbeiz
F7L1M7H9hZD0jQNSEBrbSDF3PjsCAFfsHHTR5l2Y4YlMErO/oE+d0k/puOmTr+07BazW8BDAiJM4
96WV04WQGJQmsEARQpI26nuhHDJ/Ju10pIbdYIlr05BRu6B+DD9ZyBh1ZnLhvoSQIBzwqSsH8B52
ltQZOjo+7o06lB+xVgXoH5BNgJ0sJh8Im/kFYwB5+D5Wdiom3mnmEVqQKe11qyku38XCXfBJPE7L
fqzYo9l8MTEW/jeXRi1k0vobCzU/3VXt6Tas6q471bxUtVDs7LPPgYxQGrGdnnmubzr4lJatnVV0
WpSP4rvCcyZUz0Z2RXvh8/cTpHIuDQ8mE9GeZRvJVJ9AEgbRj1Hr42dWclmxmfSIbNJ4pNbU2psr
YwsezARjXopNuLQjXnJagJwsRA5I2uX3G0/kglSQg3kQAShyQndR6es5eW9YLKbkreATRpH99ZgV
2Q+gw0erblt7K/RiPCDlAaP+iU9fljrR0Rk0kFk/OQil/aYG9XlcAd1hrNMol80pns960o1ecWMO
rAauH8Fj1dkz1syz9wEIySSkjwF4ZO6PQQj6ovydG9cSt4JErKWndeF8JvQ3tFwsy12KPyIVRqk+
olvTv+QOlIt4ayPL+cO3FXDNFmTRz487tPIXmPsSCUo9aRb3w8fc5+/TwsfxVXFcrt52cX/aflEw
Iy8mUQ1CRCYnk6xgOQ6Oo/qT06Qxvs4E+RSnVpYf/o+AX44Jfw4C4M1uuJf9pvBVnNMJbrauoDLm
bVhg3U43RrrxZ31uqbIAIAmpy7zlq0atOYOmZtfJpi2F7uRnIxhOMh+bp3kIADZTe1v5hTLbuva5
BNJWyVGmDpHIOFMrf/nbtfXQuFcycnglPPDzPAzFesZpqVx1ptsTb8A0PIfUr7tYOshc/OChb2kd
xf/0x58GH9HILQJpZJp9ljZfd/zdvm25hsCSCgVGgdR4xqnd7zP1HzrCVsRvQ0bvks/oXnY5eV/7
3Gk2laN0NL98zwHdmNlwYOqvZafTurkXFKGd0NGuI721o5xPvr6rVRlIy9LY+kOi78yg9slpMfnM
Is0KmmSrtk3SLzWOe4003U+RxoqyCeHNwPnqPFZQ+aQ82/uXsk1zp3O0rqwOT2pyoRaGOqsK/isE
8fQBjqneGFr6CwMhHv7OmpaC3NHNiR1PP2IGcqwafBh38dFOIQEK1sKc9h1WlepRpegUYv6kRpNu
JW6Ur1Fte3Vc8J5wKDmcejzLNdbaDzvEOLnaQjaL08auXX77NqXg3TZvWVQp4gF8uqRqcylc/N8C
nCtqXfUxEZ0YG8uzY0otB/3znfD6ClZSkRpZ+HyctH4cuJuB45Rer+5/ax+KE52vTyhniEEhGv8B
CAe2TQWpI9MHrSkFyYLkUrfgtFVBUzGM0uf91y+ZqphaZxm7zJMvEWFr86uuOKBhUe7yZF8iAbdF
JDJE+W1d2x3R7R//VvotoTD7kpOQa/geKJlyzVbJKGyT68fjzz+9Punok3h9MH5bZD+neaRE7Hq4
nILXikBzuN/ydp3UiBCRi0crXbVH/ADFj/5qdy6tzwfkKNc4qH0c4n79uTE4H4w5CQtcr3lsqpLe
jRJGEmOQlDx9vNVuK+UdEhYxKKY+K14+I1u8PZvUYv5EqYG1QsmXM3ZpSNdlguReW7CAYWYBbReJ
eil3s0dNEDbnDFlN8fESavt+BPypexROnBZZD1X7F8Yqoyfm6l2wmdKWJOK/ddxvT1dxIO/vKhoU
boVicWW9ty7wSSJONXyAxAI7b99vgXWzuFQAxniEgnniLrYF385WpcFf84Jip6zv0ierYpU7ElXs
1pvLUqZeG4HhzFmUs8WapVCz8CMXIHDO2O/dIxMU60SLtJgyOqb5K3eHGK0kM9SVkdV+QgBmxKjL
sFsnsDjoPyqyvxUecwivFy5VehuAijE4cFZ82eLLZN2eUh73wOoBwnrqkKdmNdUwazyIL396gliV
f4pxVpHTo6vKlo49u+1m1LAEBpWE1EvLiWTb8BtFcY9Ab5vh9EfGBAIQJVGcLPMbI4S6hN0v4ikN
CF5CUsiDIqqTh37eHu7Kljc4NwkV7k9enTybbU9RPLvTSExH2CDMaAEg1J/2Qo44aZ2HUoQLPGrc
eBvJnZTQF3zEM1FG8gqr1KdvRNNzoR2+gGaiuIItix97Pnc0DzCohWGqttae/iuEJXJSe+hM7zEc
+k964Tt/LJJK/6vH3GzCoM7bZtZiiIVAQAoRBE1fKWN2DpVz7xaUwBt2KebRoC5EDbL+ZpZ1NIwy
Hk3BOWvG8l58VfF/w/WKcMpSdCqRNRWXu8xUtZ8LRR7wDG3lCi25eVBf3cX5+Mt3lPE10hJTLwbg
kT7+CwDbsDZ+rLIV6iqS+TxKi/vlgGVrqDULYwhcgHnho5JeGzX4m48zaYPnLGTVUrimwyVZyOmk
IOq/5Bl/IwG4kurh3mNMLpW5VeP9EBYYGA2UCjS2uAxWn/KQRWELM+7yV6usibRr95W11zxIYj1B
D1exZwSmwy+p2MuQ922JZZkv5MUp/QQeT/8cQbhJr8RTd6UPtXnpzUKZZC0NZXU2+xIzOQK5Mw7V
Qjm8EMG2Tf9Y9wFo6eDQyiIWKkOjRo1kUxQMpE8bIeMtWtUix5SZCrImnxV5hsNRRY3XangIKZOn
nTg2vqbVKHz8fO9DtL25OsjSaCHjXaGuzocwtzHob2pjQHpaohixjOj/fG+JNYKy8O4xwqXPlYPQ
3VA8AfI/4Zly0AYxoFaiDnWVcx9b4L+FwWDIFCNbQn12jCXtriIdeav3/B7N2Bq7z9SccviMyeSW
nJUBwbt9Jmx+TswdOFzjcAhsL2kQCUCoqfyYKxrErpC2S/2qm2EzdSYLE0+hLdYtIaJzx7XWX3uj
tijBEh38jeNow1BPONnCZSiQyntqPRcZqdeMPF2AV8/VsEck4M3Zhk5mZgI5soROiRdIoEluBXni
YLUOjjPCYyCcYAbUeqyvhROC1512s7wbxskPtyE1PKTwK4QxofeLzdFEZbrxrHYTDpdt4mmWVqLx
MK+ppZM2rY/6jCr8MdKVBKCyJbNBB07j9vchAnEzE3aFF/6D/7xYWYB3s9SSKR20EA1Ifg4AJq84
Mv3gDJ8G+DXwuYt4O9rn7exLbRnaAraOtbhD6vcQctZzt4xXyd5cppaE5lG6J5H0KsyMz+uuNJG1
9nFuNAf4YpRqvWKdp9OBv9FQ6y/fhV9wquqlAoi6zs1WfCYmNudZfaX1/d4tSkp81sNreN7s7YAp
LRoGZAfs63YX/12C2OjYE5N3rPgEljthc18mtN79pqMeVKZvYpZ0UJqwqPJlAt1lbXX0n4qP4q5s
epWUUP/tD5QA3Q7kXZyqMtXwUOGOWrLjz/H8sX+TPxQQ2Seo/M3qAnrMfq4xrGn94Da6gQaqiba8
jGu7ZaII7KwoTa+l81WPFqFBOkZj+6AH/VdtgtAL74eHPwMo8pCfXApPcf9kIZpK2geUE4ULMBYc
sUNrg8tD98S2T7FOoc8bDszVTgU7bmkMFFn5p8Ic5NIW3s9gGQIDOmhY74eZsQbO0KkWwfZe/JnE
JSRzeLDmrxB/DXtLxSoYhU/YZ/Bxb41YFVTbwp/Y+6F9KmoPxQo86gxMJexzqFmsN0scrdoh8VRy
W2QCHylhoPnaw0Y5lOQUxsCYRMisNgDQLFLFPaoK31m0vIEsj/yjpFrkQei5CJ1BI72ZWGvbKANo
sCKLaZw3QZYe/YnjeytArj0JW8XYat0GMC4mX8MyZuGHIgRy/ctMBXKil+Zl6akgML1UeHQKBZP3
nZsKn4C6yGTUzDwdMRph7qn1rGruJBSruygHL2Zy393n13AQ0WHJRc32e0IWt1EijOQ7otcRmda9
3hPoBWToIbCHgC58ZiCrUANGSiUJ65ESKxXO2Lw0B+slGKYu5lWA2OksLZ4Wi4Nucz+lLn/uOH6+
+xcYe8OAE6NZ4kzDWpL8ZcDtSg6jgvdf5bn5yxC4gL3Iz6FnFjdWh9561Ns0Rbdhy6pBn1qQpEOu
ZJhmL5tt/pxoAGew4yKyiPC+EQPmIJgp9Hh1Qhxh1ls614p/Tn+3AMu9C/fQ70QVkU0Kq5w6RCT7
jk0L5p2fAF0xmNbhHG9dj+ywD2jdOe97hrQAfTDT24N/ekuh65UbozEk7a9oc1Qfn/i5AEhVV1Fv
mkRv4fpceQgYu6u9urW36fNcvdiOyZVeuA/Um/HTWK6WpKkD+UaC/UPXrZ8FjTNemyrVax3SpoQN
rzpgEBmjEl7fcU35UKBqj39GxCJjBC0vSMz1olO/v/2QUWntIs98dAVKaIYbq4MOtsEMEBNc22tm
TyC5+RhD2tSlJgwz/yChzOVtFR7knkLuHyZECfmuofHGqCs3u6xcwGD6frFwexd7DKZkSrf4cOw6
GTNrYPqmp+qbFgWqvpNalWd83vvi+n8A/jD9CEYI5ltGyUQBQZWoSzWZs1D6Jkjopze4cpyl87mF
W4oIWPI0KWbG5SHGeDTBpUQhMGwp0dfBy7zkiUDYhsZx8DH2QkzP4u7NXqUjCQhLb6ylnO/l+3Iq
dniyO9JfTtte2J1NaBx7HUfdlOodSPgozaUaErl1xKltsjwCTf3aH+sBM8HuLvbaFATGMGBNEpli
d4HFrpysHv5BLL/RQEzqgQR02Y48ueKg1JgeTQy+b3W2n9+lvDbWasFgNcckk/XjWcEbhwqkCeAB
6omuJkWuSzqoaCNDnLE7/OmqOrceXeXoHcNwu66NPQnptviWBnl8kvV18dndC8PyQxmz9DKdpNt7
OVJrIro7zGvGLl4RHp83EpqgUSL5q0j/pIJtzqBqjtYzsuvXzwMtRO7mP465uloG7YKwX5h9yTXP
MNa1VhZRvxuUBfgEe8nI2ZDtNBgHWYvkGzKwdpgfzC1mj34lvPatpO8xXcQtquSaXsPFLH0A2HKh
mG3I7ygIXyj8PZN/h19Kn5bQryxrhI0YZdQZTWaTaAxanw7Ol6Iu44Tj5CKjDEvsLnP8t75P4zfK
A6NOQixkp3a/j8W3NDkv+DUwrUA6BFddjw579EJx5G0t/W6Su9B7hr3s3WeZqQBJuNNn6WkVBUqI
cFp3RV1AOIzxj1lGNYjaH/aFzeGmZSD6S8iWt+xuhs+LyS6Nz/dDzWme6vaw7a8I5rOd6Yr5wIQ4
uWwSdkrU0cOnYv9TwpbPn7Ssp/ZN2upNJA19i7Hz5V6yZ+fTLyMUsV03txXDVKbNBNtzDmX/Eh1C
tgwutjT9ShiWXTWEVzmuqJFJgUMNA326UAlw6pxpLCGShcnZ5FMOx4R7PW6wlpAUgHuVYvIAK13C
FpfpDaXiPODgAVLZqA/pD6clYa/9gS+DGpyR/UnuGq9pF5NSCVMCsv4nYUUM1wJlL6BrCbmpv5R6
gpYuG1XOsNZj269j+XBFFkM3DXUfMK/DPFLTnCBq/YlkvqLyTzfz6kmug4O+3j+3XosS8jZAugdX
1giu1i8yYvxNJEDNIHbWsvfGQ2+jgytVTqMARr/cgaHKQYVfASNDDP3jpkX1tjG2DR0fCr0bJ0ed
GL+B+DJJHvVlHPPcXvC+vA2S7tISGVRhrYrjk0VB7mI9xBUZ4b7ObWss2uNbeo/4ggZZIn0Z6up/
ZLxuK5lPQphdzAGsizvU/cki0B7KmSt1qs4GoBSvKFSI9VJlV++KbdPG/z2hVe7PPbylSNi6IzHm
6pRVqed5fBpAD3EP1S3dNs3OeoXXL1L5LnOFIp0SpiJvD9PTnmbXHSuXq3rrgPUZ/FskctAwAVE/
Ow/COPSY/uwSDM//ahsbPR57+c+4W+9OGfWMPx6nvL1kpOhUYTm9QHKaHEvpxCYPGbNKLX0wiEm8
VWi4oIvpd43ZS6IvsnSIt0gE1chcObMjkROSXZn9CcyJx+2sdCNzJ8+0M+/RxDgxmXreZBw/u/hR
6o0xJ7eivXfHW7OszP5/X+wlx0dXC9bU5/GdlEEZ3gogClPxs2MsqEuMTr093xoTLigyqehgetnz
fIsQsX8GQEM5+mAJEOZtVTFmUqRaYpcBLtg8Bk3+nnc7BYK/uU3ZW4NoV05/Zbg9Llh52sXMjT5n
fCjJ55Axx35cjLoOZasUappjMchd2kodhBFkDHmOTi11A6ENAGCixkMirZ69RXtbL2uITn826PyC
d98gkOfDnovwLrU3KMmxuTSK67+sYXZrKTAw6XcPxQJovJePOxIbDFk97xSGIB0FlCQxiVTBv0nf
QiVPHa20J9otGJVXPElkp6iYw9nCm9VQyB/x1t5pVUv821Xvrt0bHWqq6rtzxdGJxTNrTb7EOUkY
faadss+6fWcPlgBaWfZQd84HtPBwcchUZyEysH4ItWSXwR86jNUURsw/+UEVD3dtTkGLmpruzJAa
2S0FVD27s+woqeAolMVkqI9hnBGDScOwum8cO4SCOFFb2E+HmajtMiGov59qvqu6aSMgm0HAfP/O
qQeTwMNj5nI5aj19nYzg94FGr88cq9ffvkfXzi37AySR66dCwvTrXmPOMMc6X0JPghevG+sDtO6k
UXzXmT3F4TAaDUib0otgdUyVEzXLrzKbam1zDrR4X+6mpYR07VBa6zj684AQa4BKCpKPKncaHNeG
SUOLXls9BkI6jIImnPdUvqxcBmcqLUxZro9/fjrbxIaptP9SBvD1WjdskyEadcQJKTXQpfyvLz18
iKpQ3yOBGdpLmLqy9w/ftr3X/vufcA5Amp4nNBzFJVr6vuwMjxpDMhTmiDuy8OKh37EzOynRkMSy
lPzCTz8SRPcQ40JBCG+KSJHMeajwk1AksAVO2ffraZjxuGSYgBpVuqbjqsPVaWL3l7KjKLKGYBEq
aDnAAWtEIq6BVVV1GS3ywvS/YgyT9u150IYupV4gsqjpfa8ulaOASD0tV/8z2qAGDpIHQ6e9qgCa
Zr23xI9a4OsTmD7X4BQvWjViR2GO5svAd1ePPATq5x4h8dEbD9QMfB+2ocF0iwjCL5YIu6hLZG7H
9I+5e4tuq0V9nmfGg3bYXh+QLZwBe9NtzuwQGjatAcpT2eUpQKOyD+qrJ+zl4/QRB92zYAn98tU6
LV6ToEP2HXnHYk8mekiKUXObucnjEfPLHAXVW84959i4rvWHW7QUMvxhxqiEEys/ZJEeWCqdTWCt
m9z6SWL15Y0XEEcf9hPl87peRRFkSt+pAHnjWtqDPBt2Tgxf8EoYuAsZBE/yCE/vK21Ec99PSlQx
1lYJmbQHfhYgTDsRFw81gV/3afwRT3Z3cc0A0/Apbm6rc5GpCJG+cZA/9BXpAJkm4E3kfHHEAYG6
77hN3AbwNQdik7roWG1NDdZkf4oQLA4lng8S3LzdGcYD3LS1yoy+O/zODNlj6pOYB8PfOa2s+Y0U
wrdtS2UNLFvHTUtD4KbfjX5lz26+ywMasKctw/PLVUHrr+Cg9P4FFgddIdcgKMcphgbgMpPBKgbp
cLwMCtOmeFY5v/TDYUxEfoQlBY/cmCJE5/snwuS+zyn1aXR0EsYMVtdtxC3EhuqxB+3S/VNhIlIF
v8WFC/qtlT1y1gL+Vun8b9gTUJDi9Xqu1E9I8aweY+YtDZB2SnticmPbS+I0GHsWTTHoDvxuBZLc
VLJ5b6DiO9OTRPR3SFHd/XY1hvyGzvEMoJUcb+K81wLHIfDS4QnfsN4NUwEP0puWlCgpcwXQoGGb
UHEMUL1cY9/J2ZxAnjZtlXVr7K3vmyHLFeDZ0UAWvaiMXS+/Tb+hCxH74wU0WDr3DL5JA/eeUwun
5YCcMvXD18XOlV3UVD1QjgbX5Z8AviJB2VEWTSyyYcsjUtB1WNyu+TK8I/MqTa/xUouTs0i7W8FG
zlNEiYzveqPOmHsDc4mEkARee0bkAdaT/R0e5CIaFxpKXPbs8com0HxOhGTSgsFXD+Hr3Sg1p/qO
dyw1ySwhwCDrsgt76HtiYauZxY+er7k4IJ4NY2J7S5dif1KcThJRAokGEJZCgvQKsaPrVCoNMBh0
H09GbCIJXLb6NzFLjGz/6/ZDF5XaPzzucqnE+hsDQHx1egUPsHDdyV/mZ7IflBZtoPyFuPthCa0Q
BvdRBmGG1MV2fZj36B6JcpwQPqhcGdEtRGNzHCgaVdFFwL1AxBb/c7UPwtvNTNSiw1z0KrF7i7rE
ZCKwiHgbU6PbtUmqht/6gwGg42vFp4ZiG9WcaLahQYRTMJIc691XDOxjp0rmthEy2wVCulevocF9
ly9fXHhyecmKxboBlYKGF+VIP9UnI2/aw6vK37UkKHBu0cm668f6H/3K86hFmCwFxy5zJ4rAK/0k
r7Zq30JALH81htcuQ1Pr6x26RakD0qGLdr0e6ga1pOJIqMIrUdPzNH8GvdbyrnXks6XxbAJ/CS7I
n2LIxWM/5KltgyhbKyq8ql06ZETSbFa7FVYy3tknVIAiTLIclGTmHUfxmV16u5J/ajO+MIQ1nama
3K3KXwEE2oeedvzBWqpRIzx6R0evSiIq31isUNzp0gW8VfYQNZQ8mbGdB/YuGLx1ZqQkXrME4PqX
XankarZwP7ootjSBN7IxzEwKpaxDZbp39oCjTrx7Y1dFfdSAHI7WTSXbRlHpLLRwqbb6ooQa7sYG
nvbvNRjS0mt72hIktgMgRZLvmMtvqVKLEazZovxNR8su/2qa87MmFyt0nkFQBxdRUtf9WXBxWoqR
WRwp3PcVWaQ4Svt9KNEj047Q/F/ADY8HTyZ+QucgCdFirVzzy9AFT478+Vk9u9H7SiTFkkrF4eyX
AcrwaoEyYVxCw2SQLzv//jqKhwXfqQCLWVeaaGZ7yUJXpioaVySD5G2x1mAiVWFxeODsjDMjs99U
TKXc7Xlw1kePYHx7LMnfMC4J6CzUCOzONCTMDezcwku0cZWEOL/7QyMeFi5vts3i1J1oE4xSef5j
KdKS0ZZJKG2Z4DdyYdzGj7D4O747djax4j7f9X3K6MeVlQ4lDDEjtXtRVNkx49EU4T1s54KGwqKE
PHBjzYqlJnOXKK3UJL8lJDNGDYdngylrfrc/UAXAu8/5h2+ON3pFIHCFpfztczWlAuXRB1no8RKq
p+mD96AxOHGexI2IED/L23nT3g1NM+GkKqtWZss8cQ5qfxBhOrccmSoP4G0daELdcpkhvV6W5vmM
2dPDXxnDK/oActipLP3CXHOY7o7mjxCwZ9WYIKfQ3QQdrX4KSpz6ysajmcWfpiKNnzq97R+EQ8+6
DL6HvdnvpTjR9AGlkgmwA9Pb6zmYF7D7cC1vi5kCRgeKXK5IdwjMJQGr+EQLKhIx2xXY5Yg0L8Kj
CisyuVSsAADlcr2TJBqMeA4oH7l0b+DQBx9toDqn+ebjwwu1J0izxEAMHFT/dXsmNc7x9o8Y5wSj
iNQrc2sQ6+I+gCRw0Q214rP3eqWWZ6QlQ6bIWV9bMI7qyGu8t/GTIh41bktBfSPOzdR8jPNMhVc3
K0F3YaDmblb3h8wM0CBmgThe6AulxYcRy0BLYhccbOU8f1cCUa3lVmpkR/Q10GMnedRj8UVLgJuf
PqS2jw1HpasEkyE+9+XJu3zIqxN6FuscQ/rOOyga74S9LbW2K284/2t1umn7uKYTGwn8FyFbOHGC
Bwis1L2tlqPPmGChD9qc2WfVZ3E4g3BzhuoknnRSGjAkk1CHC9YVHeY2KWMRJhuUgYTwOkx06nwO
iKo0woLSKkyD6eX2ZcT2/967a5IeOgBb56CQBhEkeLKoG3y2eeNb7Ztq2VrsySuVlebh+kT6xT+r
Loj+Zv3xLFfzr9UcA0uouMnkYIBI8cDxyzQX144CTjothsnr3GSvVK7ve5Sjt0DhElCj1em2aSVp
sEgJE1E1YmKlQlnf9qOq7WWpe+N5ZZCJmFaJX76nDZMjuNv0KR8flOQsZZnk7jNK4kVoCHjvh/tz
Xbr/g8/kFH4gRNkxjCBzFZHzo7nG2Zz0QgUNk0jpUcAV954UHDZu8Nn20C0tjYDPIjceS9f28MvQ
zfIDgOlzvSAn5aZbzoBauERaBSrmBA9cr8Vw99d/LNUmcvOQbe1cVACWO+8Vx1DN+TYzHBESBwlq
kW4EBVfkTPTQVVa5eDgg9psN9RJPczVD3xxTCsCFPuYozA4A7ZFxk2VPArpWQmFgFp9QwRERsJFj
Ziiw+f9YSF2gL8I3ItpPliPJToPPWwmT8j41IgKrqfo18IzEpE96k4iyywVprNvco+ZNc8RbQfW3
OqOHa5eZiSDmhj9YmWupnss26zeuLmjDbefjwWgmqYRELs9GhJUiKkwoFNElFMXOSac4VlauncJL
LZpWoMLJQuzg3X6A/tntxpQGcji60F+0j15jJBvM8nPxMa1/h3gp2NB9f5zk3OyzNoWPPM5k8V6v
v8/IxPRoeUdE5nit2Mozr4v7bd/3eJzkX6GCe8pN40WgMvRl6bAjyanrhJIVeWyIhO1EZ0lKDLis
z27TUhjF08+XhzK/DoUQ/jO3r6prfQ9C25toUfrzjsrhnhAnOP0Bxs+te6hknr+y+D9qgSAu5YMc
dTjXxvtPHEU4ilUYqwMA6I1aq9k5cZRiBn4g40NAl9W/SqTmSHvZSaMVul+eQ/UmGGGUpX+VjHs+
gUSKP9fOn9VCElZRI7VMJsUjtIWvdEZwSPIsFwuhbI6Yqnx/xtTDdpAYS7CCYcl2U1K20RmAphl7
2a9ecTmmgAElXSpmvD4TzCef484yNDLWiFGk2BGFG7EJlZeXcG7zRL2kWSz2dQB8hgtdIOUfspqu
3Dyve/EXYzf0gF2Gs8CliMTVOQse4WWDK70WSoo2njuhAedG2owH+FtdcpNDvasQ/T96++GHGJmw
1r3jubvY58xwq9XRCt/4AV2LoueMjkJxBZcMRRp3Q0jtzXqUfq46p3obNVE8JWcubQc1Ow8tqCcJ
Nvl102b+6x3C9hoeEs77y9N7WLVZpKpkJ3Sqx9sYVRQu4Im69gipSBgCkKqUEj9lQg7H/uGd1B1/
Afl6D1qGaMRRSzswQ3umD2UdXZ0KPi1au1eVtxHg7vhxjgqxjC1RFx5YhChvjWmW4W79vEnGxT3m
69GmA/PqDsOdP/wJk+Kz8etEUz7Kudfyv5WGdCuRO1kAGnzoSewjK0mmz9bDnZ5WiYQ/RdBRPF1f
6rM+qfOzeOP1jTNHSj4GSG9LoOOdT/4AR3S/zepWBw4mA5yqQnw5ded5UOdyA0eMKm5YHcqwuDf8
u8txOfFxY1BO+Qz+je+7sd3nRSU/bylxGVStWat4ASw6fV2Ux5gBLRgsFDWEMeGd4J28RfSPXMp5
MKyupKT0B1Rvh5AwB47njPt9moOAlRhErrqI6CJiiORxMmph9GkbTAGdclRsCBvjyKYBC/uIF2Ms
uNRjRgYOEw0g2DhzHVXeZOdCuBa6c2+4xScdfllVmtrVERXewDVdkN0yAhc4AR7F11aQvFs6M88I
Ifzruk5qK6BORaYlaj50rWkstVHh6IvpcbI0ZXbxMOIExjXdB9BF9JW8EpHz/eidYBNO3OGrYXLI
DhWsUU99Ndbq3BE+tcB6ywc7PO244aUJhiGWdMfWwbcFyN5pArG55bP8EDiljhctcF12RVSsbczO
ATPT8eT2kjh0NRuGkGXDTAQ1RxVFZ/P2WlHDMPnljh6AjQXc0/1f0fZMirkRM0rALmE4NON1Iwfq
Qg+c8sueVFyaAgRlHz7WlhidvfyE+y/isKf0B/VvoCWePIyv3L9k+Je60Ms6cZloa3mrykOWOH6d
QevF/k7Julb0oVpirkEzD7OZtc5hFZUcZisJ/YnNDF/Syn44TSywZ+k7NEWp+zlTs93kLairjh9O
JMr5bBYLfMpO5AhQEDHcJMpozhpIs49GFZnmP6s0Nc++eRlD0p+vXbVmhsm/C+76kr5v155uMlKI
SIDBFJPhKeLl3y8WAdC1HTjjQVR0AXms0J+MxbOjxB8qAy9+Lbh+bqasydLW9AlU8iUkCN2uG+u/
WfFPR+zWwfi2z1JZF0iO2zZ5WfA+mSIpSDjN2vVHQfWAfwjJxdNI2r9XYA7ZRxNF/qfRcDRcBdP/
Un8F3ACbG2MmA+KwjNCjtcKplwNONbLy7/B0lN1clK126aJvRGxBelElBUCDg5lBf65TNlg3dU0w
HrRq1FlEI+rESBcwPFbhiIlI0locsKIM7f3o6nyanjYL6E4sy5nCXWOT1nXtneWnc00v7SateDZI
XV7zgd2EuPGpS3hTtXPGDsOA2neF/m1Z7SaoH3XEURz0e/2/g6jy43a2S/PQvOOBAdfw+yiYiq1L
w1ajB0WwFYjMl8tibGEZPXjmN9c8nNObShYoDmjBwpJF1dq3i1jGvW3mc9qwMrPq0b+dGDkxloQy
iW+5Pe6LJrw7R1cvfxnpszkiyTLwMUzL6CvPAu8aIpazthqIPaE62VpNMpf3r95FQhZnOInl6pID
dSBVbiQjKHFP2Jde3b+uZyt/SP1tILemOc+s3juZ8pYu3XgqCUgAxPpatyviwsgkK9/IYglnJPIk
TlI/YIDIZtRdL2W3KPiqzt1DG1pXUvg8VjBHRJ+DjR2tfeTIqfpTcb+3m9jq3Mf1NqohnPPHgOwp
p/8PAgq1ePKxpdbFd8qKtEGdZM2h5/wsV2HHWt72Fuw7Bf+FUkCLgbkmIdGugfonqkWVE+0OgFch
oIXJjNFe4v2ZIQY8UUtNQtLltzwhWUNUROfEKp+YU1Ympjaz3pvDV2zk2bH9WiFkgysECwcuuvQh
wtTZs9bz+zsS5P0YYdGFJjg9wwpHXujpLInUaiVYF3xeV4swjEAGijozmLAF2i5HbZmkh4MwECXJ
W8jhT7udzUDhDkGvvz9WhTBW4RBoNlXO4DWDOIO60G41jYG4+PY8bqFOeXGH2wsqJD5AObdrQrdg
1co58GMyYaw+z3qJFuwtROG5D/PlBTBvW+TPHzFVrRz7mVyAgMNQhLihEM6RscLpJohcO7HZ+jNz
vaYwB2CRh4TlihWNFTEFr31ZmnS2Djv93LHRVS0d+zjG1mIKOoGYMjdDX8kSt6Uf54DpBdITHfw9
+ydYFgk4MprlPiYysBZukq6HcAdL84jM8bhDojKH9eQJW/QOfryBToSXLHRYnid30NL1T4QAmH1g
BWHQnhhu3IUy8rjSBH3Spn8xVSunam4N/0AP5hmZXCktyNjhDl8W3UdEUvoWaHkQMSGsGuqGCu3a
pVdEZTtYRnbiGR0olKF4xd6o6Ibwo0sn0jbkj1b8EOcp1gI9wwv8SK9Fd8PYg3RzfPFneJnBZouR
L22pAXeGLRHUP9FNODFn4FQZT67ccuq3zF5/uuvsUpLHuNAjPwTV5f8W1isXNb2J+/I4h6FI3R5U
qO2z9vWsavYm/bQG4auLUTCTtcuO7k0OY6ULpm9aumCWFgWGj5vQRHZDTQL1ejXJud5FtEQ3RWh3
oEH02K1j3Vof1Aa250ISAHxjQcngTnUcE1wh0xEhjH0m3hFMZGDa+2PnENxa903/YiTCStWy/NWw
72wj+shQudKepYmt1ULrAVUPGcZySonRfww+C9kySt7tFeX5hP2PtaTWhTj3JTR7a01D6O0uPfzd
rc9EyKVw5KigwN8XjX18suqsCSabwUyhgd+815yUFmZJgG8bebDm6lhstYFR35iYHUBNiUCnJoRW
ltkcOwgQgkJY4Q5mwVwbKCu/EgY7OFCiXdWEH3JPlmejtEGom0z5crioL6DuKgR29sSSprLmrGu9
BcdRhee0KZXY47I0H/abmn3BhxAilboufypzhZGLgIzxX3WS31c5D8TymZHEhBN8enLnaa63yy8Z
H2wl1tVopMNuiQ0RvjPMQxSBh3XB3RlqQdXpeDFCfxcoYiV1R4JkYoN2KRoLMmtV6WDjSolLf2PH
rRdxbM1jgds6Ehphki5UZGNT4HLr9rkAGOz6xceObRO7Pl24tO0RD2lPEjAsds2zIJ/5YfpDcKxO
FAjzfCkQs4tqRteIC7bgW8ybfxPLFbxfHi2b8qFj3VjX/VLc/xpJakvAkrw671Cx3FlfDagOsxWm
CPzbnim5xC8RaVu7IRVKtWfqgXGcn5vg1AnWc/DFUOAudgscduPvEABICAx6GHaGXIIVUnuFPjdX
Hosn2P8xYmqiAFzf1Xp6B4stj51uIAAXecixaWGNqTtZzfmTa9xhBwJ0ndAucqILGuISYGFDoWHx
4fO5/c0ibYYZXJwV482LCriYP46r02aueMtG1A5h87X9ycWGTeq2804b3TP7LfN0W+rtwknaK6qr
XeqbuPHnhC3o0nXWhy+6WWlRRbJewkSU1bAH4+kPjvRrtPKnmcCaNGuM0pyUZJiMDtgH4qwmsJRR
vKHCjCEJHzKm96LITCMD7VX3pVmyC0KIy4GfGZ2G0eMjgiyMxnj2zNzy9Xw9ELhvxnerFndolQpN
v1ul1YhohDQQ7iBgdbSbwIRAbJLWVfHDf69BAXuA8GrKBIDzhKquE50gbCa1+VjBau3mFLm9BoKQ
WMisXcwwjloPvjkmLOzfBXvfMk5xQfy13Fzrm9Cpb1CYG8t1+7UhT+92Gc+ZUK0DfOl/OsHJmHAw
ngYJlbBmrsYMueZevCOQTCgojB0gN53SXB3rVMFVlR9n+1SRrMeFVZf11OczM60OJqHXEUvANGVd
hkHlbjtZ2FlmVxNidr1C8hOZqb73jTWjHFoe22zDALUNpohDWddRH74UIkb9/NHw1htYXC9oUsV2
bJrLpZk1kg+JJRdOlx+PjmimV2OqX7pDJGZ0kNUe+kgIJXcOrXu6hdMVK1jiDawxDJyRvLuBskLK
5nfdLRL+7F5F4zZngA5ycSs/OCSsbpcE/1RX/vWTe1MRrC+EOTvQ5SbVdhSrhEejEOd123Ixrge0
g2SNcQk/7Jp5fw+8DGo1594XuP8aH9QB2aVedqBwG9lWboHEV6bhoMw2SKy5RkmYWiG6NMRzQSNU
fI6XqoLRzhwouzGjS1w7+IkbyICBl7AC0vWxhqR/ytANyVcL/qwUrkyh3DB8wUZAwH/yiBVk05I6
PddgO7at7TNBtxeJQSCjPouW4y5vKJAb59pHchvQ0iIWRjtIE5UsBjwQ7KB7bet+xPIUHpRs0IkF
RU+fekS8QEvvW31+OBU+EpUL1IIhDjoIfOmYzbLUku1eLq4hM0g6wngu0qc94R5RQeHAckdi7Vib
nX8+UZ2bilJY70iAYOy+UeKDFcB3mtPnr05PDui+HQCe/T134IHDw6efBj7EzI7Fvo6KtK1THMs2
W7WourRhRpc9iXXJMDQsPRClwuiX6poqpnqSYMomxFm0tvITtWvODCxK595ow6NsFhzEuxKA5cUl
/HePxNbPglHEDPvuyvBY8A8q110c7TX9Gv+mvJG452GaU2wW1Ci4fOLWrU33ShxXiDTslyg4etYC
I+Rrbk8epjE4WDQmOxbugSwF+JGDZX0TxmwHrPXL1jxU4bk0Jv9YjCCn1uswIGasYYOFSGlizrVs
a5Ev+9Qld0XgsvCiW0l+HGi+Fjv7eMhcnV/BFCluwECAAKZi9WuFY0niIjpJb6Zrdmyh4quvqAsk
9pHhSHqAIvpZAbVaoeFWRlpLewXOtPMxYIIQ0QnEIrPXwkWmyrDWimNrXrn7KfHxO+CDypLvzIzD
4lTIryghDE/jp6xySHwDI0DPvu0rJ8EBreHzMkmIB7W1XuFS6q4N1HThw3QsGBj8lPaqThOxvv6R
1uxmBgQBz38ci/nKd4Rvm3POyWXIkp2vsTcg4xmj+IGaC3a1iehb9vvGimpP2uzQSj3FJGENV15i
UlutjzR/EGcBV/osRZEnw1EO02sfJXNRyJSIrbuEfDW0G9CfKqQa1HqIP9tDugR3sENJCjbjSLLx
F+/jnZ09FOLvQKNhnWVQKarIKx1kBfOgSdAjaQP39/TgYmPkU/GFylCZCWU0pczKvE/g3juD36qD
tORGoHXI+ugQWI2/XClT95e76XomOIaKAQgCBuayF6ozmUOI1FvAmtcOdMC4zEtL48dbDIwP2LNy
5XQFB4oLbqMnl/W0gg+9Wq2BEu+odAkh33U1rDtzaJO7kwiSVO65Ty+CRn5gmbYFqBehk9gDPrnH
L6A0j6yxuFHaFelgWIpymdXU20epTSfjRGbFJ9C5b1RzSgc1jYwYupAY3aKPdORFShTk38FQXFoe
H5LJo6qmiPqRTXnaTF4+DuHAdhQOrFjD2Ae3KtKmWmIo67LiZ3kQZb8XMIjzv0AGwqSeEFZuflhR
+8w2ImfCvftlbIXFmcQE/OmdPLcL4PwVmSLVWOndbVXhaxvcTKxuTwY/GlJBg+D4AFM6xXNU6sZG
xRzRoQ0H+q2XyUEH6TDAZmTzZJWIxbfxkyjNTZvwPfyISkXlj8/d6WfCXoiCLoIrnBJXWD67FuK0
kkk3iqDbH3OmKgNOGdeUa+DGTf4fSXyQs7SOoNZon40NGXn4hQVqgyUDbFCbWOGOH/x3J+razKeW
U4p7R96Zks/M0dAJENQbX5Si934TV4iT6s36zuLNsKt0GG/89C/1uniZtQJQx1z8/y8rSE4aoNgW
uEd3lqyIoX9V2yth0unUdoqPxpI67+xMAdgUQZF8Sl0jrnaLrV80/frTOPgViptsHwFG08gTt3dj
VBM/QBbodyhjCDGiTe/qC04zsDleMtVWSU/vLFmghf3h62AEuQzTKOdofr52fLh19tM65aNiv0yH
i1X3FzThMHgXs6cXCqSVHQpWKRu3UsRO/5qM0rDiqKkSDB9iHINOgup614s5S754FL6ibrVD9hl/
c3Cw+bBpI2Vbjt8z55tk9IGt70yZ0gXVEAHg9E1/7c51CfbHkgmeAHaGrDL//G5YQR6CwUyaWfCE
QRcBwBdZ+UBhUajF+dDsRlXKNjKWD50MonUyhfxDk/6RZAjNuaedn/8z3eWXbTRkE8ijVTSjEo5r
kkPdRc0Z7HiOP/QZGPm/hBAIaFUd+UAX0CAKzatABkaHOvBoTGIEy2DXZSto5WTbi0jV2aZYWukM
/BY+BcE97Aspd/JxB5UMP9UZZ0OfKHd7NGO7XcKUxCqemWt7cucK/pXV3jXSm0ua+wOny8Kwmg6b
jtdbvbiCgEwg41ZZiNH7tu+ghbqkTQspC7towGrgA7NzBFBPSgHsjQuTR9fEwGSLrXZ62NCZ/c88
VobZ4+j9Ri+MMIysQz5A+tIP6GS7k8hollje2v4AF8yaBiQsu3XQK/wsPNWJSS0iA8Wr8JoJNss9
/MtujEnDwo9jKjYngp3tRapxzeGUjOnWRBq5ca1nsVnkaUD1TVjR79dYkPSCvx00eeX+AnqPFJZa
DoJ1yfTuXj6i/HTAwYGRdY4I5+g8f4/r8ax+qhNCsfvosTLFHtDYcvptGkH2KsnEMff2qy2MaOIM
sxYUxlvCBJPZPfozOVfHyfJ59Zw093Dg9R9/wZVCU+PXo6naGhBeqm9uxpgkGpWNIDU2WhNpVzJZ
NxpLfIwftICsWaU6D/dpMdbjdBjJOB8EnudWnN31xuMsWJcPflgJUHsYdcVibX+9DshS4QVmgbWW
amo27IPPWgnrZk3FJZbCuF+gYQ0MH1zz4UKLoH7vtCsTHjZeuJgmm+vxlRh1sU/a/KL7OFh7TpSI
aFPBe22a9BQK3nukILA+iJdkuuLeQe7u48QvI+Ei0j/hciBBVQlvTNHdj6v83V+f0lXEK4PVIGyZ
UQIbx9i9D7ErteGDca5unYvpB95JwjDB8p6BqmdrmKfJnmKOVZrPg+vgPOYVU95PsWYT0IgJpbUt
GbeJdDQwa0Oz1xgX76tQX+0bAg98uht/pfBNLT2Bgl9ENtEd04rIFN6nLGHmChTvKsZi/LeCZLCe
eiyuy/RwLcv9kqWJGwYXuQaF2DRRpBIIEmMC5Ap9Cx/NEwM3JrN7KnglA2b60ILMduz98Vd/KBoR
1e6+aHJLsaipTnXY9QVP/GEaYkWBm5Aezdl+ox3Vi2Uo2Q9jGfnc/SXRZKHFIhPNDjGpdCeeI65P
3Vte4CapqKulxnj9i9E4Y7eAxQr75Lm6oo/ZQQbWIIMNpcyq5Qd8gQ1xIYgYIeMbOR1hd9h+SzPK
YENLm8YHom7VVcdQA5SenWYgy6WrtSqBkCOVEW9KtzhEob3qcBUDS6qzdc0eWxdhswmjdKGKHE0d
5Gf1SV01cB/TjRKrqjWxBJN8miPVOoLnJFH7NtrZspwHhkJiFjOZpQA5t20xkqidqgfmc3cEiTkC
H7Ceu88Oz66gIQhuM4Oq8cbIWHHwYzpEO4qP8VbvQYgd2VgQC6gnuVmCbAGITvX09WxoYtoSuM3u
72+bCExURjbXxstR7hM3DkqcHFs7Z/hzUjTrJM7ahoxGN0CW2qXHRy52eMu65kEv9SfCxD2E4iTD
+Vr9A5lUSTT6zzdubqVsVOxc5xAZ+bK9eQGPVkI+t6Nh54JXF9ql7cCDCfbrHJSnfQEabybkAGHk
uF2zzRWX5IPyksWpsDtcJEmn0tjmatkHlAIGDuyb/jy4FnxfTlkcX5ae2N08724+fwQj6p6u0ixU
G6CJ9wfTncYsGDT7u9D/H2PumVMDShTNVGVASvfitMi8kD+HWdvrYGs0JOTGWzODX3ObU4Fbof8j
xG461BWgJSXln4J2PryNTYTxZtJdA8ol02kCtTrCNkQXLh+r1iqb77RfPhh0PcmDGDy+y3vrDaI3
JvqmsEiG19l/uS9XTdaSeDRgUADs2HZ/nr088ySFEQ5qW1AmxtwD1VlnUlp1gJcY3Oz5v1KZ9D3I
P5u2l1b7g5QYWnflu0PQ+CqqElBgbINR3qItjWahQgrXGbvjAmnNlSrSZHJNyt5w6lLOzdV7fvIC
wVVxAETug+XlLQCvIQnr5rYC6xuImMD4s8YEI8W5HW3Ao0Q+XvIAz+I2w0mjxkFIpTNxXshHIMgl
UwvNAvl3vLeLBuiSYqf4LWt+bAwIjpXCsFk9JnXblkjsq2yyJuidu7v3QDTvod6CMB//Cym9/4Jj
WjOrpk83snkzkx0IAtRK1yJOrQkQO08MFUMpUqhUJFsWsAiVoB0i5BL0VpztQFUtKLK4H3plFFJl
/iN8YNC814QWa2tuXEQKHaU/8qUiuM9TGDYXnW7HK8YpDmHnOmmplhRqFxhB5Ppa8tujyF88tV20
NsOjRpaBHf0KQE1Q20jXAwqkgnST/Q57liL6MtKNuLwfoQndLqCxmRDnxRm9fvZGN0OJjNrOLoKR
Ds71mqMSnSYdGSj78ncyUab3eGenKnM5Vw7ZiasVgvXpCUtH7FyCBHrgA/2Z+pH7da8d3QVmZAN5
abImNFFZ+jLoI9Hlw04x98HkEDzA2O5ibkIQHQjmDuMXCvJOLsnOx6SFuNr/kZHjQNbK/sJlj5gj
oxNDjQ7nEsPKHk6FGzfzTjMO838rkU2rriIWupZoDIsQpu+4Eq5OBD/vzXiqjNEEpcT0XeRXUv0l
G/WiLfqsAylWKmkGKsnEHg+IuedfMnftoeYmSPk8uM59tiGH5S+z5UrIQ9kWWv7402snmE35gtN3
D72tkPTg9cLqBlo9HzALqEI1DrBMpjegOhFVWs8ReVoraB7N5WRTiKn6NjAudc2IKm0fgkbWKXxY
m3y4kEfGsJx4TJG2IUe1ORW2LmHAjR62HI+h3rh804zafQzOUxmkv+2Fbig7mVhsSFCOueb3BbyI
tfScF4KcvBQxygOR/ziwk7T4Ub/baoOm6twOx9SstmTr3BCaWC6MusxCluLrUAanvXRYZpHXGg6q
z0jNvy2fqw2Bhu/ajHky833iwZvhCaHSN1d3xbVRd7woBbjepDsv3iQARfs6H3FdOT55eMFsHnep
/Awm2cXMm2l28NtX8c31mMa+W95gJWHP02K2mxlL4dBRHqB39NjaviKqqaUjfLOdoyyJqj6nDPW9
6XTSzhh/3PkjaOBJMr8i03v9gHOVlcvcqegzKvzUQLIivU9pCvilwM2/PVyyzEA3Vai6DEJ8YJ3I
kr2U8fbS8CCbVxfOd0OWNNfy+WG2IYXrF6xseO+znL1bqIw/DF6lbokCEqn/0yCvJ7AXztrHu9Br
lIYcHt9N5Yawcc1z2qYz8H9Ncgv1sTfHIK4hBagXfKTbBY1RTa2xTIiWPoIeK5EkpWjUEySAMLks
D68rcZksU+hlsGGfUsTdLmWgf+Ny/2DzZS5BSwfcwhpv/WGvYN2Ya7hDoCBdnezSJvrCTIduvQVH
LOQqoXQfpUiupVKWU2qrp3AWMuVtmMZoVH6SHtyTJNzH24OG7Qk5MHKwItKCCQQj19H0xhIZuzUx
1Mb4278K1TG4+kJ+JaREfhwsnc3YPyQ/y8Jliq6TefiZTPO6ycssaPwuriyaWwTSKmworWfO68G6
gv8fuu1Z7uI23chhNzea8gZkofxhrWzR7ZTy9dbeje2DRkwN7c0rcOXAmiG7QV1/0Szx2IGt9bTE
0bibgwKB2E8LcJoQZ04YSsD/4XaczeLFKz2EyC3MeVmI9N8uSxtyB4Dbmt3XExZd9oqNQFUQBQqR
QRD9KT+4NXIGGEyGI9BNOMI6QxR0bO9BqI3oZmJBkagWwwcWTAQ2tUh5b/ADRR5mwjQoU7KeoML1
QD0O3QAI93m4fMEk6/KAiYNL6LZR/eZj3RC6L8hnZ9mLWg0UiFPDi1CnIzqBsVbYJ9rOc62rJiDU
IfAW1jBWCgUXGeSVKrH1xnPtRjWtIr1WMd5LuMI9uO9Tl+P9eqPc42fRR5mGcDdpy2qEOn2/7tdc
rcdQ5m1Mn8jCKctyLKieVUzAwj9i1zMv2R/u7a/E7fvzP6axSrP8tZOBim6qRkelR4AtZodCcB92
eRQ19YExuUtb7Nd8eVCJ5eM3oRMz4Pul8/cEszJ/sYnS3jOk+Rv2lTVEDNkw6JnWA1XIOXMY3EjY
+keP/Jx89zSkhk9EnojGcnmuhpBVmLX5lqXhjcsvlX3EHKRPejYaqVGI1zDUP6Vrrf1HbNZbcx9I
gSMSwqDdstRH1j/Cu34Pj7YmX4pbKOVKp8NTTyHo6Sr7M9n82IQOXv5iYc2vRfb+uGVmdGSnlBzo
/bSLP4w+JULhT24Pgf9DHOjS8QY6LhAcRWsh1vvsuFz3mnq8KPMOjbTVB/LuoW21cZoiumsns8cj
qLd5oeelTYMt1asxDjdZ2kMqNwVjOnF24rpRGr9TVsjGJr3GYdWmgTbPVU7S3NBCCUTlKMN78/8C
9bO4Du3oS2TJIrtoRZnY//l38keSNlNpfXX/0yA5t26ASaZm9hP3RDqkrE0LV2t0buDiCL7kOVsB
iBwDEm1aaaZo72D5IO1eFia2y6n/1t26QlBE1Ejfwl67vgvVeFIiWjJ0apkJ78FNiW07gkdDL4Co
hYRwX2J2rHyp3EGJmLbmLQyyYPJr7CgmbWdIew4IHswXebVaoIIXo62F5Yd6ggcq/K7Z6jyUIL6i
IuhLgM3cecTmZgkG4Dmo/WRkh+1foiN5pjvEoQI8ssU30YIE3xXhLJJfu+yDow7gTtKaidDT0uNd
l4Hh++dlBaUkak6/1z2tUIve8u/GqMCyfwiqtXOj93zB0Og83NVDVxGIeZFgKgC71rkTHuuMcK4U
weVYkSo+rk5XT6rQBgpkKoM2mkDfqkzb7z3YaTWB4xu7kK6Ic+a5q6hkMxEMNkyCVTiCHJ+/Jt65
MOmuulz8H/EcwA7PrJ6aMj9EXOzaF0zDvlQtuxFK+IY4hfFyCEpMsgwaBeUUt7yV9MmJ/E+xU06J
JTOZwpQhrFHdyMJrugTnaQHQYQ+8EWZVxc3i1io0u+AY0Zz/Gp/gFrBiIwrYqRbxwca09M2xjPHg
IP+x2U6+CMtn456vkgims+U4O1sH4nSuFxq/nFO6o6sQl5Cpihk+C/80q5TqqR5N04qY0M++NgQ+
FsYA32bqCylXU8kYSM2h8KtQsSxIyWnPYTfsnelEHF3FdP2BirDBwiXe9Tc9BbR8lVlh0vTJzNlH
naTdI9JAwDh/YWZSgGGkLfl7bBWiM2zrVTaYx7SecmtxcVIy/qUT1I8esqOsKON4tRE1d3ZCG0Fl
NiPkWkWHSCvjmgXRrwISbZ3yr2cAqmEaDoj0dDsiEmQb4u2ga+awV8USpU3SE3mfg6LGrtMcD/6K
mCvxrDzJniprNdbJKCNZAAT50nPnxVDdoAsVQ81CwlBK0U9RepdAeJ7b5hm/UGSYjnH2HucshR+G
LysNaDnzc4kub/U8WdgcAVHRwJSKEaQkvv/vMYorCy5jx5dfM5Lwvjn4P5R7+RPXIN1vG/hfqJS+
Po9J0Zak4VOWGtVrWnrrZYUV0hcnLL3NMLxlgPptiNvKwqBhkiv24sxpCdEb9qq3wdEipzILy351
6dkY0JZsgov22E3rmB2eO5OFfkCq7FB7nvLU4aRcUwLKRqZLqiWQb3L9uHSCbHym6nmggUDAt4la
GtUWnzXJ5LtKo6Fs4L17tyypruBo9qoabzl1GNXjH1287NXS78lvov9KM2DpDGurcJ52ydw09YfI
PlDDyRcbI33C0tTYBuKKSITAUayzNfWIOpC+gSSPoiFaBxXr2FPVrybUQVt33CoIwEABxkplC8rI
5Aj+Fw7rnkBlNduTMmsTW6ht5ev19tN69GGOq20clYqPw0fsVRxIMongzlMNBnDliRGO9KoR5qKS
UxPcBv+mzsBO2HTHf6RNeo7/E4wG+j98gvXbdtdasDlNk58+41H3eUwt65GsEGnRlWkNFhoZh1Q7
QlH856UyzBzSJEcXhgn9biR20usQx8xd7D3RBs5q3vMeO/Ih7vDbkRRWh4BmVhBVflRiJRj4x4d7
nge3LPGmv30A0jpnqdljblvj4yYIWO+mbNtY9kBoval30HiGA4q9NxdRfN1rf7E94ulqHlaoTAXR
dLMJxTgwb0X01uNlksvG63n7lkXfAUf6WERQF6eSxHiC+lApm9CvXCm6N5+7MmOIrG3/P3c8pYRC
r05SMm0glDGVcjRFlUcSrjsFIwZLkrKoFIu+cszTNduowbC50x5+QWpvtMhP6B0+wFF53b6OYI+0
ADG9iuwc3G/SbpTwBjieRRz9me8jk+c6w0MVTI7MmDUZ5WMFdJOHb/5zP4bHuz5fIAZBufHm9uUX
A9f4gYu56h30CMjFdWhCHzl4LnGKwiYroGAiJ4s3pV9XPCQjJYNihWItZwqpw6ZDm/+REvl9uN5W
3WEoWA1+NHr1+HXYhJgMLmHfSLH+x9gJ6v/L/1INClC7k2hd2agxrrndFO37Ga1uNFZm4fcvv9kr
18E0UEHNCAU650OLEmxGM1lgkAdhwo+06ReXXRULTku3uroAbpGetiQywy50bEMhnXOPp4qtjTrb
VVNxNLVIcGt3Zt9vXEjoPhJpXShwlesM97rZLgye0D/pGCAvo+ZSE9yhHjcCVhmZBbOWW/DMeAPC
4r+TGtmvgb/b/OmSH9ND6wqmv6SWn8iA2g1v2L5CDyZyrskmsRDRHM2aq2VZOlBHV4hfGH0JMIxe
bD7211k0KEJ/FYMI9GkdOkdkAL+SJlJ3A3JAewu/VEA3I333OCRRngvrJIlM9YJB+MqfC4+GbPLI
OyHF5MhZsyzb66rWsjfL68KazubNjLtIHY2i+rCJxJcMh89dSl9dOJOMDwhYAGgTNsOYCbV7j1/f
ArB6DRTSCLaXyPswlPPyZ+AHDeTM1ZV7BRsACpWC6hmM6X7aSRYS3Rd4nhHFLYgD9F53JJa2OTep
i64IbBYi+Qh2zfQEmAgsycXj1tku4k2o1QCr9aM6MsMVTPUciXecu/sW1U0Pf5MlkMs3nBvKOxrS
a+rE9e3fBFO27dfbQz56p8lcmlOaVpjrYie5QL7O9IKK7TYIPsQQlO67MiL7q5Rhh794Yqo3EFU7
/MyekcB/Uqp9u5iygFxemgUMfV5cM7wmg9HSTGL4NRZ0g5qyajUn/B34RelqefuhNMSLDo8GOTfd
1oZLqqsBE3+1FtSNhBF1AJTBZvr0vzNuxwRrTUFnixLVXTZou/CGHqdSt3IGoBAAWqU18YdIqSqX
AsyZpCSSk2noh7U4MJf22b3z+asulYOUkdF2ovDOwcJph2uqR4aaQP+5E4436AxPqttYU9UBPWOJ
MIflXI4LTKFTQOVjfC8Ecrc8hNqh+eKOzujYvogk8P3jdVskKRjAcCxxi8cFXgohMfMbirEY3wJE
OKovCqBi0Ytz4cUAOFSVEP9In40CO3zh8YJ5m1QqlCW+tTSprivtQpXmhIQS546us2D16dtPU+1H
GyP34sqfj+W9APAOW2Pg3ueZ9AeWdhaeqJqivu6PiTUomwW34eRfk+kE5z+6J958OCUkLISUvvQI
hPFl1nDCaAsQC17y1gDZAtKMV4wdWXpo156Yz54d9IO00J+ANZ6XHcXi6ckovRtcKj5MUZqK770T
d64uNbvzotV9A4aMYD6LhpsgPo8qW4U8B9n+AUkPHq2HFJSfJ7LwJrlqzg9sUW+x17yatt4294Pm
orudegta4LSBf7C5UYlDcv4IZrQ9Th3Zgus8dtHKGWeOP9xWX1zaje2KQAPey9qgjaeHYtDDUARi
SFj6NV//D6NHRVXOYGq0/9qoMw/As6qnPmj8ArEpqsVvNiO0tid0XsnQcez9FonPg7oWXXdGVb6i
ycjXgnPO9X1yMy3N9c9P8+CNpVigh8fzStnKO5jSc+j937aAdEGzPVHoiDftudAjcMcJbQ74x715
ZtRrjCoH84b8zYVgLIkgnIZ0asTHM9YrVIq7Drvb5ISjh0ScT54uNgg+Pu7pNJm6X5jq8pFzMmvp
JFWsifs/gh30g3bdMs30wrijVjT5XnZzZqKghbE27lPNG/wyqylXXHHYCRvUOE7Hs4B9bYLDLcL1
29spuxMQjdkx54c3uSq253RxWYRG1X+Lp2ndufxqwLC4WDjVuH0wXfw3joAo0ZCkZYKoFyEfzhuu
pwuTSlGE0up1n4y5QUEnB1k0gkgFC47EStMC0P5F5DO+h5Ht4rFQvF94JwIdifr+3+hDKmRjjGlF
g0bRDAoqyhVYyEk0KbPAL8QYbxU8a21UQK8AjEj3aOjk/3yqAkA0wRg/3hWrvU5pi+2kRa2Isms5
EgJTFNHeSSJJafnAFlDJGXhLHKJMAQlDuesicvtHfzC14C6lEzPRATGOI1GzI74H8Yumj2JzLRP6
zgBj8S79XYZR5/skFX3ucJweX3Feaxdsh52lxJRtzP9mSXHSEyiwtddA9AE/FeQkqYtL7TCo1VIC
FPoNkY2JJiEHaCeAIEV1Nq0LMiWT4Cd6qClKRvBD+4Jfhcs8rzmdKVUZqqJKc/N30L9LPVbT2ZnQ
fuFf7J/7U1f0ncuqhMO1uycvz2zEeV3RvRo3nL/AfuDQuex91vQUBmZt+HCHn4PrU1Bn9xtaMUOW
/CMRNeKnL1geVx541d9NjWNvg5DXYhDImIcJJ1lk3Gms6FrcdfPPBYy0PFldIhqALBkoGCta8DZ7
9YNTXwKVP4uaGpn8MqUiYFz0+BzAKNv4gYbSxsau0PvoEmhXVSUyHv6tCoyqR3Mo21L0YOXdlu7W
WMSbSL2sZmzb7J5makTtwMN+D1hrkYjfKQ7LK4hWPwdZnSaJOfj2FGSU8GBk17S/2k2oJLTvnqxW
ag38RdfTmpUeBkMK2p6UHRwRfH4UEIh1Sar4wwLc3yN2M0jf4oGKwczAHsTrRmyp2R+MWbd817Px
u3EIt0gxNIdT4yWn6XenqjZkb3ytKkcXEPJmoKA84b8/KrPA0FrI3CeZszWbySOX0NgR0r+5TKEN
LYtr7Ba9IjvWKS0BZ+19sDgLxiURlaTHv+P7DSP1mKEbQ2/un1K4sRswgDSh3L24lgwI2FR0KHpM
nQXrISiubS0mk5XXwK9iae4/nsn50Ccc1TySrU04wcAdYXv8hvk7W4VBgkyXpmOotxfw60qmQ85q
oVxvoiecoZR7yZustR1LAcPThEz08HGMF9LGBGRJWBqKUBHjiTOQeLbey/ApC8xlDnFsdOly7CET
O1XW98MRDxR1TSPVZ5sqx+7TXbYE7IxBX6+2t1ukjcrOk6MaLv9ZfSP7CQ9IpTRD71cMppTHXn6i
haBsxCUuTEotIBuR0ODxpj/f28UsC6KjxzAd2nOn3EKTwY1c8OXvnoTWuMHfmta8YWiGMgwH8JZV
w2embUS/4q6gGJzJ4p5pXneTnoguJ68FtQIg5hXM2qKa/+k9EHV5OjwBldcWWr+FuS2YLW0YaE+j
Sz9s1ofUcTlwRgcqF4BjZwJIeq9bkDB3ekjsRajs8WmDfI3gGn/gGhWLf2d4hhjetMpzFz3UlR19
kMfd0evCmDtstp9anQOHvhU76q/lN/4MZ5kN0LMKiWH8YowDuoAXEzyOgvphfB9GSvgH8oaWDqbA
DgwNtQ+cqjSRChcnttu15m/BCX/RWN5+i8LrV4McDiRAugAH9UNXIFRKni1MBqWvj/jIAZrehK2x
brOxweK/y2KsMPFTeXG7tF0/+bX3PcQLpDjAQCX1duUPiF0HHFy2Srk36LPEyzGbVebPCHUg/0gf
qaUJ8JgtTZyGX4hWkHyAgOjFE6FDYqYo07qeM4kIyuGRb52ut1d+sAc9ZH4TTCxJ6zXMBYJjSB0f
ZDC82cS4qmLZeOKbXWDwSRFbMYQNN0UsKE/WtbiEqoCoS6V7CTv4ctNN+MLK9xr5X/T6Esinnz/X
n0Q1QO+HHnL0L+7tenwGgQ9cAqLWEgJhhsEwnLIjCe1z1toYFBrRXr+s5AbIEdlXKlyev8NMvPIH
DkgNt6trqAtOwzaKIbV3iiB4JF34OSBqJ5Aq9yIzy2nHBEOgyNNrc2qnA0MG/QxuGWRrC3sXvBTb
SMIw9L42XuyOpQbiNESaCiQFA4tdDOUrbV64lSc5MQO6SYGAZTEzQjEJV+AFqvqhUEuNI+9HrPac
piWBxD+RQ7srdFJWvBodni9IMa8JBItLEOjTdGl04DHzL54d/8WY6aIcyV6XtbkwHWrgIuIduhcW
az1DFdQOfTfdG5Lo+DUQ4PZX25uPgV9IgJsMPodwDj+4dh0KLC74pUPUPaf/roPvAx3Ut3K1bVNh
EK/7XpZFDAnc5fY1r1BKvByp5lFi6/M/LW0G2FPiPcOQzV5vKzEPcDllqzsS5FwZF3UFGMZ11xua
cYfxs8AyIb24JfZS84I7kUM0FnMhiGq09Bi3dAMF6GhzFwMLEsujHJdO8YUF0Hu/30oVCOsobYxx
drzlVM8aD4TcHJY5MMm1cHI+1Z91DI1iJJR7jrcJDxSlhnRKdQt/TzUI3rjAtOdFLor8Y7hxXles
+86XgDzgP8Dr2BOH5x83+nmo0ctL/5ufWEniAvgfGP6NL5ke7gBEzzQkhquQVNkQUgc5xfYIEwIc
v3gUbCT0G0+s+z16isTOF7nFGXR7RijAEDJ92LvtpdWHLFcc/qzJCNGjo3+9bsVJ9ynAnjoo7vEX
kgRE1KfmjSVaXstxo7xhbzeSoox09vPvrfp8hCP6M5rlXhvqJDtZX7XdQVOwWb2dlGMfrOzryakP
I3noOtNai/fjZGM9rRcI3+3tBvQIu+igrMoSTbY6hpny/PiI7piS/oPTB4u1y0hM0Mb6BWhJtvBR
jy/ZA1TUStUxlOnm9d9xzByqgsaPx7HFh2X5S0Gqb/TPMh5SMA/g1r0mhATKfPwzVwEmyEbvKaLa
aYt5u7qTCGVKo1kipfCMx0EwiHqSlCgEj9uHE1/n7G5MQy6MQDcTlpdvOp+ULohdAL/pbnSc/tpF
SoIpbdh/SdLIkKhjCKnDJM7wgSeghR847Wy4Na/XaagXO1zWrvjooTjaXmM5axB/+ALoOwe+m9VQ
EEgyR+qpl3qoqwREzmt3YNyV6t8n4MRl6CTFB1IUGuBTVaaJMBdakPAK5hwCzcYGZ4ZR9911OK2Q
w+6zdWRvgM4CYw2OAU3jH0m6fFY71dWSe2OF0liGinOund0Pi0dpZb3aLBV3N5wqH62Pm/JfK2uN
GLx+hRoSoLXqmzOSjtvc1c9/F9Q1gaA34cyndK9L6N4XTbyu3z/zKVSfHoqBQn4iVObAtLl3h8Nq
2nOLZia4jhg6fWMvLY6U5IYORnpYayLO8Hyj8qxbXV4C+2/BABkjBrWBhB+5iby82P3G08rCtH58
rlqX3NdVc0o/XvpoD9rqluauMmSDcrJ9kd/VBJ6MMQpNM0nRk/om0Tzk6Xw73sJ7s0n2sTntCOCB
GWdvPlogyIXnbS1kKDpp68Ccpvc1dQftQ81rGqWf2vam+HQO3ME1bSEepVHLPyEwZ1RvBB6+2+5I
A+2cJZRGBSI7zqFgqXWieMCkXBqho95uiM51iZ3yeXTOml7GH73vaFg0SvBNNVAxPBfbacuLh4NH
LQn0rzKS+GqEwRNIV251RYjv4n3oKazek3pgi/N8trNIwfmsXuVqDbJdztddckBujTc6fMcOkzFv
ARU4/9VwVdqEG+kCzqIA7dyKZSkeYflhlaZCbMqjiY9nthaOwc+YSkCV9foaNUOBFTr8mbAFmHLu
xTNZjRnlg8ZQ/+WQzccR1W/xkFNLjLXeiKK7oalowytm7ynPuwEQQcqqdh5+Yz4IVt8P5gSC9oRV
oVyrp9+T+yh8mR98w4WGa4gMpskRBqomRuaNDnRGNGtTm/lLwk9BsY6uhf1oQ77MlKDRy5fAyc3F
f5vKrErEu/iu3NYbPjkdsO0OfiFbAhGF5y7FIIeFwJQlHNKxRFAN67/82n1UjSEj4G/DHav0RxyN
xiGZXkCKz0evQ/UVCuVF8EdHF4FRoOWaXUqIsfpvELuJubvdzIh7dT4CzfP7/rlNDKx+D3NhOrMe
K4uHtPvNi8hk4xn6/8bE3uD3msGaayZeOGWpZXQhwCg/mAOlQSuvarjgm1toPvp9g9w9lRaGIf77
jm2Rq46DMwEEe683yV22vMSqSKS0WEamza4xSrPit4MyaU+xxTTgEJtQhT8k7bjuE7GgfN35Oj+T
sg2lv9urfYZw4n2cewp0xzKtBCEzM9qOYBluPsz48xlscVCvsvIFUKTjHFJR3p6d1BBVopQ8Bbir
SfmHEvH6kx+P2xxyXdQEdowcPv/Egb/EpI9yFHGELbGzRNZsS6fsIrqYMmF0KpV7H8E/pst/8FXT
IkX0g0jKqg1TF10GaC2dZdRG76uLzc8a+GVPKPdxioK+qwb8OHTKn64nXjClvH4VQtMVYw1Ar5wn
60FUTYRFOJ3cGqPI20jJy6az+EodCUtCZswc8RwBPm0c2r+1FgIlpNmoHXgd/As96b6jmYPN2yk0
Dq7bz/AZ79zmjgWe797CPWynShClPm7uBGHbqYoK8z4ZZnguGVJsRCoDjcjVmoCZuczg6/u+GGm2
br3d6YHX1/4G2Lurj3SwFV6SCSnj87awts0wc0zUC1m0cFNJNhyzpZ3SuDj1/9ovzDZNDjuV93pe
0ty2Bzk7x8KTqGhHcy/kdgAfiYNnhGnfX2aNL7gXPSZ7s5ZTY22o0ASIMrJL5xvsn2tf3fT0uBxu
yqZ18EccYp1bEG0RKmaP41KkX5ot+j4gaRtPW1lblvErv5m/Wd/TvdDoNKiyg8JkCZjsaVFuhjuS
e/Gtnv5KhBWhnS13azVUv6qmYy1drgfTv72LB+hHX+eGX5fRryipjnNb5eg3PDQWEr/Sq/RV54Mt
KFDfsq3yvhYOdsq5A2BkIXx1XED2qxXSFu0O/orzQ5FtqAlzo8pze+8dh5kxaUCtZ0mgOSpNiOE9
2n6N44vzSZ/8uAQsDSKBrjTQzo5LL1/ncpOSm4gtiTlZE7THxfpD3JD37cbeUF70uCM+tLFb2EQi
mkYySYQZieM/pWxpNBw9LCQsVCzUosA6Jyo02PCRExXyZ8X4FtvhK43LekJqUSkY3L6EOsVgweim
PchjQCjk5IIUZ9MHg4swSa/nswgdYJ6U7zM7sJisnVo9L04be++nVQzcPj+ufxQiflEsQIb6Eh+H
czvJaEL4GDpox9lUg+eNBY18CrctLit9N7YQdeSRC/MWxT8jXY1rcjZqcQg97ADL4qPOKShxkUxG
tb3MKtnDkeGiTEzMZ76D1srG8+xHeqJbrvBBP9PC+O7hjXhz/3BIksgv1VqcuB0kAUfelVhWI4uy
7ouvyGcHPj9w1bJJ3fOCfi2e02jBJjU0K0RghT/RV7RAin2K0o0arPn9eC1tANqpSf1uY/Qv81nJ
wpxzA51RICVcl0lRseUDweJ49CJcmCSOaxuyJl0zNMjx0fklXg4+2ikilEOLot3lhS8hJ2QFxZQG
pJOkPK2JHqAN1GONjRV+BS8DRzFmB+1GRUSw+5HrDWahri016MuzfNMG1QPKe1kSI8jByzkUwXH8
jyu1ZHcpZOzm2PBxBpY+hMQLeNhaN5XHIE98WDaFDjYsYNV0WuLMtShnbPI/CYfDOU/3ObmTm6Ts
i9ZLaDp7SCadKEz2qJSEUFIqdY5bVin+tMzVrYirowONzuWQ2DZ7Dl4rD9Ip/1MzYdrWheIN6VeM
teXphFimadySW+RCgiLuieaC+EES9dEXhO3tuxe5zQQsg5/pDoBqmkLvgN84FRRgQKRpdw1+qiOw
Nu0cUUmWC8bsXhlmTveoRywUooOAC9EIPZnvTW3D6/hu6HUpo3EFouKZr0zTvrCDfe8Sd03uf74H
wIuU/qIIIUV23UQ9N3XVRm0SR1SpoqKiddwY5wBk6Vp4KPamySEMUEiPFsZyFyUUbiHNMIM6MpCU
ALS2YGb/pELEvdm70jIbEdlxtHwzH/ZuMCoicN4ESboXZwPHN1PnMsFT08lD4uhFhJHnTNEjdwdX
8V8+rN12B49CvQwlO5Qjrm4RTvRbRTmineHfWpT9MbLVeLbxUjpamjtKP65hTjimrfFx140dgN0u
H8cgxmMh0hrf+Rz1SPSjmh+KEuXjrcgBTU51mvZPMK9CJHlfYrlLD3dhU6UPxx6hxF5vJOfrfMUG
I+BseFoqHaO93XDPRV2Ss+ZmXI0/x1IpMvvNBDMLN0oAl16G2hmQ63ROTcKWAtI0UtG3OFN/KqVt
D0Fbl2LWvfSXuozgX/W1BdzgUOhKfVOIEw/iTu3CnHNQckHgYLT1nqHw/zHF/DR4x4/OVXNLCMOT
LPtrhtq4eXFIVRXOLu/9uRJonzimQnqcBmxzzlDqG6MyR890Q0b01yRBCwgZ4JbSe9ZE+vk643Le
9k9Cjyeyofhu6eJ3qNF9HwtNd2i5qrstL1zOOP2EVg1elAQryRou6NvaB3/fAG/idQA1BRkmCVMD
m3bbnDkMlhF07CUysb3gzrR4765bFy/fcBU/Ezt/u8aMRiwIamin6mqHYa4hJ6XB4gPMd/StqsBi
iuGS5dsOSEZXxKjmZI0mSFoVWD6gy6i4bnhm9ghKZ4G9QsOFtGcjXCWExEJXGrBgajig9ctxKFbq
AJv6COw7mbp4HN17yB1yk9SimeY6+zm2o5ko+FLxRw90S1TCNrj9M4pqEiKwCBeVYab9vog4n3TB
UPnJRfje0CGYXwyrkLLBHfEtvVhqdWEWlwVEB5nBWJDEmE5ckrBeTD0q4ma/TIzdn7NGNIJvmdnj
0TNv8/Sm6a0cbK2gZjTPKZIVWgdqAnoTBFuoWDHBDuTezHocQznmW8MzPlbp/oNOK1e5bkYnSRTF
HZA935UIrE0CVzZZ7x7vPBnHeXWJ6ADIVIzZqvSeOrjN4kOOXOiut3UZeUlfkyKGgcsQBprAdXmc
UhFo+v2eNHvyzcxaT6vCU63fD194cQkSMx2jvwpslvVpqSJya48/HWK7fA46TZpoULC6gC/KD9dk
0uwVPKwidC2yYIfHp4CZ6ORuzyfeknOWvuSmsZyhWFUuaPO0R7MKtLyH9wnoK9DZ3mhyGuQUVhqg
GWrm2dNnlYPgvWXtbdK75QKQlqqNHnWn7dxHXKzHzWQAYfV/vVf7gcXvOgmr25xIxGmNl2Pq0PGt
8DS+r/5z4Afy7HCKpwTDOa3Yn06k/2IAFiWDshTQlIqQFeKn7gpnVdTN8/S/NjxH6uVsLOMcLUkf
wxQAO3SS6UpqY5HslrXrNwWTw++mTX3SuQHE0rl9leE/LpZ/5dvkbb1wLeCdNkd5njmIoy5cGC1I
8Q5Ahjr79eOFpnhZx0GnLJK1nD7KariK1GNONlCb4XR0oxcYfMX0DLK89Rs+5n5fER87PHZH8uz1
KuauzdQeXHpRGJphhe5e0RjxIpgapoXHv9CmzBhFEDpJH5wPkF7KtfCkpemBsb4TIKHnfKJO2xqz
7HBaxScgCoFmBXyzlAY/PBqxk05MMTP1aDosBHSbkHkc3covSg3gjib1sBgDXUYq6u8u2wgSMfDA
GuipDEjd1HXCNEux/qDAGcY020YriEBe/7NZgiNrYe/dh97I4Fmd4bq6+raS/wOQHwbsTzBIO7OA
1JSUup/VZQHZOqr5JqPaCew6IkOhmKSE4Hw9jfQPH8I9W/rgjMrI8v2VG5NxjkXvT3PrFP730DfW
tbN2coLOuq8PzSbfZpe38MVlBfFOq8gdkMci7alCluQOe1VGTmvi0GQeUe5tATwTFoit2NfcuF6k
zJlSlvnchLcBFQpPuypR32ORPg0LAG6BY8hbDafDKTMjCZbgt+0PuaH7BX/glTdbKLCEgXkZH4gE
NLvDglYzXwlJCfYphxJprA9t+E8BTSvsUHD8fR+EhOlCgPiagaoF674n9GX2yrJnGZdyu7LealD6
0hqTk1QumC/mqH7KwNWUYAPVrv7niuKQwW8clPw00SKHXgwBPB2v4xMarJniq5nrLe2vLUEssAhK
DkriicL3KHhXcJJEKi4McjBzCfGQsQ5Xivd5mHRthXSZWpruaa0pVB0+hxZFCRplCHmHubxwDPQQ
3pv9ExNEP5QmzeJ6hOvjY1luxcRSdCnr/Kxe4D2JwnCYXhDfUVJu9AymlFWMGFw/29YgNQhcwvl1
rhPUGfLefM8Q1B/ijgMYlMjyo+9EvOiuqON1f12tSwAp2zecjAbsTfz2ljg42pHPO3cbN8h0Scjd
akjyybPFwMm1jEW7L22AswrEFwhQFwj5iENnyb69b/1pbHOObzgC6Ockg57bvV0ymTumASFzQzXa
UMNE2IgCW2iS9dpRgY1oeP0vG4ch/ocBOXcz7Y0ERIjwzPYzC2EAH4TzVFbvzp0jAi4r6ZXgyGEq
gXifAIcNKNW98jtIxl8wrN5nD8mw72xJLcZVswIsfn9qlvkCWM2rlGhvVPcGdehU2obxm/sZJWWS
amqAHNmJ966OiLFFZFpYyGHOiGGNz5cVJYLlFAb2NHxHpH6/QDJIYJvb2pvngoH2S6nKVOfkAiXy
wvC5cfcfc368mRopFMehD25GH8taxjYU16UszUg5a8FgEuiz5aFld+lHAYosaOECN/ynbpPNA1SG
2xlgMoBfuGq3GbrpdKV/wvcgnpvfqQyQnUNxB/aSrowntpn9llVD7A4LcvmyUJ025H7EksCmpylS
70/fU+Ah5ItEzcDXo6HguFIfKcY4p3gwJdW3/gQRxxWy1PDhlSAlVORx5eYXltI3R1boC5ucfFTL
IJmNgrgWzAJWkgMHHlRdbcPrmxXkT/HxBWKcuYu40ALMIf7hGVSl22uuay/XGXVm5DB3COqBSEip
sLSxsGeDoF6T9SOHFdV9986BqdjSfayPyLO5jruWLeRbtcr+dM3WGAVG0vY8K0SAyRkWHdnwvR5I
jrzENZ8dCtmQtJboYvpobxcuvHpd5LYjbOlBgUnyS62wmfxhg2u8qIQM+YXAoGhlzpmBlyAU8U9z
xfQv+FV/DYtjYtfb5+64spl5j7Et8q7+Obb7LIiRWEpj76ocytg1e/aUSqfGFhIUYMzQukfDB068
bU/mHnU05DYyYZeJvr/sNgn8ioZcZ0/CfHY2wA5vfQ/u76mmbtC+1TFtZplIxSQ6xF0VIzMHC/Ud
CGmJPUW69gbxuqhdaDIQi+13u12Tnzkp1IUEeCoRC5JABkE/XEcdwivCbL3xSUWRRscqxh4XBWaX
kvnUTBp8iLilowltp9fIzhgNeLixPRppQ/CRD4CI6vu5zdbMeOMpMBhRFM6zf8CtSwUmO7rOIVMt
ciZS8YNOl16HGgb3Fu4Uz1w/gmQ3JWwFeJ1NwRNjfSjnISsV+O/Us8QOeKV0xWLb2KzOTBuKSTRx
Q88KYnYwHXzeIiy9ASAbyTLIMqUyMZZtYWDSp0dYjEgNYMQXNHjRTw4QGBwND2g+t1qpENvKriy/
1MVSQo05xlwMO+IeGGLgt2YMi+GLoOGekoZll+rYXePXUV70uCCVxHIm2XY3ZxSuJiOKOcDOAWRo
JzPt1jOfSr/SIn6F96pVCHMrOxamxAe/9l50ar6h+hHmAoZe2thAyGRNFlG9+CmMKh6rg0O3bBS2
iH8rUVGKs1IOF+VJl7Q3NVPHJyOoCK/S7ifC4qBspbwUXL5jiCBgIC93mLyFCJfyuJeG18IH1qsp
Zt1zhfp2Kcr5h/neceVLpo2MOXUG3Cr0YcWlO/C8zmpixmQ8+V+NJWAlm4PszT2ZyLciQL3LSN2Z
dp8087ZzUjLzBw3ueSzZIrnINxb92rzS6mc2PSDTtNRPgofxdeStbCO7Y5I10AWyKnPKr9ymjdqf
dk/llVqYQsbU9RM5At/tN0DaJS69c88T2K82BVEwKyt5Faw2o0+oEYfxRWWB4kXWwYWmsk7/yLod
txvodItzCEAvZ2gmI6CinDfZh156SdNi/LYoryVPET5i7aARpDi84MNj1KMw/EmRlPvkUMd1qr9Z
GI8ME1MGrMKYWkEcVNkiZFqyjYoAzcr6HztriZ6zi5k35qY4Jy9YCVQPXOuG/SjlgixwPOb+2F9S
NGYzCqgeDApiDrS/qD3ZHMYtCBM2z3/1v3f//I9BlRoHx5+ziJom1/4xrDpTkYMaADmCAAUkm9Rg
T+JfmA4Y4jKkkIWwAlWIosBWlrqPhllBATdHDR65HuG0yWnbg1C5bsV273dqtCEJKQZ5mQ/vLMiv
RTqSJq5fK6B7y1XxEOFjiLdjSiEbyzRig2TcdeBcMXK260S7IDDBLY3tydX3Jfs9n94vUpgzI9Za
ly3tdEKw3Pc1xLrVOnD2YKd40C0Wk5e/Pt2Y19+BcMRA9tpE4h49hB6AofjpSSj+gyZCvTemfXFu
ukDCYJSQ9+Rq67N+QW6Q9BWsH7l/iMAy0Iebl1RhnZQTtQSWNv/x2z5nI0J55L5fm2OWFSTCCewi
0+aIRGTwvMlg3bfZWNPW+IWgj2cnvLGO7demQ3lFn6+mxgbyvfnBoktEmogNlK+2U42a9NVJweJa
N9L0DjEeeeUXLsN2V8Js0Lt9dro2vM/yLRNqEqJY69WTbBcDTIElnVYGPanZRHaBeVu0+c1olJuW
U5J58REjok53S8bdjN7kUQVB7KU8wZxFGE40R0a/mdXoFf75bNgOnSo80v31Um4Xgl54ViIccAq4
CVb7oxcw/3Hea1FLj/dij+gGPkG8R2K9C76fFJZ6AC01sXzlTeXVYdDUad86CSKOibPkhDfmdvpJ
S+uWq3qvd/AJ08M2exm1zXUpMhibk1wp5GZsw2T7j8w9/wE6/eR+Ghi6PtMK43KbxoSDlWPiGL3c
kYIYeRTwubWniLbHvjLW/feav580YFBOMV+TbqGJ3OSgFxRZIQ85Jol4ZDjzN95j8bTJWbm1EG8+
NnRMslw1JrO/dreb4GyDtMPEUqAvdHuPoOvhLK38G7TjUafdF/fqtYLylyGwyaoFH08xzD4gQsdY
xgSGo1R4UCgJKjIn3SC3AhXXipfiPsXpQ6oyM4ZYKgwQZIn2p9dfcrkHC6aP/sZ19WAlwM5tj+/S
IqyTR1mxuS2TKO6umdbaqFh6ASPVgcW/QAVLGVEdFIprl0zVhiysMfBB7zJbHDEFSNqiQU0Pz3/n
rtSa5ha9JBSf4+lbVPOSBXR6FK4lwD325PWqyi3ZnErk18kOPvprzwi5DgJPG8bxZjP3Omzhcx11
Q0hbkf6QDhQOpDoe+O4Dl6Ucw21ZeWAT6T0iW9I6tkdtO0hLstqO/0EXkiVCKW4ZGHmv4bXG2Yhq
89K3qfi6S0Tv7GTLYX9jjMa+0AKf585CZdjuYG68uGsBe3deox3sCKbFBl1KOomrNhNUw13MxlPZ
f7UHGZt1Y1zobU+ckISwKZxDP/yzIEt64H51m6k9Z//t0Xe6Nxlo9Imjgy5WCKFn14NdBqac6DEh
JeO26xsCzFj8J4HLoZtet4Ta5EyDO4P1BVlhqk+PYrsHHLn0FTRr7XH69MG38TyVzaHP5He7dCma
OD2xTn+Is7DGayt9IboKBvQTbr641ifTKWZFnONwmaAuuJ4NhWXgXwoeqjnGcLC6h6PGtLk7BllZ
1kE0cpOkGBE92p/J+si3VTzCForbC/sPb5UjGoEnqmQvRARGWjZuw11dTEarrsTVhBgF2SKJrjfO
3Ek0yysHRdV0+rQIKkfgforU9SWP3UnO2Zphs5ToqpBpAuCIKmnLkAip08HBVQpzzvro6/lRMRaZ
rXBxP14NbJaDp0JS/ownLA1T8tZ1cc2mTnUVtbGjvU6u3lStK9SwDXc44CaY0PQ2f2b60kASt1AC
euMcz64Pejlo+szK7NcPg/gcAKdqAqnqruByBj0vU/bdBRB3woS9lahowQwHnKEEgmz9pKKD/0ca
XSIXMFJbARCyvuEyedbKOSOWEIL1dbVqZYnsRN59c7E9921VFmFC/VfwFp/VA9Kqj1lyDGzdLXhn
v+RV0WlPc3rPN0kERt0CJxfG0NI19ebcbY2KVVysfxOjnOy2kMQVFUaP2JEQBlhb6nhp348YwRNW
dDPxPUIOKPxI2TaqnZdsBQQpWKro5T4hJXb4x8Osphzi44BbgtVnw+ZAHHixi7JxAFtAsnqzOjy1
SHtx9VZ0AuSpFE/UUr6FuLuz//gyaKtD2p2wWCE5GH2gl+0uu7CISbJ70h5mOkpbZFYlxhwh2hN/
/ucxci503x0Qbau7SpK/HgybNO+dVCH7HQsW16MyIIDJ4BkxIH+hNcMqjTCxYRootQR9NofAzUrm
zS68HLOpt/B/vARXvdyEMLFpweYUFABGRC/vYKpcxnYUjfxES2C/NOmEsPqvjZ1kygKQ61tbH9pP
n439SuNIkJ3S2t9aNAXkG2LAptefq27heNYD6ezm9qqaSjG4jvdSCQTG6c2gIBOaweTJ9+CBVEce
19of26AwqMh7HBoKPA+DStS1Zo3Ku2/g4u/alRe1yFUEi6Q6vvJLBbl8/Gbe/0DXXimBOA2B5FaJ
g3kAeQBKyq/lPHbZE+D8w+sV1livoP5GTspq1649xDdQ7QxbrXpQLNM1HRldX4wgo1X2vJdLpv2+
317qA1vhVZF58aRT+pNwXB+fD/LkYW0uqbLlsN5m1yfDzQnuGEP6AnJzkWvxCFJTx7EJMNCf/R/0
m+ej/iM3ay0slBk70kPVkaa3msf8buhJylgROfDs/Gt3v9HhPmK+cpUUn+HFsvKJYCTFLf75zMG2
cJBB3DdSN3LHLr4p2YzhiylSsxrAf2zPuyfqu/NYe0lXa7a8BWN5PUle/YCPP4Xzmull2woGseN9
sImy9N6o+JUFFjS6tJGfYwnL6ugy7JHPBBdHh5c4QHEjm2D7Kce61aJ4uuBpiVFp1qfBcDB+LMX/
FgL703MWt+YxUxC1mEJlMmW1sK0nlk1RjTab7GW8WMIpgqK6fRL8x+4AMOPLWtDrCwXPowg6ajkl
4xli191TAPv8P2VSmwBPtGpTZT0OuT5Ngi0N0cPm0z31FDU6EATfUA4dDbbiF/fMFMrm3wDIEUYX
n2fdWrFIgcvjEIfLkPGJGTvOSZs8rwfld6n43ObRg9Az+JEtLUw6TR45U8vi6RGl79K88xxzhryX
MG51gTi9XaTRHu675OfKJDTlJoVI+E0smNMZn3PjkkglxE5Wquq447HSHRspzSGMqOv5SkVSlnhE
7PAozGKbCrWFEPvZWgg7CP0OxsgdTC21QnIUe4Uy+ISpqIoLB5L9kR0OW788nOU3ZJu+w61Ytzu6
291ppU2/nGAvOX2B02PntfUXPDvZ85+QELZeUALh8IrdRPh3QIDOzoKG6VGHS3qtkGQV0Z2L63Ra
z3kXRlN1as5tlGlr4C0atEQRKB8S2wiiU1cWPdyEyaxituoHBuZdAKgQ/iueqM1EOkOVJL54s2xi
o9UkrTeOni76Dzxk8o/T3Fzxz5yyYafdTbkPqq4jaHatODctNyPqN628fOEnl050ybqBxdh5a5bc
HLmpm/QNaTqbj5XFwtXfUCr7nBpy12hJaLEnh9qSoOtY3YT4WWIzhC0i5W6X5o04m8slkPTmLr6g
RHI0ivN3V7aI5Sa65/AuCMXarQ7V7D+EzCD3z1jTCCOGEIr12JvhLRGFftMjZvCXpTOFIKnI32nx
mZSvwx99POymjUo9JxZ62o9dV/QDc+9210QbGmUt3rULvr/ZU5DVvlXvoZbGmkIwGikcpEMtr4Tz
TyXeodI/n8eX9G3Jdvu1n+YEep2hoxnEvE7bxT49+tAV4jXDZyLs4pTQWl+S82AMts01Z1+4sSiR
ADBWRpFojIu7V+jgVspztXfV8CCAYmQgl/EnR9zYtPUMWL9HmAoaxmwApl2ecO6uCGolNkaYqh8J
nrNC2522qNn4zOpB2e/ojSX2EcRgcpCgQT9QGFrk4bZ3fHDLI/J4ft16lZMkuhCn5wlNinnxicwB
v8aebtGB2A1GF1/iEZBLKpJHGCSgbX/6oNRvdTYh24WhwovYOFmwUhJHBGfzIwbwn3AimtZOJAPd
sTrWDT+evIbqjMiZKE3H1DHKmz5xLmgRz3pLcx1wD2Fo5d+gdOh1++fCnZ5p/67YGMK8TOVt3mVn
7QrItS2eig9vNYQTKBfqT/WfQ+63/OT3HHRlBPilsO6KYqditTF66Z4folBEjXPuZReiqPtAsy5i
4mZpd2Sany7ne6oZwrP4/TCS/zszDfPyJWfc8qzMfy2gB1ljuh1i9eZt3goGK9m6Wndm5ZMnYIED
rru8f+tMhjzWWU94RjYkLxPbJGd5+GK6GuiWfS8AMwgtbtYJxw9U5Ur0+KhyAwZ4bfKDyPIOZuYP
YjQl71/cDHPftO3W8jbuaxWq+82wq+LLw0gXKhbkYU1auMQVTNBLMoaLVf0ShwYoxoN0aVlyy62h
K8XWzbKpYz+nLIo+KZhK4Y4OHyJgONgKMzWHetser+fADB00dFMuscfTr/7HF5DtMxOpMXGEI1aU
T0eNURzT9JCiSjY0MAE6s/SV3TgESKHKVPWBSM4RUsmozbXbXlu739Pzw58ESWA2JC7cJ5+ZIE5b
72BrhvFq5bdP1BW+IKSUVLt6u7VJMOFxXWlakPAMn6O/WXBKrItF3ZIvH15j0Ntpo8z/VOjTESir
17H4SC78xl5CGGHr6JUjxKq5s4zgqsUXzQrSZMjxCljusU+sCNbOTOPbwKxM5XbGVd7TmuS/qCmo
qfYCg8RsqJR/5YprO7IUW6nt70Rz41RkqkTux62TPeq7OCNI9rBJ1A2ek+xKCvtFFO68oJ+b13GR
k+A2ssLK4OdChHmLq/mst8IlIhfWAbBAexD+eQXUXpnnMxUjooeegfHvtdHoS8P4DWV5cgzm82LW
81IGQfJtwxUHLi7I1DMMBRyeZdCHu/zGp01ukIMiXMDRiHCAayi+74k1R89/LFwlbSSrq+Qf71uh
18DWyFeQWEsO//vJtyA4ALgN+K7ttkp8ZX7fNoTNTx5bkItH47C97xhdR2e+NmPMryU8IIBk7hex
xz6j0t5RvaXxN563b6MZpv6k9fWJHRVynq3Sh+HciH7jSMF8F7Wb+b9yf4jgOmpGSSvo7/5CAvG/
wpnLvJd/VPZ7VaXoaTxAzXxcSoDa5t71dR27DmqGI0R/Lj59Fs1AUxMzc13fXw9mdSsom1+fE2Ft
0uIIv8okeuTQZgNDA4bBoLXkURR83xXOaxUEeIgnFla3JR4w/eKY8hXqOY/caKmFrL/B08DGDzaq
oGlmp6BaqxhQlHswBoCacBJE4/fuzmNv0eQfeLqXfBp2nv7T9nHPSvj3HsFEPeQkwpVlV2+Z6GNq
2sQ6ojaadjhMXV1bAH8TkTPp+EnFBM5RQvcjUqHOZ0Rcffki5wdhA31NXwBnDW53K6aPm4OkRy4l
f66v3iSvnzRPKAIrN69Ig65eqct8oCLTJDGqKPWzpof5BA7SfIfEpzf6AJkpkdIYhV9laMwl7M+U
p7zcSRq/KoiuwRLfOzS1HIM9yCe+q7+pAUMUnbCWV+yjOWljdK2n0TpELcOXd8trM6bkWmdyVtPG
GAY8kvev1XEPXlpmSAQXiDsj7gCGlWaAm8EYwggA7PwpYGrgGSZhcVmzISta5irt8zas0EzinwNg
MGIPB6/fs1m7QOTGNYJ/avQXKtTIn0qB7fZ9JYZcgA5sZdoSrxMursSFoiV/BY4OB7Kdie7Fu2pv
it6xffcd2q95gp0M9cyTmeCQwyuti4TA4bxLG4Da72DSyUbtcQLpUbUxc7paTlb1qvE3wYGz/bzN
iqpZ/PrZAS8/V7k9lNoAb1hYmxy3+q9J2NxULSrz6ixYVLIkTo9GgJ9Ad8BfPRFWOQ0XKeIV/zFc
1l3PoaHW014+NxHmcuXMQRSfg3QcQYSDfjaBzpgdXw3DWM+aJ/9qGwDXEm/yM3VLOS/bYJyrpLFT
f1vNO4iF9XVDtO9nNowQGDHbHyELSraKCDZWe138jnLduztZhd9JUF0B8ob7233R0HcpFv/4kMuo
qgKE8oqXlk09U7YPO2TA4AnP1/5ERQFBN2Pp2LFNmDioA32Iu9UcMg42pCwQwZP+PfaczqrXi8es
nas9RUiGcOxDJHgHtPyCeNt4dsQmTs7oX7a9fesvJp8rrAmFRAXLje8IygJ3srjw5OVrU1i1/O0Q
Ua7ylwIl1ok2unT7tNcB6PeEkSOjPZ5NUnJhkuK6Gky+d0gBcCNeCMHqyWH3yyRdwmxVElHPq6gM
scu00fWlW7RhMjjmwf8WRWF2XP8nLva5QnWpcmfH7ChsgYIBwpTBr6VGo8svyIdXj0ipP3bWReGv
clcVtQO9UXgyv2fPv21OcDl6NludXiSkiDPb/CMY2tRYSBAsEfMPXftGjCCrJhT4pp7pW500to8v
s0ale7uZSbhdLmP0ETXk2bhdumcJEun9wMByCpLvP9yMB0fDvSBcBgt7tSsXtZMQ8S5cdZAIKOro
TckJb0DN+3WUQIJ4toAhYFnxvG2rjB0M+Foe6tyVQdVNlWjUUe6elQb2jqRsZE0ZKcASq9oUvdej
Ip1OsHIpndol5AH9YpUChc67k3kYQ43hJ4TiQQkGtFzxNiYgjfCx3VFaBf945OnHbMIlTLxqjjYF
CpLnbZuPR3hGnaitGbBgfzPjxKqRZIqawFjCNKKexuQk4zyGKAKWwZBvpSlEePcCOFlnK6OVVlIJ
nQVT39Y9g5rjlHA6kKVZ8mUGcJSa+dkuI92sAQg1D47d0GLmXZ3wAy8n6Ssqzo9Wh0+Y0LqgP+5L
O5MlD4P5+FxYT1AzO2+KWUAGOLbhb4WcnclsHUXtEXY6Vk/1uJJqjFHLjU4IEOx9806xCLCi0RpN
jI12IK+cE1vSSWBgF2e2lBorXRm0F34RRk/LPLOQMEeeskN1Cnlnbhx8DfbTctq1shmrPRiOwPJe
ezfhBnhWWzHQb1t90Lw9CoBc4JcuXc7opzzRFWfObu2Q2edCE1+S6aefZBgmhgDlFJa7qlwzTGzx
DuhzkFi1shOv/nKyV2FQYZyQjYWDJoNZRgqxOGH7vt1KXNZRq5CDdMsGDChvJheQPlv6SMyRHrSx
LjYScM2g698EhK1231ebSWVmeTRvBXmIzddiolgR4p/3jZ8mukxp8VKPQoMSHlJ+9Y8bCGdNg54r
qcLN5NPMvq31ZGRY+C/rkwlximTotnPFqAG3aUn02f61DYPwR8ULVrUj/bS8McefXb5P0BATuWyZ
+4hEyWDHSMFOuf+cRBOI5LHQuaC3rl9+WipSZwrP9ziHg7MW3qeE6T/ONJ3EXSEIPNuiYWyyNzxM
J2mxrtW7YvtYxibrEVZiu12StrjP7y21ojzYdiK0QZ3kg8m3tgw3QuILOt3B3xVaKP2HNRILcByw
dB+ldA/SL2nBPun0DfnOYEsRToh8DJOiA38b2TpZkBvw4qIuzoEqp/WyeLbxW8oESpTIOgdLVv5n
yipl/Zsfee6Avmy804bCFuE4KPQ0cOD3y6ydw4oSMB4HD/vcEP18pkWUh7sIz8VVmISpzjr7PMsD
/ns3MrJcnFOictU4JlyCyF+JON4oAiGsPsDPOVhTSjEojWNw7oKiUV7z/ZI5wWIsEageVbu0Mg9g
SJoET/kh7bDdua/eJry2E3kYYe4gkEhW2txt+rLBqftEHAxft8+0BWCUrDDT6cdF2qObvil5xWeG
8IhoxOqGuSO8F0AhUU1hVKeN1GriXoFptBMKi7/Xp8Q5bSWlcFf2uRcVlW7DYkiCY1IDiVvV91fJ
oylsMSRGipobFP563tstx/0rpBDJiUvUR1Jcsao1/KydDpkXee6AJQO6TUnQ7h1d5FS4bei4tL02
Z5ySa8wzQLOl1JnLLgELPQEnnUqqLZ8o+m0Z9OneihNPm7kCVpIL7ItDwf/gw03bTrqRi6FrSwtV
i0jri51I/fFXEiQWdW+JP3kNM7nGIUuoLCVUR6hgVVYQOSzf935ZHpw5FYBvZWbdEtoZmA3WxGdW
tJ6XrTj6TAMv+sWhk7At8fjRrzw4H0+hQo8BoTulmSLRW4UYsi2dnk5yOPFkjZNvxoJyL06Ro7rB
H8Vaqxfm5SLrDv5l4dVpRmde+vMxwH7zjOQ3ExOMabqoVglGAJyFphljbgKItJxraHualnXjD3vS
zqExpPsp6hUy18Kg7rktOfzCW38vEduAIbUo4a1uuo8xL8ALkWrnmBjRaB1AH4CYryDS+ktpZvO3
iXqVLyiVvrJEYT8y3l2snkxQF8CEVLp5xmKwNQ1VnImYHyXmpaQBOCcLoNo6tiCIMyCTrX5+41WH
MnFcouL05O4gb3iSysI0FYGXQd+rL8wK4R8Kzrddf8MYJXD0d9zEHyIv7uewH6h+ddaqrkum2cE/
wBkxBgcjHLTin0EhqmF7vmx57HisOOskqwq0bwS1IOwllKqHPts/p7C6wyKx2qw1Ppb5Dh0TY8OM
g9CySAbVjILUOaQVFeuBOvxIuhJOfuYVjWaMv1KYpZ8y3GArVswGKRxe+yHKJ571e06CHIqBR3EZ
yQamBfVMJQLVwKGTLO58vEodqux2ZCKf8/8CHTR4HglmhBB3+xblPyjmPaQK9JNeV++K47Pw+k/z
WOAmdcpn5E6XIOnbH227FMnXWZc6qUjST9NRHoP6kwxHRbM3nKET9DHjxYMz/d0nnOD46oXuzidH
VWfpoNobIWQf4VWZfksWTVxQbAcRCZSXsYt9tzPnNsmvY63uEH17XQk7b0b5BWMa0MmImemJx/qx
Tz2FG34NQc2kr5hub0VgqmcU93y4tA8wzCtb+6XY5jnkuz9HmCrmBet5cALj+tJEJLl82EwfmJ6d
UommhXHShfrLoZncY8hvylMFpDLjoYdHNfRio/DqWlA95ofPtuUeXM3yxLF5LGawEApqsBWlpsLV
p06ulNDX6M0UZ7eRyFH9bNNSJ98rY9YtaHzz0GayaCl5AL/6BBHmuvvkpKGZjV3CyWDNZ5A80PDJ
twwJFiqBTfHlTWZcnd+EdBBnYDkdcJPAmvVk1vUFEHJT9b8x2VIF+QPq169y5J0H10A9aF3kLq3w
QODrYaiTf9MpVIYsjut2nfmi1szoOtHH+4ooo88NCjlBQwnyY8AG0DaSR8O2s4UxzpVhUYsPUK7i
84F8PIN4M18W8yX/F8Jpjjh+o6wVvXGkuWEgjZlnLwmfeHiL6XsdQ97CpXHQrwk5+YW8uyq3AwpS
4Ouee9I4o3Qfvekr1KKAwo2etujSOYTSVFvcDZXK3KtDAKyWFd166FsLlUK33L1DEzp9sIhIUGDp
+8l2tvE/f9dqpebClI69FtZXr9OL0Hu9BX7LKFdzYzu+rDRFOCmcrVatW+j54ZlabgS97waYNLTc
zpnyKG9gIuBx9nNevIsvm9vHAOhckGKlSCwd7gns5jYpgqfZoDYldV78E6QiT0ljY/aneI4qrbft
cbN3xiE0uQufzP0TKVlpDqts1I3JTl3RutQg23eFSvxxZCB4lCk0bW3DRCLu/Mnqayz7cx84H2rQ
VB8Qx03llnn8UmwpsGEgH/99jdP7QHhgrq0ZQKJyjEIsHM0YXsDAtcCjCCwjQ+TYOoxT0tkXzn+a
0RC605LxBdm7PAUFWC52z4wr52XSUl0doy3rwQCnbjjDDnRkHFmQi588iddvHDILUWXTTMnTyIuP
9dQEyvQ4IVnC+loQOW1r9EKvgftfgZjPW6eHG7FzuIhQLrAz8jGIHV6kEPQBdEGaxkmtXnDj1ZhP
Y4J53rUnJAtiSw0zGPDAQkdHNBIbBr4862WkcIXwwsgBDTNlef1BEDsmKeHgswwBZXQ5en2KMI+E
KOqaUZs/HiJT9E9xFzjBLCzk9+qTEeq5kHpPY/zTKrwUC0WPY4D5k22+vNiJZnQY/pY6nrva+wcz
3ADFN9s2Z8U66/rzCPhuegl2JTIjouaeVZUM1cOwm4sij0rERtY8r06VjVvU8pCfQdLOut0KA0VH
aotUmdKOCh5q/7WdpMhWTtguAk1RAy99RrorIQW6u5nE9VZn3iHCuypOefq1wKtoT8TnaXv8ZJzB
lGRCNufe7svZW5MTgCM2cNq3PrlGzKRLHy1xCeRAN5p9/QUwkEHG/+uABKp5s3B3xCASzXQ/hccu
wTbEh/OspvzKJmLMv2bvYS4Ljt+175ITn1P5BGmrZEMi/YrAg93ZvukgkrVMOIm7Q97UT9I55wef
CXbWCkGNofaK5D+LpifdtSGUT03g35rLwJLNdJ6imSbFrT9/qc7YTvPu9h8gXHRfkD/aq/PHob8/
m1FuyxQdTSbU05JfZhtE24brpZ27xSygVEMpgHTUTQvD+TuoS0qgCVZOSWz11T6qgWDULkZO1bOJ
0iavxVvGVBEBNBlhypaNM2riKE2Olg2RmWBTFDVcm8O5emiRAWEaEdRSLT4py+Ro1UkK3PKvhdWH
D9kCpe79Fe557qTNHZSF5eLpGpZC3Az57qWylio/inKGApMYxCqpmEvz2UEmxxspU3UkhAfe08jl
mCamOSi0lcIcsDa/xABUI8LYpXi73hS6ZGWNI6Wa9txru9YLcwZjlyPJi0CEXCK/UNKBbpMC+U1U
5tSIpGLESb5huNoZsZQkwwCa0L6yqHdrEWl1557a8IUbhOChAs+6copR6NCoLhSysjcCv87Wt1+9
YiyabsUFk7qWYqMnzd9bjP3mHy1Tfotx//qFzLlaN94VCvV1Nx8UdRzUSzuxGNERWQR63RdBGrpC
EzHUHSDdGYoAzsfY3bMDkBMhxwoH3wn8xsI8eAquae86PK/cuDHQVt5idDy3MB3ts+w21HkcWunG
Oevr+XHkaFkShIw8W+CvvG4TNGFavj+AaUxvT81QY8GHFq6Wcq5dxIAWAnFZEwVnyP30g++lZEPP
GH04ioTdzi3397iHcyaGMwPnzXU6UofpSo6W+fgJt+Gv744XS0pJWAcjx7AgeXQVTgV98c4rXIbz
S+aRPkezSPjGf9aKqtveRpYwFi8TOMGml6PRvn4qJO7crCfeFCqWh6aczlGrhlyvbHtpheti2VL1
KXDF93h4ve6eHliI+wcpXDc0XJ4aGLO1w7PT07hOic8sF9ZbC/CzjtUeYqhhXqPys/Rp4OaqE0t9
3H64SaxOycCjB80uKKRa5jDH7RVC6HqAYov7eryH5fZgERy+6pgpsMEQDVDJB5JHucSZURa+s/Yc
vWRw2mz1BdQKJobih+a/xZgO14mgjpWZ+wlCxN9M29eZZ0ec34qILTjMSlEwAHiuz7lUU+SaBPXv
13Z1rE3Z+dmiNBYubXJNZBjkWZmjC7tODlqHbt7MBaza7MKxec7uvfoRkP443avtC6go3y4+jvJg
XgeK2tE9Z0ErZgZ9+/jpJvSAHIgrCsDzQ52bJojbu6oEaEJenhmpqY8f2YxlMZ0zhzIkS4Te0lMK
NoR/14oFT6vLg05SgIjiMqmrMa9wjhJrfCIB2RwnyOPU11aj9UJT+38yFHA4PkCs6E/GEVCWTpLk
q0Jq5GknjqEUvc4bhbhfhV0RHwwMwtW3dWSYO3YyqnUDn3k1RUCUB6+DsO1zvca8lRNz+HlbZ9BP
7iERcOPWDKQjwVY7I4/2iujkk/Q92BcZLS0QO+UhAQzwlEh8grXp2g5q9ozXeETczWQpZ5aJIl8w
+7mqqPT2CVWQLhDKNsrF+TA0aH2cTA4TbA3Qv0yM7awAJ8xKw2wbCbwrNOSuoDBiZCH6Ttnb0Wk9
IV9x5VoAs/i/VftBLk33lCoz7OxOQIB8maTIKtZU5/AmSD0s8dCKWX1tXutgwpAQZZYzChv625gG
mAPHkPbOqt6lo6dsyboB4HNnq+mUQvGdE4VfetM4etpTbfh7BVZjcXz3re32xXEBlHiLDWpIcYYa
HE6eRv+SOr+mk3SBKyGlzF3Ikdf8Ugkmm8iqJoFK30BU/sxA6N4sDF8cHHzj27l4ZLYKieJMzMB5
cBK+lydK7D//xOpNWPFKCorYddvai+J1YMxlliqOKsYk49s9eRJv+VKZP18lXCmhdE11do6BRTRU
qaAMVYK9pmFhlT6zxCgJgi64lAU+PIEWJ864WlZ/kKL8Hbx89UDaMwI5baD2csmryUSbCjRzlzrs
cDZKKpVcnlkIUhQgqMOF3lEg8DvaBqvlt9UXTiRl4US34TYsCYqIA3CE7s7WqI9Z7W5kXsYt6VV/
z8UIEoDqJdM3G8LcCLthMgD4vbwOfnI8BmvYzZNzGb54Ta8q9KnWciFF8ADj9vE3ucVffUBtby0J
/8VE7g8We0jgvypA2FSkn4EQSqhz7hEsfIkKliW0pw0bHQLtlYBIldhUVppGiSfojKJmJehZh0+U
4q2hy0QXSf3uAYFVgEWkJbeU9WpinLP+yl5vbIjtukuC/ra0+zsPOHigga/yg/KnYTMHsN30hAyC
FcRWChBIhlfaocRKu2l/AGXQBM71yvTKcWqvIbqTldCjXahT8NMU8Q5fO83LaH+cGvTMeWnD/zQy
/i0+ICZN4tYuMxi/30iF4/wDRxmt+usXIf7z95YK6qn7vdybJ2Wul10al1DirWuDlWkkEQZbqM28
VssF3cBFacTCr24/PUw1p9dcE2UJAEDu3cQ69g1DYdkjw1NYv4MvZp5sPPmLR/1/bzkesJpId8Ow
6bCpZFZnalo5p7WCKTs9V4K9mo/h8R8lWg7uIAiO40y0dqbwoXaGJo/7mQTkTUBgUJgzHY3NVMk2
JL86zaaLShsk2vY7uzv4QrY4TJNbDsyUkB588SCXF8CBZbRjEcFpSL6i1qFnluAyhKcQ+TdaPCOJ
933Z/ferAu1TcPyGQmDRHJYF9HJMKcQVLi7V/H0rOSoMUJmKeohOX9HCPnLwtboorLMxiff2xNfy
oqjtpzwTfcC0kzVr7pnnjn8UXFXPzX+Ep1qhvtblp4fvr59+7DiRkBOG74Yl0PltUni5Ps/80Waf
0tC3EJTkTtlxmtw68A2AErcEUn70PUjQVsU9xGdRJEU+vTpL393rTrq1Vlxwqo3CifJBMdOes81F
+/mhZbeJnYXjZa65yPawdhBXjp/DDDUywipdjoVOGv0gE8lQD2vO0X54s4V8YPlB4SLYDBT6Xtit
KY0atczq1ekP+g/VMbro9FTdBUTH7LYOqfmmYe8IJW0fJEXRTOeTytuG1h4SIogHe2Tp6Zx7ic38
AulmRy78LYYiEzKNfLzsiHx+5OVk5UjUeDmrRFzf5pjsIIXEtvRUy4Ukm7mzue7sHlS4xFivyjKH
gDWhKNBQ7Orlq5gLT0T7gnXLEGFGemg+PeT8skuqlGob1a9h/TrOGEGmNwLP6nSJf6E9P+wPtvCq
OAM/6To49nF1H9qCrKgB3K9Dwje8b1XMXzUCdzf5aIhssN6uK63qNm/pjcENPk4J0CBvnpvBcACh
av/slbmuhfUvuyskTk9KpRFIRqOPT1LAxgttRAv7JNXT8pw12HeSphJ+h7NTbj7c1yngJr1zUSdD
A2GjWgg3mjdQkxADHJaSYKhbaqDiJVXbiJ7Hpm5FqLt/DbG5qGai1zM2Ea8bDSPqgLkjcfA4kBvL
nWEl3Uy5TpvNG9mHwsZTzgL7LiY5Jztr48R81RDkjozelmBY2jZu+z7sFPaltbs7Mf88zztGkPf0
LlkcVSRXyk7mtIbdLSXdDk99MczkPKjb1/qhdOPQGCw7lErU3ycedmmuoA7Dh+3qfPUDg7TA9w4K
CremoDGlRtzocHunZz7URMP1/JT2oKXCaV3oO9G+yALmsQiFoD1fN+Yb5g9/e8prf1UR7OGRHnq4
VSGCBs8U2gXmM6lMz0guHu7jMNTnR7h0EOJYRp5w45VC7qY9p5Nm0G72wYnXBhs/HdTfflp9pcPw
ABPI8ntq+ayP/TfoznAV+Kx4OuYoOpxL0Cxi0IjfQ9m9DaET+pg637JeSaVCxa5znuvUbQZiaM3n
+uD4lEkjafx2inRmPLnSi0aGSkG8uNX+u48mXf9oswqgVvH1lXyU9OhIw75746rs/vTQcY/pIk/Q
oocNTB/HRvBOUM2100ztWG9EKocEYSuHNxlU/OW7mFPcUft8S1X4HhHG2hwaNJpo1qYAUnZ8AwOU
QRAUVU8RoIwjP6Kmt2tTRc/vys8JmVCnZ1+j67Mp34aPDuORu+nBceQ4Y3WdlS9vKyyzSGqPVRKG
/feqVGuJ9MixgLW1NY74NCm2aWKoniVN8K6pwWKT7mvKy2JOpvdKAptlFwqLcSAW6O2Tzaq0hmGU
lxwWEAac2Byk4FqbvJ0PolF4FVWFjdBeDuzrT+UOBELoBThACCbIwLVowE3BuV/FavO+fVS7uU3P
/bJuiuNG9eys9gm5ej069La0I+YZlOUwDMOnAA2J+fvRzqJKFGqFpWuws8OumjUh2WaARfvBNINo
XDMa/e+/dQmLflCs4LASPsNWjchyuc7Xi9z4dL9js0jLlR0BelvKkHozmYiJy1N5wHA0GYdLf69Y
ARQj/EgkxOhPwaB9MEyKJAakQddpIDcMk5iqEvZLJujFwvarAFcxx2dyES8U3hUnud8K44dUStU8
/KzJ3oV16IfADdqGvhPDGEGzu0rs8PUNnTlSbU/D0+ggPDfp7xeojgwHFcy2sOI2joBlcPjqPNN3
++sQ+8MRZ9VHJhq94eDN3BLZPNl5gU9yz8kFPFhz0qKqTfzxHdfNrwxUNGkd74E0BqJxu5Jqg/Im
/twsvgRIboKxnj4fM0VF32gsCnpRMfDFeFh9EbV9ikZ1urPn1W6BztAq/zuCxUFufSRUVBMq3cDY
4R4vgz45x0hS/Jj8UowrSjGQ1Imt2b3jddPdFMqerHw5y6QN1KuR7V8ppR9E1QksNlpKmlg4KnV3
2J4WEuHK2ZJaPEjqrMB/GxwdpgVzf264O+segk13AVt2gT5BUwTT0cttbVOTnhyh2x1AcvA3xl3V
txUISRRXdTg6+7Q1WKkG5OIcxMb7iT+cn4Z1AYWb2t42ItbrDfB2dZiowX52vPxRIOc5j+EjDS5G
9xCfMPOzJC23Z9ls8VxzRsSkzhaSQOHyXMT7W5LjMv+tf/9xO66FqZJDWDmQkBAAHS9f+wA0xOmN
9uQdNOhAAAAofkzN4RvTOAugAXOgGiuMHTmOi7XABgYIbxDpHM4CICAdJqRkd4iLfEr1+ljJJuH4
iXVfo56KCruP0o3IjyVWmiLhUcYX0zU0nbmloGgmhMUVsPQzDiGtKhgNyCFyC6RKipTELbpRfLno
63dC8devLN5Bk++Mm31GZpFMhN9l8+hpu4ZAfra6m7yU5aMw2cVI19s1F8SnlfoN/jcNRq4BfvZs
+DbTgAZBqtfrR76Pt0NAazGsJuhObTbYD1C9IrAFXp5NNFj4KnM5GmCgm/vjyapSF7cDcPZDjaXA
gI0h8tk2eL6wons5WAB8QnO8CBei8DDXaSKMBjgDX5ldGzuCADgR83A3VIvCHbvd23Wk0AgO86NY
RIY7imlxGDUcCGP2ln4XVAODWXaJfr7xRxmdAgFedKDDBM4vJM8D1PZ7J4O+jK0f0Ka3SarfjmM1
aYVh1RSNyi13mi0XgFTe0B95uRz/k8hIhKGErKR2fLuHlzg8T1cit89cG8kZU/bq1IYXc9TWp1hf
vHVglgdqFlPYrTPuNd15lQiEE6u2mP4HljS55DZO1I5+tMzpPAptKkNKhwZcHqpiSxqUqjqWrhbl
RWfWImVMdme2Wzu3PUHfr8uXDFIJNDB++1Tgnc2KsLSTiByYaMZv4zHw3vLj3VUDVaN9B1ISgP4H
Lk1ZaNEVB9gRoOOrrCgbq/vWhLeodTYNdYqeSVg3jFhf8AKw0yfZxoReIhSYQpJ2J6jSXWE1S4AQ
yqn0eaxsDNDKSpPyqVDMS2RCAQfo03ntgqhkmiXxUNUZpre4pDsvl63FvuF5LQfJZKvzKSjPjtjh
yNpFcdF+nPepBfT2FB+s8JIn+QTg2a61x+G2nK4yzvmixtDIRhtXvxf2AKbQB1xtneFcPGrJer3y
8z1H6C1SiVjGdEG3vqYwjX68a0EdNqppJ/nR52IuqFwH/5lwEY/c9Rg6UKQBAGXx6CnSJ1QPYlqa
YA5hVBFWbAGh+VcWa3St82UzNVPXhz+1siBOkLrGt/ttvdno7iZVTWYb9yEPYzIS3/qmk9cbmwu8
clM44MdYFX9EYZYTcIZh55r78Iu1KgsHBDI5zQ+m0GDmHw8oOCYLIXOy4uSsmIbhSAq/6zxaB8Ms
6aYhEQIP+y6sFi/HCEXpf52PKymz+XVXHpmWOIMPH7RgSoeXirFQgNUdvVbkS7dnS3xly0kxn5t+
n3J3efre8yYoXrqvzb+nt0shXCQEAXGdyEpBl6NtGqWL8LVosWqRrUsTFs19hH+X9F2y4hcfmZmJ
jXM0IsdfERWr3RcFr2s3LygbCJAOcwmsaGUPECeV/3Mf8ONE/ZVha46nxmZWhG6I1E8jTSihH58h
hxzczulCPtLARwZ6t833si3i+XNtXk7KpuFWS9scbgy7nZMW4t0O99ffcYM5bGKCkVMPHFixOiC5
WgJAk9hcLg567thJG0YTg68Qs9H2c1PeeQw/FaNYx46+VFncOyq2elpJqTHtDA/PPf/MCGaURyBG
VUxaA732hHJM2DOhojUGhYaYxI9p3TFjqBwOVFwdE9Zvgnlk5VXnD5eKCcKC/GrbgEt4Nmkp8GtX
VFezRVs8ApMYQRTtNGiC0Zo3/vZXMieqBWHadk5sk6ImMjaYlWgZ7TjSKNYgVJ1TgKrVkJDhwDHz
0/TLnnKyt0xahVqUFQi9xHbfklcvmWGOzGLPo7fxswXwYH1e+x080tyrlfdMzW8odxK3S7U6+KhQ
cq08iXCJk/oPOGv17fixKRoqFrTNg4dKaCkXlz0RiRorALRpbOqRl39TqFOjh6Hfot/zNeZkYxE2
W2VQ26m/ixqktWIQCDeRP4OUtHPbTc8w0PpNwoWj7oqQ/nnkh5lt5Hn7IhugHzAuHs0U3HsUMqEe
uWQzuTPXeL9qXAXjv4/XOaT40M7xJlhCxn5ORGHcDnKpI1pabm136uaj1xpUrhIsZN/slx4pufNg
AXRUb779r8+8ewWXLpSMwP57YOps6XMc8/NBvmuQ3KVJ2Mj39SIflcgFSVFJiqC9puLGa4SpyFNt
4NPcHD/Bsqg2ZQDVspmhLGDpw/piVJub5Th8cKWAq2VUeKo5U7KVbrQ+eJ5YqSA+g72ANId0FaWP
bI3HOuFPAH2Mnh4Y3ZuVFCNOvlZwaAkMc8zzYY1gXzVKgcnXIauJkbBg+lMES7u2c55rNRgDBUMN
oYFeIzvacVHZ1Cl3DYkU2oP4540V+WZt5AuP54tVy1jNuTVfJ46XhL5fxxBVtpeOjCoHh6TNGYRx
6sHEjwdDGw8C15/hsP4WEJOoyJYhp90WfmNPPgMDDtY4yiEa/wYnYppRzg6vmKFJCM6zC1tfgP5T
J59t71Tt7kjiSqJjkdhLZKeMhxyxrCycgLTAVk4lkNjq2OaCAMkkmk1ZHfTJuoQXHDHQrlplUF0H
2KgTlkcIt6G1MmTYPHy5qR9/ASvfRE3nLzKFJRvHxDaGs3jP2vLrOkPZp+wIJrqXWqRHkXWZNEPw
+JMcJFzd7jX6KQyNfPLQVrVsK12OW5skOmYbCv3LZ3NAJwS6kiSA0vWQPC0xStUrEyQz6noP9F1R
P+Kb1nOYWruqYDm0GT1v5+rWixY6HtnBuzJ32cW7CyX1q9HSkKJDK2CmkutvgiTr39ZLX2fmupFg
UnBgqySoZQWgPv87m69Gk4s+Q/CnAt9qj+W13lq1jQ/cAMRWQRKs5Lf0KMXhG4kDVOeIssxhCu0x
PYNn9RdGINAFIKnX8MDUtGk3P+aFDPq/OXkM9zSS4n3ekieInoK9dxKDUppQutUSiUVxMx6x0H6T
qXUQj8Z2HEr3HQK6CDktnvGieqGqJfbI+aLFNqt4WyD4BlD9xyJ+gxL1u704YGudEyDFf2EEWItG
EY3h+T24Xf0Xe+3lDv02IRmInqUKlQ0NwRbgmIxwwdh2gvJQ2re2SW+DGZzrCJ1DW9KO4arogXwL
YA4RScDan1WA+09NgpgmwLhe3DKwPIwbFzFEcH0Rsh0i/UE9I36voPr1lD0U2U/y5nSsFcbN1HWO
jl9JJCd0pG5rrOLeTTUCSvFHPNGV/wTgDz2c90sBe7pO1bt1gaNqBZvovSPVBzROUSumD39Q6fDP
BarlD66C99lFDzqGWiq2thWpUfFVgsdchv9LR5XXp8iWKErXdukNroZLVg8Sl1SYtjsSqAh4hZmJ
Xa8macrvVLnC+sJvkpJw+QRKPKesXn4FgiOYSygWs2Dn5VlHNI2TSTL3KaGpCMq2uDQ5gazG2Y8x
0saiG7mHliwmUmaMZYbUsu3bf+tGYtDg0b2cbTvdiSVtEF803Ww9ju04iuLoLJD5Q1UakyHauKSI
BnxyfV3r/zhNJ1RtGLp3fhnUh99bF95hytwJwpHlYiWOKTyHp4AZ0iaxdLMgK8rVfMPm4QanDjPX
AN0H780Cr7Rl1JmCAo0g03sPd7RFGsYPA3DCR8NCfZ+hJiteVaGh1PE/+EGJEk37GGcdVtA3AHPS
jeZzwOr0K9CGxF0wHIzeuOgtKN//LlNdOE4HZV00XNwLDdlycFf7YAqGwM0oxJkEzM/tVVCqC067
jAG8a704KLGEuuAFvDVqAkeSJkiifKrF9Wz5f06hNDWGXxsch1UhMLsa1yYdg2DLrTFASuI/ztAj
/jyrHzOQVByDc7dyhLoqUecf14TvvgrUSNX2nguwvNbSnkkcyaTjJoWWBnYcXZQl3opkOj69Tdsn
cpdraeBHvIEAD3ksZkAm0evF0B/jGEHkhPbQKglVcvbuXeU6koaxqmDFTmm3JxAmXBGFpF6mhCpM
MpyGdnS9n2WB0lYc6GAzEa+D1BgApL/5cydgh7PSapHUCEf/roPXEExRyJEj4NIe34Vri2Q0wUik
Pv92FUR4rDv6uYrf//6HmNJJJJO9o33wgrG/89/A/c6lmBMa6BtFhSEFAgh30RFyZkbWeWSrwGUr
TQ+fDPrmUvArXbUeIrw8whStCr+MHBa8v4DtIBJBxg5MQ+q3w4zqTrRhpKmsYc6cgqqH5+Ix+Ifn
Ds4hhWJWbOjU1KtGraI0tKr+zN+Emj9iIju6Jq4NU3QzM5gAzcEn575hEWpVvgHfPIxXrko6VQXN
mwg1mw7tqL8FMvlxhkCcr4a7EffpO7bvtevZwPzdGFk248wj2fjqIUKLza9Aa4tED+tMKmidcHQt
i+TGKsDJV5dlnwS3lZeCRT69L5kxRp+eFyKbTn3ELw3A4Edh7V7SylH4aDgTbfF+whbgJY+9ghbI
YPpnIQMWKqDwy5JaCtNrkjnLi4bojmtWflK7wwSS693ZYXNri4K5q1hWZGZ3la4ScZCeLQzx5x/A
ZUJyrcxy8F/NylIgPCbQIWDc1PVvY9ifliEZw5JZPofW904Ekz8Et5q/U9LpVfpbhQfgUROXEWRD
IK4jmTrYsH4TxMHBKy0L+XyhUq2aSIZobNS5VCK9teJ20RJvAJIgpnwI8MDFcLlr66MXZID2aqZn
txaVJTGI8auQf0c2nbb99T4k1sThgrKO3DzFXC3TLZnpDwlaVesYOliU5mjVEGoJkELva+qi7zHO
BYzLaUeZ4qHDyvik0vKDqVvejUfqp5XntNj4NLmouZJ9cGT9YgbFXOn+5PP73z3tWPalAQvZhvJo
R4sXFsNNGm6Ow8WuX6Crw2LKisAC1Om6lqDfGQAHMrAuNylws95nZUQFgBKYk8vc5Cp1DjKpb4rZ
rocXNC+/MouxhElLfpQwQnYHVCsc/Mdi7Vbvk6WmbfGDxx3EVsxS+fENHx8nIvJrARUAa/5aGl8e
nsjts+GthFoGMb8yZXULEkgogHhf/XUI5muYVRrBMZ5KDSbsNK/ocDQfknRoQKR96PicZTAW6430
pyrUZqxu+Ta1NlBpXnBS72SrYVx9Stad4oEnIwUc2bkR/l6T/6GzWlNQzMcScEccsd6MTtazlmEP
jVLN0tBr8sJ9nc8Eufc5lOkjD9eOEk3AC/TBGlBGo18xavn5ErenICrZrf3w1QnaY2Auxfq/15O9
JxoxjkiWGAhBF7nunSf6lBGZu3/Pnz32E8//fCzp70h68fZTPQc9JkZ6ytcCyOp5KpSosHgpvvPW
GLznNF9pw5lj1HVhzL8OAJHF7gxGOEnpnSXZiTH8yqJ8jXLZDJxmqFSDcx7qHQeJnnefX+00jOuB
a/I4bo26rwspXdUt28Sc3b3hNy0JPJD0f3d9r4VVzbv0kvz6yobKH9DmlGtnmMoFIwwYENlMlNMa
04Gi9w/Gjy0MTFGKCKIplFefkUrXNPBygi43k64AQZePC+m5cxb/7meaTz/lnDyZ+s8PNhUcyUXB
LLVnevH5Y/OlN3ynhgaRJJPdmi2/ZNISW4D6YBx6AQK5Ih3WaMBfq5xbg+g5jrxYCUeLJ8Vfgl27
W+6vhBKWTfLZzu2cpkz2KDc9fT5IjFZZLJuHX6bRX3yBb8hhL4Y6ZG03jDuUeAmEOR776A2POKXl
nFx2NYTJZu30O1uXRXPxQA6BCFqqeHFow2MbRvm/Y+VZlmtlQS6Yg/zn9ci+jpsxuwhQRDaAM8B+
VkjMwk6tUJi3ojcQvfxEcqnKbU+aEOYTf23ij/w6BhOMfv3bNlL85UtmTFUyvZ3Ju358SfPIkuZQ
tCg3sNGyawA+IovPynmEK+IdgQpGKko/4Gjws+jpRpQugStmWaHgdEQDvP9gJoxLfi2GLIZw0CfV
9bCkjEB2ti61FMsFDhGJLpM1iiX7FNkP/rEft/qASsM5vMJW0JG6Cs8fsa7ik5vCAnp1LDO5+G80
jGD18DAr718ts1XvHpx6a9u6zLEkRv6dJe4PKl4EXRzHI6G3fkyF72WJfgAytZBq8ncIeGG7CSJj
VpWKEJQu9HHhk1e2E8fzo7QhOJswIb8HBpXAbKBAyNUYF1Rhh/bD174JFL9iI+9e1YzttJQEqHKV
xyvJ8swODViZLooRhwVWPWvh5rBrAALL+kUekAu5sQWNm4tFTjr3Sj0bHA5MVdUibQpK720ysZUM
yKXEaaJpQ5ZiXoUl+3IPttlA4cZLEFi3syKwj/58hZ90PsxuRhThCQK2M6WtiENno1zdG4o5vRyS
5wKPIKpwvDei+Ixopvd42s8XFy49g7CCkIhBfyXYOEgXkR4aAX7wsIcEOzJVs/A7Xq68fkrOcM3N
uCLVXcYA+Itzjz637IGZS12qmPdDneAojIsI+6OfIIT7nePf2Rd64ec7UD8IMaEB2fUqnXza+PuC
E2rbZiHTIC+WSy0SXG+j68XjoPgMAe2PePLpJIevqcohNxzGVjaLQe4NAHrrjSYLdPJRSOfxAH4I
nKVrxtQJAH08VHMpmH7zsrvvTRgWpx0Ge5Baxq4zS/IeXSvuieG/pLFPSScVUXCBeSEENxZS/qZR
uuJsFHkdgzaPF9jITmCNbnq22cO/KztrZLzhv+dtfZRTFs0mh+wOAyCUsMoqbx3NGogSoND6gMCk
guDAi2xnjYUM51zbchrI5WA/DhQcrNEUrn9oy9MHkITL+JRDmG9DYwklnK/OKD7ZGowfrT34390b
9PIYkDVbpGQhfoog/rWBIhiPOQ58O6pwzOok2QYo3dOnUbyVZKdWV4POPePieviWwOcF4P5QHlWg
tH0qI0honauWTTWpCSqhjjEpP5n5jxi6ZuX+aZgJWvFycybqBayW3CZXgtPBhFg0q/rn2WgJif2S
deusmlNg5DV49ufqx9PCIrV/AvdMbzsZeYPCHZmMM2qOzaZu4V/IkgnhDxvyqjP4rmhbCx3bb4hL
uEZS7xu4bjhdEWVJoa3KtBcuHcx2uFAMq01+qnbIaPDcrMCxgOcoCAase+6d8Lm9VeIm2SyAGgKM
0V0xrEc2AqfbwhJt4flr23NxShK8faydmRk7/4fh2ZSijNnv5auWL59VAPiSeQFmeTj8iHA2u5D2
l5au6WXjOprVUG9ljwxs7WxSZ1+EcnBWTg/jtH1vVJBFzDN9xl6/a616In2ZJ6DT867Q1VYE5f0p
EyPnz0ANpaanSmuF8/Pb+QLNiHuExngax9oMhH5IqO7LxHi5bTAaYjEgwYJEHfQkhEXHYGlQm6c8
SQQnS4yn9gJw8lAh94mRAI1E28OkKab6Pp+s00hJJe/DJcP1DsA65HbOs/r4mhvA9VVwxojpQjiM
zp0nZplQ9OUInmSKdvtrD3v5uFX3vhkl36FdRkWgdY4eMGMtAqeUXOjYilPH2d5gQ7Tazx7uSjhu
LtkWnev+Qvvt9NhlRLOt28rZpdXLH/QlHjA/Oyo+KdB7F0pegmCzJKr8aKJ9Xd7i0FReCtKt1Ntd
LMFezoD/uNl1GnYLdC3axXiNXjn23AY7+Tv6zoUUBln6rcEHMYZWpEnC6XBbNKQNM8Bb0lBNpVt4
31KNnXIhqWS3cmRmg8I1TVAyi9Y7GCwSMO7/nmmuHSyykvWHual3V98uIZYjPCi4qZ8ILiGHOago
VddlKabrdCpew//bjXr6sN4i2SriE1iR6Vjc6UjDItU+At46GN1DkuYfsWNbWrHsE7aVk5RtEb1A
hJp7fdhoABbTLtddE8cCR1LDxgLdHDtjV+Le7Df8MznQWn8vFpUF53OgXa9vBxnfvCx9+miHWc77
vhkQTxxn83LDQVKawhyxBs7EHG6CKGKgL8D7W+ymMDBad8pP5668CFb1WTEWhQVAJZeLR8wKR/2L
d5rv+AdriD8R0XI/LfBOEbbZSjly6+aqUBFoj5mQ9iAURNYY0utNivd0TQmvg6Yz9eDtXXKH5ys3
LL/KDmQdHn0uEyMyXnqqlazv/MQWCEX5cH4rrgsA4G6o/Czc74SCmx1JRnxYZGT5YZcud9HgVTK3
6SDRmlu6qsAxIhsBJ/ToUja4NnyFTLPW4PxqS94CyCRjErLsKVLgUcj69HNbW44mtCrKKAQDxWP5
q5YEBZWYR/GDeZSLTeFm1+GhV30tGaYEg6ui4yEVZY6nSH0nO257fGCnu8N0sR937uHvUFpRk4XP
weq43XanI8LBBW/D9GcUl8sAg6orIMZUBJ86B8KXRFov2QE/8EcTStUg8CIXV0Dqn8EaTj1akjsQ
libqM1ybLOBCh6+UISDrr1gFxtyC9YjhS/GMEcLRVdLTRlsr4NVaS6+6eAvT5lU7amzIUJLGbE4D
Akl+cAp0o2LrHpUTNu6vjib+1CDrmgHzY4Vl96D1gSko2WOvlvGWs7qz2w0WIIrCQxwHswxt684P
7n02VZu9YElOJcHkA4eTqM7pQekSGwEOg+0lJWyEnBC+Yf3xzMWg+nUwks6iVzXE23/jw9Ivl0ob
gAFxa9IjeWF5WK2Umj78I7tSudhRAaPbVGUzeAp88af0vuwBfZS4UwDzTUC0VHiyK1GgNwZbmxKu
lMOOrJH8E6QSYkXBpiq0yOQn8ltXs+d1784f9Rdm67NfpNzMRQzY3H0qRXBvSUvk8pJlXUPWEOpg
WOfgE3COCHigdcjrD7xOEMfjYkHdK0LM3816+YmuPT6r/gvg8glGgdeFdw+I9ztvalhehuC4GVAD
WDzoi2E2Ugb0JR/kF+iOvqhfYJb7QINoSrS/OOCO3mHXusB+AX6VTb53vpe6Mq3B6ljs4gbUGgvV
CpZEmYx05S7DejGxglysEvTfLqSkNkqp3nkMrUfHimFSaOd3VW5QK6rEge3Ig7USJndHOjf+RjTE
MhBl+eF1i4uKkoSTNioKtThQc1Pjq4rC9EpHpwFhh01r7iOB3wDu8sbjWT+vE5A7WOPTqk1FA18g
JRdheh+SiWeEhdBlsriwYxdk3dI/K8hVHz2jtgOtIEemOY3tac6XYsXhc3ZLOpmixmmM11fcSVV9
2bfpSX2nayc5T1PGFXfG/AfHqgiQyBxuy0VKehSAWrPlQcjbcFvc7hVGuSGyiKqYSmx26nhdk2p4
gi/wfoHRz71/mTC3aqI8AiJ9cThFnCGmucVUwSWiZtLiQYah4LSDPH1KDwrP90MjxbQAyeEo7K5N
7gGOVJ81cHYJ03Cbcj++lW7Xu1nmSeMwXN1iN0zKsZYcxs3EuQJGgmKJzuQ4ADFn9TK1UuJwxZ7Y
H+MA8WcWyLEgavE7s5BRNK7g+XIpl4hFrAfj3Db6GSm7Fvt2utr5zvFVcsfIbDG9H2fUjgavnn0C
Sfw7x6OWJuwklG3RGzOHF0n2e0wKuZOFlik34Sgxd/f+ciT4clS3p65q0UnUbnoXTFwwtrLnqODG
u5MEfcX+NA7Pp5Ic20x1+NGyyMIkWLdVrUs5RIuTaHzUxTvx1vIuEeuIrBsk1/0/qhKTuiUevM0v
NHQXq8LyLwdY7oFO6UjnwfdCPss2NF0yryAgC2orPlg996+5oKF6wYbNbx6YMAa7IRuiNTVAqKf5
GLCVynhedafyIkvJIl6Wb//tKqccZDubunftB3/l/5La6CsnKBmbQ8Wjr5lt0YIr7B8yQwgue/0t
cdOW55unKwwjyRSRhNeSkA7roPaEK9UUvXo3H2xy9ZSJjKs3rIdeeBRwlUn58ufRlXagRvz3K3HA
qwyrqaEhGNZBnUX791FmpfYLmWOjekD5wIpX/s7R4N+hcP1bBCvziZbHZB4stxvrPRPgCfKi+yZL
t0B6rt+nVCDlUx4xd9l4gMmELr2nHR35LlJ8W7jS42+hQHnQRl3r0GN0Sx+Vel5Y5umerZlILNdZ
d08iXbGOA1pLpj5TuajhG2imYZdOAdbwv7MBJjBANAejiSdeQX1wq7Q29ayVlahVMd6PUoly2h9P
DjMwTuxEnO+zHEblP4Qn4izI9IrJFJLSiBSQl3FhH+euJpxTCxhvU4b6kY5/2DhxItDdx593OQ/R
valR/dGFHdl3r48RiMyjvTbQW/nhpn1dz08wvJ4J+eUZffGOqIaZdmW+cZ0SMgi1sdflEEn4uYTz
05Em4Fb1LWoJ+Pej9krIlPU997dQDfaLG25lHCYRtLGIbnYnw/JBD5Bl10ZxakWJxwseCcO+GaSi
wIHUiBdl7bX2/4qPNb7FRU+XqzITxpjv4vZH0JPIVDscCbZg0oQV/Nzpq2RWEya2l1obSwviFu9Q
vPQbRMDbjoMfx791wCbcu2T8MXC5t8BZUOLGUtvCnXW9sZgKEkgs5pLTo7AAgqnsEWxgIhQ1o3EQ
Ly1whVMTa6I/r5xcXJHp32M3iCDfkQ4D/xK/CVq8baL+ev78feJbtJppXsg4o8Td4VduutO7sUSe
MRzWkbbrmr9B16HDbAhpBwIFRKDjB3B0WkkB8nuzvNLE/sTcWMyzqpowTrYE+0DF/k2TjNZhJqdk
ey4ALmEuF5mQJZ0CBypIbrQ6xj4vXShz7k6v+P3f8kV5LTVKaVXf1FssWqnGjxx12tkipZ6MJ2CO
7QT4/9WQMWnM4HY/oFC0uKRDDjJq61vCkn5UU1uI4BtOJhcXlU1LOL+qvdqNyGR6fz11uWlNjfnW
9EAs9+rI2SoHKZasL31pPgTmsACc6r5A3SBYq5c3PqNx3s3j7NwxO9kBd02d/v+PgkW55WIykDPH
mxoA7Wv0/aKlsrGviMTw2KknTsOnAGADF/wbV2CYMGyu1CSR8uXty8/zhX7kRdlePbgSIFogO8pK
uxCzovG1+6UWestVeuwPFJET1WzMbcLw/u6I0uz479Y+VBTnhPCx8rCAdyTdbX0EW9dGx5YsteS8
nXlGyPKhfmzds30b8b95T+/A3vPYaJcPIM6iqDg2oe0fcN6tIWWOxGsjwr3O+gb1kfADJ5FAIwMR
wh3GiR3+JD/0fDtqJ5GG4IAzZhahHM7MOaNahmL17/4O/90ouQimXjWuXwBo1JSvFkcJ2yVVzBRD
fxxEUMzLsq6vddgAycAU+yFeNvk3Dcdl//9LUDrefuXTJ0JShogoVxOO/S+Eel0Nyu6/6bjclOx4
tQxmX2KowOEGecLlwFStrwmwq8bgGlbrKLRbRNJeFGjl3jZ9iR1/DD1cwJk4VFi9EmgHyFb6dua+
VN1stjPzZTPbQGwUPNfhI+RvPyDtxQCrwJxHp2K7Z8OrG7oi8Oki4Yq9FLNwhrERJ+vaxPs/3YLS
UaCB+mYQc4rlQ58cdQlc0AU3IiGkntAnhW0KfNoh/wscwVTtyKM72SJwmDbOcXPxGLBuEqPoGq+v
1thHCaiTJnUpyyngQnXFZCf0tZyqxj0zJkjhuRnu8my07RCSDZrSIidYA5nfz1zm/FQIykaknJ/r
KS5aYXPyakURpDrJ9rqm1T+f9XN6vWjmzA/gVXtFVtqig0XDGuuueR5/yS14yx/PKMyyd4xS0GcD
6thQpFpuoJKu96jWix13TTc6oA1titTjEA2TA8VTtyTO5k9/dDTqYqIEAXBQWR+lV1mulln9O3cb
pe9mfx0brjpnt2kp0C7AoyEH6P+hIeQa3F1mK4VCqJj+PO0ARGvGILP49yNlQqi7AKoZE+chck1J
uf+y5wrrons4B0GB0zTu/a8RvaEn2dqeT3fQu433g4D++IkoinEDBRdItVCMzWLmzh+tQt4FQ8N1
60YKfTPe9mX0i7mWO6FHy03ECJo+Dx7g7oXA9GYP0A/g3RYo2bpMvIUPtG4JnAvbb9tKhrxF39Wl
3MZj/qSKzag11K/XWjFIpnBzqlXR/CDfewxQQMRzbHua16Nk6QJnaoo7QRn/M9LfIHE5I3U28v0B
0GuN1d+qLOsUHArYaPm4ic9JsbK64JCjBbuRA0pCXFDiTqZxoP7yHNyk1J8cfggv5uttTjvqiyCL
adUr3YloS3BeUnnMoymcKoRgoCSBBD91lkH9qGkOf02T2XAlVR352abIj9GF37M/aSX25LD67MXV
zNjPDp7dq2FNTfCUkt5+njo2SHQqT190g6y2CUdPEXTmEokx1y63MosWKnl4/bN8/L29WJwqY+7X
bouHETK07qc/SZV5Tx9V3SA6kMN7rLQ7nQO24LD3Z9NwuZDu7ZnZtcTl1K3xf3HLNalikesvxRLY
tTE51wL9Qt0A54spgALHcHw2t3HFRRimMCUViohLaJiI3wK8VqYZCpNocXrK59nMqJZGaO2yrKvS
+sSYXf+MXbC1lLW5Fl3/EbftC3+qBbq+zPPniY+kiNDNrcTz0ItXN/JQPuqfM9aGXDNdheEgh9uh
YdyOZwbxz378KxUcaTHjDbiOKvXYxsc67E4wbvQRuHFecJK/rCP1eVcudIYBDEjkuC0YABdSCb+0
2a/trwZt6uzc8+QBa6nbBQESoS7/YuAOqs5yj6UK6DuR//f8EBYOval6/v2vOGMX+1QeO6xquWUI
AqJimq21heQ/by2coQYLTpRlLsnI4j3H87zQmfGtoC0afiBrQ5JeXw9y00GRupRmsdi7BHesO90r
ueh8j6X587/DMTBlupug1p/R92/3dAqJ3eAt5Tz6ybWH0eCWK8wDrFoddB7q0f49FUh0dlzx87EQ
tkgSo6NMXozZL2JaxDdl25C24sXRQvoVk7IdFGMiqp34C9vZIg2/V4B3+dVI4UmV85zGIrkUSwoP
QpJrTnCwZ72ko63jvc9cCTuzNEopa0+kdVXvvGto4mWo3W30R1Ui0gHG0ovqMvDkl3HCbqWic0ED
a3jVISruZD0oPWIWruUcYAID7Xma5XjahmsJBFpMOA8NmOGfz4/1BPax4mfcZa6YhjL7CCl9mXOb
LjXQtEUeIrk0WuvoL0ngClPmAvdhRpbDFdxas5pAP5mtsWdh/L0OM0lJniOtXIEgdIyemt/JqEmC
dlOeCHvUyLA7JQtxUgw+1fJH12Q4a9BtB4LNr9GnBQAD5ljPat5mURVasRMHWZKinrtyX5SF3D1c
ZBR1OqRPC5Iihh41vNVcO1ut3nx2qocedmkuz0yt37yuvomJuVM5Z5LcsgsVyy0gPKWTXtXEKO1+
zkN7V5LZiydwkZTsLEB1lMDx9/qk36o8Tyal5oYSLZNVYCy9VHTzE4l5iUcckB8yXyA571MhI69V
BUgHqY2HoGsUiXKMAmFZm2sKGfvihH1/J0W6LAN1btgCjWitlB5fYMk1cO2NaBZQpfeq/V+PVyUF
KUBoULDzuHF5TThYji02zsug3ZdN7r7MMhQh2V1rP6B6nU+I2d5JbRw3eK4lRRnjW7TpoqZaiuUR
E23snv55fjtphHDzZRiWM/AYXUrdGiHspSfQSWXiPtJEVP90zauB3bAbkwTLfE5FPY1XA++wn9ah
EhZwLz2RNWQsLdylnpfS0OwsSa+Jl4w4xnHU+oC95EqE/1t4lcFM1AOSEHHg916rHBdFe7CGSslv
7aVaxnQLV+Wc3nOxQy8LEu+kZKuw1G38m86XTRmxlwY7thOysMicBIYkyoYI6O13ixgkqU5cLhY4
smP0mzFY5Yjy9Q0BuK6i7da88PxOu6zP+LdwhzP/D4P0TKATA0I8qdDxUP2IxD6j5/cb8+bEPdoC
q/DplY5v07/k7OhE1r8n78g9VFYrDYAX0s+omE+I3NfcpQ0lYnQKtQstFseJBIWxawKQdU7xAyJM
JIaHuvoeIujIgD41e49icizLBThIHxTIL39oeAcGhE07wLWl5kE1X/dcBGg8drk7VOsOGtz6UYsK
seScLnwbcyOwzlsEKychjustx4Fv29U7U++0ehFNkPZmpxbsT8kH599StF40futc6bBoTaZ+ceQJ
Y5L/yPpubQu3NSvtagHJ7Ohodoo2Md3F+rjqbSplOxF8nMjm1yOejoKAefrJwhSbTfKVqEGjoyn/
IHYS56Cg10b2a/1N9IAP3UxHbi68Jio6d8jZx4J2GaYuXMktFFYiqk7xXBBUgh4jwNQTR90ROn02
tS50q5YImdHi7Jqxo+uolU/po2JTjzOd1bCK8qHqZXTxgOqNlIvxUA+KbK5615E99P9eKv4qPkUx
alafMQn07Ow4wQBAm/huDaSBF1RuluMQFL4+wnJ8zOmV/SOl4JrhzMeOoCtsHY2dWJ/2OV/jy3fs
Z7lq7nsVaEjW1kQ7vQCfNjp0WTCWWOZfR047ioI0gfNK56e7Mze5xmoi9QrcuLen9RZAx9aIyLVm
dMQnFP3mH608LifX76beGfQU6BstORLuQloyu5jmo5BYsjnIBipOKmLSBeGhZGy6MCgW3crlPfpP
tAZdT/8R8qxBz9e2URkpAb1fvumAnG9dwS5MAk2sacJGi3Dlqo8La0Fw50xSdCS2cmI3e7fOjKMI
pz6UQUHRHjvpbvvFSUqyI3LshxtbhlvDWWCuygSuRG7n35SI1LMihQE0P/mpkJ2HpnxTvSIiDu3z
kE6HqbLBREDJqJsOWd1zEr2RaLCOIftO8WagyApEODS6nFPgekmPozqPAV4KvzcnJiKDdkDFFeWt
9QR4JfCg4b80tlv0oAUtXmWs8VpZt+l4Wrqp+05y59ba7tn/IXDGfogBE5Q0Ka6bWxKKnc8bdfGp
8MNjVOf3oqHQPUjKiNhXfIW9m3Xx7f41oJqu/oOXUkfz3XVenwycvxY9RCECWsEZzMBUAWr6AmWd
bMp0cDewdaoG22ROIEu41iGwmYFnUujtu1B3pAm/6LkbpLSUyhlNdkb21wlU62aqe5QBTpG6oLkh
ZpLtUr7ByBgeEgYps5pXbumv9o4rBT8R6A7oMfdhcKLXabZ00qgYal6dYlkIx9FzH7gUgpufC0M+
9eMPcTnkLv2B3QiupeRnipDncQNkHP4FNCvjAkYIJOTz1U5XW0fNGYzl4UUln5y9iquATgIFofZb
IEChBWCpvlSGVXc1QCG0Vt1Fe7fskCGKRgMlapFKLrXjjBwHw6ID9kR+W/q8R6klqv2GWtx7xKLG
kvC05crh/zbMiulY3x/Ncq/mqj4VN2k6tR4QL+lP8QC9VZVTOQOKcUVhSlaot8nlN54qtdiNfmIp
IIJA0cwfOYhjSesIeUHevgacIo7SYJQWRsw72/S4p1uFGAxA/pNWQ5njSRALDhPoeapX5OCgHMUB
Yt0WNY/rTxp14DG2QVZjyK2qrvKUoJX5pdx8rmZwGdpmwyF/q/Kk+9tSRs/RhVd7b6jvtb7rjThV
x0Q8wwzO6NfwrH5AgsoPAjUDJVSmID/29c9qsgCNxeiW0FTXsIyqlI6cm3RvF50kUBpCul+iIcbs
7Bm3ddpq35MocwB6Vb43k6YCvl0QL/vOmgZVgc9dR77IwAiu1AhdB1LDnQ7Qvdb0Ci+kge71amOK
c98K7q0OoYF70UHMcfw7UEzs/dtFvVnBn6m7cYoT6S6npwBfKiRgnbx2jQQTJOKWwwttlC9eGKX+
Q7UDfICYCv03VvNVaXSu5KbnCgXvRnebwftgL50RU1YdRGtYnGHU6grrGta4CiUN62NE4+0NjM/V
wrB5ug0KsGvrKkOfphp/hpgGI3dh0dOPKBu4DnjeQEDRWVsm/Kn0MDVoLenXwMPGx5gssV+Q1Ns2
t6eC30M0n9niKwPb5nicpQPW0ICmjiRkPFi393KyztjPb1D8gn6uTZF2Kxa1b1gyjb0EQDNVWl1v
Ana3lfB5HLv7QuaOPmjTqelwD1FbDwqrvqZTe/kM2jyPsNLqdquJMID7FmItMncDZejVCOkTwjg0
+KAotN4t1urvrJwzU+CbSNzj8gLTugNYZR+Z+QE4oOjfDdzYK47TWeRbuSj6kk7kW/R19ChJqyKB
zRkwuwNmG7rzrph5Nj677n/H7NaR82uR2o00I9wYfCBzSKhUI8jmSmeaGL+lIH0xRYJX8spSqVt+
58txw6bupviTO/+ntndWwoQvxeED+eco8yTOUKJBYO8xYhCghtdyNoYwup6INylsNUnL/4lWbA1E
E25ZJv0o4lDOZdtYHUU8ZHvwsexk/PCpTru0GTMgBiU9+0ciiUuXRWrSsUYmRvAzjB7Zjp4cNGi/
6gj8S5dPhVgQ7K49VC9+pt9IusQ2abKCfetnPihRjoL0omQGkVibtosMD4tReiA4TctY2MJ2lkAC
BiKTw2nXuFHKh9vSv8xW/BfhyTuaQGZPnyK6U84ImhDXrHSLMa+iWbH/knJ69PJxfNXvZMemEkfh
2axRPDbAVvYga6tNxi5jHeRZ/Ub8WjTwwHs/XMRAHw+3Jo0G2jhYHZMFK0X9QCmU3LARi36FbbgK
GkDKd4n3n4eyKUe7KHjVrvYTf598OwUB6jJPPBbxzP3hRghRYwELFV90uattge0BhhpnL23ftXDr
jlJRk3nqN2I6GCvDXmYDuBgPxSBoPmmhINkbadALXxis7WdVC2kmH26sFVzqt4INWU0oZetWR91m
GyEE8nclgh15fejKeBV3+6kvg6sUeBcqOypm3B+g7kDcGzKEM5D254G++CBMd4vgmEhlvH1/IXIl
p0IWaYM13wnmw/MZolUooxlEhYGJgDzjeQS6h8tp9Y5IRuVU9bfs9XzRh4BeemA+RXLa9F0feomW
OHPWG8qQ8NRyrmSb6vGHs3lB6KHXRdAXQK9zOyz1x0oD07ueRTvZZfQgwmNpewnZEuhh4ZyNs16r
U+bJBCvQm4t6PagIO2uOqhc3RuVzYzxXLUn4j+kUXpXZl7ej1ugF+m/HL2qh9AXJj/CaUiBDdMfl
VeTMERc6/Ed+uVmuPYr8mkC2O1BPlSCREHga1uYqy8cxPHj8940T6RUPCTwQHXEOLnemTIkUxf+0
cOGpZGPvwE4xBwzGyO+qa8Agx/Jt90mxJwc4YIIBALfhfXjx71KP7ASZmiub0LBm2oLgL5EkixW4
G7vnEaxW93+ZzSGfstBgwurauAIJc1i8E247B0tFdyP1ybXDarU8RXLTUcTVnlgExA04ZrgH8eiI
Y4Bl+OnkadKBDGGYQFffTH31NUhDmt9/9HZdPzkDYB8cMn4scOP2OXesgfkjCiwd1C8H3nldPDts
YX42fyNZjj/QTze+4Q+D7JhEj6YLA998URZMrlOY3lnDqOPNlQ7FYkT3G3l2FqNzQ1/yCuUsSwYw
EGQchlhQzDikuPCOd5WG5Z0ii71pn6JewfvEYBworohKVWuSORrIcnmO8SojjI+DV90+3Ce7I0Hu
uyUaeeptyVo/xhuuQFKiHrLI6qQMTIbvcNsX6WuA5Uf4dnepqd3+2u0UL0fkTZUBhRng+rU7NOYF
7oCske58C6zcEGrYPtvMalYJfoUSrQRJ453n6EXs9bQe6qcoRyAq62JDGMovIYKPWf4tmUkRMu9+
Q011drjiV2k0nTodhsNY8QtPNnmWk6FSWPu+iMVLsp+YhZzkf5gZJa53NeTEOj34WonT+yDwXNlj
unPBGVNGD3wXW1WYRjNjZqlLZ+5JEjxNbwKjwzqDtfRxXvNcKBTrq9go8dIb89HABCMY7pMyK9jW
BVa3/SQEIvne+b0UdyyvmMiXFBjsn/pHlB2W7SPUrntr5wCLbslu70TlF9PhQp24ZZ7yFhCLPGfc
qyx3KeqA9fSg1kH5NE2nf8GeHvOfd4CDm097xfIFlcak/WZ9nSCq4z2FWaYbyaOiTZQ/v0gKJ9/z
WAxzHPZgrLYi3WfEtEli2At6peLO4s7sslvlvmtyc8OTVtXvC6CBdzbc0axxFW145eJpR/6DLOt0
WzDYmTtPS/RgJxs7jOTOmttsFxvrbmT7ICeMlKF/z6w98FE6xtQOUYEMQQYJFJ9HDeH/Bd96rRCh
hDkOMRNX3iWVAFZIYTmVpYo1cFjJjaU+1NUyvmmBpB5PYJV7HULjrWMoUGXjN6N0aPki8AUl2Ddn
kwh4rOJ12SEaf5t8yjbtJqCp+yMQTNladCB3ycvUY0f//U8IjZK4STkzIgU7QAzwvovo9edJs1tQ
SOTITatLbv6WCfGcAU6uTH2ShXl/KtqlyiIynuMvCNRru/thMBoNBOZoP0FFCUsaYQfNcxzaHoep
if+UseZBLTNqcoI3lpX0RFJa8GSEZ7zeirnFTjhkH62j9dBGjdh3z6x8pyfoHdEJU9GKyJ1+Remf
gL48Re7Nu2PAUTJ4ASr/XVTwH5dRolFxD3K53F1UESj3/Cw2VT+hXgi0Y2/Bnox6RbaBIYCCps4z
lrnL0SLhWOVeHwakoRJOIYnYJYJYCELKDgjPWoIf/WRkI1PGEGHRkggX6bNypkmCfBDGFda4hKkj
wkK6VN7HKmrcFcnvtGpCMGKn4jgOfYZswJq32g4psdCaxpaXfUK5oxAoI6ZK/+BsYxKQIIIrE/56
AH/n0xm8USBtseqhzxV+oI8u4jjinzGqHCezc5+Bm9X1xOkpC6/HPJXctQXSpBYonRYqL+398eTu
QSgW0X5tb301OR96DEdrNwVZl5qqy++gIq31agJY5f9BIlZ5GXU3c4RkoPphXLd8l95xIJqp8Ik6
c8F9R5BxfRvt+PfF/dk4xrA7I/jaMS5NJsQNal0QueGoreHRXrJeelfJ1rwFm+CqzbuKLfAJTFBH
kH8EiwwOUSdXv/tkn9Hh2mur7npNUJDg5JNKh0qCR9KBZcpdb+tuGPQbXwI/7FX1eTZETTIGzynU
coNwLbWTugQw4RW6FG3DCwZ1eUlFdj4REQlYcNwiIlIQk4Meuq7DNPjkQxSDSdE6poYtnmsvJyNK
qc6Orj4RRz3H3wBTdnIHmoMWFh/x/BFUnbt+pyE/M2YEmPzxEQ5IoOxMMkwdGn8dskNXNNG0VZOl
Z2DfOK2hDQf0HFEaqEzDpFRoO+RzpRSW3/HrMs7/sDKmRWdQqei0ucDHKkLmqY4OJ8r+Go2SwvtA
V+06Q2ItY+X7Xzfg6PX/h7IrPdwCcvXWOy0Fl/kobiV+kcwWdbdt3IzVJgdVEPsvfp3WQJZLJqch
A/3ppMS4shPuAOxdlSqMSJhDlZuKBFjsxbQU3RRTYv2itSFy70uJQz46ZxhgmV5XIN1kkgje53xo
one0vWPl7DRQuIDvOgAnbgS681XQoXIKX92CEyHypyFyRFZ74NgBZ2dtxNS0GqLpf2woFrueWQ6Q
z5e+ypmsL+KyWUAOdXHaG8iJI/U/TykjO3hIodTPRf/cFax1IO0ygJSOsAaBvSEPQFH/vNl9H6eG
CVOxeFoEcy/h1V/Mr5AfHAdi0TxWz/gWkFeH7SNBSeACVE2kbTYUNz8wmYmzVcBy3CEVkuKDRrT4
DgZHk2mv9OYmri3RD07VzrFvZUzqkmMSok8FMMF120j52aFrB68BCyPjXoeQooEiUdR38/7dDq9C
zOR2ZF7jgFWV5ojpr4lZch6Py0DmJusGbw/W+k1L/yozsKEsAXuB1MN8hNRX9yU0MpW5a0i23E06
zw/cmGBh0GkkKmi5ZvxgEJxbguttjX3MDJiRxjxDyKwvqWhN5HVTwlDOYMxud6W35sN5ciKgfUz1
mJwRG9Tzx71xSJaAMFSmmgtSJIZ0wgAfRVTkeF/Q297WSKWbgaDef8nxABsQ7PVRm4i2OYOkXcQd
YLzpLrwcSrTnI5Qe3RJS8qbr/0iljzTNsUTVKpi7kXao4JCsnT1Cu9v7CxcZhoZUaF9xF7texkfY
ATvcXp0tGwWm7Z0ZKUcM1n/J8HEeP/sn7rU6/RD+sYlVypss6/wio2r2duH13u2Oa+fhuQVX925f
S8BiaqIDBvawygwYndnBC6Ri0Alg289IB/gnlVeiq0lSnN3Ubz3TnVPH39Jx0DAtBpVPSvXxy+4L
gcDTRazUXRvS31qkURmMEZt0IsyA5aqS0C2ksV4FMpCLzjTKpcZBaUOeYGja7ZTv2r6D9Ku/LQaG
7SKifBEo2ms/H2o89ptzK2vrpxDmSrM921OnEQ+fnhgaOBpZYbFapCA2MYRo6OKzbS3ENOwogN95
2E6GW1qvjgKwD8/S/n/U63M72lu9lEYV7gQD51LW4Ii7w0//4GH9YuhPMTeHgQQgeNWzjDTTjXZP
zL+OmXbPbVV2JE9q9GSCujc4N0dABEbbPbcT39JLi4yc7YBD25Uf1jg+LC7Uuf8QnsjS1tWLvzth
BE1OUEzFbZrQEUlIXbQcKPrkGc6pPZY04d3bsh4TLyr+93ANs4zmyHASp+wPrPmxYuslyHu25Nqx
qBRzpit4OWQGknO2xkHcvenCPO6icEg4baWlmryy37qRmvEeNDA8xuUS9zOtdQZ4v8c5oLi9jyl9
bhhmw+YKmURcW/4+FGg58+GmM7ZRrZsSocxgNv2Vlr/GojixACtkuvPKV5nJ4c5EIdcTePDs9D8M
jHLExxZm740EqIm4I+pLy44Is6wCoheg/XzUtCtnrWHy/X+9sH743OU7DJLYMSKxbKUKgNpfpcWs
+Qa65fdFEjjVhgxxkAZZ3y2pPj52KKX0JhsGw7GhJZojnkPgmgrUCrZojofVMH0NVAJoF2aV/iTr
18SXVM8YvAAuXjAHz83Kc/whMLz63ZhkEvidzyyrL/6sY6uhdSyZ2tRd2vDLh4BrYINYZM1BGzKD
22mypZo84UG9eKhZn6RDq5gjSjW6sV9kegGzd9AElcIM7oKI+7le5goewQ9rFD3IHoMn3227FlYU
CQGznUw7farpcst8TrI4XX0tn+7Gw59rpaVurk98NMLkenzJko8bRyu5qBzSdHn27sadsMiXr4ef
tNWu6+MNO0qn2fkRBNb3GioHYrL1clAo8xPs7QkRZrLIUYxUdL/AyH6uHrKjHzuUt4C0EjCxUWRn
FF2Dc577cytdujVQsBwcwPa/F9KmaswPudtdJiX0u+u/TW5vHCZEiPa17CKB4Fmh15SRFp/87v9n
1v9XLzRHuijVvm8sxyq43U7+o334P3tJbf6Yy0USi+WONF8kuxgTZmhkj8AJbZBAQKMQuPwq59+3
7wvKEZgDc6PjbO+Dly9Lj3G9nMsMa5BnJmOKugHf0mpPKyqSp7VO78DsIPpTPghxdJ+kAkkAuhie
sDbCYgc+TZzMonojTthWnwHGiLYs+fbcoAJD81KJP5nIouC8nbZNxy7Lmdqg2BBS+IZJJe0UESdV
n124zaOYzb/o60dlRgel4xtWmqKvzfR6ScjItWe80WA2rAQyMMISJNGjfjAZlgPOS2hFQXYppgrO
1/CV69ChmVg1puxgKnbdyRMG+S4lmehV6JgRsKQo/4Fhi4g0WGMboYLfO/pIKg7tfzPKLrKBnqS4
OsLPD1IZmt2SaNaERx/y/B4jCduhzaj34MsDvP0kMSHwRtE855J75o+wM/Wv5TPEfcMqzlQpn5Wx
+lBJGUQJOezBibS0SpzxEDQBrYoDowc9plcJWz6W8l01Idy7u9w2HV8HbmPMDlhaLAUxUUWujtiO
eGUj5OzD/Y1Ud3oJvvz+qgLmhHRSFChsjio+tPEYKpE32gTXh/L27FjsqRvojhXAw7CkVSq2Xizv
/2poc6I8HltSkLqelxlA8KXR0bhz7uHDLykGBjwyTCQIsvU7sTZGhA4wBR9mQNIcw4ykDKqaQ1HN
xNLKfaxz4W21iGGAC3MTKXArky6klN83LZtJPxy2O50Y+D4FlOSR5+OcRPURP5Z8oe0SLcAOi1My
IXPq0lKOGTTTXiKGfj0nDfJE4TJ5XJXws5/SmGLmz+3rUSn4agyGCn5laTtsjQUnGLvuWDc0gRmu
+xJwtBBZIHhs0XxnTxukU66tDnPdwKyy2AEt0aPX9hLWNJoJL1sNYqX9+YHpj5Tcz62Wwalj8FmN
pK01jvilhclU1qPtkKeJWctJqipcoO/Qgj8esAOXHQh8FQ79cTsyJdVNgb0MEy1/H/qfqIQCI2gd
mMAXEvFUj1h62JgMk5zvVYxZklKooRBuIDvD3r1TSJZSvfPMYjqoqp3vcTzn5vr/KneR+cEdrbzc
PNLOU7KJTxI9v9Irr//ZyPaOXN0dWERF9ta+tEVMPIuNFV3tTo4hjOyrJWeGSNcKGELI5BgwND5i
8IVQbhKfWQ5qOkOmU5uWTnG81YytDZ//0eLMzm7DRTLm+5sO67NsL3fSqq/gZCGNOLKTtATZwMzC
MYAvtqsQbiJpqqIZ3UTLkhKKAYC+Mbq+FTMB0Z6ovshU4m95mBhuY1KrgQ6Msn/AUONBaU75GHPF
XZvS5ZD+Ik/4bdkvH8+oWDs7cRLYFJBgvLXoxzsqfCBkNr+FFzi3BQllTslhMx8+VvOvbkOpJaKS
7quNO+EY/EjT6rYLd/STQEFgpvTVjOqz/1YrSbxtYa3WxBXAbyMsbpI9ruabZW1G85TrcG+mptAQ
kPIaOlZNC9sLuHo3nehBV7G/scfsIanyr5tu5X8KHr5iyoo+mB/KrXPXkTXOej3TznxkyNkyEa2k
s5OrXhsElQ30G5yzNwNsZSXTweXQ2l2WH/mKbd0Aqk8/fgyw7Bxso66Vfh8tEtKCRoZoKl1Lam3b
12E5vLgneyZq8khfyLSSq5CKQ8AMr5XseGboOuYwi1+1cqP+uLYJo4M7l3P7/n3+2TUoBBxewDy3
NI+tRMH16kMXpIgSuJIRyN0b/uPhwRbOph5R3LwXrycoEVGdcz3qpT6GTOtcz/uKJoL7zk8Dax5D
+60Oq3QU+ltOQlUII7eOyBm5RuxYqRriqBzRe4WfrK9bMsIaEcIM0PGdNKpRCzP88vQwKX8fCmb4
UdQaLh4PLMTIz4fK64qapBju5UC8z1J4f7Fjb1NfTynGH7zMQXTNUj7rTtnmxTz2w2CNJLJcz4l7
yT8GriGadAdxxzF8tEcDQvvUebb3U5bDKWkY3YlF83yBKaT90VaUd3Y1sQahB9Ft4nTO3o/KvMPO
lMzIues56WfEqY7nq7Go+KocUaBlVuyBsJLu80JGUz83CHbgEAlSUf+KcDS/D4ORcYUYSJNV6+8+
I8tt/3TvyaHifmoypAjWkYUGnRaWCma0tFO1I/DRwudXJTEMOB1HY315PP/J2vyV2YgqQWXOKN7u
bYy5p+Ae+GOmqwYkUFOJJV4Bbo3stoKXA2iHIG5PIsWvIwAawa+sXRweEFhjvjrKUUGtEUCp2GF2
dx3qeaCtjdhFFba41oa8zIvb6z+uKJBDYjXwdGEaeS9xBiv12ka17Y+1mS6yyCtGw/ulhiQuPguP
V6nAAncin6tNuzwZQJRFq9QzpL6Yt1wMXUUt0m57Qm05vAhROzpZ1NJp0FhAr3Izz1fSIPDXrgys
Fd0GcBxAz79ijPjHUx+oP1jPDcGUXGPHDRgGwf+eu3ZKA5d+sEVcvvaxgutzVM1Xzrxvn75sIeex
1JjdUh2t1zbKeGi6YbYCttVxwWVkuFZu7E+0lqUzUu/AyDeJVmTtQlp8f1aJ2SGww5BfbaGMqUmK
NjagzXe53KhCRQkIou+bPuy4vUtKZ7ue3rdD0yLS93T4AuRNPn+v1yP781O1dXthYsohvCU2bJWH
/hlq+GaiQs9C/Gc1r1wUKhxkI6c8B44OKuoY2tkQ8ySWJM6izN4a/B1kgtURQM+EqiCRSjVbk4aO
QIans7Nc2KmRhtCGEU5eJLRTsR9qvFzswIN+pNhF4cMNudAmmXSudXUGS9dxgZzi+Vzw5yKmuIfN
/qmTe9kNa4FWZk+3e064I4nI5Ucg/uHvJ6EIWWQGAc+WAWutLHgyOj04oXyNqCmKYW5GFBezo17j
unXd5aT12KuETmKoK1r3mn571+8s92ZT2bdQtt4B6DId2HbxhZBiKJLQFUTaDK9dP0hnxApzCgvR
eulZ3Ks5y1hccCA6FxeXDlS53BVRZF2zPHcvJTzfoYdnwdEtcV08L6TBaM6VY6aQUTgaBph7quom
7mzupsnHN/YHuGq6Fy16StPf0W6pDj4j3OKcAF8VzwuIVSxtgS0MToJG0N40Bp2OBxCpLr+fwXK4
aLxElMNC5qTzUagY9c8FThLuJaCw/c5RdG6513cRBDg/LNNlyPune9sKb6MDO7IKFD0jxy5sGQrr
oonCylzzfZa1OpK96ctqXqDAciaAzqyjpOiu7E+x0HbMHVUiL+Cb2Wt33k/jxY2okf8dBXDhTF0Y
xCdJWOiUITMRyUOCwKp7n8PGKJEQr1/U03rqjlzf22JDHyYvfK2BozeTBB2WC70QLAmMstBlDJer
R+xKzaE//ETzr4yP3jfzsUA8no8Vw6I5EUdDcdQlXmO+DhI0q/UiX00PPpRd98jwQNMy1dGzxAAP
RDC91fWDwGpkPI0Zs6gOSGRc1cWh1i9suQFzfgD39aA5BLg3evtkycDDj+HNkS4jBlKjdxf5RFwg
EjyEElZA5ICKg5e7HdOKttGFFAbOg0ZzTFDHq0QhxTpez3OB6x4dGwjow1g4J1p0Bd3C7Qk97BxL
tzASsoG3s6f+bDM7jJBfOHVlQVUo3DaAE8bLGHEMTB6VeBA7iWkBWVGVuKgk9q0DFDzK2MNCluqx
7IAtLiKECTyAtVlPHD7cK8ZbcWDN8FEbyCR3AH2rc6GMTVCoOq7cY9cPPuNH3kQCkuvFJwqQLxvx
ccKK/YvqiKWvF06E/DlU/nPtZCo2Yidjclt4Tw/yznhMVivRFlkc4bjD65ahx9QbqdtWi996aVGY
TtAa9bSVoXZV3U10tXgyFSOweCx77JUX/RrU7JAAysPYaP+ifwuR0UEgOL1UUpIv+k3v4I3WtssG
mr/TCWH4oq0+voF1EjbrgZNJlEx/ruA81yxp0bmvJ+TDLy2HlM8m59UhipBSMsZykDpI1e/8RJwa
pmUCuXeevNuJwVOht6nvvWzvp3O6KGgQ1DR9ZzsIDujedvBSOxKV+RDL+BJhGRB0ixpBiYjxFRTL
f4pY7crwXrlYzm3NLRC9pUWQAPCpvIsv88d9sEeLJ8IDbcbp8tKxtseE/ZnEBf2D2bRetlX5furV
gdlT7ZggraotNGhK8sRqBrHihFygx4/W0Yp+y8QmAA4kqPaWcn5Oo8J8kgTvTdDxk6uwoq1ECfn7
Gr5LNFpVCaK4rVNWdcIYuPh9jYGVwB/2IX1or6ruX8s9zJL9pYVPi/Pz5H47YNj35hi5Reju9AlU
sc05A7MzqRuiIqH3xvdzabb7y3H4n6rLSHqOKf/vsW3Tll5F9aH4tgxzUXlSKyEPxKDYqMyQ7XKh
lX4VQeZ6BPiumksCQF1UknMFSm1CqHj75M7WP0z9F4faMMTyghYnQrm+yHQgjfgGubfAWO2HDHWD
yFks81C2yHk2wv7pY5kWxezGTIZoRM7T4c0AlAciBS2jpSirv5gcFpVem71bPBBVFtGMD0a80uZa
p8iCvNQFSfKRAGV+hDgg/JcpKajZ0CLI/0Y23DL9vhcHzaoilfJuOmCyTA7faXqFivdnANJk+pg0
DttuYxOiQvyCF9XSr4jvD6vsJgjt7XGzGR1vhBxSdodWDgLWtrLAB0H7J5P21i/NW6ZApmDZW3Zn
OfSqYhvaeOQFjRi8T4jEoZUpx32QZt9hGDgUw05gRveFborZn66pYdLmoeke4mMtf5vduk80QwN2
ZbbN6N0Yr4UIW6lN/zApdR+GMhwZTLbrccoWVZCRQu5qPgf280zPSiQtgfsY1yukseLtyGIg9+H9
E4efdLVy211SPlQ5qkAzHix4oMHtviXhsC5wDRd8wXFh9xiv+4ZSLWyMoB5ELYfsvJgwjNpp2gT+
yB8RrPq9izgoDb9X1e+ZwrGT1L8COE2l9u5nEr4ETDo2a//D3Th6G2j2m1DJe4vPBQ4HPD++x4S/
RxB7a+NaDetzTrQ4WLgq4TGNp32OZ8dec+2S/hHrY+6/mjtxU5f8RCdIE/4pjNjlsiXGEXZS/JS/
yMRut/71Iua1I3XK+dna7HXDct2AEiSQ5f8oj5YFrdZq/CGowOmW4HKhwt9xWPRF6cNOcFLiwbKb
LJ31miOgYsSOLJ/rxupult6PP8ZXr5D3GSmbJugiMXNptzU+MbpW6vGHG+0FMXPYsXbbilkeoqJz
GO11C1OBIbf4/ouKnp3E0Wz5ErKV/juB3WDfCFFcBJbB32b+qJsWATgfOUCAiC04QhD7BtegToFN
K0BRyVHOnGvTfPu2SRGHk3y57E+K8hR3DU7/1wRwIMZfKwMHiKPdgI1M+ydOyEjmrs5hU7HHx0FO
FYsry6ogrcomw7cjkRopRAAUf9A2mYk9xVcC4y1eVESHU4xUgl/a0rTYQU1hVm5PNSmJUn0X9e+1
8Cuy+AftTtP35oRyOamnvw1pX4YxYXwMLv8ZgA74JaxUZjtNCGykleMSjgs82evL/NCXgURh9tsW
2cO4K19FUUCbU0cUtwp7mu6RacJOeen1FhAfy3InE263ew9Q1TRjbnnT0C2WMnlwIGdSsTvhNR3b
5R7K/TFThlA/z+6cj2ary/i6xbQq6J2bmTAulO4x4Qy5mBoIt835IleYsX/guyClw44yVDzvsdYX
5MbLywAXIz/ibM34ZhyFCG59ul8cvgTag1Baz/De6b717CWclK5ise6B79HlH3P46Q5EJTsjs95J
AYSPHUPPrg9MPArzyyOO7DOWfHsf5AG9GtCvddtLFXooqZWnazrPIJfZzWkO45Xr6/9dEd8ov4ow
+z5fkjUYsA4tHpzd/dfFT1+26LgQRgNvP2C7VuAABAtftARuYHApFxw94Tw+K1EnCPfE3IpFORzs
1gOusBJKC0c8Z1OKFNCKvtuqXJmvKFzIk2Gg8wA9EoOOqqP+IZ0PI04mwUW9aM6MfXmk/vlQt+L1
M49gnoYV9axnacAqA+xX8m0RUmUj1+z+q/tieXs9VA+oIx+/6/Ahs6ajhnJighGC3wkB+LxpaRF4
94T5p8HwoVP7IoSfhPo+Se1LJmZp/2KyM3tHoUpeZZr+MtZBEUHaxJaTxArfhx1E0Uar+rkIVMqR
bfqox7xuJVAm2B8rk7t0iOOYF0MhCtNtUkUraAQTC047RCEi+wKbmnXBVA+Cu41sgZTGOuHDIIX6
hFJxg9SBamgOBddqKtftghTnaWyL0t7OA/FxVBflM869c6q18GdvKQX0K34CA91UL1OQRMoUMCdq
OwvoxzOSKQ+MvggLjVkowze8xsK08rlNd0TP0aW816F3o45J7A/vYBoPBwvDdNqmJf6yd0fjn7SL
Y7Ux8BRrSCi9mOz5iNk9nx8KUsX6Rpxb28xLU3mPEpN+k/jJEgsEWtAjDPQtFWJYiNSuUIeQSfVQ
EJ+KHcgFkaJkzE9UFD+HN1Qmiux1HZo9fzT6Erk9g9PtsysNgWWJnRVIUBwDdq4BFzU8F9jphzMT
4Nes0j3ssKbX3p0YO3Q5IULj0vrXkFq6/osfG5pAXkgi502RfI5hVSAc6nwO11PUglpgFLWBkmOd
5FWi9UbgHkmai9ILKslFs+cGN5PI9wbWmgUaw9xqknyJ+EihczgYbn3GzyZJ2wROIw4inmvaZ+Nk
7//Qf+7yvqi46MWfImp/PjuxLsWFyBhjacCj9nmXulim3TDcX0wwhXhzxDW2sXVvRMv60fW5WJ4a
zl5WQy581IoJx+Kkbw1934+jVovUJWr/TvXw54NeTkAYPvQriiOyBpUIvk8iweK7jpJ/THNFw4or
a+b9lm8jQaq2lsWTs9HOCGhtdXcvTJgv+7hoqy9uHOTMDu+4CZQmDBSq2zdf+HAq4geriVLLkJUv
rCyiVtgO17R3R7Arh1DnOR0pqTGigoaDEPU/qhjc1GnGjT/8MJLwxpn2md7omV9t9YT2JzW/7Hgd
obPU/t6lqN8k4JAOo9fo55PV7+nbqI/4+lYPI3JKAFqBHNdmcwrVXa/UA+BArqt3iUvV/xzBJs2l
1aZmi4x1IPhet6WGtfCvmasM09dTxEojHhX85IfmyDFwReEMveh5o3pCX54YnDVkZyiRfuSCq7O2
DIBByiQ0pe4g54TXzY3osLRL+tH6M6v4LxjqCYipPUyZbhcJsKu8ThmO44J+yxVj0M11/lx7e1l/
DOol5ICz66Y1392lz/8qGTuSbfbF8ExYw4Cm96l6If6GveJ0OnJgPeKvy71tsDcuyQBRP6+/zx/T
G1Y2VdxpgdgKHjeAvJ645bI47Hq4vgq8MFTP2xBlISPQvfHjROkkQutG1NHMFDohi0fRakPboJ1H
FOV4tRh2RQCqZP0fl1in0T+emJATWs9wzoAv5cnXe2POl1vUhoNzVku7m2MdiILvOy4ICgi38Qb5
agkPgjBoqmM+Kio1kluepT+clEOQhhAnosjv/8RFwFnmCp0A6tk5/wYF4RkBuslpnzgLaIUnmAEf
yudF5QSc+FweUJE0JGTj4Rp995yvbJcEl12NPrWx75x7aSt9Eg9GTkBRfLkPGHl6g7TrZnbeQWvE
xAAaz1Skfv6owz8jqsaCpILf34DEXGxY0TEyZxiQBPhtrNCyxZqFbqhExzfwmJOkrW7LgS3FqM/0
8OjQA5ue1qKpnBHAGu6vyRVq0PbKmVyrMtektzokNY4K8jyQzM5CRL6L/MZ/aosX+RorYLbDz0eP
Gya/ftOGITvf7t31EDjr/Py13+o3eFen+VuXDJIfTLMz2hsbzmrrxapnaCJK9V1053lAC+JZri5N
MmMBxnj2VCiPpXQmHNB2aDb4ttcxZkX3xUynqR95pPV4DW4XPVtpob/YFFBG8lrb9nIZTfnwXPOg
IbIR8RzOZz2R7aHJwmCB1G1vmiP8QP7sx44t1j1J5gbGxcHA7UbkYzFy1ypYwKUPs2RKJ7y/ip/a
YJO9gUfW3CtgtzkaGC8trtP4Nz726pvV2TWERB7xPhfue2S7vaP+wbMhQugC8La/iJDjmG3BY1qo
x1TFc0DK/a42n+pk+PP/fUvEuKAehLC0TBANzWi+l6LfU9Vx25Y0+R/uq+CRT9QnuQWsJQveOmTf
ybnGYWzElZ+ijFDGtg+o08U7XKYfZWdh7P3KckRHsx0SXN/clkXzrm94vJGepcLCBs/ao3+cstj7
hOjE73Ccgqw7QmaEC6El/VvySSr85XJfWfhMaeb5a55uQ5290JvQav8EydKkaZn6FzucID1VfHU5
epRlpyjLNwvo3WnjOGttvfDj5ax9IivvofqtW7sl20TKUtYB2ieO3XhOadFlFUjyXV4cdem+SigR
g1fhj5sZwjYEpJFB+bnCb37NQv39JsM62xdp10qdNLOXEgpPv/zSSkGUzDaxZPk0hoS9YeGnUeS8
blJR9pC/RuTkqmf9F+DBjvfx1EdOfYFm0JdF7kPbC7OejyZr4onqkLLv+exwCujXeiMJk6NDJJFq
RCjvL405rsmujmgsG8FQC4BA/d4mkKWEbQZmJvXY6vSele8MWBOkkbC24OjdyEhXXX02H4J/SW7e
75rBzUGBdaeWf0zCTSIJ3775tFgG/8QOUIHowY29vz7Itfy50JCtk/kID7iufqFPZ/pmoUlnKCca
P8fp9/DhXojOQGL6xR9TE8LIZ5r/BUGz5RNDOptfDSCqemKL7Uwn3OAho/vzAsiTh3PuSYbYqqJl
crKLUbvLk5fHTBXXOzWdVsNIVke2H/4RaNdKV/OuC5029muAgaUGosc6luwySgbpy+bwPhfkH5sf
cNCsnhaY5Z2WtDfA16FqCJaO+64myxIs8vuPc98kNrj8+S+IeU9efV2ldk4J6bi08af+qgOCPsHK
RoDpPdiPj3nUAu/qqkOueWx99U7c1o5Io/CbfbFpOWerqD1a2HwAEHMxGeA8baz2CY568yByqsdY
CKtWOKjWkS8nXXq3vI7QTxQCNsCdETm4JZwRDSuBV9IioDBpB42gN98adg1NRobs0z4uULzL4VQ6
iEpuyzcNuz/ToamO8hPa3qNZTa/5t3sQOlElNw3qLPq2/yW/gVF6TpxizoZzuglmydHVkYSzdEoG
Dyi2mLGsHWFdRC6JhXKS3FIrniZtxLrYp8E7QS/rB7c1QzQJ6F4zANRAF9EIAlm9fAk/U8hgC+fl
AS+rC/RlDda8OFNuWVTWibdfHnsWlfkKxudSTIx8L9FMgeTb0CpEBdSLgAzM6fk6rTWiUtaHjte7
TV8UPDATnAINT62or0Iul0cb05srblRzUl+Om/vCGrFLweQt+vHHYh9c0Vj+JBzM1oxMDhN5G/A0
+a67qihClADZcmYXS4i8py5s7OfACcSzZlVjC2EqrifKOcWlwsRzhhg6C2ZqnOV+fiLTyTPfWrNz
EJVFvQ5TRcqgdxt6wyo5nRgWPyGQUEvbCGatYCO574Lm9XWJs8In+rJngniu0jLsAswnEciFGGoD
q/LTyvmBYx9DoCyZThCm1AXFx7VhRIbxaQ5ShGeeJ+32jolxXHXHbdHbYTg4DCvbHr0u53E6nrWu
d1Ykma+2w5U/D6Lv7QcH+W3t6LooAlqlcQGdcYZWxpacNgkHiWR3prebc1s++vsaMsVmEWXeeNY7
liwwl/+Y/u6B6K0RSrA3mVu1RstW5bxfoAQc4z5jg4C8Lmdx8Xn1iIho8XiWtt2Tuv+RidbZ02LK
DPbp9axTvMJLB2ZZue0bLjFkpPnPpqSd1Uou0on7vgYPtWuMkbNokSgZ48B8Dw8jpdYcngjJaj8O
rwMUG/b5ADEiEg8pPUg+RoDv9Isg1Ddum7U2rolA34CGRUUyVc/ot+rgl4zivArJoV/Oud3bSGBL
BbZCj8+rtM0Tu0NDJn//wmSddVES3S/rIkdG4UZpLHIsJmuU9qD6OoLCTecq0eNlaFwltKbRbOKk
WZa0W7ir0unN3Gxp5uZ5dqd2NBKup2xdxHKMuuKRIDe+PykOaerOhwqP9gXdb7xxuYWfntAnidLU
EnVN4D/ngIWuV+hzr/Aa4XuylMPNyKO/HY17+AuYzp+IKzuAq//ZmBfIczAcC8JcUyS34cXzfXVh
zqX5ZOaWjs9RelaLQofHwFBPnNj5SW8+chasskXy5z3V4iwxl/9IDvBtyCUM1FVXBy6SXzd2WSX7
5FruS20f4FzmTbl8rEWccT1tuIuE8RiLNgldlJsG9X0YEIzOcdtXavy4tPUY4yHP1RMjAlf6o8jv
eqPSiMsCirNIaiql+qH+3Ff6d/gGckp5rdyCwB4bpCooY40AkOYsyGkA58Ghe98JcnUnSZtApeW8
i+Vyd+WUUHUZnS93yMYjrulgWCjG+oDEqnD/O1VQvOO0Qg+11U66uPfvC+ETOXfcdP/kv1TTl/8W
gI2Fe/qfut8lEnCkva8lwQQXH3KTwsr+8Jne30ayorE6duSQHM1QMQbTMmKUpS9UEiUY1AW7yWIK
QlDwg9Q372xkmOynWAzHNrjT9uEW4U2tOleqYTRH80HhWZcF55hrB0nbYwz09/vLT0xL2CFQwGLM
QTSGD5rDiQJFD4Yz1yeWaBNL9demJzM+RZYfqG3Fxdhb6n0U49J1WGHY89Rk+5gFQnpoFtkGIbMV
5hE0x7paBtYVw5xNNX+iY/ORRgYHCkJs/WG74GkaGKVlI8rVt3Uo5Jl6y7THJvRm5qAmtmq685ub
kKOEuzmvbsHJDnRGa3JZufNbVTVYQhf/zsXfGKxtmwz19LOn7di7ZrliAtDsW3DVw3nqtAvrvBo6
Z1vNTK2xYC5EWLe3CgG+7b5fmvBcEp7vxFE0XaHuEZMUHBYPZTN9qJ1IDEFAcvvdygnJd0QDOMeF
Ka7eNHZ8BPhzBrNyy8dh+tJ22Z8HkYkauLM7xLmaFQga5Zzhv0VpxodLjQdvfXbOTwBxlZ5/ReSD
RFlTIQ3RLBb8zqfFeYLyWoAGUQXoY2OLAHHfZPCaUudDcQJ/tQnVC+y8iGzLocHVG/dWc0r7qBI0
+euaN1FRMs4cxi03dSTgfi+DaYl0s58vbFtqdzGOS2nT4q1aWesCPr/cYmA69aDe4UwCrS9in2sV
NtXjbgwflDhmVInHPauTsejtM0iVGMKpCbwed/9hbLQT8GNA70gydIRD2sGAPZqANpb+TJo2DUVA
PSrB03yyxQXtryr4Oz+LHr3D7jeqbTadHUo9nuNyyr5A8O+byLMhR3YvzRyNrCHhbRAe8PrgP0iq
UM3HgpBGXmJKmA2fdZg/qOW5fL/W9c5xV/43xqZbidrkHI9HVaxyaotw4sF9S/S5mBXOnQ1xR1Ct
y4DvefEm9+2Nz3CFFkFnbvV409/2vCuZp+QcJKIyEs4YFE2HtYoNLmjDGNscPFo5oDRxHwaAzm0X
uoH6fHkVsYqgHwF7Q/xLQiSajUT7NAM6FGvl8mZ/w14kbZV5gKq81mX0cDvlcG4Nsv9fDH0C5G65
IrUmefaAzoV0Hul78k/cyJswH/0U8L0oM2AddbqHwm86uq6fVHd9nQ08pthLwRs18clL1n1S8zh5
oRjeZB41mVtQ13sR+3gGGoljZG6NCMprxaqewqoQw7/ble4lSb5r/whxD2dBQfSQKlyLfwKSpaLq
R2iXLrtr/T82gGy2nD90G618d6s+xGd9OFgg9c57a26EotpRCAFn9/rJ4hAm6zDG+zzqOdFTjHIL
/mD2AcienvNckZVw83CQwMWaV4L3IU7wNFwYTg9+ZHSvwquhJcjUoBEVAmmoYgzsFGx2zyDZydPV
lIWqq9HPtVIf4UXZjBcFg3KCayO7FIoqxQYWuj/vxGDEXIemvwgr2KIXMtNf3ujyC1Y0xZVnXd+X
GqOAjW8NuJIK3B62U/d5DDtp586qv/C5aq5LvXaoPAf8wQC1rqX6ixElqBx+q0hn6lISOyXjmu39
pklW/SwjLcbe/w22J8bDah6Z6bzPqQPfKJjgop/IoUr18XUbB2P00IPW1aCr9AOCmc9ZSo8wRoXb
GLzwy4DkgZExRYa4jx6kXKuO65Ht9UcEh/ONweCl+fSi3ZQE014CwmWGzuc7DyB6Un4D95cm6llp
7DHmTvjco17xktJiCMvRsIIt8bMCZbU6xOUyMR3LLcHls+xUM/l0HE763qJcSREdTfgdabpQRxyk
1WN1MCli8vZ94fV7+2vmZlsr+x7qR3JiqLD8skbR2ynQWXu3bN4Tuixh65KTjtNLCUs4yXdd/Fw/
s1tU/pHAWY/AbKwguE3CRGH2APyu6+OXkpgHSHNYIMku0a5mc7qvnlEO+vZN6OK9mM0iX8ARS3ri
a+YVhJWRcSFIaKL0J+hB/fc0yl9hmMB/Heq4zlsAuZK6nxf0pl0rNHyyOWKtvjQRqbOy4dxhmsxh
cEvz2qIrD+yw25l5U3iOBVfjJQpuAV/iXDRx6dU1MrfAgXp2I2dBE8Vo+qAEXThzHwjplOdiSYOw
VUoKfoMDQhhe/+4RQ5zs8VRANfTTZebCMXT44aCk7tF/CD25DwP+U9UMSi+yJaStSms/4m+Q9CPt
z66j2WF93SMElp7YvVlXWlO+mW0S/CMo/cgpyNkyymDPNryf/Hl0tNv7ohownjW0Jbq78+CHPFMW
+wLp5mR0jWWTwgWXCclfa7RosVvx/ZX04RAX9CzMKpbnKZnzUQlGh4W+Zk6xH+QvXqx+w+j//4Qy
7An6bhWBg+i0530YQh1b+jaLcOdJmVDlEFtflEKSTiRuZJQatT8zvcrrEnDcunR5DbacTBiBOnF4
9CTcxPzXEO0ktYcejuJxgDuhufj78l0AZ1nnQ/PNgg5PgS8mJ2wPYYPZJi4XKWbX417MI7AsE89M
6qOH4JWYYDtcY/zdTkkVn3tKc0Z2uZ2okwSEG2Ej9vD5PMGaM9Ffg4+ewGpRfDqdpr5RbOxcoZbS
sWjyWJKizX18hTjh9Iz2K/jt9HkyJflUFDN+shv34OYm+1SbjlTGyJacJwbEK+jUbKTwvdUHDnTX
LYvCre7pyPq38yWunKMXEJYfBVbbbkyOyf8fqMFD9B7gY8RGX5Z3BzuQC/YpS/GsK1UlgG820RSQ
1XbjIakoSHvS4PD6AMObUNaMyfohKnxGk6Jq0A6zTvYwkKSILtH+UCh1Nnf8HTaB0zUpD5BmwmMi
t8VIX16HHrtiAaqWqupO/K0qyIH1jVd8c0wMfW1hdb1uNhAYhqEUoEoFR7fCn4V4+8CxbVwMy4jm
zBQ83HgO/ynRD8hCT6uH+H2sfcXll7V3Z6nykQQ+WZDsqG3Y+EoGLkqjFysr8InJlvh3ia/1RrD/
5HxtWVznxThgXyXTEhkn/1UlmgqAdKLOzAjWu6+ubwV3EgPepryohXQUPDG9iEaDyJyzyyKN2/PK
zXTaAMfJzcqbltLKOw9THd+52heRk5IMYlTtX2v+LyGSg/V7n6b3UPhHMHqnp1XUX8WchjWBqknq
KAr73bZqCyZRUX+MD1HRXPz7IDBxczRPuvIgGGJYc5Zb9tYhK4pcJITxy95Fet7r7IN8ZCdz4/Vq
/fPtWJwAubsFstng7A8oI/NsT+HaiEjXNufKUw/69T4I6+6zn51dlqDKMSwwEgasyDBeX0tnzLPk
qIEiFi2vYaC2DnNwx4c5oci+dFaWZq3gs+GHbnU8xoouPbcsbYW1Njfj7E7+invH0jTv4dny/fyY
ZbjxLMKw5oEA/a+iNXKzClqTYzqcLT4W8sTcsFl+8HF7NdtAJ2NJhoEMcd5BaDNTYx7xvywTaz9M
NDpyS1xqufNBym6dHPxCUGf4be+gzYLI+SZwLfgULI9lwEdBpdhUs8vs9RUNf06bxYTwg2YumEXU
yU36MRX6iAhRp096/BE70m37vKRUXDmsntDKPS1/s/dsHgeNCUhyjeuojoHJaY/SI48ae1Fs0Z/N
fzkJSCvArQhBQZPaA9EkIY5it4lO/Q1FBcDQwo3cUTtlRJ5ls8G6fQgaEsKnt2U1TdPKge7JjlkZ
0avaisDjLZC1FjrFrqS/Qa4Jv6LF61B5ZKdMbEDerMBel3SF0OA8UhQBw47C/n5u5sytgLACqJPb
6qhQLn9QTS30hswh5W0ldhFCmj+huuy9uc8oUq2FTXBHtiQPH7RumG/bkGZN1GtLr2feMbicm3Ru
KAAYxrlfJu/CoiiNH/83TEvJruQusKqgSendrBnIu/aWhFhb/YgriPHiWuoeoi69as1iov5L2s9V
ln7FiTqHQhUR14CSLi//J8l1wtKI+Ocqh3moijrpbgQhxFxxDdOJY1fjS9yshOjXAOf9gmtUUyFQ
5cRJVJWIP4a7ep4YuCac9QufCYkDmxf/uO4irSXtP38Cr1lBKrdQlPsAvJs+W+VWE6LMFDofjYE+
y9abf6wN2MbJ8fGgZdG3tIIuolLNRyQL3Q0047Hux0vOWFBuop8uqm6p5DF99dsQhgPTyVI0vFzW
LsC+/EozrRzjQwFbEsA9ir2ErNHnMh7ZhGKdT44EGVzLwkAcxr/80m2+MEieXru1/2hcFxrq285m
jK1kSThXltMpLUSQ7EkKo07KweEHaVNb2gJzWJ6dulXm+HPGum+ovok/Q4Cx1BvCkLK2HHnLbETN
SzXlQctfdKavT8Fig5+hakvjg8dXoufJR0PFVZe/kaXaW0KaopNFiPNtPJ8QwBcRAcwF7CIDYhvy
tqzYP6bCwHOP6OMxeITuQ3WNbX4TIHNJGLizWlw0w/tWNA3kwjQ2qZh9t6TEhhpoyevcUR9q7QTM
zJjT9pISOxurVCGVGT8IHI2Xeswcu/FXd+ap3IT08F5VaRIMB/d91PxiCcYCNsNSdfYeqKKkl3wU
ApRcbtzLQmAsO8itOw+Ie3UIpGZlj/TCe6HKjDwx4IgUPXO5CVL+YHlNk/rS7h8vMls9j/pFlpCS
DyyEYXZ5kYg4U0meLR2p8Uty+oDgwFx7AAZ0HMfFcYU8hq5D1m6ZnK3nGKhEplBSyhWO4Tef9Jo+
gSoXKHPOFtU1FQGZhTw1XhlA669h7DNlIyEvcFGK8Qv+amLs1LzuBBHDcBKbb3KqIeIIK3tpXLWJ
XKSwQ5BHJH4bF896WdD1T0ZhOz7YtKwuu5gzwKQi4Oar8sLUPLZNLgha/l+NrOzMiW7TjJWbMflz
zHkY8lRr+8bcXl/zr/HbelQNxP9eJ0d3UScVxOTivis52/6yFs8EG8jwpqHg9jE/m6tP+hCVj6r1
AY0ESjnFdHfi0I189CZZYV3+W55eEvQSxok25dHhi1+BDCoTo6GJi+vvHW+2OojJhdyJOrPdgo9u
K92l3/FHz+C7/5EsjTE3Mo/HAZ1M3m6cZKT2ASku2xqPxmjXavMSpep3DA2h2HQc9GHy4dUiBQTr
FFYms8ec84BFG2DlCv92kx3foXg4+Fka2bKckx048W3gqHQMcmLujhbat3hgFqa6TWVwtj56ZFrj
inu9UaNDRYCk6cMYZe3Y7CrTfbrL7JD25N//Z/6KkrPrLvzWPamyEDeW+J9G8UaVGAZwPdxF0geH
YhIEwfopMufeqlSks3UWV9s3g3o7Waqdg+1He7sPZcHpIxknw2V9qUt3nrMm9ZjJFoGuRGFtTeU1
12IZZElziIGHzoxlY+OwAdfLWKd5FG0R3qPtrzeHcDo1sUnNkJLMmjJ/GYAY1g/QzonqdISKGSgc
PzMktRFDhU3EfNGMo8pBk41cNHvAJRRp/bZnxE2wXr+fr2I0nRiYc8OCXPfwoS5VemqUAATuvWqn
uQlEYC2KAx7rOX3NpLum/7+zyOjs6WeOwdx0OXgvGJ215j+Y3XHUzKw6AetiXjqTXLEdMIgRFY2j
btah0DOqYcaLFEPbJW164iHBF24hU29+/20ejmPL8jQqoBifdvQFEbJjKpk4b7ERyVc63BR/uFpQ
gAu/OPw1EL7NjtAwy7smTCxe2Axif0Mpmb6Kz0KJL0VuPcKzPO42U6O5HTewsJuNcp0P3UeOK3SF
cwle2qlBQctRyvII7R+z9gldcBr5yfzCjTmrfP6ugf1oh/JCYsJ8KyCXv6fdgOFXpBQKN+j85/OB
Qld4ybDgrPdScXV7EzLsabxcwTzIXWsT0Pej0GB01HJQn0s/fpI7Cf+49fWPKdLM0jIbkT7sq5gQ
/JVY/rqVwujjS9U2UzeK0K3ATycGDJLVK5qh946hYPflObitdEEf2zCnHYm7hjkiJRIszZYAAcU2
7Oltb0onRHb8N6NfoqqrKnATklpFiUzuV9Up4nuwpkfRpxe6gRye85ympHOWIK0QbsD80uhd/6qP
djgE7fujAu+UmD5rdG129CMhAvwtGMyl/gklepHscsKBT5ByBRq83U/7ycrqO4JoRUfZsP5RV2dh
b4JtYWOwGdymmwPUJhekHSO+nDDLW//FUBBG3aVL48BtKftYXTWOtpjECysLnIi0IL6ZSL1eb6EI
8x6HEqTMhbs/Ob6sjvLTDgq18zpnnbsOL3OWTa79vZA1H3RHiht1luwEsxEuSYIISO6a56XWWuNT
SqoDyiVGDzTnPHPUAdO8ndUdjOM8+TyB3t1X9J5WRZhxRxaSUMZSqNsc6SEOoEqHuSEOsiKm2KI0
yLcR8wriSAWR3r70H1Gdu7lTiP9blxDZE3tCiaEdy4ltmUXIRGXW9FEcrp/+ykHfwlJwOOm7gEQ0
5I3nyHE/4ISwja4aD71TiJecKbRIg/4qPsAPxra4J04klF85ZXialn4+O10hpqZ1vZmgViTArGpu
USamOxbYUMZipbsNuZxaDW+VAnPNQ6xq2f0wZ7asAdaXTopgVLP/t9ogfJohWtAV1yLp9R2XQOzC
nPhvMxFLxcSUqRdD3Dx+ymtqBygjgNTgTBGnevaLqaI6+WOosPcJNNMJYhk6GqmEXEVftymxX5jD
mTP9vvW5+Raonlkr8XHO4jU8YBf2tzVouvlPVxOV90r6o5T1Xs8Agr3HhXj1PHpQ6gJ0A49w30KQ
P03k7MhYFVHu/fTELFvo1+0DMedCUi0udTzh15IXSisExwlKE/C5ZzKFp17AinhDqbdi5BoLzl3i
TBJtNhABkF+1WhQFmpHQrAeT0W/HxzWcFyR4yxR14B6IYjQM+RYBmv3JGQtTdtPj0xQkzLoMMm8x
p4Yut2Zz/mQHaaPm4kGIxlT+QOUgX1wElZX3m+zy//AD9iZwG+0LTv7on0STSg7sRoImQINEhqP6
KaqFPb56YuguU6XTyIPynBNGoGIlSb91Ued27HeRFUaAgNqOOYnwEvA0mgZ3CkRcpiVCKpHoWRo1
gLKPVN6s1rT3Gs+ywOMvJDbEJXUyAgsx+ZVaGvPnJx81dHFRuGlvKhJ31GD+WYBQ/C4+hOmTk6F/
a7dVXuQGfJo3klwnA/DweNvjAqh+/TJcvMl/Sy5sRtqlEJYwSa84ktQhY065m9ophKebwy9sMLpg
CmG0f5TwNMIwPtkZtDbfoRGiXjtRLRDsgxFL3Wf70boAInoFVNBUGgY7uv93lPPACZIZAxb4ByCr
aQ2cRWcLIOThZGGwhUQ8M3yxHNfiYSXwcBt7rh81GMs3KbS3LQXbs+f3h9HYqC6GM0qjIlCX2L0I
qzDmTcifWKl0gc7kbhePy4gcQRYfmMumVk/bsMZWKOyA7gV3OT9J+c1Iv9KDhbW8mbqDadzKYolF
XRvFzz3FL7hdOhO8JG+e+avw4Il8xhisWyKqE3w2sELM5vhMb7MdG/pNK75X14o9zWw7mEKlB7B/
RoNI+6SC2qEQSJrG9ooeWeuu/USZ+6NMbBCqYu+Qx8+PDaSxOnViMmEvW+/38mGHE7J1l+UgZnd1
jEK1bViIydKfkllKyrUTGue2rLHAjkkua7HGN09+4Q0ffGulHgDQLlFvIqyDwNzb3Rnk/YFi3ksi
KfqAa2dy64XoZZyBE9/x/dEwvlBN1GhNyTph1skNT29Mvvgp+pmpDRyy24YMaHB7yFoH7IzZL+BK
nfCRFh8w1ZSUysJsv7vYF/44zHFvj4mbfCoSM+bKXcp3pfoY3oNsU3FPpGFa3HeGaxWMQeGnQ+Dr
qUKW1AbRY7UbPtNgarUidA6o50kWjG+yUFaCCBidD3V4OWxJHPRrgxaFsNzYVLLqUK7x8/wRQm9J
SL7oUiSBTy0X7JrpRjtRf8DaidXDN+nFv8+q3pjQx/g3f5bnC5WV5JL+sd2hucs6nInzjGh5OYYK
SsoW7KRtq5vhDcIJp9KO7uhHI1OqRMlo11CGKtQQIyOo/5Dw/+2nVNQY11xWzS9YjK+qjMna+m7l
jd+KIgZ7jJLVtYWVrebLq45a6lBDkbJElnhEgbNGS2c5MKVbA3GbJylZ5qI3U/juZ/xDsYMKbxnk
eJM6vC5brB+nM9ZH+yEBdsITCfWk5kpBI2mu7eEF11JihTYxMwhkIoKqCw5X44T8QBsNcF0duTFX
7n9F4MJ1qp9JDgKopTPhNxjyiWA/jZC/nQwkz/Td/LkXCrCvbypXUpTeyS/tCnNaUthRcJodDsdY
Jw5MmwAt1Jvz9793/THg0EBr6uGvjkqchTBKcwbBX3bVVGvKOVJGmRNSK57IAxl8Iwv0gM9Q0O6I
M6CMQCHUNzJ+/gnRnwF+mmgXM2yA4myNQlxPpOHxbWd5iBWEZtTyULJJblpE8wWFc768NDewTlXe
3VC40L/VWsyyo9jXYWNbMn6JSXo2vytIZNZoiZaN5ERSXIpi81OSLO/NWvzcKCETaNq28cP9PyV2
8gTBz6LXbeNPRq8McDxtjG6KJKkU+Q+/7T5xrl1Th3hz6h76dWvwW8ZYJaa02Ie5jEflwMCpRo+9
pjGM8JczhDMsvvO7dpROlGE7GvL4fcAeNAOD6Rxr5SNPsRhamNHbQSX0o6BcjXm43g8ziAF/xZ9/
k0AJkfj+HmQa/bL/jIp2wNqtMLr2q5eD3/eRZ4IlEk59+ZjGbs4t9xXygiN1GqAyCa5mkUz0eEI0
fCcb5oWVYXeDIU0w1Uba5GDng5NNZKiwQyK91PTmwjiGWttpyplk1Z+1ac+W+F39ZBwfnTcPhTVZ
yiIQs9RID2W7s0hDU5ayrTM1UPxsd2z09IC/Fcyygx/GD+msd6xjGSAwdVvvwsQhbrSd6fVwtyS+
zhbPiREzgj6rKPWIyBZx7RbtQAxt40Q3J+mgyJ56l9KXdPzG9wrDsYYVPvasuQxB6imJ7BDhPJzR
yeuLqvEA5zr33Kzwau0IvJpj+uOHTRpUQjxLNtH+OYe0o/Ha5kfO8eeCbPHrug1vJOq7xTD7WdxY
YqpqRaPdSdeH+Jhqx2SySH3G+WxGuLcsTOJ1PQbUHdzltyJRrWn1lS2pRYP0vW5AZU5web8hkbpg
fVy5fDVdD/jMfAVAMkWbmd8AL0PnnJj7Q8cRRKoXM89psWCHlUgz1/CCdl6lrcLIou29OXnrTL3F
WAhrM4WcDLu4agDTKidC6PwZZwG7GCARB+vQJcmZTwmEJkHXBie2PwXPHGSRa4yIDPJJk4711eod
ZL6RyzJxRmR7FQ9vXcgZ+1/cB5m/Pxn/7brvwleQN4Iqmtzjh5K9+BA0zovmAbbU3mOsTNpfdttD
nNw5fTALbRBd8h/fgss4e66o6c0OnJpgL0PoiSznfrNDZ4IrDC0EabGj1bSfT11B1AebSdAQ8hDF
Rdl428Apu//LIX8CW3CidT+9kDr9XTTgPPFo00p4jtcQ8XXCM3oMT+5787zgZf22BxVfo/J+ZwGO
+6UBjyTh0+uVHPseILxXasiYV5ZycCXAVP+3/jgq/7dIF/vRJ3Fkvtg3QydvvhNWBxyyRk2e1X/i
LnQCGDAaUFfvLQfXDBXZZSc681yCkLNgThxpc9A5rq6MQNukMS+sb0GdFOjW9PebcQbq59/FhDK+
ViNKnpcUR+tkHfrwIA5HVaUL3a1ki5077V/oyVQJMk31ALtO3mw4lslHDJKHPRnGKAPzmXmRmaIO
5s+Tm+5vMAuEgjVmxuzvrBoWpsDg6O9R+w+/4C/ylLSKFuA6SNaykR13RPEVcRgM6LcKB5rfjbCK
s7XaZ7ZtUH0cWwK+ySkM9bTq9vKRK9y+A/jVYoI5F53OfMlekldmxJkDZyywlAZegOnAkCgc6L7w
g8WxMOkabvtHn96xLZbSejoTrjzkippBK04weqAhE80YA7R5BKvmeHupQTBd6Ba6IZUbRCX9gDQX
QsliTuMmIDxNsWmysRN4Bry4N0177ZmmD575A2GI6ObZ9kk6DFSdoVn2SsMnd4TioROqsR53LStm
BgO+V0n/yvMF7zOYzo0vFbvDP6+tyeoOi03MXUM7IlcLP59/SaRtyr65zthQWjXIei4y+SvyDmd1
CwppIPtetOxRg2TWcv6x2gBTjG50BIYxxydOIiKHP4FaEI0beXpVIi4tru1KgGMJKQdtiDALae6w
DQYCewcfNRfUPI6U53slxqYkhwMPbmYSptRQ4SOchHlO7bk/RE1PqfsYzuHo1ZfXyGGDFxDlVObI
3G1FI3D3dtPtSKGzZSFEXxA5tjmFTE9NboqdXgDYQbkSbi6loihuBb4NOP157R1CzNGM7JWwfs7T
13m4MYOsewyAGSD76Pg+WxJKSv3DvyoVcpGz+zf67GXBdnDtTvLa41rezU23jipVzhhGfShuxeWi
537/CW92n7p4L31ya5YLU3l1uu38Z/xkFw8U8w5xYyXbyJ3FGD4j6guD/StMY3w9MWxAyWvtRaGo
nE17jobPN+SIeh0O2TaMiVILMjr1bnrgMHDdjBgW2Qth5J4nQ68j3K8G+/E+tJWboJt1ppTfldwG
6qu4NBRyO8TyOE+FqhtUFeAaKXRrwzT6hJB0PAnLAOwvPYflYAQPJ+IzZQr2F6gbAsXpd0InYCZI
FncJuYhM4HqiamkbFKQtlwspEQ6GSI9UjPdILDjpe5tQ33eBes3J2LSSoc/sAHpND/FtuRCVkII8
ZaPuxCYEZvFG9OxjuMYBzyprYB/+oOaZHoaxo7GOzzFO6UqwM6HOJpQaoeVGZ2FjN1uyXNIJQNpN
2zcOVfxXRbg73Efm3gzI0V8eNTW6ljgS61Ys3VBOix9i347EDA7VHxBcH2uaJaqB6d1ry0b4JjdH
4JCX56pd+VBUG9znWAGXPo+vamvSevaGQwpjJzjLj3zighD9ZY0aa96/CKibDu15sh2WnWUXEo15
Jmwv1Sum+gxt4eJr1lFuLLvq3R9XGpmjwtKz9U9oE5ie+UX78ItLdgzhR+UeyfxxAaRvsFgIRQl8
84jnGtesSnYJmXcdhL+faOlBkUHp3+b1SDkYgSX2ymtlcmp+4FQGXsycco4iJZFHz1rFIC8H3t3i
x2KwH8fvOydXvlad6c6WdObzHh5zADuXrs5mVL9qW1+ZI7HDl/glur1i07g4Wnj3yJJYIVlS9l2y
fWUqHq1MzjmQaOLXm0DrDy66DM4+D/IE8LidUJtsT8rVaZKMCcy5lv3SuP4MQ2n5J1fNwHCbFPI4
84+8/PK3GOe/ZrRBFOAI82kht0IIJaYDqGS9c5bUNXKKOHK4fvZWy6M/f4GJfQquk2fLC6uQkhBS
xrsIpgY9IL5DmOUOtddcN1LJhHbYxoBalojb6PJOihysS8yYBCbreI4S4xXURPSZ/XePwfs5B84q
GPNCUHSbcRLQ1Kk5HwbTF6M5YcCmWGVqPOoTWfPviiNALfWSolP3sWZnk0nIff7iys3yLjeDQwCq
f6CmQvOgw/byscst7H0K+5f+Y1IGavydwpSN+E7ecCItErinEbvjxLsf2n8CCEnZFqFULVDgVbxi
3VCQ4tMSHEOFYZAOg7Iccw/jIcYRolLGZBpjyLKM/fbuXfDYU2fNZdkDWfLzTXLHvSRNuJq59TQ0
z7m/8i3qASK8pb8VsfVxSG44rYVjHHUju4E7UIf1PKDfM1RKUKP0/i89cvzlsJ5msu6/LZvqIO09
ecrwOz2sXt1Fl/aCsRxoH0YHJiqfvkG9CjvfO2bncKZJuNRyrM/D7dxyfYvE1ZHtQhoQVh8nErHm
M9dImbJezj56a/3TgujQ4C03SGeu6wTbhPd2fniDNocXZH1oPYcdaNPV5KkGlMDrp4tGUqcGZG6v
V6PvJ0IdCrPHGmB7ADW+vj91QWpKecdSmr8V/Bo4F+cOZYrejxOvMWvDlkj6ce/gf4hfnA+Gkb/h
qQwd3SMIuO1byfD2ThOQKpO0gJIm4pP0j2EirbaLQT0NJ/dqrDkzGISKIH2EBeDEHnuX77NojDe6
WDh61e1JALnfyxIbsxrKS7OXXxhNuWF1k4Q4MPPz28ZE3cxLjHwhi6SbdDqCZeRgBAxhCpO3yKZO
8TnGOY3rzA+pqMAGaK/oY+pVX2rBu0k/UWM9CpXMtFxHOTSSx7gwa27Mzg9IrZQnBNJtf71HeBZW
ayvl/VAyqlnrCuNvt6w50JQRbzqu1mLZ5f//7Aro599vMTTOSOPqh4QKaPujVF0rH9nz9mfa5OYW
8iR5LQ+NsR+zemZDp9Ba5g2LDV37eZLcfRdfM/zWuV5Gk+cT1BW0u68Ndi92fRVLe4fHM38XPHyn
P6ZDDq7Hj5mScBA0PmzumrEEuWwaJWJwMKiesEBSQADh5c6BABdJ2zsgLcz4yuNJ1PeBbuvQPUdi
4Cla7NiYD+ak49tqvep5RqPPwRG3jMs7eDd4T5J/oDTGrcGID2qKK73KNepTX8IwHVlI5mKprbe/
Vg3A8dypG3TF1iu21ef+Iru+aRLtdJ45EUzVd5dWqG0RYjHgHsw1umOSlfh98BOSI94jrXfg2YpB
a6lhwDNDXUpyQrUAQw3Lm57qlzmuMD1vewp1Lw6bMrAygnsOzNbx2qp4zTYWn2Qzmg2XZEZzQ0oK
10W+P0rn+hgFNd0r0d7c5otI4omcYZcOBmaXt3MyV0hPd+WB6bLFUa+zgP1/RycFLYae6ehAyIuj
gRplxvT7gTMJmriNPlvWwA+jXdZntQqoPSX9B/goHDWx3MiBJHYj8F+rpxXP8jTjO1nC4D10Y2US
lGvaGHr08OZutN0MGKF1u9IduNTQa/FaBGZ+N63lb9qddHvegj0Zx3DdrMkv+zUcMcw+qoMdwIVQ
GPHCHhb/ODZV+Za09r+Px0X5k0pMfZTSKA+c+FPKlor0gKS3Sb9n2iQ3eZNt2s/JwJb9/HF71haF
nDoA6m41HR2SR4NUawMBQji8fMFBj3GLtRlaLZBzzRpgsuCkuL5aHRoUs9WGt5TeOgWysB238/EX
8yFfcn+rXx+iY42sfis1vjQsqEX3VpPpHYO7DNaB11lK7KqCifmO1ml2z7bGGRBKeeCc7wE7ui4k
ejY8+XRta8VWkGvE/kfJkePZh9oZ/LlrKHx2FCGO4vbEwa6On/2PVaj+/HCREnHAgqXieXLpv2T1
FB/sO4Ftz3WyhHZIFao98ZSvLp6++yUrOU2ebLK2mGdnGVBz6PSCTka5XlTtjDeXoE873cyMSrkz
LNMGg+MBfyUdL09oWgm9S2yzKJle2WPE2ZNt6sshe8AWKtJzdd7rxY2h9oW9+KxBc/vJF81+g4Yz
GO42T8sw46XhA6DUe3hDywiPNCAO09SN1TfBOBZwP5ZpR6UIIgbU9DhyxXSk4Xs9PeLV+oF3E9by
Edh8yV+SoBLEAiCGbcl+LxpWxggujueZggc+9ju5Rs2x+Z9dgYJFTN6VYjublgP3iTO71lqPRUDX
2pGG7tKDJkcdC4meeXqCbSK3XcTpqx9nZVLTMs6oIO2H4QHDNuL6jxz/tQUwBqHqtjm4OGO97qyj
6lcSJ/iZxt5UbUbKzJP0d2WzSuxlOReRLgrVfwhduF7InAER0th2QLh+6Kj2L8vb9aHNicDzFiZq
6PGGQ511OkP68bYn1WApjMBMxbPu/j7ka8/ztG9XzW6iBNECi4TTOLwT0RQhBv75CESwAIvMe3kk
ElMOeCMhiH67DBUp2r26FbBz3K62aYg2fJGeSdysA3pUq/ciGpzzUTWr5nlCkC/d3tqfjsDT2PV4
SDFpEF3HvSCKqoGORIqOob9QzKf2DDUoyxyAeSN5mWPaLgGNWcBh8AhREWqnBHQSkaBbgfxit9Tw
39huEKG24dUjhQaWUQ6ELBXfP+7mr3ouDs67Iluw7bSqM9VYtEq1sIYziyFs77Z6fykZKyb51Afk
vglxzWkp0nNr7xR3QkntwiS8zZpT2jDy2H+KcFWFdgQQoOitaQUWREf8gasiRLkwcpGNvM3mHxDC
eKQoDuLkBChLCCXNZwYw6d5aBy19z2/RcuBr6vCNiYxpojZ0czCBM1fgyupU+DyxENp0NwYvgmBq
hRftVh4HfErT6YJr0V7dwbpfqT3oHP90luN9HVEbpP/amZXH9Q8sPp8Y9maT/td3H0yJoD+SSdJg
NFaeNe2i4XkuM9QtMjo3rgxmwenHFUyfS4+2sLRrxFGXd6lbwGJ/ltkZ5vvbDEier9qdoj6Ox19j
q2ovi8TujutgI1kG/DjCOBKk44DLMdMfC57kMJyJkHjHmgM/wVBVPeBRxZwKx4scPurBZwuNrSLt
3VdljGt2RuHvzxYU7pcH1FPwhh+JHhgz0xFxDNZ+Fpt62iHb9ur9KwgHVargftzrqZ/PMDgv25Gi
cmmf/cDcP+TvDEuix54z0gnwzVe+uI+fWQl1i5rGHwtPfwqc5Eo5oiYty6sXSWqyR1i5RSQz+Fmx
UVCI3aRpqLhLfpQUGTzhYftFb8PDfgXnnnIXRCu2mLUd6Pi0jkyYbd/uBde4jjMT6NznvqCXq7hI
cAyNeOEvA2nI4YAQJfK5e3lLVNtyYAj7atsH2ypZ4W3LTMt9HWWuZ9HKsiWfh4A20JYNPHiI5w3H
/JMwIvPoCUHvg9afxhLemVr3eoKTwh2TfbSXTi9lhk1ipySm8+jw95ZzCd9f2HBnUkvhkRZQc9ei
22qbd/g3jdXO5TRhpuhtC2EFWeRBx3CIdkzz2w87RHk2YH8bhySeigleh4flqj9y9W2rFkvf0+ZK
DRBmAJieL3JJJsD4ZA/KP63oSsbuq+dB94DL47KYEcbDnlkRxs7cL3wvFlM4wlFP31idiOaJs9rk
laZl3l6L4YAlkj8m4Ucnc7Ey/ClykupRk47Wi2RpCh6qlkdvgi2WVI4zu/8YKpkDTBvY+mV7k6zt
xmH2T0STo5hzyA3i4wJJz8VljwgUYaBudwcdrcTfVCryp9LBuZeO1qD/grxjfmeYHKsdmWi32v1+
qWmcLKkdFhH+JLtc7qCUxVohlwgBBurfs/3Mm1AK6Gw7hznFn89ooVc+D7dR0/nfO/PoX6LLl6er
mohEd2CbKQ52agk1ROu9D7oondQX7As2Ge8LT4vJq3scVhnXuGK7sTsQYiUtN8leVcRfzM0P+0tO
kIJYTQFj7dzI6Da2LNPTwWRL7p/TK2m7yoq9ACzMAqGtzmB7sAj5ifxMoQ+k8f2vb2wu8sAosgp0
AOmr4DS8lV542jXynx99kBksvSjFkgv7Us+tnWFW93i/ca5Wq3Dux8253bXIzeLLZlhUCVrcKTga
RWx9t3fV+RuSQ+00ode3TJfnMW5rXz5oEm7aoI6BL7y4zpxIkWc6QTG9yNAk+jZy/dCwZSrI2TvM
4hMUk2RfsfAJfHWCZ63bFoRiB6hVm+DXLZTLPsdpa6gr38g2HGIhwsTx/r2oUQDRTfgnGbVUGImY
oAd73qd5jlqdJPDhMYrvE11UmrDOSKrmn1sqX8o+BV7T3lpjvuD6QuK/SBUnTq4x8X0eRfS/vi97
s2Ebx/M1zjz8/wguiCYejwIBK8DjTi3GxNhtgrtt5msRfLwn10EHZhc0dRW6YX6uL3AKS+WxIx/r
OGTijkcN0sJNlOXTHm84UgICbo1DTvEXC4clMAGUDuJoop/pZm+x8WVzcG/KkwNcA4nr6UM7VnGf
Ab0Joz9q+lPbU1+V258EJJoL6nS2IKgDWuu65wEwL1sHxIe8ExgR4/Gxu6V+mpyfqu1wvFN3cet1
DJSsZY21JYOBIZ9vqEilGOrEb8IZHMynGNuYgmVpHGbC9bkZLjP8svg2dj2Asmlhs7ay5IJ6Qj2s
3u1CI8NvFJxKKp5b7g9rSFys7Ol8Zxz1w6Nc9pnyi55k1dfnDeLJFn0CvSJBqDhc+T18sOkvZIBf
9yIXb/oppEEq50VE4LhdjHSPT7uSO38bXSa7PcuG4z/gt/1IdDsjjgd23IydO3vGu6rPAEGUywOj
q0WRFQCp2Au6pZn+EkeQv/yol9n53P9auDKfNFIDjECqZdIr21kBnKt5SAQPXNg5AE0C5Y6cNS11
Es8O4L58UfFqu5i0CRyFaDWsKch4xnXbpjXw158CewEa3FzZSY+mMZsgT8pdYCSve6clhvatMD/u
OaiIGrrlheP55+IwqgkewARFd8rOqSZgtH4jyrA2r+02uo1gcFA5SCiBm6fb6mIGNvhfCaXWeUfb
7QXWBGuL76Lx7Gx53hHE5jOe4iHczB+bMaTjUJ48c5SaCfod/4ZJJ4zFR3r28alhXSX29kDtHMTg
RNNlablf/hf6/R1oznGLp2PhjdseJY3U/W2ZaQMhUeLZ31bDrABQvyzRwHCBkg7Z18gwx+DRL6z1
yACYpNn1bzWfdeuxrCWvPca9/ERTZZKWO5PY7E3r5bO7da3WRDcRRCtoJZLS1QaTyhVTb8hBLIc5
qFBbNZ2HdOFG1obAmTBPho970wvMqpifU3yBr4dwUX0dfayFHAdesW45mZVprU0cO0CWsqsNsgD0
6DmdmZaedoT9hQOXpXrb7ypsyQRfCUKd556dR8tVXxVv892/nLc9GA7X44FbxS/03mL+CM9lWfEE
ZWyVh2zdhVlfKob0+NGjGRuUgkDwkrNgmeS2hEMRN159CyYLd9tyiUvK/XdvOXCUmXstWlZ9Ko2Y
MWVBZo/ELr6H3ZR4VphTh/h1y0xhhTVGGrLume+Hhblt4O0Ijs5bBaEGRUbeLRQaabL97N2XDavP
v/tca4vCHO0mypsJX8d3UOxd0/7NJr6bEnWH78G4UqqbGYvh5bHq1RoKwatUUNZiBdmAJp15l2F1
YeaB+kcha1X/RYTbTLYb35PXkfTmAt2TlIQ1Ganc1WuRcvHrRGsiWHkVODc0k3/eV8ftl2xdhGUP
8ltlIFg4K5QrEJCAD63vFliaNdQ//ESgPmLTkC435ML/PBce644hzhRRqIMzM5YXydyK9sZu0qoC
O7aOXhUgzUmqbGaRdQBaJkXwqBPaFbhE2cDXDvUc7SvME4InUKpO1PxGQA99QjZpMsyZ8JC5cdyw
KIgj7zy2ryvLDHH8/ufOJ98yXsObbpBT7MnyVGcSJGzB0mrr4KiIQOpwDYD09EEUUc2uNR8EHwy4
UiyK6ldGFxoLKE3fZwu/wjhERBax0m83RS0AzT7MX9KoQovFZjhJT4sQi0o9HkZhqOKp1AfsoY5Y
/VozIeqZd+SSIs+BepyuPUp6msEk1aOAh0N/zLzIvn5bnIa847PwAp1YuMqErDlsCSDXfwO87cNa
pzAoO83QQ1AjmlX90/7kOAy2siD5NsLT8QWutL7P95Tw9AOOLTJDDI/fPMt11tqsAwiK6p8ZiXNh
ly7oMPBVWzo+e/PvbKbErHXrE6WjbBT2ZjMLgTgN+4uQpAG6eL9ajEC7BhaC+uIBIY3ItNXr1T+p
KXcS81Z1Sw/b2LplTaEEmFcpZ3TMzDV6vRaSNiSlTXod84cbi/tKmeB+jNpYBVZl0HOFTarT2LDb
jMHlttEcSdbqcR9g4Y+J8GvRM/qV+Sv3g+1iVxYyJFr/I2b7d3Nfs/F18h1RVz9c2iUGd2TIkubj
cL41knxqNvnifr+zmAkLCfMa1m6Piw69bC6c3Si4G8dx24Bs8gWX8ys/dRWuOfVFaeeVjnqS697W
dmXN/88kVJi9GXog2hJIoCqriRmvKnHNzUb7UCl4lb43x7uEBv/NRr4NBqJileoFe0jBouuwSxYp
gAMGE2DDwyPURd3JYju7Dx8fszyp2EtMRsRMcaavr9SqFUp5U9z+ljmbJCD75HFrxbhpcI8+L5At
vH1nenJRUvDMNybeRCuoU1XTyDqpJ/YOWz+fXARxlgi0qawwjuANzAVQm+CIzGz+aurCoqx6MTOt
lETnB7RTARMht96ZXzC6/H53Znob2SzfBZz7lpl3qvJoAIjOp0MhZdXVw5PaVRdMomhkFJlT1rng
puWiO261R0qQMx0uPPYcqfs27VEBXCzwwdcky5HR0Pf5DlZ+tek4SLHVz71DeGgXAW0+eO8Ufh4I
P+j4FtHF1WV7+hLachSUa+PSREdB8D+AstCh/thEs7BPM1ZIHnBgnGcSk8xvUykJWwjkRZattJ1u
QISh3uekZssLeKtblDrQjXkh6Zx/a3q05uPP6wLk08m3gVpMYLQ07CKoIY1RaS6PnKsCHsJnw7B3
/qWTlxLExp+Mng9uB2DheMsSfxAjixuo4VZHuW61YKTxZuQzfeBSAYeDRsKhIxa4lean4F86SPt0
dBcJdCqpYNvEYNc2yeJNUeFz1VugnUUNkL+YqHSxSA0iewjXmXMxDpVS/WSj5TEwTS+cqHL4Llbx
DYk4UgKsdHmD/zsolyGcJP4P3Pm6pHkchybdSjZzmb5KFSHvVDpqtTXfgRTp1rV9mHGYcKBjlm0l
woxCPy38Ne6IW6eEiXoRLvK5w29/ul6D191qbDb8Fmq1KqMfwVidLn2GpG4HeejfHs30aGgASqxW
h4i6o+yk8SvF9EDBd223gzqPVUiKZ39WFs4jtIZAT4wfQWjjOzzxEVbUUSsXDc2rti/BibSLSOID
N/ABJiGGC3T5qTYIL0KNFQzjLWe4tUHenbxEypZUp4+j+rO+7ojRr2uh07mDhZrFfg6lkBbxgMFu
JjzSLauQG1Y4stX6k6dRU6j/dBvm0WZRyxno7/RmSeSwo894CZlyiqj2n8F3yJMyGcUlcMVZhyEo
nVgAI8yePR+d639fbmzWI3hx8g5Z9niZ8a48D6xKNtiRpVgcSlV63mGUk52337RbzZ4S0J0snGyH
iJicrSzcshJ/0o8HyGPV/Qc2JmlglYbwV7FZKecJ67PGBvWURybwTW5K/+7v8KMJhjl1O5CXBsS0
TnP7u5P8+Utv/4SYF+SHLzq6UaXlnRnFCcoMrijrUQ6Pele/0WtEgKg3NyxeXvEjugg3usxdquDf
g6pYXJytTkTXXHws3nvqxEUaI2qM6WSZ5YganpU8rYIfFt4petRapoGlURtl8bv1zxxylRIq2IG9
tiJy8u9KEcINSfMxytxQYsXs0gkuEyZnvzt4iUcoGjBsXresVHfehMaMDJn2NxbWKGw61E03mB6y
YtH2Gwm9Q/MkTBrCLRz9tWgMOFiPrSkFx0MN/83P1X6XCgmH+6BsK+IvzhyxlILUh9RNKN0+NrgK
Jx0hAi/czp8bdC0rjzf3QZH9sOFedQ/H7OSsttLds4DBa70bCdDuApy6dB7HvecERODGvIuRlxml
lV7glkjyDIRG+PFk1gAC3WeCb3l5tpqeM0a9tGKfVHa0rajt/O3TgVmPHf7ME/F64Sfi55YFUBOU
Eh8wD8DjtiGDZbnJlLx9Jc7XeF+MMafyoItISIhwArJruLBBGDT3IlASSUwkir2Pf6U62rXKETsR
UWIC/Ami5TxeRC4ovYRuaS1uc6nkIiiM2FmQ9Ao/euTfjdbIhA3CD+EsC0peMAKjTUZJTjTP2YkI
zjNPxBCWZYr6J22r+wlJaVsDj4BrUKdH8sT3PDmKXqCCmRavDKpe9/yWiA9MEoKSsOMIm3gtGFVX
dcC5u1Iy2VMkGzc2QXJ6pGl8x6U6ZPoNRUYMvwwZshkHLii6Z0kI5M3kTCIMLoKeA9mA/RJL8iqB
Oke/gBSt6q34H0C4Q1RtNF4wSh0WMPa7yFpbDABo6T7NpH4rSSnAMceAzyNzV4zIUNA5x6dkmCmj
dxRRSEdddinxLPcmrbXN5fcv6FXtX/OP5EARa2pYZeQzm4nyhFMz7XnRPm4THNpdocTLNi6PnNjS
x/A4j+w3WnSLpDMagUfY50QLulY/JLbI4RJSrep8Rwuo0caU1IFoo0hSL7k0qtlg+6LqbXDQV1oB
wOPksnPkVy3RgwY7Q1EzFb10mWXLfpffABWqtnmEq8VidmIugKsyIjT5+lEr+yLArAG5D1AtKYxz
irFUncDbKpn2Jt2sJ9aEzjWX535v7qRb9gOk7AJ09g+ihRsWRGOQqfx98t7JDAOycyZyYHDiTPj/
64m0/MhtMV8ft2UvArmIgLDffvUE9vjhz4i/zDC14sL00zm+ykbY0Vhe9AdIYhq8NmX8Cz2WXSNr
Eocv+T4jCFNcHcjUE9Yof1PWm+B4Oyvdqc52VVtwB7HMOZVzoRAFvWD5eHiVUOmcSc4/MUq4onDW
JpVT9EDNmlFD6gN7ovvZNKlb36kIHEgc9xnXT59ZlpFaVfuKXfc0o2yvvfNiRu8aujOrEGAlXzFI
VaZRJ32zN/3V6uPyLuxhOPR4vI4RraxVcRg1HPReQTw+tyzUTQcGk4b7bz2bfQShPjeAEZSe7bWk
a/5GpgZ8elz4gDtjwVWrOHGsdSa3XMnRw8NRKDt9as7TbUEaWRiC2HVG63EwnBYx/AxW7R8u/fKQ
+NbSP7zGaj6DPVKXJx7pjN+bjPtEnQEKpJGZryuGuiPQcMZgXs6Er50yRVbEkciPbqEB8fON09QG
DzfWipoOIi481GZg7W4T/y+3DuX7KVjq11UKkxDXXfOQ1KDlMIuMhmbZo2S/Z1HyxWZg4dRbP3tR
IcEsvnndb3F+dce0+csv/sFsEzABSkcsh5t4EhI35U60Brb3xq97VZxn8bZT/S4SdvazxBUlzwlv
ll9tqxSH8NW2nU53V2BqJn84418V2wVr/tRRNl5bwMA5gMUNaSaU+ihO3RUH/KhttacmSh8BRnwy
E0RSUHbYyudyUYsVR1E0ZrS0cHbBQL5QApFBb+0nph2Ai9lsS4cyZyYVA1poDrZNB+CGaogsaJPU
0nJhJ+ezIK2yZePA7EFtFGpAKxE2sl6cKwj9cv6VDrWYBosVuCueJ5QERx3TM2/we6lkJqHkiRLD
XRXnVGj9D4K7jk2iu2KmoJk+Pbk6kHEj3g3GMVK8i6jJ4+ZIfkg5WRBcq9aaJMgUq1vyHNzEo8A1
m1iO5y1tVlUJRqDXCzeHmC7vda4Y5sh0xt3b9PzVVgGnebxt7Wf2JbRVDZ3FqDy8bOZEJsf1pcFQ
TklqfiqEMu7U+PLatSanDG2wBRtjJCaAJDSbX338VNXrvbO/TWHPMCHZcOCnQiYOkt0kcscmNxJX
JA5c3WPOWbINnWOvJHS6K5HYXQmwz+enr0VYrKQCtC9Vni76Tebzwpaux4KygGiFcw4h4qZTfpCB
7YxRuVrOaM1IaCfe6Kwp+D68mbhPHth+3RFt6fDkLUgWQyoAF+erV/fHGWp8cMxh4IKKKDYQZC+A
bezQIF5cVN/TSPVv4wZfkHp3sjuubbBc6SRgGwCOum6JUAiLwycojEZqx0zfeUCiZlFmTuQmigLy
vzFPw1ldg9gmcj/zn/lj7Zh6Z+oEz7xbXJghR7kVfhqcyV5yZwJTLnYOejeAx84xrSo4uUAMWFbZ
Nbj+K+p6pWH4bFnZCMybINylVLYq3kApjYu7/whhs+/gVI6QEPiC939srnsd4Y2wZZHOm79H4Ki3
4cLQbMhA4e0oEmN+Uc6vCbglEoSu4j6J48hEpUwZNF2LMQBh9yl3YZHik3G/o4BtJdJPPYmqEKtt
IO0WPu8BiSP5eQ/VcmmG9wkvC0j2KfiOJIqZpbF1bQXmQ2+5XIZPn/2J7vMaiPB6gHQ+2ATooA4s
FkUOoKz0WVGWBuHf7qriJENI8sx/qRihBpqhEwATxzDTSZwmhqzSyuat3wUgUJXonro16/PuBBgP
S2ghRkxgQ4ziYk+I9eOBRJDKC9C1VYaEdadD19ho+uyNhOst8qX+oqSnKrtuDHOfeJxmOjIEk28a
NBnrVRuQQOiI6gQgKLPir54k4+n0+q6KCIFVJZ4Bf7StJFuuTOLot/Yk/bugNRvMqckaj756VJqr
UFNOKbXL0snNT+reqTY2UpYuvIRR48UyqJj1g37fJLsR8R8GpKTdKZ5lev/NQZqmzkxzukfJwfpu
8IZQeRuffrv5PCaPxE5/sXzBOHqpuF1HxPJMayqBzGmHDLwMqiu6F/kclz1/O7w4HKm9XhlFzDfW
SY2aIggIPTon95FYRd8lTSNUcLxH+I3t/szsaUEH0Kfh3C6FHJ99aP0qnV0vfGZ3NDnZBysahxCR
yBT5HePayKyw96lAd3EEzXaDSUWn8ATQ5YdLi8qOb7PfvtfQrkAvEyiRmYSCGBl2T2sg7g/FeKeW
haATJYP1EyMCTTnel55daIQi9e0lkv1PhQo3GxxaPz1qqzVP2b/RULLl+IzIpuoGq3AqSIz1UX5u
LKW3WK7vHKj8SbJx8n4wio4ZBNFAP5a2yGXAjggCMtXCWI80XdIVlEKWgy8E49XJdE/wbcmyuDjB
vjWbuL6qkqSZBmHOE2fK774MpIa1BwPFISQv5CWbtX4vf2tgrzqoyUgzIlxyxOWACj9ENzlf7pWJ
uXq1T//l2eY7nRGOKcjasDuPMqFWsqFPASio7DTs/IaYS/bcBJ9MEZkmI4KAuk6EDLVu+mbdEUAZ
TMRk9YM1jMxQ7rcLR2cVrp0ul1S/BCM1MPjorfdH3hyXjMVSKKXJGLudS3HPDT6usXsVVqsaLt7G
hexLy3xb28dj/LvyrEbEN4QiQn5Z1LvKgyLocvaI+ndpQ6vU/Y+/vBVfzRuECp+P+BOPUvU7CG5a
ISgvdeeLdPat3KgCaRKuW4iT9Fw/DZEYDOAQ1iF8a1gHuxOxg/t/M9tM6hnFr0aZYP20kAuSH5mK
+itNcaqFJIrtLqEfZAfeJ6CRE6ilU5BwlDx2RipWoUlBPPlwY/9ed6tXHe00x5fuCLDc5ZWCT1cc
h5xIN6pkM0V9PFFV1CPZwHoUYpth8rsrODf2BZYDg3e8oUfI0uleqAqeAyme4DPpQPt87wM3w2V0
Z/WitwdhFvBLqJ7l5WWSg+A5kWujzeGkaUgWzAtlOM9omIYIyUT/d2ktfBHXjjjVTOOZCPkn8kpY
v7kY3Cbwc8E1zwRoahThhmh6ikybNJNTl7upDYWQ7N7w+1cqp7ZY6Yfiov9T9FMnRmIpsl8mj0KN
e+6EUV6wDFiPhTryy38wZPEzbzCtYWoe3vFqCRi0wgK9jR7gRTGcXFxym1Gx2fN2p+O5ZjL9W8v2
BRim4pJLcCg4TFWO6qytaYjU7xMG7MK7G1sNWE/lKyqs9NRgQmOATZOKF1xs+VWbrAhbwfb12dDn
pWsiI85IgCkiWAEpc4cQoN/6gzs4o/BJcd5AHNP4lHSWXLp91any7NeQFkmOUMldXnLtz6llg9F5
SdS8GIcaqLREC/7hMLPrF/duR/ttu3D1UyKNLXzgdvoWHE6RqY7vzD5xYhJ2aUHgkvQcd4PXEk66
x9qOy3SlaE8K5C7/RSzBsLEm/CRzddmQCwnkC+RWubnXEsoca1Yb71d6MKS9vcnHPoNStfk1o7+A
HkwGQXMfxBKrj7aqjRqbICMg7ssWdKM12+12Flfm473HE98p4qHtwFmF25YdjgbCvsbblsfTfKXN
IwCTxZN0Q+BpbmrY3aPOz0HogeRMtjOrNkXeTcKESZt8d27D6FFs4DJn2EqJdBAKjbBHUZCCvwSC
VUmWq3gVrjIT6jcCEu2+JLdIMkDYu6a3yTjx37lh4NqPuvXQtFyp7pClW0nHokiSZLvmm7BbK7/4
ipSKNTSk9hGg1qW+W5+QLaDSaNXPGzqyAoG+ev95uXR7fIRJPeFPI43XQsZy1riHnV4+wEOZNxPj
uP1UqvGuMVLQK7qH7va7o/JU9yFArmPZln4KTqd2CasLsGc7Dy3+n4mgSieEF9OWBvgjBtisnFvj
XDASBsj1D7OYIQwPga2ulDD7PLuOaBalLDniMg+skShjD0eEw73AzTi2ckeFCNZJklxFmg13n6p0
TItfsu4ye/WRGG2d/zQ5fAuvDvnm/8MXwnFQOT0gH7aYrxhEZxc7QsOtw4l+RaOwhxw+I1IbJMHN
poUqJ9BhKSmp21YhbxJN+pFvrpj6LQ9xReTIDcCegKdEY6dKz95QLsKrj7WHQS4rGbrToaj1tRyB
TtI0PWVcElQtsV59qlX5OxoLgpjC+98Y8ZoMsFbwt62VXykVPzbvAFM29UBTKg9lwVT6fBQ2HIWx
CkLIWO5jnYEkSy35mebv1OQvBPf+9YpZQDOhVKt9nFV8X8McGZbDSWWGZ18VwtEvDhToxEz/X33P
tKz52RtU9sJl0NA7TaMGsFetM+thtTEEn+jgpubcBsKs8al5vwfoXPXZ+DggmXOVKTG8aLC6rN0w
dlCpDlNJsZ29FXhah1j+nufi8ZsGmtU8pxepBlTTXHrHzOOJCuz/SinkyMseB2Y8+5icDQeqU0yH
GOCTtqmXihl4vOBuontvicH1xvN4E2rkzgsBOOVz6nm47S3rmm5LBdoRhO+wUwgVQtNjViFA680A
kYS5+8Asbfw6ExBBjnKvBCRYn5yKgucREnFUVoEIq9crdd6GRRRrNpCFDsL0zGghcrWJea3pbF4z
zxpjGHnQEGmgdTGICkoj1dlFjhbeNCT14LBxafsInUKbSC0lMNRdSXysqn+YKpV+MTKAK45y4RMa
ZqnUhV1CYr4gdU4X+uLc4tjZFRZ7qVyUQGYY03NxtUDn7HYT/wTIAk+5SraiJfDToIn3AajX6Iur
8nNpIri6vtMO1bnwOpDb+NRPrNHgaz6kDhiY9yFNnoj3oBxZ8MLyiTlNWaeukZqi7ftZQO9GQsuO
NkCIEXnFV4MQ53GkIferbCkiv1HdtGWa6jTXDH056ZMAwf6c8eudjD8X9Dd5ZniZ30Fpqw94gLji
g2PUsRNYemZ5RygtRJmnwliNwsdzmZ+uhkeLam8mPQbVu5qC+8/NcGmUuzTt+4nSDa6gZ9BGDiao
NqjWLNo2Ke5oDj1qSBX9R167TQOU0HDIgNBTCjTEpcY5nWKfE7vAir4Go7/K5AjJBJvsC4MuM5Wk
5iXXdi16xUjz6ecCfbznNi72dhKdF6RJXwfg4KC2ELf/sF1h9CAJumd1pq3uEJPcePIhH1gSrKXx
QSbjUhA7Mxb61wijiEykAoK4+akIfT2PePUKBRn0ynB2ON+cazM8UCVgZk0ZV/6dW2Fs1HXCOMW2
2pEzrxOWdaQBrOHHgyAuc4ZYE21NpgYkk4k7vzBdscN4+b33cEWnZVnLFbFJHVssAo6VqIRLBUJu
DzOY41l/lfEclHYzFZGDvcAqHSJAvvF7rUZTDffyz+SbKeNvDlAf0CQvFIFMFyuCFGN6Uh7nL/4u
VLZJQZSIAms6wDIUz1mr6P7eYKmlldUqAiE/CnU6L6jzpNQM7K9luOKyF8BXK8S9OqkEQBH8E3zD
uEu09eSQO+Udunt8VtQ+HvByFTGtej55Uh4chvzCsRuGhNeB3l1wFDkQuoMviIQvx/5foMZ3xTGd
dgBVHNQrj8QNkBoS8A42EP+4JlKCS15Z93HEGaGfUBhfy2KMIwpwhI5ZXp9Ssva/53ecb7JrcQCC
mgbOMZUgarUhm4uUfh3WtcT/m82Oah5k+Lp0grjfjBFRw6ZWEOg0R78XONNzslg6CzOD0fClbF1K
YSi10RrtrWn8hEbcrASoR+VdmKws21BI1dp4JrfQsF8UyxwX+ZRKRtHX2RWXIUfdflCeMBOFeY5x
c9RBM1+DHua25m56Adn/vfxo5D/Os8y0WIC35Y5aq9cLrafWMv80E8W/EFbtCK0Fl7e4NBlkDmKY
BBtlWhG/wxoexEF37OyM7RXDaxhIZnqv7nyu9usNJQBTAx4m8Y0bxv2UXYe8YfmWFP3PXhnSuSFp
kmKRjye5347SYUHYafxdFroBlif/S4HzJg3Q/Lv2CSf7rVEEXb1yqMAXwxrgEhUQBuUkMFK6iUhJ
3L1xLg0E4IvtxXSc9VZQPJgvJYyevCS4fn+/SOFO56x8Y2h6HxmrYi7vOWK1fgzdTKSWOw+cgZow
m08d8daENWYBRXU9sexGGIvQ5aNAWDrT9N8GXAbDJFGsTdZRyKdulOGaE1/gq2KpFW79HweTn9X7
M5VvXWOLF5OHnW30hmeDke9vmvUg6C1rUi0MlSnb81MW5GWCCpah/eEqXdNA3ZHjqUVnfWIdXwKx
yi8mONj2aIdAJsY0krcKWxj3DL5lK8MhLXiW3go+EAylXjSa+PUBEWIGXqS/SL4JRpHwvaUJHJTJ
1DRuyvKsWVHn50kdBM/xrzgtpufzxuMxlKTKyjkfuD34fxNId+Ad+LKP/eLwypk8QjXZaettHVV3
2S4YIafBhWdd+hOIIkZpxQVnwxKFAJxN+wLIjYWep+jYnvO3xaVhwEpIxbUXMKX3QwOv8hDcqhOG
xlCdIxqZVbFnqsC46RgX5oRygGNY0lS3JmCjyZ8LbBnYILuUFoxRZIf6pG4x6YIUzHsAgfv+9qAk
9N0jG8U90PWGumlCgoMzDoV10TZRW1GQ5klCAacETgM9aTxSM2uCFF9ekmtWEPr8X/5JDa309bsr
yyBL4b4dLuDEjabyzHeIDl1iPFDTMb7YkOJzjtqFIxrZhZgxbL07rRqGVc8bWT/ArKtFtf1ttONC
eu7zWQOa7220RmBd/B2LS4UMBDkDHDnMwvctKRgv5auUi2FWuPBMFe/DYXNqzlR9usT2pbPiw3XM
6CC2amO6QTj1FxxL2CyEZnielCSCU6ndQh1Z4WdcC6cQZxOLdBkV2S5n4dozKUhAcjqKHkPUWPXS
E5SAUK+NRwZjyYdZ9bVHzm6viFeifmLcbCL0rWYbSmm49gUHcFK+89tkpA4VszCUeJAuVaCdI/zT
IYx1MoHqbCZ3TRDShCejhcV999SLDn66FelHOMH1B2fp5jM8vUhEDh9FDhPrO8ZEeaU1ipn4kb27
dJGpL/B1wk+CqkMPtCJGGBLhLZ5h9NPCdnMlL8FuC9ixr8ZsgkMHvJpyFBVOP9KY2wla6QbupNxh
Udo/pDxckOwNYxsRcoDyoO0im0gJtEIyTqcsSIr2+QNCGxmSmpZtlkAiq8T0gU9FQS2Avg6KRAi+
LTPo7bszW1esG/74p3b5UjsTORB3gBvApLIxnd+RxUz8UfYK+xirKr6M3Qp5KuCu4ls1K1foJcOR
7MH+csgCaM+hgrsSd2NwAcD7EvHwRX4BqX8pDVLqOHk6CgmpWeLSdZUSePcvIishXaxb3/PQS8v0
W6zTvpjO4L4PQnSXS9CZQrxLlgz/CeSplairrvnbxPfE0L5TJvRX3dZl7jNicuV54vhCHGrJTAjr
R0daVbDyvIxMtnM3+VcOKcAnV7NnQri4N8eLQyKlSFJUO7r0EBNzfEkwFPX1sGpK5FYAQGgj1ud2
Iw+IFPQ3VgQG+nvQsH0vQKqP39Yw5gVUY61cQJJxOTFO0pgxZ1bws43TG6pXNBg6cpgJn9PJygrw
Yqk/x4bt0M8Kyop3PN4ZJlxyp8oV4g+4IqfTGyRLYvr+r7IhVmnrgFntqP80K3LKvMhlF9bxJvsU
4wYcC6IjMSVfG8mxrt+wcdYXxHbu+HaCHx2tsfq9swqMd18xtlF633bQ9fq9tTD9NQP4y8Vzn7sc
5ziaD9BW2vDtkU1dQjuKOgYDs8EZWSS//q4DqTIEIk45c7NxF+U4CTSdjc27prU1QhJkRuc0715J
S6OoDKzcqyMG0r8a3Z4GYhoaD+VfKKWHvkqzyxpJ52lAQG0gosC/clrvjqb6DB/doYO90+QLNxq8
HECsBmgeGQR57KEHDlZc9dOlHHkiMfWu+ZbkJEn0kGYe5rIR2AFqdpul/t95Ia9YKS1znhudch2T
vhh1rwlfGyt/ZkrFgAx1vMykbF6GjlzYeOmBUBh1COjJtMLAxnZ8HqqGjq3VWY8AzblV9Y/DpN3q
15Tb3jOod6AJZCteolLLU4jbH3UT1c2DtbGprtz7fLULcyoGK8YhX1d8pE2ZIIRiYydQIyhL2/rk
/2uhyHW15SLg9chkgwTsj8cbMtFsLrsNPvO9A3bRR0e2aUcw4N9HcXnVn1wtVJ5HoO6Epi8iSIHc
b6Eyf5gKloyPFe1gXpVJu/AAXi2sAAw1dadLm/6AQCQgvO00FAOgyumtX54zwABpJhn7ae7AReHE
K8PabdcbO4J6pG/wIdgALvTTt+tQ2/gcoWkk/6pY7VnqarIGO6kBgR9WxfHW1x1VvGRbBmcKNoey
43uKJj2Vn4JqJwE56hjQL+pkKcKg4pQrE1CKXiEPcDZv+m8Ey3BwkRjqp9Y9168szJNFmijg+Uaw
Yx2wKM63DgAsjmUn24NGfRy1aKHVEmMeJlyiJw8l/Rk0I+AY+/MxA9R/AnJ6E+hm8mKThyyHCLrB
R2KomhME3+ga+j+ognbjEO73dzs/PPrHirkmrKCZMM7hwsu2kBiCJTdA3hjzZe9Y+ZNDZyiWOd5+
rzIyJh1I2lFyDYaR+shZ0rU4ouYBGu4MnI3AhefnrKLdUvDXiyYpBwa+uoEaqMLqPKGGXHBmcCex
4rYqe1IoDaaO/0yUBY+DgZol2VnTrPoHa8IG1F3h6fvW8auMMWvNRwFmwotfCvVu5/k9V222uALb
0fcrtb3v03KpzHHlboG07LpBBT/r2sX8DXPHHBLEPGxdb1yfrT2HhuxlRWYi3GzUobuiBsXZHrxk
qF+8RE0fyznC0umCz4eUL67yVkcmMqfsrdP+jCRA/P0WHdCbMT4wi906FiMZmLUYT8dcdAC2Cw9p
0J188imEUnaiOPg5cphuRJNbH7C0Xmt1Tqpc+g1VgM+DhUcpGuGZl5xE3nt+NjgHMjWiDGQkoAgh
//B/PwQb9GM84lAGXUV+agbv+yqYdvseupz4uM6HwIxoZiyiuarX7HIJPRXbjnkWH/QVB7cZgIx6
Bph9dt/8CtC7wDcXzwO4gnpQsGcuKU8ab9Q7/vWP8uYrfDfMEoXmPjbb++Uk8kX087hDNRFI6ahO
xDqk+atIw3IWXfdaluq/0Gam8+FMXd0vBj+YgHN8DOtYReaCrSNtEICcGFoF1OtXt3s7Pd3G9B9E
LryaOAfDqedkI6ND9sIH6mSVm6FCbJHwCXjKUUM4O5mpc3ICc1GnwFhQbgdiFZE5yx1OvkK5PoeA
Xs6E88p41XmpWWbGdtQQBNgvXamN50vFG30tzn7ABl67cbY0IUiOWMcVBoBdbjKAiYESn6vPubBo
FuBDs0ttYjGK7VgGKJvZRjlcJA+/4YWwc9jcB1JNWMVuKTi7kYl7KMOh+swvIDY35vFusvFsqdoD
DweRFmGIHz9YU3xYJyi1H3hs+sYOs05iqsQcqqyqXNsY0qGIlUX1nTHSTIXg2wk3ZyT0BmcQ6zhx
HFrClfoVyIqkxxuAoxg4Da6etrHhUVTkIKe3TOJ3i9KGapjRTjkVwmi4CCDHthjXH+hAcdjZa3KB
McW0yEz+Qbcosw4Y8e8LkGSlAl4uLo3P5BH3dgZ78i+mCv/zcEc3cgY4CqH3iT6FtyvLOQQ+jC7x
4B1zvgGNBHJ4lsS4P1fI9GN4S4wU5JW1lVH4aXpm2Mpid4XNi9SqZE5jCQgN4CYf8x0JVNMVd6JJ
T3lAD+TyR8i97vp706xCfGUEKxZiNwUBAeD5T2UndOXTEXZHO4FWRDhQVg3c+aV7L/nRiQnHCN2y
jydTZjH935xgF9e5NNLQyt+kZwMOBYR6v+/NPSW9yLMphjea7cthPB+cw3pkaNtR0QRjRThcf47f
fF+EuvepF65llX545oNxmzceoxL744NiRGPV9eUiCyLGgHAt35gdKc3kSPv2uxtsUT3f5gL3gFgi
9kcc442y8V5+wOuwdfj0sqMoCEAObqGfAV1z4cU8C5tjUngMDNbCtspAwIiFtDnEn6szRQt+9/mw
HBlH3IMraq1EaWtUzLFDIHnoWrt1vjHwxf5kp9n3yv2zsWqKwAUJ4wzKF+mJjsux0AAL0ehAZje4
pXNw1k9czkuznC2xEcT+UOqM0rX4QTwbHYzb1cHra1rSjCeJLFutvMr/Sd96qxoW/Bra7xgEJl4J
5VvQxBWyup9GBtR5qY3RfWutkgm5r8nCu1hv1D07V5O/XJkgjxuqL1ezUR/n6cQYyesrOFrS42t5
6utvYpUmsNlNU7+ordSakLFLMOwY2IAhV+PMm/orSDjf7qIhzkPJOX4uLKXp20Bjpd2UZ77zJdVr
jqFUk4bzvwOUmYxloNzDytxY4VYvcXEg7voWDcHVH7kPKUiCrQST0/P/MeK/O9xbKryyGmXxvwWI
s2n1ulM65TEAzYZV0ZnC0yzNJCg2fV4OCh9afBRJmPNY9ceCOpJ1abzPjmg/st0m0qu6gqO6qPjn
2JBYs/lOTGE3mVgIdiImXwdWGl2PNaYZaKVaxZkuf1sqKOs6psLDI4c9GxjlOLkYA43z4KXW9Nby
zDs1aTDyPS32X1UPSD5J/wPN3bY25UhVBzaG2QJqpEHAxNpZ9A4xiB642QnROJ76opg2KSQDPvp/
v0sRC8zgR+kkja75Cm2orWw5M+XXEo9Fi/VacQYTgn8jSKvK4M9udCgafkM66DHThNzDP9664psf
BJ8qDio/5G6CfKrZ/YaZc5G9nC7i+i6YYuWI9SBFvcQ3SEI5/4WyODbfEJ0p+BL3AFWwwtSX4KMm
Ci1wicv+v1XGfhBjgJEw7AX/fmaplflC1D0zxfupAZ/E+LtCbFs8YdhU8meQKR+vJKEtVRljYsm1
SLrtrIXvvOWNK6yEbj1qGHIXjDvlfEhQi4PRHzunVGVkFagVmRQzqK6R9hOwRHS1lcMRsYsPNndU
1emfLgb4A0EvsS+bWA9GQkEb16fj67CKLoZm063upM3BaXwvk9YEEoHN1owhdncgbt6xUtdWqmES
JCLzNV5NFOrlyyciAzUnioUXK29Xf2QY3v3+Lw6JAkHbydX4hualaE5hy3S2jHLGZh2h6Vdio0cS
PVaCx9qu59cDcIPpKAvV/96M8ajWt+DsYTV5Iy/kpgU9h3Q0QuCK/i1dwQAO/g9EBcXPpzuatxJu
R4ahSNWRXWOIVptlUKicaTrfkGEMmDKrnG0tsjcRJE9c9w34Szj6GSVMmkKERIIq4IoxSrYje2pX
5Yn5vz7mM0QxNK3Xz9VaCMmjuTuaFGGtUNAGie+Q5jZD5vKy0s+PqTJj3GCgsMWzM5Jo1yc621iv
hpwASaBTje7F138sFWV9Bb1nuhPBjYdRabFzM4OR43c+gJtKW8pxza0R6VIA/NrcKegXrp3LxKbE
8bgrPeuKQBHjcJYlQluFlWFZhs+SFkbkHP2hBWBt0LrMKwrB+WcGU9qEAd7iknAz3vjI68aZ7/Vw
rh2dlCf/GS49WtcPOkMr773uDUuzYUd04dvt0TBSg3Tz+0XnQX3g/X+vV4Wg8HzAPBuUsPqpeadk
mWv42iagYnqIHwE0VAstXJ9xOY8Ixf1Kj1VNmZX8O3dlZT4cce6zzrNbtIui+ywKCFQJR54YNxU/
J88pBHEc9dLfafEIagkflH5+KVhKUgpNYw7fNkGXqPipeBoL1BLkmr3Jrm2uq0vlCz4itXlM7XNE
/oU9qQpMuJM1NkVe6eBAaGrwxhuM5q+hhWSnhBYAFoXIs2msqJt2vhvIMQl2UGhH6jXw3lMPIT8h
IfRCVAG/ZuEzGMrGtVEQ8dIg32pagRtAFudGGJN/Ln6As3BIbyuJ1IVQZqCSPKa2SxSdMbJMZ8Ij
KQoPpLWFjZSJDaAEcEJMFts1IWaHnKLOiUjb/2RaLlYLXHdQ3IkV2jIl2sCPIzOoaR7olPiB8Jeo
yqx8mdQU/Y29Y45+X+DDQqKq33qdGMTjsrd3GnarQ1GfdEROLQSdHhT1HsoSAiHMy4zWlLUseONK
atckWNtuOkcjYOk40XKcx8xRBAinpXN1qQjfqLRgsePmm1boWkqPPpl7OewNXsGV02oTVTcVrLGS
4Xy6dbGAorD6yWRGGPj7JFqx+U21XB1fn5o6CbcpR6aQIPOfMkrTEjdeais2etlsqiB7U3QAE8Dp
R5qpB9yOOv0i78gWjJUJem1a/xQuja5VJQeHkDFeCo4MEx4PgfQP3IhJTvVjM1E1IVtMrUjyJDrj
nDF/PrdJlQAfObMO23diUU807yON4V7QfbvLRtx7c117DCyR0x5dFIewB4/U7bV2/Se4SqhVPOiN
290TFu5jCOqFTI8AGIrrTTf3D9vuYfYvccUDTr3hBhqRf1/huCu6bGeT8MvP7pJ0zz+hGkUn/MV6
UXb7tRTBlJGKwC6RfwdYr6lBe9FE6/IKYhGo6bLd6YBuxeWxGTx8ky4XoIxqLqiqRskwck5QbCqK
SdA+AtGgDgQNFl4acuLQasp3zTcNtnVtNX25xBqRRXr6Af1bfuOCZj2N+UbgWKOzNJOQJrmkPtWt
toNQOSuqrQmc54vIs6sslNWHQ8eYcu458SAeYqru/PbWR4u0MgHKqmeiAH8uw53WhIugyN8dO0tU
0wNFwR7+eOd1frjfjV0dUuDkvQkG05JGdd16aTdJ6vZ1lR8uNEl8FbDTyqc+wiKmGkTZ0SwOqm9X
o5GwNYPnig5FAQvFQTfQVmnKmqMMdTflHSX+JRaBwXSdw6hFtmP+WzZt4BFClfScxunG4aBVOcFC
wqP4AHwHth6++ru6k5DKbX1u9WHMZlKYztzEG0zeZZE97OOojElqMjgh6v/9/2qVTtvTG2SDW4iG
5JkHQE+F7K+6pjP3blzZhAHH+wW8bB+ESGsYHemn+0P6MP9jSfdQJAtcfItlODPbOlMyR5et6uUV
jdXZYhpWLzssCtXiVIg1VKt+C9hALHjdo18Rwu70MeWq2f9jieDIqxDBVMtFZkv4lYytJMVV6QFS
gXamJxQJySFwiS4keQlIjMVyox69z3sCSGPQtlyF8fyA/ySS+KtlueVG3ICyYz0RnerKFuc9QPB3
u239fWuzWx2bkJbiMFM+lnEZXmHzSmsZHdSIpI/Oy93BItRqTTnfy11yl+RvEe3Bnd+4HlSMmaQH
/G5+zMsn0zWwmGIZvYX1KjofvbG+alUSRTtLGEQYi9WmBsoYV3yJmt2hLJMA+tbcIQtpBWwjQH/g
5g+JvgJNF3lXCQ2B89/OreKelUqhY148RCYzZYqlTPpHl9Irg7C2IHdRwwyabp3EhPu5HPKl4g8X
kQdPf2KneXBgQoSIJKvGj7NGwcRkwEbjdrtSR4df5ZFBMZIBWQOa4oXaclSjNguY+Z6i6D/HrIXM
mwrKh3ysB7iUevd3Ys+8VR6AJVC1bO3/sViAx/NhZMzPnlqem9ge+Qx3+pgnsiXw4ozEqlIK5PHo
WPCEx0PGqMr3DAQwl74Cc6albA899G8kr4bpK9POa8F8juHSWum9rDEFaj4q80h6G2HQYjmXN1IP
71++ZVMGTcG/Pl/w81utsGxapOQYtBCHsuibyRNFkze2ujKheUPhW83gzojwI2xJB34e0bY2zNik
WZ4jnt4TfdD7XroXudpoGnmHEnLBXQuR75f7I4HeA40B0buJT1d4BSXcl8ujIgvt8iH9udyv3pyt
kVj4jLYuCGpo/an/Nl+zX1wUzKiEsEPSEYvhYpc1nfakTwzxIpnXAt2eZPcygrw/ClmfyZ7dVA45
Hp/iICJXKBZEpVWcNqa375n5qZL19YgzdtrIsKYue+lPMNf2/Qq5MJjLSDQyBOdjWnAnaryJZL31
a7X3iLSRfD9sMw1SAyibDwACm9WgLykWCVQWzfOUWl5Wc0cP4MGoKm6EDn9pkyP6rP18W0IRwowh
XPyhjVUBcfCyMlcCYF34mMwjzBcFmVux2Co6eAFXDQvgKioUe815ilpDB2vxuC5BxD5dvrJNfd0Z
3V/coIiHvA7CBHJMNS73lCBUUtQccB+IRGaRLe2e5oUPDSQptDysuQBxgKnqrjEnDspK3Pf6mKPI
1IkVamnkqj9DQvXGfggmGVXayvZGBUH40FPhyLvFqgZVbYCf6jUBTP6TtqOYTOnMh9r/Loy8daIu
fl2Rn12dFmirKE/ydyJmU+MbSNf0hDlbLbMNxdqWGvmI+xQ0GbuUDSPufZkRIjnHI0n+4RiNwnE3
7x6AR9KuoTTkNIBlT3L70F7Tn9vRKFR2zRwEjeL/bw/cx/8zFU3W4tm0tJXZWxP146wDzYYPwEXF
ihnU8M5xgKMdOs7xJYhd+MKBBZ43PuBIqwPf2cC2Wn9CxII7MV1JGDSofXxe/vuHMtT3R6V6ks1A
guCB5TathZ4zjd1IpTm9JK7eSeKGuHzP1ujvkJ+QLX+QvNs/uplR8ykLRtysxkCh+uq+SB8CmrNk
UWdozHSXZf+o6PwF1qGOxNeVJayHtXKp8QGHmVbEkToQK6qd1VH49ni+DEH/c4TxH1R+VXX1k3W3
5jbGPAHSDmamRSfSkKP+h3FyH3+tQo+jdEE7LbNrfFFuX6AL+oj7DDgdHscReXJtMppZnwCExoe0
4QQPl2eL5Qtv3eZnT5U9Ky1AaG7c++rzt7FMsyOoGvi2MB/ESJn2UOkMLIxISv6mEfJdOJNdKgNl
Rb6CyQBhq2q5FvrJibEDoNpEMftt/QQ3zNQKY0yFeSryJn8FoRO0uPfsC86Kn/enCj5EZQpUnVaU
AQK47Mx+q1mCB8EWyQT1dtYXbAWuDjplXfVkL/VPYcZgvuo0Y8qI4iRNg1DZtrpjxQh3QotKVQHn
Tkhlj16EIRqlKLLkasmjjTrz3Ud81pIlPkVqa6rguxl1bIvyWzyXy2Krn8Pn19Gfxs1Id3ETr4sN
n0dpjRvDnAoFhVG5aQa9G9mM/Ci/nFXnBMTyzzreqfPdiBgRwFT2t9TJw1t2Y/mgyaSsiWFBknrH
Ld+m1DDRMLsXSolZPqq+FHf8E6DBw2soSipL6LNYKIA+24lCMd7ZAPxOVRJq+214MDf/aWC7t0F6
3dskmIV4sPxzx14ClypLZkfcD8HgO8FMPBpUFZkLclJyjZo4Q1J+tpSCBXXNpB5STOFMq4h6mYgI
IaOrY19HcZan9HM/m9/zSiVjjs/gi8a30ACwVvjA/VoGj60JRbJrjU4n6F4j4EcJ2NAkKtAFuSjk
xDfbNG7QgpbrAh2Uv0gfa6WcypX7z8QQeo+rEocYCg5nbgdBYekJa/Qa9adlF5CyoCwMKtTXLVwY
Of0iYYTlll6rNJuENZj9We0pn2qQx/X3ZRI2onJq/1yDU3CarGLRBSSx3xhx+oVUp8da7TfNbQpP
F+STHn0gi+j3LMvxWH+xoRMkDCEScQw3l0VitvZV4D0Mk3aRM7gQDN9QMldXETMLLsp6jv61jy0h
+RLod50EnwBpAcr48cW9Ba3YzSyluP4WEYbwL/DhcOARF9KA4dgE4w4xalHfECcn6FuS2dX/g2Tf
Hdfr+hV8SJMsYdNGg22uQAb/WlOPvu31OO6siP5qyP9GxzWS0q1g5g3q1KHcf1V3RsOs9zlSAuNj
MZCjQrC/V1MNZPRmM2HAWyorLVDvD9gy1agG513hE+xXrk7WXwqwtC5qts5y2tcfAlajdTauTnHV
iJupaVNuPoCu7Ua2adTPEHL9EyC1iWHRrxxCgPYv6XBbvaOWhcF3DfC2wM87H16sNP0gfDaxRPsR
Uue8dUohBMf0ukh9dZ0GtVsjaBIREBcaiVr4Aj6NojGdTjy+UAMcdxr+aEldBf9Aw0R7voVcjUKc
b8NFA+uTA3bzJfn8gMRc2fkx6zCI73OUPunN6i5jD2nI/pgRLDF8gNhMA243CJCjLnZSZyFkdXjL
PHzdmiRdYz3DDFeAVvkc9lTm6Vf7ity900Wlf092jHFOO2Ace2AiLqiQ28aGGNj0JoMK8K0ph6D0
B7V3vLEXqwe4tUYUy0v9G83rA672Dd6wdF+DahAuf3H6W5UWTi4gJWAxHYwLvFhxUVi4N866dHjn
Etlno4ggmIfYurntMZiCvVXpZeTV9hKNx96UW2c41E958QRuvrduayHfpRtwjrZfrz9v5T6Vk3Td
a6q2u4YAng5RvMbDd9ZvVzAXA+znXLaNYGJ+8ON3XomI6qx92U2B99cqQl0Drs9a+A2dTELjL6Pb
rQHVIiW/o202xWVvzBvQ2jzPlEen6iSHUkUkqocJItXPsP+NokDIyADFd5UgNF1UrIO6Gl+yVeDF
AMycbWrX30kqMbeTocXE+OfIBv2GpLlWvJsNP6VxavRqtjY6z1tXH1FqYMfEJHgkqSHJI3xxsR4g
y8srRNHY5d25ilkARA1rBKhwMh1XhatHSuxWSMfQaBadcxbGpdj6CLrPZDFzaz5KcM+qZdrDCcH6
ir/WbIdrtmA87DXiv8Ewa7RVbcQ9TePQHg4nAPpSFfCLizYxn+jrOC2Bzffzii9Pm5KjjGgT7gHq
29pjnJpioLo48DMBx8uLjmuXTfFt/dFLoxoydiLUkGFHUR38mSz4oJk6OZNr3wdnRhcZ0I6xuUZC
MO52LpX9+BIcSWW4GgmwQk0S36YcV5FH+CUJhhGsZVfPWxY8kZ26vO6ZWV4az0zj0j6sHnDV68vy
yfD37j++fVgfBSvfbqyXZcHzBf6gVCkyfP18urv9CEvecJbBRNXvXFA94+L95ZRWh9JtWX2iRhE3
7wBFIvWXaytNQbcaFCPfcwHCyV2+geExMMGX8FqWSm+LbKCsDKl2MLu0PAyPqrJlF3RAOV3X5MZx
STyj2z4RLDj2oKdibRPXkVEuYL7xZRu0FsxVeP9WbSdfZaKFhjKIT/qI8VffXILMz+14y047d9R7
X78oB2tn+3NaeeOFSx7SSpHTCRleYoFZkpLXqoh+Oh5bLri3UvRmFigpDQo4hf+TEPKf+GJLSR9E
Ky4Tvm+wKfVoiRW5lqyl9zUUBAa3CcNlaZLJPIzVcnKqKuBcKM0C+1X9OicULErqs96csqtXXMBb
FhpPPOZHov27wkdoCjOc+TZvnBm2Nl0njQfC1VkQootpfa2kwdeUVKhLnNAt9uwUhDsMXb/TtQtm
H5Da5lXCPPaI8dmPNpaXOLNmprV1C9KfrufO89t7JORZYKOAZpVV9DTTqxLP9Ehoz/E3aKRvt8HW
2MxTmkAewOZJADv7ACvGliIBdhIgUPc/7kMU4fDP4CVbNkzGrUWDf3EvKjNxDd5lDUrhVbSrx/m3
ehOgqhiDUwtScyOxGl++Z/UcTqhSzc66Jw/D/mihZP1FPEPynaP04JTmL5P+ihFgvk9FOZH2xa1r
v3wiYOxhURbcgBY3TG4H2rK8T1E/ZJWVU5yNE+DUWW6P49xeJgBKsjswNuFqcewpZoBvYQaf7A28
ECNePmaYLYKuPwG8zrFEM/dny7WmUHcED4OVwMC49PDn4dLGf3ZTep0weNOshxtDCN5fzJa+gaLI
5qhVCV53ZkErF1KT63MU7dm4aOmrPt7vQQEgw0x+SxqFwPHphrfsZ07qkvVHiJQ+sx/IKCcV5eut
0CON5jVnbgUF2ddE5190dSqHrl/BXgVJ5OmqVbsb/NiSIAbqAT0Dyv4uPINxGnRBm54dwXmG+QK0
/Ynrf1PSOltkXWlpeoO3NmYjm5RKIWeGSiHPHmHJvfJBATPyXwoX9Ujsal7DtCOoPnYqJK6W7ULv
Iun12WOwsF492XigqIm65yfj4CmDBpAgvJ2kov4ZQ/xHKiff+TR4AytO/FWG1RmsMYcyq/h4yUJI
48G5s1WLIlvmRxzmYxlG277x6fFcsLCD8A/6akrsB1hC4Twc72cGUQdSOUz4nSrrIQcplbxXh223
lULWJMbXBcBi6MMt7WK952bxaxmc6YXDe0emoi9jI+jgHrMmxJxXhW7psFUu6fFtgm8rrCFstR7B
iyBqblldZ3NyF6PGNFut3SGsU+oARZSShdM5HAUkF5gBsWKzwDvRg4Y7/+4un82V/ZDp4kV9pW05
MzW6SMqaOhS+Vdw7asZ9VxxXK3cs8GjpumEm2Fi/fnTfk0wqG82HZ6QADyL8VkY6yimhG58k9/VR
1B2WWmr+MZH4LJ/mxhHvfhebKHTFDSiDp6m45ZtkrBk4R64vQCVN7kRARx6O1DI1CH7m4mPshMbg
/eD3wGajg+O6pMk+43qgNxsrBDVs/Mz4DPVkP6iSQ0cc/JZXtxAuPjz0mK8urfnz/zS8RkGH2Ixq
pqCk6fnrEylHjM2KRlSPLf4MpYLJO7+OQMl5nyxQqQkDr6wwQE5jHBVAOy0bCSMojRCdCVNXPGRn
NFRKg2YVmMeAw5iIpe24FZGDBZ9DvfcZ2WZisYJI3PFHLbTaiP8966qCOluZJAKFsN5BahLUo0+N
BIRb1+6ye4WLojJ+lQanB97fvvrA/VRYNJ5PSfmIKwx8eCFcNpncsKQqiQtGlR6o58RPRz5fYZu3
sVA8iWK4UJHXxT+FwqP9CMzmY0Pi8bPtQgAOKkd6q9N0jREIyEKEfnzbEy8fkGKUXDkwVBihWsOK
IGsFNRXhvclze41BTMbTZ3dlvKSfl8LkVAyloeeq+0v90wF0m8bBArMf9zZQlzWSELYgUJ+qj7hc
Z8t8Uz/QPDWa/shdbrOnua80Adfq7pzO+75ppLVyb30iQKYqSjDLqMUmEu1ZsHLBlxWAMUTbrGnD
vO0EcQYJ0ID91ez0Z/XmSIKKwB1DugdJcTrl97mVS4zyR3wdgsjn5IFGPQCvRDQuSv0lBoEwfLjc
hk4ezoorO2Tw4FsZIq0xNigcR9Oemf4lYyL0fd01bUTrFQIttp4XgjlBsQwyLHT54DIrCbi/dIh9
SDkdU+fMWbsPfo2GD5zYYY0sLm6qkyirW7uDTK/B1SN8pIVepkAjal/TjZ30QDGPAvR9+Q7RqkWJ
5MMc4ENV5zsrp2RXXQqXQtfTK1oSUrMr0PwPEzZXfi2o/gGkzvRZLexmUgF/58o5nIrDBSQNBnlF
XXCElthd+BNlZZRZPJmx9O3IyreD9/uLaihjkvvgLI53eZMrz0nVA/opH8JJjW4p8wZnRCmkei6s
hx7ilT86oE7GQWUH9mCoEf3WGF5BZRIkTRUWihOzfcLtb4cwSJvh9FG6JWEVwuZzSO7rTfV2q1xT
q8KnHu7quC1JdzYGeQ6v7qBR8IsQfq27iq5pO8Na/qoR0vzKUcZfHb8ebz/DnAMALL3EeekKiwOE
4K7HYb03FKKV8eAy/GiAtvubBt5GfZMHPKPlf3f8eQDNVT1FCEMyqJzvQMY4lwBGrsc6lDoUjSQg
6KZ7TElNAdDelkfz5m807Q3D4LIVbsTBpNh7W94uR7c8nfSgP4SYPBiCSjQ5JMa4PEPENNwHbBIr
YD8JPjeab0um57lp2YVFCPoYiWDdqCxgnq3EzYl9KEQZl9E8GlpNDOqT5w4eiBIDcHKvX5ta1IRX
uSy42c+GQDvq91yQMxO1klqczExGfOZ1BKAECRwKmE6VdYoZvZERtjIFgjp2oIeikgqoT3h7xmGN
X4WoSOa/ahBtGenoCySk9bTD9VSuVkhqedP8jxQIrkmFZ6DFBO3D8mv05ovQeaaD3HKKYWRnAgmx
gLyv99fuJzCaedPaP+hmsCyaNYlquz81+2cIDqQuSBpYR+0yJr1jvr8+Q2YCkBxppfiX2hlgWgru
fSIrnUIoVPcnbRUyErUa5Vu7FXjcuSs4gwZB+tMtltoa2jNDv7/vCrmUCCAewWQCex+WkuLZ7g/4
n6qL6JW0p0HQY6UbirQz7i6dlRh6udj8NM3qPwtbdjfARICyEB379pwN6Z8eeCPGlDarPnRzIJ/G
XB8TY1Vj6bjRph3b4jUfjc8kyiRX86h/sg4C8OZgpfBjcHu0vohhE9n55UGpt+SeHmOeddwUTWo9
OcfOPJ232twFePrQkyjwnggw5OYrNxKCi6AQcB+neWt+pBQ7/3EzKgGsK8bbcXrLBmvYo6TSv+RO
fcdjyIshd0sZwVCrg2liQhZf+Q7bsHW6eERDlMDnnaE1RHw0CvIEF0hzJk8S1duU9rJNclTVoIky
K218kVyKnhkxtKVy6YnjDQXMpiRMfBPghWB3F4fQwTPVKBRKePkeP9A7XI1t+sXo18CNaZS1aC7z
Rziczd6dFB31YbKBCICGl2HCN7akDH4iB3YXU+WXjRCgWtk3D13T71Zz/WNgeidC14iWiqzITEo0
OjMCHPFRNKhwslaG7jXF4uUoFHvI+phZtpZdFSLXRw2R7AVkeVPKZyckUwAxMtxK6fhRYKyqPWb5
Om2tZzPjlFczrWfETLKwjLuf4ez+3gfd+rK5ZwhYuLmcxs1XMAGBn1Pro4i8nYCBOTVo/2TXaSxC
aYSlT5YC3zQh78CL0gmG7MzXt3A6IzdHzj22ipLaqn4PRQ8fzZL7hWjYZvlBHS4DmWKO2uX1dhqc
TZgvNaBMiUXVsEbVG7e0DviHxH7zxi1Wz0wde72y0ok3OyLwlFFm0YDlQyhatZw7teDefLEiAdp9
r7azt4JH1e1l9EtANZum5fYCTL3TUzySczjLNgqmTKXFF5P5RvqIG3hWQXuUmFrpyj+OKVQENDKK
65L090OwCMGlBtBjYgyEkXAKRtFefLTCCYmn66XDlmrj99vHMxW2xM+E7/edODI0qck1bJXOJ2Dg
i9hVeDcEGJJ9tQ347thxcsqWJfT+AsbXnNAkl/EXCpWNs2L3hr8owRC9H6ClKFrMrCxiivMvEJp2
b2Ob2zR04rYRtPc6JJyhfjLIcp2H9hvuNy47PLd4NltpIPF9yk+jaAREIDStNZkkgX2ZZJHmX/oC
PYfXieQNO+54D6xfH2LjSYd1wUPMzOdHDGv+ASTpDIf+1wK+37vR9caY3bdyoCtRL+1bANZYM+iZ
kr3M5Ua9Ch3HpKkNy2Idzg5KCnjtOi9Bxp03DkKfCeLLYm7JBVzW27BwYxU0yW4voi8Cu0TeUKi0
xUckIEG/vanvsRe1bqaVLlsQeYyamMieWFKSdEh5JvTiTku7Ksi5J58mmZtcuMsUw1QajXhvZWPI
s4qyy9adURWeJmz4PLrd70bZkHb9e02hpsqbdldOnUR3qxIudSeIPjaNvb396IzrH2K7fDQkKPt8
Yx3SilpQ8Z1O24Vn8wl6tZ6Xv5HcNFI/J1V1muF38kakXY6rJsMXRBZsvYJRzHgVxBmtKaOTtg4b
pkVMjZhldbDw5xRXfxNuS3H1g7NjTmEbpByQNwqJdbx1AaUaKNvJlkNHzGKKtv/XUMRzSMKDczCc
U1/OEwstpaBXnpimPxc41GrC5Nj4oNcQ2Vn5DXog17N9F3iF1oHH28g4H/v1GSDwkxA6PYQLDhdq
YOTq5jbOqfzZzcmVHX+g+BiU2EHVPlnsdiH7lsYty1DwbX+93upW7EsxIjhmzLjUG3XwssIJKB0u
bixsri522493xgrxt/9nTd3EzYlfCG6/XHOoobTx0keJhRK2IiYqAar56jJXGOsq8MoaNrKx5FsT
LHw1T83/9HSa7K4SsNCa4AYtEfBTdyTITDQtCi2c3WzIauHYBvgP8QJEwH9FsyNIIe+fwL/BctEN
GAATn4AcnM+GLS6pXkf3wJDRSM36wuG68NJcfqYinxved8sNQLtNtVKHk4yTKWn24wzpCT23AQEO
JzSUhuyYNEbfpVIPyRNkXp3tkmnSPmcRahisiJISScAwsCgwtAOKFBiQCplrAp82yC0yCHinrLWt
2GETzPU5bldr3p+9j7Yqe7ZhvjoAR2OO/o9cToazdI0SXZSo37oX8rjy+hyCG8DeROiwfjup79hU
sQN5Ok2l7zW9w+pV0VwJbj7ZlQtsurIiZcbgs76jiboTlSWdF0IlmaECXi0zgRNCdF90NpOz8c5j
oO1mW84pZ1G8Ijvw6MyRCJVZOABWOQAfp6KOsJ6N8nowVAIa1/ZYS+63fAPOfPGvY/yLEPUx1LKU
WBcNapnXT0VwOd+efvIZuiSRv9MZTjA2D2p1O5VM+2mj+pO6PonlJbAws/I/8DMN4QO+Q3i7yBDq
RzqwNS8jD6XM2x6q5SKtbVD63q+wcCFfii3miMRuuO2s7gQW9/gL33W4gwXUI04bLfj50FtYdmyV
+4d+8Rb8p2vBAqVp+WPRx0sFx0u3gDUedUnfvCKUvjLw9mZZJYr96+oBcUipK5Rvs4L0kxYC888a
8rA1pr97jh0rCQOEghg+OJXFYF5mrbRPCz4wRPx46Mh8IExzKx/ALnISQ9X5VxKzEDguu6Ts+fov
jQ9P7HZW02pFR1JdSipFupnG3Quyze0QWNjXTfXSf+v4leAJY7hv0cK2J/QuMr5Ee2TReYwr9eH6
5UHbRZjBreeLVhIMUse/KyCPw0MxV3/32ipnE4TiMOdFleNiOYTq/9VcrUfd07da3d0XzjgZHKCG
7JOViu0yuJ7pIqzI2y+vmaQ2aCadZ/imRk5sjp+kpNTfpBI3/YE9KgoszpZivPVhBzzFjbpoPZPY
+9c8Kdt6VBYuW3k6t+CvPCWmw+sWdBMyqVaaQSP8y9Hxc8TIPG1yOucBcUtmjdYC9iq3P2K2R+cw
8wF9YmGthAswP1QfDReMgxONvAQOi76uAGi2jawVX2wFxpifI2oKv30A0jY5URtatlDXSKo97Bfv
ujMgxAEYQbuhyz6whM0W1pZwOhsYYzJwoo9Xvc/143XgUMThe4DM9uoDQwucAJbD2wopx68+l5zM
zolN3hO3PnnWmiawLtQXjNl0qzmCDanl1Xj8Z/9fPBcauwtwVsjQJmxa1Qcr9Xql3D20/ihknm9I
TCNcWj/PGm04M1PA5JWkKl2KEkC9WjpnU2QRuFm8Kxox+wC1FPrE2WAz5bSedgQO0uwT2Eu9HoNR
qAFHGx4Mw/oSs/76DblvQC2qxADFFIlGNsDRebKKvEpu8lyId67676byg3XtAf9TrJW3/ARwDyGH
+6tekCgHX5wskVXPnbkouNqlPOQa6RPEBdqogCVJaxRPRqLXVMLQ3dWRILpthzXX5YofAvkR2YkI
79GP/5pReLxwB5oaY9p5vpl639o31QJn07t916yoyj4QW1PEkrbJCzZ9JBNfpstJn9OvfPDqEt1B
NSJ6cvqYbNZX+Doq2mD2YRwM+QZalbTYvs/7FU1l/LZ4rbm9EgjRLgE8pQztQBRthUHlV7CNRWv4
reeA5ZUJLsbb2ik8R1PDpu1qMGFzITTfhMcsJiAX+a9Q93buE9SKP+SJcbZbTX9+zhw4dPymuNiV
3ZKfzbHK8xmh5oNaNW88eOAdF9EHBdU799qwwdjmS3GI1WnBDozvCgBRdf5xl81FyrAVeJhju5oY
EbEL3WLzei8TW9ut/PS1tVoyJdFNweCZtfQINLFnGH4lGEZ8W+jamJToFpMjcylRXwk/RYnH2eJB
qkEdbVp3vWc++3oKOZtyuF50RcOreItdxsN6Btbji85GoKk/ml9IseW3iyCzjE3y5aAyk2aA5kvj
b/xiiEvPuTX9oIaFiEjAFgHtdP6tN66XFaIK43VfdNQqk1MJMZExKbRBXAJ6BvU+W1rycPqSjfdf
voj4cYSYktmlGH2idhf7xf4ML4Ii5JsBxrow3MwWEAoLBrmyED2gr+cdre2BGCxRktSgfcVsTNw/
0cb0pVXkUV37t5bSb6+0sMNwaXzN9aScXO2+yncPYsWZW+1OEnUVo1IoWlCcz4iiI1sWQ8uNjh4V
Irk2xgG2iyjny40VJfiI2rnmv7n4tHdo68uRx7Oc3bDNqAuxVEuDmMLeS4vWMu1m57gmfvWOeS/G
op1jmq+bSGxtoMfkJFoBwFmPSCYvM2Bmt3196OuyxEm4dn3viKPlAfCcnok5wM+63GEFHLY2DfDR
t9hNntDMQzgysuJaPPK6IcwJKIJxTr644NO424jCwsePpoIW4Vaorjft5bbU6m86Ablqws8KEBJV
S1aex+IZ/3alWAM6Ob4Teq5hnFHYSFnGfH/hr8kV00dLK+hbWkKw0bO11S1JoVitHU0b1Wk4rY91
1hHjUnxlGRUu9j5vJuq/FoQLsyfgXS/a4cJb7k06F0dtHDkB1O9ZG/ivr7jNhOGjk9MGKTxbbmGb
6OFeaMXYKDCR2cVZaNd/YnI1mWr8fM/OkcKMRvIYt0XVV95zSMMjJDhaxEHIiaBx3uMHqWlZFepE
jHpbS28IextlRSDnFX+jPbmGu58K0U3eO8OO9egVvGOiONcLoqqzGE7M9xjXj90NBE37pejDhxkG
GKlRBa5VS53xXhtxuKFyvqv/KgWgKMwcMH8RqdrExkFbexa+USR5wEMXrZJHPUh4DE61f0jbDL5f
eQZugNPMzTkBkMufGRay4UseKB4PK5B8zmMbMfHiWqINS9Olory4A0hBRh3qqBqAwUQdDKSseuKt
pT9Hu7hGa/bC9ZtQxDy6uuCDyo5w0/XCnVHqTQZri3y20ptXHcMojOT5u99sPuzfYADdKUflnxpa
YoAVSv+U6gxrsD7MPJepoyZdkuYjwTYKiL/zstZZgqkGQsUq/uvhIkx/uFZby9oYJ4L8zdXQzn6v
GYGcyfze6jJontCfAJrhEyjvNdVHkBs5ZO5zPlLFfVQT/pVN5opGxFUWDzXJdsnRdlHX2va2UbCk
03jCtseRdlidDsjsH0ruLLxBOb3BFnJjM4CipJE4OSIcjXp4yWBNuqRn3j5R9WJiCFx+k8kfKfko
+yhyhI/UujmDSVCNRHGaxc1CRN6nfX3ph9iMn3cENznmQDMG/xziQkNIkkXKOQ1O/rHke6KiJHmi
kGOInKF2hAZfoNpKY36N9YhEoo9mt0E3Hf32RiB6GRTMYE3Xg18pkSdXBJmbm7uOTIuTrBrkzHz9
k4ivcyoTUaEf9JlbUsZr0/3Py0g4q0dPsXritVdx7C1jZvrG9aOS9kV/OuhwLFihuwoFZOjZuBge
92XyVk2Z2slESyf6xxAAM7F7RRiPQyLdnp7SQdz/oO4vTELGFBWXmRavXMpXCj7ESz0iULteDl6N
OpaICUJoHy15EtiJ1kxH3RnVIkboKteehEJP9CbC60duETm29b9gO8g1AbnfyT2gF9Hx/MgE51Rk
7l/w9BZUz6keyZc6/n0YWLrCcuV33xjVnWFDHFE6N91Vbf/7oyiHz2s3ugw3ZuSezf9aoVkVSjK+
HVohzgTuXCcpSdT6mp9E9uq10N6foyJPwr3BE3Uq7I/zIvZDZ1n2iDSfzWURTYGtc6bZ/3Yqh/3q
t9/WMr19/RpwLOaPh/VmnBCSTgG/Xf2tBFEVQBK6ZuSMc3Y0xZbETMdRTUxKcTPeqYBICWHG0z+n
0lOx9FkllchI3sSVdE6MetpK42vbeTr8xMSpzVFiUFi1DaYDULODe+mCTlTfCg6+1bsQ8cJKUEMn
dyiRsVqmDJK2l0thKkpIABu8r0US4Z8n8XxWJ6SfwyRqUPxwK9lRtNIOBvM5UJibK78AnYjL1LDm
6Uf+D1ns6gzEKphApPzRmAUJb+jcglqkqyPHAwA+h8fpYEGS5Zdm+Le4+a+BpBP8tAfYTAA5cj2a
DG4RMPOJyqE3bXI2K8cHZRph+e6onpMtaOeBKdxszSDNWgg0XjG4GhYjqzjGzTer5fN1UB6/IYKG
smS/vI6Bjx9Ul1Ns9VRdVno5GmrtZ/LiAQMgzFNkA3StbfhkBEvINyXQywx0VcrQgaPgw4ot7vO8
OCGy8W2oqM0Wd0//w44/wLD/YLJ9cepD5Eip5dThQXvNVA9stKbv07GrThCM9J++BOfGoFiBxabr
pbYFNINaLgf4DuSiokX2ewIjMcZ6w2BKlbtMQZTARPWFp4FISdg7249VpAXwRbuve5J3V8AgN4I/
a+Y0fivyFmiMWDfQQ8+vtpwGnh2/+OmL3O84HBZn1rlQ3TewGyeEPH9mAvoR9MNQCyUzQaftOXwn
TFvlwVOrummIyb64rTqxOIfP9LYb4jSQWlhVmANdWfYGjAuurx8fUuIKz7wxCM7HxzPkg9m09ux0
UToevycVKwOZtqMPHCDyaS/n87iSajSig4T4i3Kn9dwD1FIUqwnwlTlGl5e/PxUlb+bFv097OWqn
mTSua+peZ/Rgjx+OCpir/TquD499Bn+EwSOu6plehUvFfEdrzjTfMbXMXBpQaD/7edwky6IfsRBW
QkLa1yuQFwaWGKZuknq1VhHs2k5C8KYsL7mL0+2UPwaHUCwyt3TJzmC+KTsdto84F5U+Th4S7ZHO
41WeOGUWuG5WpdMTqVPxjyKwcaBRMt5oU2uFkEX9LAWlcZKTpLxtuLMMvj35H9pAi2nZe0e5djjZ
ZerPS4GcuAWICuThd0UTWaDbcZ6/ineibXz92Do7UnK+os2z6psjYgihkvrx6uI+xb6BkYCNQkif
0Y3f7FbZziHXg0lexP5ZjbxiamJvvPg5ZRj0kEtD/weoYdPlwRIeLM/4o0b73WGi/ZprhfxbTUAZ
hPdwGF3Vs7dzWoYXEYkQA7nwVJfiEMyZhSFtIZAgnJICxCKrF3ynfJDEzo9HJG4dxT1vLHeqw+ho
U2qIHi24ClzcOPzXcmYMoxlLB0oBGDHoF6WF70lSh1ZbHCcjUpcIgr571SPbB2Vu3TrEvXbyh7e0
rag/AlfeCzVAK94BxntvgqzZIZOjOdHDo/UZkrr+gUMH9BtsjhUC6LOxNgUj45eFOoe7ymyRqsNG
UmIglHu49dDwta542Bt/OPpgeSCv5+gfge+MFWx6y+tMcv+3ZkwPU6oPU7rf1cSkCP7uPgT5gx+U
1JQ9f/mDtBVt3duxUmkpCHDVvaWIPAsli1t/muiSfogcUDGqrm/AWGOyegGRQLJNQSYcF0Ek0jev
7vQaFOGgSkML5EeK8VJ2TlxhhUOxnX03H3zThmYRdQ/qwdJj2dH8Fw55OgyI9kTZS9DFGXjyQYSz
YcfbAAi9MHY6N/HmnVbtygN+iG4aw+tDWitOa29iuVs8dyJeCR50n483sTstA9GpUA2Gk0P+pYaJ
XI5SKLretYJhrZKkjq8fgCLJ9JFoODksaSAu2lBqdEgGA1qRr0nMIK3wCKZ/A+vziPYOLakf26FF
NEwSDgy7Fg0lGiMdGt8uKtnzg2KvZwbqyjL2eNArvZuh76WgBfc0towXrZTRUXva1GKqJSJvvbTt
I3vTNKsRvIEe/CZcpCzqut6fxxuTgA834NSDEz3zspX8SgIHt5t0Ju0xC+WqIKlktjnv9pEEBQxM
MFNOnKYcK8gs9x2nImYmiJEsqJ1ZNJ8DPx7aiSSPd7p2hPz1qDfurp/+Vxvfia+Jeeim0qniPWhv
lx6Mv51GKi9eprthByHCDQnsT3f7xlRU5tnXv2wgApv1jy65aDA0mnQSmI0jDWTwyKdkt4Uqcg9b
C02UYjjrAPftwJ6GTl58DwLZFQ5pBPBSDF8FsfnPDxhaauAUdkRZpSG/kfzGVF1UOvsIA8nOqE+Z
H7EXdgfrsP30gDEo+J4YKCWMZbtT9AUzqjSWkCINZDv6ZvRSMzkCNMAEMXeqESFb8ZXKphyHCh1W
ifvKEjfxpKKUVqA5OzUShDUkESBQ3hCtSWnQXJ0DRkC3yGatsSBJfFO4Z3J+c2tpH5uC8+svyruM
rpf4Itpcqu2sCPVHWmLOqSSCsrOT9+/BT/5j0njuX5uQNWqH48uyecJj7fJt7aeLNg1LMQ6GkstE
Cpash5vGE7fjmfPwnJX/hvHPQuTjWz3nGvnPgIYrzXn8fDoTtdGEkjdaBF7yL8Tpm2hCtrzqIiKh
tkSudRC7iPdJTfHMaagLRAMcumurK7qlled4sIfOJJmlWLVnPkAgRI+3x4Z1p5qZP5gpRAaes/RP
uSgNhOdrA7QwtRbE4UTLQfBYCSLhfYfeKOkk0SSArobNq96DoQSerBtpKSCDAaHgNhkD+Ezc22kp
HbIa4a5KLNrbmo/ekxlyzKDu2ndhgC92qaTAKKhvrund5lk1ZXtsLM+xzrFGp6TPqZQPwGVq2Xg3
dgPZBltnYslmE0BHOTFtJavxesOOULDrM1Rdpgm81YF5aC+B+jFxmX4h/JVhdn3vb5uLUxgdtBQk
nAxKNmZ0H5byOB5WwRqdfPRD7b6IyY3UvTpOfTfHvGw3bVcwRlgpTEBgfRfQu99/BbwMW1n63MEx
2Hp/ro5ckqHjxtVIA3fijybUH42UUxxzzE4mLzhQzrn181bpbDSNHmhzjhGrhzoOZZ4Xdy9DAx+w
k04RYeyenR8oHrkpYnoqb91P3rrRo8U8qOHou08bzzlgkt4ohjJR6cRMCIIRt+Q0pX/eEAp1ph36
/ktFThu02TNQqti5W9ZDMHd2IP26lIgSRyExso+I0rjhPkkjjnVHBnMmH58qYZBa7fbXFOgG6LuP
1ys7jwoM5TK/LbzKts9hDuKvkGiRR378vgD/lgn/O6708307dBBf99Ntp8ycWAbuah4MYM50kJFz
brH+vlJ+CsB18Jg1+b5Ihmo1LvYeMESWsJbxldODmZrZc+sKq/M6yGvvKQ+nGvLQI3+Aj+l+frVB
cMNppyFMPaDYcbqaFaXzaVdhzKgnxMaUWISbSDKapRWR0PgTV2r/bBKVEmjayA2VYcEE/0KgGAVj
ajPV+ATRZ2pEhxBctdKp/zo4iuPtUnagyj1Mf6DXUaqK6mH39XHwjSFGYkAmCagny0dgDfvitHY2
lxgMjBieNwWMktnjG3gCsy9y48daBJdvk4mtQMMSSUPQvIT1kkN8UxnyW3YeQxbBfWfJFsPn0XWm
vVa/AhWb1xTpk8hrJWiEdoFuAnkgUXssC4Gr2f7lYxOlzgf48y6aa5xr9xze6S77Y5ysOeI67EG8
Ppjckvapd9Am1THYOF5fLCmq7JNv8jWBBpBy6BRarQxrQQ5VbCdlPZAYQtpyMMZEAlwdnYNvbQgl
YYkKGuw0ZJ5jZTvHQ+Em9AVfvz37yQWR33FMzrxSaEf9pnoJVocL77xvUPD6M4mGlfaRIC8MJ33D
3xqrvYcAvR+xGGa0i7kZuzvWayczM4y7YVt2yZTh/ggS4nJ663Y8Z2E5x7nf7aSbZOZ+UxJMH5jO
kUk3IWmSE4gUzLjAjIYtd0Px6DNgbosWPUBx4Naqo2LPeoFUuPqjSbpKga0ym2LB2batbvuxLOdo
SeEiZcMSJ+OaeNDn2RV2dxxiVi2l19oey2AYtIxrIH38BPcSNKSkg8Jgwnh4nIlQ2SnujeobL3uP
mM2PNKptirczR1evqvk94dllLD5gBHYJeiHH8IQLarGLWns61NJOhIUMez/JFiSZYfjEVK4iywv7
g2MKXmFQV/twUJ991J1mPwHy//XaA8gmZChW692/jKmE6ZE7GN9FIEefr1B1+yTP/arMEvit3YY2
cbGvGA22JHU/GvNc9XR5YcXawyV+Cfxqg9TsBhyAl6s7TGtuurTzCM1DQkA8EdC/goMvBDe2SPqy
lt7e1Aq5nDaaxxJA6eqiQrBDJY+o/1ts5QzlLaFwcTlPOieR44oX/wotIdgHi2evXnQP9Ib71+XG
SkGVxjuRNLMN6MK7SEbRc2IzZd25KlSrR4punMrI/KVa4SfeqI6a7/BIkwUcwcIbM/Ga1njZFXo1
YhN8LU/WLWrJljqecMaTr7Pa9S7xGgFdi3xgoEM20cHsqE7nAydxx6bCjGz7tGx6xy8NMgB6uyKY
PO4LM4T62F8HIgpyavw0uJPT+iOydkbScE0upkJp73tFFZ5yPcDu84hy2R+FxgkCD6ybhkD4e7bk
hEoGN/+d/vOyWetzKUe29j0PkejWBZ7qOrwKwzCZEFXbsDTvtncO7QCT8Tkhw1iI7kxTyYKPfGfT
A9gteeXEnQQ9joCeeXCC4BfiphMmh/ImjfVytMmGvJ9zMZ0YHah/9d4ArODFbzy1V3Ll6AjWBfnr
JqkWr/afTlt5LW9L8ZbU2p1ycaUyF5OiqHZ4IFqjHWbOR82oO8idU9Aa317vKXR8C1aHg1XCwtqn
iCrnQzTg+mGmRuhRqxP/aYw3Ror7QUCpkdmTVEhTl5isIFC3vOEV5nZS/JCGHpSk7E2WzorfHgVz
HZCJviIQuZaixULT9pN0NbwVeXcZ9iZgBF9vkp+4eOUuRJwoNIWG7nKBH7s2tqF2YTXXYYukkRo2
aKtFd7W+YZwdVRQBHoTiKPmtHCc92ajSNq6L3gQRcs8NQqi4TyZjeuuJ/TyQMJXQvGFBQ59CU9s4
Wx4/lzoI890Y8mc3VxMvriKI/DG28uWVZHq7Pb0KljxcpsormW+3eVLGXpjeqpUilGfAXQ5S2kTj
s38ASoATQtPO1F7WAz9o15Aa9NxMX9pSVojLy8pXxN+ExVWm2yen0uvetmsaYndnAKBhbO/74d3Q
6L5gLZL/c4ZDXytP4VFTvPhb2GuTEeCFbfoYRD6JSdZl2H307ymlqKOYR/59w5cI7NlXsXsXaPHQ
VhRlTsd+aEZBz186h0FiS9W4iPYGzl+YhJKPnbwLH/nPqkjJh2mugbxDHQv2+j7ZWfEQM6QX0lXa
b12Sdm27cPy90x73MYvL8jPum1IWLW8vAdRljIf/xng4A+TwcoDgifrvW83tprHb/NZ7k1Xc2EKx
2gA0dIB86s4O4gWgAiThWCppAOR8PWGSDsZ5/NvK/BER76XbJofLTPEQTYO+3ky6fGc8S6cOetff
55YH10xgaC04IQjgQfpmWVxI1FNVvT+ifvuzWe58MXQHt9oFbNu6DZ6Cki0+ZkYXjiGq/B59LGoD
W+GK8fwXAbU/p9adj024E4VisTOoT9WwgiQPArENx8jKnzyr/+bqX2QOLR2xcFdemgk/k7YORBK4
s/3sre3McXtOtsE2gdR0DUpmF/2LfzVLhgoK6L94vVdnWBWHvik8DjJTciR8H4XzZdBk9dhNrtfl
Zw7NsVjJ1FHpwvmiUmLPk+2zmm2t9dQX0kdfuRqmzSSNrV78NrB8LhwiMa2RuBL9JufAHy6HGDDJ
/oGqOTDNiOxgWLGX70M9iKlIdZkaP/hKSyzQO+TAkNe9okyylpjyw6qDRVAXO///jPuKsVmWZ2hH
jWk3Lp9SUMPQZzKkWaOSwJG31X9OLgYxKosyz72fQHQW1ObAddLU0RQXBZxEmZeiyYm+Lk4mrhDq
WV+W6zi6Bo1r/HNA4Al6MtsLyGPzUjrUTdcRRJqdjko6mL1/Nz+peF5qiPXf8oPJ6Zs4M5BkkZOu
gsnY7AFWgUSoLZzmeAI5k5b0eUTwJ2ERH9gM/wCVMIUVcdKF8Th82gDra9c1RtF4Ai7MhonYL0ZG
fWVfcKIiUw6LOYijZk84o5rLE623du4WTP+dZmuBlMuXWXU0kq0ZOHgQbcckI4qZDJgL/BqUw9YA
4wajkmpVP7EcQheFxSfDh/PTAn8u7QLvM4ShiS4XWD3t+R0AmLV3hDW6543S86XJ304ss+ZLaTvw
xxPwtP16GoyJn2zYtPW377/m9atxQGsxcFak980Zormdf28LT8kDi1Hfo5nOI2yeEH7Tvqa7VDpe
Thrn1Y+LNSQ49ZJCvX9Ios6CV+tc4S2kYE41oUKBTybhAZtioBLeE55LTKtuVMEzLwgOg0dmPlPG
F3lpCvajFdvWN8Ifjn15oNAK0xuxWV3q/HHi+T6zQgh/Alq+Z84WMbRGJIqppBDaZbc+fcjCG7Rr
U8zUFo3UaVDKSEwBzJE6jQp+TUj+mVMPoLNCIrX5yJLDQEiGb0vgrhIUq+87rghmOD4FlXUvaXrl
uTQeB2w3hmnJde6/coE8HMyLy0QAjz77NBoYPNmuJNWXL/eOzO27j3ievc1ZqV9pHAaZrsjFHAf7
kj6ksVFSY/Hb3dHSKePEmdpyYMQPUfZoyEOmAjA+UU/uH8iGOcWrhcJPAVpozoPLN3+yIqZbNIiK
WDAGBs84TA/o/E+wO0SUh+IZR8lu5HWYn63EqHCwnz0ng1ZMcfrJP0BZe4JvL4ySYjIyE3/Scu4k
4fz6kD374Ty2XilEs7dGTMbz6bIazrmfivHFV7scGIfXLsrzRuEVXb+QUrgPtg8oVyPVX2NxdaoR
ZZnZGXk3ShiYsmYSNrDlRNI8WNhlEPlj2mYjm2T+j2niEgjhIxnmXZwxPAeDEY/jbaN0hD01aH5r
bdxyiKpQhI1j63cnUaQZbXwigmRiMZ+kvM/bTgv+XqUk8JvXHYPVR1iPt7aqlevYhXWArR28ht9k
2XQ8qceJxAtkxQQzcCsXNjhKq10IRMe5GbED4yRQax2P4XqfaBmbw3PD7M6qfb1Dksp5asfHLLPR
jIzQcw02Z022nBbGUV3d8eGobC09DNQ0ldn23MyqZpV4kSifJ4gwvFERp30f3CRfsU0xbd178RVr
BnizMrzlhlQvBcOU4JeHpnqdluyxZnFIRDU+GlW5p5q+TOTpXKuuSSLctoVYpkpW5k72o4OGZKjr
muYHbxzWHS9UXxt9h9pZ0Q8G0J4/enljr1EL6DVOpy2rFurEfhYpAT4WYpCmF5qE6/iTcDA9GjTY
IyLKYYWOfTc+wQa5Pj7Il9MkMn8NFLkhu/M/32MZK37DcFzwKQK3EYN7eeU1qf8J0622WSOFJpLS
ivV68H1pq3u9nl0KYwtGC3Oy3V48A/geir4Iv73bljPR4PgEx/ChLlnpMToB8FP21ROzFOzK/pCH
iLa9F+HiUnuJvvz9Ab9nHIXrrdRg/6qawLpFNTRr1DpdloqLFTQVpFMh9YmVL5Rj3BgKY9PB6azK
f74uvBHZIDXkZOHjnRbFC6x6y32NwhqWxuxYotd2Az5z/fbrl0VwF+9La1fSG9bPxFJmi4UYuDhu
oWwczE3+a9hE4+skPNh9AQSFAQ8y0a4E3AhhulZ2fHoTwppyA+SLyKcpa6zvZDMC8coylISjlGxo
0q7F9W428IqV6yV/Tx2xKh4+92uGg6a1prAhdfAPvJRYgx08fGJvDgMurq9VQsAGk3MD0zQINxrC
ytLJEEpoyQHCL7Awy1lamggvpKLq+qiv1UjUPnrjSSAuhb65iQHHCmQxyNenQ801emXf+H+x+Jom
kUGJZavzKzuolLqaT52/0Uh932vBJP9cVi241lSclFX8nDZf5AJ5c8c5Q/RqT+xQscKdjynvovBc
cVVaIINJ7VfMzd3H60lnButw2rxrcLCh60LKMyP9QAfAFmzmReWk//kHcbIoGGmE1Di5euxvhxWg
8M/zmNGMKuj7vp7SuHmQhw7me4kNzOaaKQSb/+x4GlmsyFl2GmtmRPJW+3iBDu4jH3z1AjsoX6yK
LgRkn7FWw+lBCONHD2K29UVz5OXe70iFjPuPAVSiIh/kEwK/MkFcDjC2aEAs/iWjPWkLyPQvQdmt
RBK6ASQtr551LHiE1BeVQZFsTt43tCpdQvPA64gchx/nx/1BpOhUOkbaiktfLR57HITTcSTFfuJ8
8nnePVIaBVoajSdVAxB8n3iT6cAAcZw9MOVgs9XnCbQ4ipWigZKvpNnEUJRtsLlm1ZtQDgX34paf
lHlFMHsz3GlSMEvvNFMQ7snP91iVAngyALyPAydqa4njZL9hCktJorV5weEQKUAbT9Ns/+iTVUjI
w18Ix2VzJm1E+a/udlQAFcXr2Mn04RTn2FimTxrq2Us/D73WjJGHQC6/Edu0iekM/d30yQzon241
lu/OasRbAj3K7zH4uvNiOP1Nk4PTDboYZoXGcJTwVcVqTBZYD9N1z5m6AJmyhd9VAt5TTDIMr3BT
eDTXcttO/4rHegHywkoawDhGFEmh4AuZFYH7nxMbFNq9b5kNguUeZCUhCJfQd9F4fcIqTN4s+rah
OT9mKs+oFMSbUWkzaPS4BsX90rFbIvU5eDofHLQu4pgFJtaBDpF0Sci3HCCM0hkfQ6Ev/ODyOf0B
U4nm26tdzze4T5rAzCvJ8hzQWgRPr+GseIfVkXhxJ6oYd1i79mJvaYrYVOOQ/ZODUTkTXEIO2ed5
uJO0Mc8zBKdg0t9ky/SqD77wdJQYrWKfsLXbl69QlcIOpKEHquzqk8P9O0gMAqvnJUj8Dlq9kMKP
PXHwDzDXWj7J+ziCpZ9DseRsqYalXfuR1jWV/0lu4zWTi1IbrO9vUC6ModTOXQi/TBFDhl0wHlkz
EVuIfP2Lc9sCSBp4sVnjxWyBJE7lc2Bkd9caJXRhki7RxidUnS83ersCOT0QR3TuMIkBy9h+2Sjn
OBkw83PwrzIecO0JRJ0Jk/MU/RbeuJoqRS+qaoozDaw1a2YWYwmV+RA69BmrIQRBXv0yT6tLDVNI
b9VSegws0Tr+FRuGkzCiX850bVVh9k6BGdC536ebeyXQo0FbE2FEVlUZ77nKiFsuI6sFeU8WRTWE
KDMbDZJ1vOycm9KEcxybN8bSPHZ5CcYzII63vQdKmCo1nxklm3gmXr3MTZU7akBafz2KKL//vt0n
064GRnEd0xFkNyMAqsAuBtnGXz1xlgLPhvhL9ItFa98wZQzdLEN3TVN5t/cipAjBGbLBp1ohacfB
Q6z5xpu24XGCXSsLMD0P07n1r36sEk5aUGH24kOF1hJF6Ucl5r49VA7z7CEiOcpsBPT2qiqwFrU/
7hm6t4PGZ6O82mIX/zNowVMAkZ/FZkqdwn2yOvt3cTg7gZx9Zy4QMhesBLe9CPPGgQvv/j4UbuCq
UarqbdyvOPV+V0EgEVhD0ixheaN/+Y6j5BYaPHP5pZJqXX1RJ7lkzSmTHpHsM8RC6SQYCpWOLLZ4
RxreleLCkxyY9OZnKb6nojAPmhxD5Xff5pNDjjEQOuR5vSJ0B417baNVc6BL2JMmwUk2PLciAttP
SpDOSDjtE5Yly5ftsTS/6XVCVqsZOxvZGbcClBsQp/8nZ/BV2hfjIgSQv7L9bEBamrioRmQaC/u6
0vOjV2tu5xQaOs7zxi/bTzewBUdpvyk51t37N19GrJ8ASpGlWTW3gn7RrBYQwBsFdHq29ZODb6Y5
QUjpC1V/MG7y6Z9nJLOOVFdHrsiVa9jL3UnEbcBIiGzUFb0KHh7NrvpjHgbsMdD+sI2e+GUorYd1
Qr9c2mjI4Hl+bf0TwuuUSgfb1M/pKx2CNGfR5pGIBlVVDwxkhmCVb14VzaV1LroJ6oeRYVyZhHRE
7cISOwH1Fy5BL5m3htSQBq8Ny8dy0MOu/RH+4QUHRPigDW+AFPGpkcSTXiarsnctiZHe5SikKF5x
po3Zd03DCYOTndJ7EHKbp5fzUETJhkkrePY345J1pFT62EDBFI3LGYocVyPxCikv0hWCMW+kP8nw
BY4xorUktPy8FC3pK4Lt8IchYr8ipFLUtrEffkEgRsx+s0rznRkHTFybLLJZ7+ELfp6QyNbhc2sE
czrO+naLezsGJnRCUu2p+1osUo2LAu8qtLlez41IADglRhw658Dog83h4UavL+nguPMwAWqU7Kcl
syml9covKdaT6fKVPyxsY1eSQ5LxFfabhPxTZbCOiROFGZ1zDKsS+ewQAeD9QY7M8KiGqM7rfotH
9aGEw77lZExcAe78aL5nRA46KiGmt51FwsWBRUJrr1gq8Q4nuJWNPpNoFtMcSFbcHEkg4tlJwRdH
Dylfi18NKu9fm4bo3ImegnGVmrIlMCjDRDqK20d8TgWO5oDrnY6by4F8F+lxse02Xy01Y9HSiPMA
dXGQR5hQkeBqn1qih3HCwcmoqn134W2tNZgGpefCcKtd/gP/iLsg4u+DgjFVi4s7wAI6jKLHCfwd
itqI5obgKk3DvexLQgjU1PEa/8D17ZWFnR7s43MVQcAQ1adrGKNdG9C1trOXAL9iV93w+cqAtLl/
7OStNTLegKRz09qLAQxbhWkbcm0GL9kLrlVN3mBDqLr7jnOOAy0Fbad+mcOdDv3E+7vG8Vvv7whZ
qK3Dq/0NDYuVONCtCASjKlInzGh6YITbbVNFCdDG5DAdz5tteSCXsBzDXtMWSi70mrgGHBMnvFBC
hHcq1d9E0cN8nYEcZc3QVqs05islTpuQHpXg1HqMC8jj7c2LG+QqSE3yQ+z1mn+UxQeKXycs4hfw
xYxgB/EWtm26JaqHd0RwZdgnswLXCBU7IyfEwtd9cyvaUI8JmnDB1aStprI4JTnkZwgQClI45OWM
xwmhpc1ldlyCSzDzxa7UZJg0flLKRWTMGLGQLYglNwB12Zlx9zgUgL2VOC2k0xuTIllsaV2sYCHK
zribzOonERZHLQDodmCeaxvDDLe4Mj3b+GGMCHF4mf09oPbK+gY8YU4+jGqOSm7Gx+Y7KVGaQqIi
osKfWENZl+SPkDf0SsGVo6FFNqWW1TGBEPZV0eVfJwrVrYFeiv0DVSMUYK9bLl0dOIUK5gpNh7jX
3AjTlTB/jWunLBvjGEl04IOC9aOFqXlvIn6hYnm6pk0wpOkXo801FH1dTs4BVJ1ixDqw1hQqCuU2
Yf+N7bfapoiLUCxa2Dnq8/vnZ+01qz1Jz2BsGaAOQaLhtbcqfaWxKnJZALXMt0QOrhsWFTDWH3qj
jIX9+pcximOd9siMhYgy44J0+Z94yIc1TXr5FEQGx0bCI0/zt0sfLCePrRyL3G0spJ6BgzT59n7J
VVsFHjBrkSqgZSOP0WuLBN2MJGPmKY+I9umViE7q4WKp8ikLo2lNF4Y1T9M9fFNW9VVXOqavfWvW
SrdG+24EaLL8QS0wyZVzUDp1DB30Y9Q5nnrNY6vDqAstHsbH6NbtC3W82+RmuoaJFHSMlBL1PgC8
gvdWR2ntonU7a02Ix+7kcjhOg0LGdr2MrCdMzVHEUD5SJa0DWfYvyrQZvhQCyXoy/DQsBnIFp19Y
qVOypRILpajg87IRKlewxoyuLSbVLIEZPI/1fl7wxwXhbpv+QrY628krbD1hJUx0euhTKLwR9qUt
gmf9YfESNtxxWOQSRTeMJ3hwPcwUukZcwbBhj4Ajf3Y5yn6A86Ey8Fr2ji/aPneB3z+JnK/Bcg0n
yXC/u8IV00jILkyMI65Mn8XMnjjCmzKQn57o2cEgStWvkUNTH1GMhez6EN1geVIdyKafMDrw6COX
JLb0w681iGVZaGG97sSM4yrE7NJUWjWr+fLto6uKax32yxAUxKeRbqiHq8m+mWBPVJrq1y/HkARg
aSPYi2jpo55FOuodc+rlAMEW4RaVXtqcS41Id+xiwGgP9DEI2A2eMPF9tBc63a5D0xfe7ol6JlzI
UtD4ZkcioYYJGSVumCu6EgLi1k3VhOFf9ttrm2ms1zrRW0Txvk6m2loA/CcIr+DJloFRg6/LLwB0
ZnhT//vmWKDqkqe1rmvNHm6u6NsV9RKE2jBOM9y7GKtAEtpijHQ7dz/gtKPFgdisnMq3j9OlzSdl
nuSojD3rFdfuXBx8CeEPFBjIDauLNTLkCUhFMgJNQDVpepkAcCZB2oe/FOYD0S35gbrcJr618Yeo
LWUtgxiWpW7O6lA2Ti0xViNQ8taRfc5KtsulET8iNx6ggtYTlrV9x+HV41M+o+/374qLvIOv8qVN
6duvrumoqgK0iG5Ak7dYH/Zlw4WPPAdy5HLDQQeV8n6NaN+IG96Am+exVYG2y0i0UyfBy0OzuiVZ
6Gigoxe0jgfstrfKXOt34QTKeEta5/BuiWHMdbP6TiiDL5NCRBaqluM+l7RV95GfBeh+Qw+KAvHD
/MgKG7+3sk8OYnn8yugFEcfn6v0J1dEF1kJv+3fsyhSikuhn1JRnxOIjNg3yBDo/1yFM2x0GZsAY
zz7YWEPYKTsaM/E0jDh6VLSZhjeyA6pqUlWbq9D1vWr4fzEa2IUaJRZ9X+/RQH0tWNPHtzJJA29N
jKWl0vmOPgNFQuEZCixS9u7+yDezKjOH6gWmYgYcC4wWZ89nlI21LuorG3UYoyvRQZGwJQS4fxhm
0KNf5rDFBDSqSeNmYY8efD9ldFEploRgskzgtebO1tGT6PpKZNW4o8ncnxQ9tT40rEvRCFr3yoAf
7h8QcWsYUgaotFirfX/naKcqbHGKTCdhHAxIYcOx0hQ4ryXSwFkYwu2fazvSNZp+mvkJ5cXWIhdr
ROdEnGp/kBQnjiQ4a9tByVRT/1/rLlZLtNMRhX/cAsN1XnaqxTUXehKUbGSmU72aup1ZAV93YEfQ
ht7Ol0kWc9tf6drV1zXh0NT9xRXqa3fnYukYk4PzTfRk3urNgl+aoh3RERexEeyXW4wMTfcpK17S
Hv6pY/iWI9ZNXvXeBXUplgNqhjM7UvKAj0UkGoiY65eoBDxZX0dYf861QF1xh8JK3jOCM396iApf
A/Ne+IWpMxHBrOqWNByVDpZqiJZSJfZivAchuFQUO8NUapU3SWLMujBEUooonmvtuF0Q3udPpU5k
QXGeewO3IKbmCKwdSueY1qcOO5C0tcAU3iLVgVy6uQdj/KptXC+irGyBsgTkZfT+PUjpacagP/pd
GHRUlUTGhC/NIGaOh/v+Pz6llcYtlKCM4EAK0M4/p0vw6VFl5s7Bt4BxjKnclhEirbdmpqys7SGi
1EO3Ljap27hC2Gcsqa8CJdz0Rrf8ro+Z3gKZBwweN/sqbSV7b5q4ilxEH8ct9uSHdgPVP9pwTmf6
tjPAOadRHN0VlphcCnaPnd1KB//7R0gxKveBmEHqkJYpvMsLhpj8W3CaZ+UbxT2uypDfTQ8FUFpe
1rI965HfvLmZKFxIqgkM5Uei5ifcIDRaZnGmloVvMV2LgzHkIckLezQa6bMJ3i57hwQ07hPSfVq1
7iBBGuwuPIO18PPQTqoWisu38JRaylJ+2bJsuaCMkWJPYhuxpryBXtTRK6iq0JtqEzwHxPSL0Vfh
a5ACvvl4y2phbnhMIE/XJms+QC5IFslXrfIBAwfwqGXj+Vmw/MKglseN3ISZAEUDxW7iYLZEdEGd
oo0nuK/221sNaSA5/k7zNrwwqb1EvI8skwTloFsPi6q09I8Tm/HqG4d4eRrfrmtGOCqeVGs9EYMb
jFtyHcKI/VPdpicTQ2Epl7js9NKHdP5xfWoZsCTmCaroaQhoKpIRPhtG8E3xD5A/zxo5rTswW4tr
aLuPkTZBfpFNDtKs8P2HpeXTPcGMU9HKL0OSJ1S/Q8TmeUP6MO/OfXPzhXNEZFz5R/KCzlkXAAkt
fPLO+Nd65jXW7HbXYF88MRrsO0fK/aCvZhXU24zKa7dYX7QnL8EoEEiCn1hkQA1wTHMj1jw8irDN
2KxVvDRINqE0/KBp5JBTA+DkBqjn3BaB6KlQfUnATJaKsJLR5Q94P68UQ/pR1k0KsROVNAX3ppUY
9BBH+HGPkoPqtcGPMuzvMWD4z3PgSEbpkOFRLmJy3o19SkH27k4OaGZGKkCkokwY1UAxd7PVdxj4
/nOCYm7Ex0xjGJUtk05qhtRSCCAiAimFNzbpsxQFg+mgAbyXPyim2gi8FPjTzzNvwBtuRNo+Z/Hv
MzfWWTIS7LqFJVKcN7vKg1glDUd54s6/+P9dz4vmw/gehatiG1m+1Ys7ZzPBGaZhYvNGWyOfmhO6
UGh019HsBu4IaDpoLFt1lZMEhhJB7ngTfXDjD5C+TGWb3zeIspLwrUPcSL+ugtDxw9IsUZGdlIna
sDCKmpMTw/JzNmpQnLtMjgg7rTzru+K/LUX8V3q4N33WUtYfkRoUlFXyWba/7XgtzWRLIX2Dx7N3
xWYk9ayFgpDydpxYwP/W3pFsfuLsCTi0cAyEVa6nR4OfIJWz63YO3y1M8Mj+sfyONWwjFTC+HlCf
0t2XiSjpjWFskDRPocNnIFNFJduV1mISlK3/k88yL0Ul+VJW6+0BnjIli/9yn1lJkaUJ+kOHOjIM
Q+oizRP8IS3nB183qpAzHoT/nHV5cFV/jWJ4ZuP/vHnUYJ+KzdK04o94QAxr57XkVEuP+O1G6nau
wmmP8A/+VSzA65L7P0AitQYKUmoQI9KFSltjekqAp0gckoGvCkysf6aaJieHugVH4Z/njU5xSGhC
wgml9gCYP3wonqMdSUXWSUzDej3m2FYQdq8wZDQnusZ0UvMiedNCoFkCtCIEA0gs+fBsQ26K/LjG
a4bRxw9EdS7QxTNdYLo53fo2J2/dV00ULino7tf8f5oD9rANutixUVi1X6N1luKOQdW5zIeZUDyr
Fg8ADiHfLaw+tbq5fEMHx2TPWEQ7X8phvt+/GzavmUTgwe7/ziPgpMc5hIvjSNw3pnaWVgeKIh79
Tr0JCucr15knI0PS6s3E1J9XlvKp+nG3BnHuowKBnFmPx9ZE0u/zQgSQZ+ZCvYppTM6UqRo6/raa
drj4V1zlfgHAbFylHO5ViZ7JJJFiBszPIKMUjPcKv3l6CD4DS4Z+WzTF75CdeQD2kPZkPG9q7584
3+6KbkqlWpLM3WUqfq7srI/BYDF7eEnGb53DisKnA8ylPkm4AQqwupv2FVURgbxOOf5mOIoet77p
EVDUo0HpQFwIgN2bKRcLc/8OxgDkil76D275FJuQl4ple4/ClszWkL3VeiE7oZcTd6aUdmA5rhRD
V8Dgcs2gO7hBsY8wPsa8UrCf6C5pyHMEDuBm9qj0tFfeSaqmAt8+PksZN7sFz7QPyg8UbdBDUA2l
A7qzKieSaAQFNc7bArDw6YMJVNyBGhejtVnOTDvsey4wVdgJgKKDenuk4v4XAGy5PFu7zdDaGlT1
kCdKVclfI2M5arD/yIuINhEqRgIOMUU4rJWnvV1O0AsMm7XcvNagft+bWbLCKxoe+CK8T39QckWm
1NOp8CbLaR/EyRto4MD+oaF6GajjB92itI2uoxyS70/4YLakgcpwGj50ygfA9IRJzX5ApniITGPI
McIA2Mkzm+1V5amWeYCP7q6vvvpM5tmKXECLFxp8SGKON2kYxcWW4dZaL0/wjcthp9IJYZUl4CwU
ODkgNEL4MmKZskdhN3rV5zE/FopckWvboj78eLVnlHfYzuFXY3KoSDxL2N0LC/Dlf5cEicPO/2tg
IJdaFZpsFRR+SkxtFiORA8ULyB1zy+0HzUb8B3BVors4t8Altj9eqXM/PjdZbyLAEPd+CCZHLA0k
+3vWQ2reliHXcbM3uQWMB5QUCVP7VUh6nZwe2HKXclUIQY1UNtr/YTyF/P3dcJCyNt7ZoO37Pbtb
M2HEK+TWcIg19H9KBsh4C5CRJ8lVfYQy5yu9VkqutqJg5ye8cabL6CqIbMy+Hfucf1G2smb5KEC9
0+9tEyBRO0l+LpSAZfElvLBeYFVQQ68wNOERYypOndJkQiglFw860cOk7C9QVXwkeX8yoDM5Hw6T
suErHT6k/rNKAfx/bmxFOC5RLtW+BTfVEjJvznbC0rTXC/cZYoWN0RdS3luO4ulhlJb/jbWMtC1L
4MLwtAmGTQBpTqWRyZnyNknLOH2/abM1BJS6Hdo5CfKnQW0CMHEUxf8g3E1kHtAqVMw0VP/ixxff
Q3YAo+qFsWXqKZ/fQM2qblwgjM0+gHlaT45PTlSICMUaDukQ7C2orO6mBKToPi33Pi+cqX/Iidej
ju/5SmWEf0pH/opZhifuZdJc+8mBs1DDYHejpw23NIfZ9hM04LwK1uT2SO2hnY8D0rh2Vhu1xwTo
DT7zUX5gDlzABwJP5NcIRuMedEJKMoxs8pVwoqtBU9mn0ctbCT92hdZ9U6a/4rvm0NfXK8wM3IAG
QojNnc6BGhj9pQX8RTlN5UdykRlWdSg4378UVJdvvbMkCd7VI6oh+7eusw7IYad0a/2XkCcUlV8f
ATya6k0J0tVr3ikgiJju1nnTdhA7zMqjcqd8OoCPYv59o7Tp6aAcZK0ku2E0ZXzYyM8DaPtLzsJW
j+zL3q1kkFI0LW66l1n1aEe/+NDnw9pDjRnUXNO6laF5MHxRTh6yis3u3JvySEuPaFWk4C7eKgGO
RV6OBqcRXmXJDksEFyTWwkja7Uofm7/c1/1MHRNihm6KiFF0JM2jFVxPEYJUqUeUpZK+1tJgVsou
Zn86SxN4g8FZ3b5O0ARIU35IWzznNgoy6xCpsTsD6Mipduar7IQme0TFvZt3JTHl/gctFZCsuJ+B
NJtaoACt/4UPIjun+3arqMHLAt3Pz5xW6bO1XWjpTdJSjzuVaj4+QhjpxXhDARipwv1pZUDBYcnJ
xQ3YNwVKPSC1scMibBbo6nGSEozRKlEF17Ig+AnnJjntGOoqcQBsaCykSVixbjfAT9/2A35Cn8SK
tAny8FYomC1bkVJsiSNe2kHChV4xZGaqOkia3erAXk4jAMJIs5VO8qvXlNrYF3RQ19SzqiAEzPup
Zv6GRxZcIg7zn8pshFKOCltQec90WSWhL85/cIPxaF1Gq+SUjLtXcPcyfR14StwA/3yBTskor9+8
89poYD3lgdPNrJp7Tho59NlpFMHmEfyr1eNvYd7fn+KnllcYt9k+jFrEL/XU4b6GSMVKQwJ9Lf8o
3j11KO7aNxms/f4QfQUbMYy7hi3p6XzF2wXfjDCJgyAHYO3C9r3jUlfTEBpJmj2seu1GNQ9p7EIA
ZeBShrgbV92tfuIxguLzWvJ+kw2jL7LPJwuJ6rXhB+808mn+E0MmkX6M01X32dC83++G1yTm3JpS
wSdsGZsWu79H3DndttREdiinizvKp3HIeIO2nmC/VK+55T+PATH7sc6ifGRa8oHG31qtZGPPICP4
BpzagYQCNDISaZlEiV4Y1DaBxjKDSRytJcF2WUPwy89lC3opwUFiwuNM+vYQH2melSPGyCWZrszM
aePm09GqqKoe4C+L2M8CH6zPuHwVSQRQuRsGU8QsaWyYN9nbK+LwOtLpqJK0KqUZYw/S+eKspbpJ
ZLsn+EAF0YBmwPHvdDxkjXnFbrFRZR80o99r5S3+dd7Wfgusy1a0MYTbLRlsW08uPC6uCnlcCTTJ
A0dz6HuztX+sQf9d4kis0e9gswRx3IEDeaushBb4Pu6qguPEy/lJyRr+6NVO+S514EBMcncL62Qt
egoP3psLi1sx0kOEpynwoggzzYKLDnNdE8IO0HKKVCWMlLil7idBYVUqag2XKfeo/9IlkCdYdHzY
o89m6woNKI0Q10w+/GYoppAbTm+oQ7+3BjLGu6pUs+bANU8jbfGNJ2HNvaOWHFo5Hsuc7oXsWFK4
UYBP8K2uUbG6u5DznUcRzJgh+GNQR8hboDXjAGHNwoBqiTn1tw3t6e4f/fewjhZcQJRpRPPQliUK
yvAHRmuX/0xwwvAgqvU16ItkvxH7i9mWYdDxJSsXlfYsHTNeb78QYrmi4PQ6+44Q0jkw1fiRDmCW
DVAEFMKfct/b2cm5d+4/r6iuj23k2kkzj1PXaBKFRUszIYGeL9SeLnyfnS1s65kjmRk0oIRdWWUF
8oUNBznSOZFNJ022XO8KvjgnTFY3tGpNFfPklo4NBHwxohRMqb8v4rUUcSZ2DpvOByuo8WrJ3W1n
+kRusXSWgO606fKCaojtBRjo5HjDjBtPkaXLWFSQbyI5CMDAQQ1zw/FrLzKs8yTBvNd9FgZTXOQW
/dzKFGuDlczXyM4dwDVQt+tCd2jdKPUleSgL8h/qQ/tmw+Duzz+t4VfehqMWlt86Uf5/aJ96Ub7b
3d8UliquTb5Jp8prQ8rmT0QaEU/T/CGnDr7T1rff/BjeqkoWzijtpwDFXcxC5QX/mOR6Gg5NK7KU
rg6PUuwSC5MgBB0q/uWAZOQqBBujAnSfMa5bFp18iC5alQPfTYh8SS45I3KrD5xq7e+CtCKzceVr
f9uA6XzqBVcZs26kh2pX5H03sM3552elWSPWOMzKK1cUiHxrTBfPXIeC1tV8Mtiv6GUdIx3TX/d0
z0XKD3bkaOpcUPJSGL6lCGwupXxEHoVNZL9Yugoc0OEje7W1+40UA6AO/KbkDeLbuURbaqVVAZCD
fnT5G3T5erXxkdhwcg1vC4CNuqnj7vJfu+kQDnBu+M17KjxMSnBWd3fmD8AzVPMbEBQ9hNkUtQq+
Cl92BN383Jvn0r/uTMohn24jJczQZCvzD+9aGhTJ3Jg+Hjjsm8dnEYG8w9FB30je4Ry8s5t2MKQs
RYe92UsqqTwmUD4clIzRJw93vKBlcv7ffTnhJv3l/lFlkeC3/P3hNCSL1fw5ijFOPfd4x+/g+mKE
RyihJrYnJ+RH82+23zMWG90+E9lOSHXc43hU5tZLjzVFtDz21Il9Zl2SWcXTNi5NfwpOeutuxF8G
ihE+7g9cY/4LjNqQUIeflPxcEGLP/C37g1pbQab5ZEr25I/LMG67N4f7LjdmprSJSaMRevoTDjOS
a+6IgWOr9nWAZmd8FLJZcxgQm1Q0OIYizFAopF1dl0zIxAaq3YL3i8UzfTtdfGdMIku9EEfppvpW
jm2jgKrZN9uYiMpOsJTOxmIul4JmrENzIpRNydQDGz+YN19HlOD89UUyNh2nVb2UvuPOfIpxWshk
Mmm7+Kx/6jz7T6A6DoBYsMug8Ydvw26RnFhAKe9pfacgbU12GaCkw8hXAj7gAfqO8koFSE1jup6q
TjJI929gCQJ8ie5LrcP75vQX6eRW04+LI4MEZFxaHyohE+2q2A7GYgWDutJ6ff1Q2ocmNJ/clnMm
fSKKZW7jP3pVuazRWEDmbT3MOK1vS+aSmj2PXj414n8pUqVjXaZqW53Axw28Rxxxa3BE82wZkenm
Nr8uOV8jfWAV0QMoO6Y9vZk9nujUkhkrCCZJXcrmBoaWjn3bIDa/VONABpTw669JqiOTM8ZIaMQ4
V6yL7b7YQ2QabWJBL6YWGXCU5uvQ96vx1+ovT+Wvmn6I4M1z4e0IFfqa9FJWCApII8ZqQU497W3B
KaWhK+12aVi10xfne+kamX2zrKUa4T8mzrVvA+G4U4dkaSewPG2UTd7DhxPfHPMiJlgUsoacCMmy
uIMT/bfex6+VOevGcj8wVmolkX3/0Pi/UaYCMb4yAQnHinE/ma6tHysxFkimtvmCzSOfUxVhIO4h
k2GsX2eWdfvR5j/N5DxlgA5NPC6fsAth1R5Bn9MqcO6rAkScEUNkaBks3H9WFCsR+gEgP/wXkH7j
w034s7Bg1uMvOEdZcgznizWzDO5f2whjbuXXIncZYhVvLCioYJFNvpZEwqCpV8jAx27iZ9ZsGbRa
wHEXSIYjHHy7VTeEPWw8RElvN/NeglFeB4tJ3njEDiLeMLujPBIWMDq+MANxpg7lzmYjJRSciDqn
xHBK8a6oO6RUtWfnx5qzkoWm3i5dx5ZOVvGJFzy/C7hdsAoq4lO6i8KTQZm/GfRiw7Bk3g5W1FP4
EYFS4GbLtB4QuxpuYF6U/XYlS2aNfw+qGRGQUu+ktOBMDBYuHzKL/Dol3KGDNmFiGi+Oc+v7S8Yr
Z/EOXZqu5ywz3tTz/oUCn836ZtZWAXK5iK7h1nJj76JAgHOTVnq3U7O11RZT93TCP/bs8P9jaaiL
VA7VTUoFP/uoLsxOU+BhYTvQHNdwA+n9qCgFUuyYFw1k5OhwaKDb5AHzeuyA3gr7H4jgths00rWf
dk5bmRyogiCQWC9mvtS8EQ2W+s2WU7FZRRVa/ZW5Y1j1kMKVX5bivmPiigUmmVPhYSjimm84ztWM
BNRgSRrX50vXEKYJLuJU3STF1FjUxSMFF6/Jl+eGHWlOirAWE31PvvhRLCvlgtfXGtYRzJ7cCHch
kR0UGgBuG/kMj9/NS5kvl2TCek9xX2qlOwpDBRJXhCKlxYtSN9Vl+TfV6qkefUg+7De6zruOAh7l
bQPSSMBj2woz4GOGiOB/sCiTo/oVToqv2ypiH2MWCVsYRPBwmiPUwYA4FlFrvUbLKCnM9cqNasE1
fy+NsGDC6V/y89FTyU7brKpw2vDsznk0KEtPDJAtLzi9zQ+MjpC+KnV00lrjCeybyDds4KeXcGEd
ONLGCu8x/tSc0LffYA7Qu5nQbYbNQkDQ6CDPiRBn9EcRfvx3lS5FNRkPD2admUXheWCGGE+QBZ1n
xfKHLkTNPx76zSl4kg/n9j+tbTdhyFxPaUjAPB0HMF2Ka6D5IPItXfeKJZnry9HcyvEl+WnGFZvc
4cHbAnlBRrFIZzNKYDUf1r/fMKbBIwq930ITR+Q0vZ/LnF9HWxZAz4irrG6FSIZ9i0g/hlZLZPj+
EWM7mhKp7xbg2rUKaak8y+ZmcK3StquQbRF0lHefd2PO8BNy5cK8OpbCBaHsvPZHqTgq9uJfIQWg
nrSKLbBwe+jf1i7rzttWtwzPojowurTTF4haBwB2U7gd2cjFWabXPa6C2n4todTzdfE1lHOS0tNs
mLb6dEmRdRcmkX11K5lvZkaLY7DTobriibAC6vCKx0N/NbwRx4ZaukRebGSa55BwTW53Nyq1rWgQ
rihmIjYmgqBB/5tqOJcNsDvGLWdDooyNssMXLeyIOp0+hkWtzS0CB4WFdtUyTnU2WrI4HYaEk4Cn
lIMSEm7zF1bb5ECftyWrg8rkxlxFqXUvqjUlIyvapYwQTzhNVePdrqOROazrBElPptRxnfbpmIjh
mXZwWSnV5MAZNH50m8lCR+xCtXnQ2FzkK+9oPOxRp+1FU1seczt8biod/M9xtU6EYb7udbLjTzAG
K1xtg9WypOr0Qpf2FmU1Gsnk/V4pWoEIgGoGTHT4Xg1cQ3AqdHUjkon57NxsHZOuZadmsJcTJNLf
MSZQAhwROb/jodlKIlpVX7m+Goo0KjBi6ECSRtw1B4cK4zDGVu2Y0LdxX4eob2YX1F0XmUzLWAyk
UGwn3MQAFEuuZJPgc6IGr1ZjBMQA6bz9VFoMkFqkRNpr8FzKjYps+miDiced9iQth3LOstbsbYKU
MjxiQ4V0mRKoX/YJRnTvz7YMVapJj+tjivFD45dEa41U1/j1YGfKRV2HFro32a9iZiQYHRyIBHbr
2MEuMSUdI6EBJi0DOtO7BgjtNBi1vUcg0tEUOjfz19vV9A0KC2IDLPgFjd1Paq6bkc1KoJsO/1WV
scb/5cjwSIbhl01DiS/LW6VxkGmVwcI2GwOG0vxm+hsF9/qdGj4yMJv4qQqBbX0Vy79jy15RRG4g
y8JzL44b61GZzgPySPpl6BEKZ4zusQcb6UuyjTpR798h5fWW2JvYJ5BYz5IhyuRS5zGojFQmh90W
KNhZdn1Uuu4q9NuCwUtZMg8bUufv7IOdVPkA6MV/7+D1DsChLxvsnlT9tA4LaSRCPdIsftppP0OU
M396sIPrpC2D3HT32Wx5CST/0YulalAC12D48AhgqD7bpCp/MKC9M3wuL1CCEr/1Bi7/yWIjmbEq
uQWCIrTs7s28XUKE5KDTvLhUpR+6KgoXlJyyuth8SGBoaXp7TE9ZIliTjee/ISywPymVbZM5ot59
Onwa//TQ+K6zX3sQlmqlcDmCmIw+P99auK3nMl8b42US3mzuly8ydsX5WF6gMFJUqKKVU7vDy6r0
A8biaRMxwmJZ1dM+RqtFWYe23xyTF3JHWCBoSoj9UypQ4qC2xr/E2fnSFwJFGnS5buf8Q+tghQDW
OKhZ/uSeTiyJvLHwksNopCZ2MYsHy8AwJBfBBGPT09ju+HXAPnXgNDrFHZq6omkMquE0pOk8Ctxk
heNNydxp+ZYesLSbSnHtKc8W0YwSrpx8XoTbmJVFbvPaXSiX0jMjAP1YA86gNnbKuOTrNZYt17SA
EqtdqZgnjt6fJaadvi1UF90//bqknJZEnB3gyuWq/jLMFOBtN/Huu8Qwem+46wxul7FdSl6vqfST
kRBdxQX9THdZfhEyNXghnt7aF15NpACPDgA8fAudDUgOG81fy8nODWLcWF+NAznWeFgzLm0BViNI
m6rEiuwqXpeKkn1kXQQRdzostD9H4BjnmS8y7A2buB+TtKvTn8YdVbMK5Me+kTSnMnpntpDN/M38
tcqDJ13ZzNnnaWwPL8opCD0UePUyjB7RYrOJsUUCq0rd766KVOqmMOpsrP7yMpRvuSdCM2d+ojI6
sVba2mWwHOAryJ8QV8LjEDYf9UmfURGXrvdjw7CFwWyNk0srOjsD5+1WLngS84JE2hHy3C10xDHd
1VTF9Lw/Vm4TRLNEYTW7iqxSVudLAyj+iyPeLtJcAfZRMtasuNvBwJ+NhCoT8cod2sKOuCeEWgqa
5/WxjxqQqHaI1knNQnD61DNXqmpoG6Vz/xG1eYJT72r/AKyaBGwZPIKYJmW6otyhshDls7Vyz4Jy
BT07Xafqitmw4aCv9DNz5xxT5p0itkMPoB8Ims8eRyZKzx97Y/Xqz9ylpUsIC39TtRfLI0gmG3ti
HS9rE3y8qn4jXlvAn1msS8l2DCazjI4aEkLSxJCf2cpwHORoVK6ELrZkfsAzhuu1XnnmLFjU8W0u
2UhdbbnLNHe2ASrKy8Dx73PJG/67IgoYwdOAeqExvw+sZjQiFGnbTE6J4MRUkJ8ikDsCVj09sWbN
zoqZCRecpUP0p7NFpClKFRbCC0rsLeWlnKrme/lrYICWRnreccFDNQWJwz/3Zi0YbTf1fUaoqtwh
I77wJZvZsi77P6dW/qJmvosDg/eof1zjPsfMkJQFZDYHPvfRPJ+IPYGl62Faav2pA1yTcYiw65uF
S/WwKbEYJDYpD8C+fOafu2Mp0+KW56XDsO6nuWS7ZgO9ZUwhrgCQTtiD9lEid8hcTqbNqmCX4gS2
RmoeTV7uJmyYi3eYJLHa7r/khOaFbXDTEux+GtBN+Vs5XDo4AdxefL8fskinCWjFYVo3EGrSxp66
JIqJ0izEnC78Q7p/tcmJu0XpsET8Zwq6/oRGWTYRA5KRRZV2XrF8CVl7dFdSn/qQM3xVTrDnhsKu
yfbvtr3MXMUaNRnA9PF64R2gKM8CLod0pAmoR/+nPQO8oeMRyl35b25YqVKT3J/V0onm9rm6brWB
pJVDT/LewLLyAp5LxgDmWF8fLEcmgOiFzunkn/AspMO3tDddqoD1vxdmdQ5/L8rhClGh2aMvcOFW
8FbAXYdFwaXGAyEh9cU8fz7M4EvmmRog3nhSKb0deLQrz1GYiJSg1eWgZ9Q9cicGY2SzvqS3MefK
EGO7ik8U27m+YbxdYIg+PKFPikt3s2Ou6hAwhvBtqji90pifFxWoGgdW/fBIsUEAyRfdkauKDmWx
85emuO36VczXUyOZLkc82eEcL0aPiD4QStIZ4XnEoBfy9tQUxgJdLafCmSw75TMOPl7kcaLxG7fs
LPU3pAHwej5P0uERKxwDhAWaY7LKUXMGfc85eabZS8VrYrUF/GboQCnY9Civ+SpP3MY7EIDWiFMK
+3WIoaUUuljlQijgniHNeBixBYmaSTg1AVfEEhkj8Djv/gdq7GtvjjNfH6OKqsqSzfjK22oLWGBI
3bL6mHmekUgTjY21xSTFzN8WviX+sQGGdxP1eFIVrizmKceSj1w95BbemnYM+QLbzz4F59gRQ6TP
cDSYZtaG7RfoDKrHWajrciIpc4/qfHJueufGuQF4zoDWsYFChrTl7jXq6b8/HlvZ3gW60/9UgHvI
1LFwCJLCtZCZOz8z1RweAmJ4TeoeJtrH4DDVBn6+BhS5AvUL7vHldlF55RzdZwasArrIokwwjitu
A2be7yfMmeEoCms2CDGgos71dcSy7M5w6B1g2H79MEbubWWHp9X0UfDA1bKb2Svz2/DXdbWgSRjC
u4HJ4weekW3LArE/VmopvozEywNInwgNuyje9WqB+Nv5PvAWIthHce/ph8B08zCqqCbvrehARO2s
0/u9Uru5df1ifQsZoC/308y4JP1tHETn9CqJw6O6gpIjrvRoORhb+1ef5K9tvqphNpJkiCITmPMo
Lg5us4fHCjZd4VSu5Ld/iPv96kTTWonvYoN9WMDLtCK5J+Jmo+atgwwECDRI6JGRhUKn1iVVZVpY
/2jlbkKeEvRpjoTKOKnDHqyIUdLXt2wVF8MXnvChUrTaH4oRZB/Ik+2cMZAF+CLiQaahxMu3aXlW
YjhwNC5sF0kqNPkQe8P7zgTI///X6Xx68b7pC+iy3ENHLikEENg/cUwb7zCKv3mpuM/8zsbT7iF2
ErX4DuksVZiiMkQit6gQii+IcIvg/0YGpxjZcpgnpAW5CecPlb7b3SZxnp35digNUce70AaoatXb
vWRL4lc2VZkXnCqUKEaFjmz+aWhEg/l4PJHfNra0UW1c7Zsumr1D6yNFUAjzUTiqXVWjQo2eiTgE
3O8sljwJWN7h8sKwf72/jEiw5ea0OcEo9tpuZsk27KG6xOskFqNFLZYylOAU5lmPG/L4jauN2HBL
TY3VZFXHgDyIGXA8NgtJ0VY49xtqTnkI/8qIymDJGdxwEwtDWX9deQCkv5NJ6cffRZu+a+4Q6QXo
t1oIIRpt6mdJ+Pxk1mGM/DqUEcHob4rNV3iQxk69/xr1pcjvKyudPXObLz6LluTQnHwrWA7A1ExL
ZzyLTBaPfQvsIvXUYD5NMEI/dpZJLbFLMWhDssUJWt6DyPWeo02mDG6eqmW+wui2JjVX8fjF5U6Z
3soGPmQsFVxzO45XRdb3kpHPvNogG7i5KXHnpjzmPgwTTwB415tEuGS47rDGDdlMvD9+huMYa+MT
L3c/LeE0tz2kwIgn/vf2znRfkcD1fK2+ByDDm6nDTPV3OY7nJWVzhZuUkykS7QEEeeAMnhrpXJAh
VBWpdPLWx9XuUaHbiUcS7+XM2CKpg5R7yyXze1UHV2eDRGNYFWJR9BCTNzJi8iB8mTuBaZpdXtIC
e/EF9CjVYtWoh+LVDN4R0POWXtlhKpkOOlk1fx89HaEp3g2jTe2wRBgtGzQHIfWOUS1L84GDKl34
xObFiZFnAC4vRBuOefBGRL1yW/BVLlBcbGA6xoY/fNlYe27sItxHAp155QEkvobli60tNDUhUvgk
joaZ4BGoM3ca31+6gbPWndKIpn57hW+FgwTWDhl3+lUSTGwmQRrASezy2InLzESMivljweQ17VrU
vt6WsyeE6Lic75gYrxdPasmA3tmE6fXvOKxc1qi3mps6EKByWRDKz6ehmXFNRyfSh/2LwBbmu1zS
ep4lfykO/slueLTWd9zn3DXvR+lIL1fN3R8YkCD2iA8MTW3aTAs3nCcXA9Dj9//iPnbFKKEmZoBP
hmmrDRHWMnsImxxc648uDlQgO8BP205bVVBYcafEer6cO6hdOpiznvem8nL9JMlS22DJEn707k/G
6ul3mPG9gyUH/zvTjG0feDsbAY3UHZITLpvjLjOpRP3ZM5zeIStSD3xXQS6TA2Q4HBS3EofS1P6p
OzKMskpkSGefVaXjbMhzEsyw168UiwZb/yZU9tPvdX6YIuYvkq7ZPRKNxReNqTK77qUEAXxcrIFq
2K3V/cqt/A5KjKtUwhEAsA0GGP+0JU+3DA0evCYghaJc6Jv98JK79v0RwXSF7220c7evJRuxMJxi
qS0MPfsHAer9Fp3JJ5DzZ2zKA7sgG5Tf2TV5/db/8bM1nOB2LMJ5rCFCN2bymBWK6t6wib8LBYcn
eO8VIupr0c0nyioCNaoOusfiXNUOHqePM+Thkjxv27e165B7uHtkQO4Y6iHPpCZ1dHIT8pk7hrdl
gyQYC3k3ab9nQ4U+Wegm4ioCs3J5kZskUBg3tNzOE5sKiuwuaFtGkP+8vZ7gvxbsmCwFVFsRw/xX
Tc5O4AUEpVHGEBTIpLGP5hUC7pqhH1IZxj1eT8Po+hgsdlz+0jgfJva0HGZtHfZO2KCDtSUfHukl
RGUrE87Gek6R/sI3n6SerHXLw5C/v+jOm5yLE2nfmFM3YVpfYaYPm0OyxelyiuRK/UwuFLRWhmoE
fp0UqA29jbeRWVkuh9qacBeFY1eUfh/VuYpZkaW+l2Wt/K1G/1eiDPSWgOqbWNDSMTP0eBxDrafk
ztY1wbOvqFUeVGveIWmf2p6Hp6lyG8Y8x8ni0pKLRpfHSviJVRf1GM923wAofOlMxA3K3SzIKjO3
h+Qh20s5AJHx58eZhEYaDOWdww6T5wUe8fKhk6cA7PldEh1MB0ZA2prkWn4nzwtHzhfmquUBW4ty
fTn5xcdT9ppYJvKT/+yFJ4H9pdLwtWWI5s6wkeyP1JsakxDM0MeUUPEICcZ2v3ev2Tor3ZwDiza7
ZFqnGicez18fQfaxzATgdU12n0h3IJrxq3vjspvegxbX3g5XzRy9i9GH3QZwEtdXWj5n9ZYgk7hj
KgMXAhyeJBjFXNBtijw0V7sih71XMyE+bK+rt8HOxQuiS/xUGqC+RBAv/UDCR8bPhOc84UTmOsTH
GfhJL0xp01NS571VQ2FGUiaTIfM9FAN2LcDAyOd8SuajcT42Tn1LKBfYseJEbXQ1lZHQGIvDDn4C
fcG5PmLt1XH2gns5Pi2Zu6W7fJAaTy5PbU9Z7K0DFLUrAAa3t/7cBBnPTjfQHuQY2PJUQUQ9kQwD
RPbwoiyHh31czOl6MASQtsG35FRJtfDJ4o6hZpI8lTHy9V+demNBrVALkNMW4bkvkShKXrjC28Ms
NuAsqXLig50YuKyDmcKqBeRA058zUKFF4TnaS3dIAstBK+RJr4xyuMFtfZiOjfn1RsbBSXI9mdZs
HeoFpbn8Iuy4KPQ6mEzsbLuoobC6+Mf4+ICzM6+zmrTutpH7k1xaQVzN0gFEaOxmgLxTP40kVISX
G+YIcSvgyNpM+h3hnBWflOuDx4FIHNhHqSnScLRjygoE77oXdqecXPFMeGQClJbN+1JbTv4AjrHb
QkCc/v5tvU5PJtneZ9ELn6YY1PtrDU6g/xXIaPXoh05M9vxt7al8E2GFja4fDIO6PkTTATC6NyZt
ovBAZICn09QmXHc8QpMS66hIirMJepXAFSViLgDZMxZUX6k1yRwL4ZRZtXrnnsY3kROhVbinxGSu
hdRNfsRxSGYw0UoMUjoOpTd34Q6gJwgbHK9i+oBoGBG4ym2NSSjMRV+O/NSXJjhfTbhDjP8H/8o1
yaSRDXKCAfSKa7wB0XUOUzahIk9kzBLHJZul10EPffDRohRGI7FC2a0CnERG3JcXHG80ZWqS6LPz
ZiRgVaydL1DCJC7dNijiXTEjI/sEGjW7Rv5zG5orWdshy2iip7cJlI9OLrJ0fxcDrHYgvQJULnvd
nls36m70OWL50tQsGEhvnbi/AO9NjxNBXug8saYG+QUxtpNrGxTFnVhf/nbWdy5IwnsVsIwlnuqy
2l/OqBPIz4iTq9irmtVJjYZ9Amw+r/50pd0lhk4SpLL6OAFSGH07PYTWpzOsOD/krUqR7Yrahsw6
oZxodgFMp68vwEyrNjr9t4yE662QPuspFH9lXkVhIIZ18IqFsj6MzTP3vTro2DxJXopSo9aXj+SA
RKJuQN7PL+eGI6TQDmmSkEz+7V2SxgfMVJ4mprrnwLES3UrO8qiV2MILy/bYKYV4/TtEHXiMjMFU
Kjv/WSisoCXHV3HSTSie2zPDcBcjXiIK26x/rX/TEPYqnPczhP08fK0IBrKlnHHhPAzxGD5oSfQD
J8+9V9uqnSXzdT7S9gnzVI+bZQhQAS//w8ZC3Uda/WhjJoR8N+2rUptCX9RAHXgOS/stYubWW4ej
FxqVtWYM2ZjjUpNKInn23UWjdfFJ5v00YFKlVbrVFMNsBCXlE8iC9W0bw6SOtDs5m1TG9ockc6Kl
FQ65kV6dYMHkWNrtWxD87eun5KYtBXYfqR0ZNEeYnpyuuh8x6mvrRwRJJt3t6zANWS78vS7sT+YU
CBuL6FskJyUdv9cXRtVGv47hNipO2X/INN8z3U8HpinTzeW00ogpzkVyJB1GtDM93g0UdOGMUpZC
tK4XTsqtO4tOfF1DrUTrlAyjLCnj5tp1dVpI6iV12i5dhl32+3UGPp90QFB2d3Fa9RJUi11juWNI
+zomFv/YFsJBXpLC239/zEz9lLf5Kt3QHChyO3IAcse9iylnxmSb/U03iRDSu12KGiVZYuPVaN4s
FljSI8qXTdld/W7pgsiJji8GSbYd+q/OwjN9VbPOCo8xeptTkwcyOklyTtE1h2qK9OvWisuPM8qg
qtK3LOKrl/HOocYHpfpEiZAufobRB5E84V3++je+XhVQiz98mAJl/GOh81CJjYIztBvBMDxGSIZ1
BIklvVBtPwc3AykXkJJHo3zWIZWKhlsWIQAZhS/zaJ8L/EM46GX3etcFXiEziJPfJJ03ALl8yIXT
Y5UaEfZlwZ0VAezsX020umwWORn2wAtoHIN8Qz0m22nub9IY1AHixT2ta43bQnsFYvTITAJfaIS6
KkdYDIsGU/6SXdJ0D2FsV5sR2dHFDSMG9rsisNI2Aj83y40Sj9kulmQml0O41daZBG5WbNbLLoau
83iKz3ebpHUi29/wtK3KTy6IEwelfn3MjcAQH1bsurFb+s+zvhdjlVHeDjZt+OxqY14FdcqA9pY8
6ULaGVcDmjEp8zLBMLS7iBeHC50RguJEKdbO3JRDKM6sEXRsamK5tJxJJe1eC7BSzvZ+XdPhIngl
A9cBD+UOdF69giyJ2rHhKwrxTjoVQbAb2MfcxRdsb+mgG8tsiuZTzqGDqUkLm/korZerskOPwnv6
6fvs+yXsevKqFEgEYQVtQCgFcRWv+y0YEnIfZ9K+SWe4veiguYjlNVxd44UECHhUHv9xtTH0944p
Gb3x0uY4UHy5DHn6Meg83yiqkGRpjE1CKsIAgZn0UB3ELRZQeHwP7SQ5y9hoEf5om5BSnv93N6eX
q29bjU9VEuanDa9KIl8ueic3HgWtpxY3x/UGAkL2D5NcyE1EaA9GRi2iWDM/YgzcyZgAjZUqzHmb
Soifs1DbXVBf7DkkZcfecq3i7qEnVU/nxbPug8Z9vewQGQHIDN/q47kWTIaKf3uFECLJrpOwXFCq
olVCrFtMkZoDa7zcqX8Dk181/HSbTBn8qbTKb7TWxSgEjklprI9ZVA8lhVwdemH3QmVJ1smyJNoN
DSwXEl2kDHXcBT/1WP9Aeorp0N9Swz/YIManTwdtR2tVqnKXBQEKgogNopJ4W1XgO12QC9rtKZeL
pXQXeh8SzkwBwnkvSkG6aM+gua3zVlobiygrd+dc0H4uObxDWqWl/0X0C0gCTT/6mECOev/jeb8D
6TgXofi+GrusUDHbcgymXe/GPo+/hVgGIZzLwMkDTqdNCM9lvgbWDRyJySxoJIRUMa5Qy6DNI+aI
bFFfQxvo0KV0099ANWv+RXopRYcS0J+icS9OKmUXkFEXCbICcXaz4hCy8kQKnB+Ff9f/CvQ4W4Ll
hhy+ya47sWEUatcD8nc/YsyZfyJiM6+QzyIp8Zz2L+5uQy9v/g+GM7s4KbeJc+5LcoAGQGSi58Kk
oQKqwkrTVUpK9J8Ll5PnCz6fNkURKCsWT8fdU/PPXXpaotTCEQ5kTBoSbBFIj2dQj6kA3N5U2SYg
7jAylgpsIbXIuTG8qAS6+ocOw07S+VGO2HaoiL0xvsYVyNbzyL4tEmnyry4DS/1yuMA6FeilcwEw
sPg/c3+K5PC5L65OSw5LnjPQ0HccQv1XjMFnbjdpNEqFDRkG7ppomb3Vsl1uSf1XEOFRYVOkYzMr
pYboHNlqyMvkaD3E1mo7/WdkCwgoiZQbCzLCRPY2zUI8/t2b118A0O2mrodMLfWyo16ly27CqQqM
rwE+rNYIb1Fl0atkJoorJs0q7RyrLj0LY4yqQgN8sQNx/ege4lf9m7P5hMs+hofd3eYqHM17Ua/6
YGst2OKsnpwxIoK1jHnVYkQ9KB/jUVdttFT8BRu9qldtf/NZWavEEoC+8xYYiKvYIs5oB2ou4eJo
Z0xpt2VbFD3U6+u6uknFtegZExS6pYkiwlMLuBCxgiml5kRDBnke6vd0gW2Q0Njnfhwq1Z9EkuSI
ETy85NLw67/E26S+3lEK2lXIZrar5QG0LhEYq4Lple0z/a6zQ9BsmWlbUlAC0jODMEK9dC+X9+cR
zpynVjpCaIrEU4wPMtrn0vA3HzVzBh8ZKXhhmCDXJXd8FF/EU/eBc7CLVYtH3nYWLBAewfXraQ+a
LjYukkpq3uuAMBcqdb4NoQ91hmp9KD3b338aVasupQnmUpJ1FVN+CjhoP2mgGb1JTs/Esipewe6X
wEn5VcF0/EpwtDTrbfTiBKYShiFqskSpvxqf1xbDQyy6knOnGklsNg/SSE44t7ZUrfQCLvpnfZ83
atR43r2y+1rB2+uV3co4vf+1zR+U80aN5hn7+gYG/LbKySPBoAsSF0q8D1KB8HBc999LEz0knro8
foAN1oOqfi6bLHr+hmle5S7io1gHx8xzPbpv5fyZ7LlmYKIHNKaK4rdqVIX/7qjIiznAbDehKxHC
dxkOunPysdAclurp6lTGxYvAok7LjqraGcLAoSKZvWyQ95OHFJZzUFpU4F/oE/is/NKoOSKMyr2V
RhcWGhuyalI8yGHb3frE3SSNoeSL+far6mlwVIsz6f4vai8WvkVnTtMVArvRrUtS8iKlZUYr7wRg
Wl1NRrxxruKhb2mf5axi+ssVuQbf10pLM7Q1Iv98c3JRdTEsfDEZXI7xV3rz9QskBiyXH5r9Yu7g
eglsCppzyhe3mvit1EjMDqOZIlFr19t5cBGkkIB856BiAH4hov7OyY6u/3z4SqiIgiq/sBZy7P1i
bYHzO/NTsrHgS2WO0RnaoqnHGBkSEplFBG1lqHtA4JmgPqf39rDur97Fw9dL/1D8nEBBScztvcGq
LftMtEoyjuvoy+9+v4VobidqfOsRmDi7Md41Ql2ETVAj+IEIsVIsL8bWCyUf1ZcRYRrRMUlWlni/
MrYWfM6AEL1326mBvwK5HNuc2kWewrQfoQ5P/V/hW3H+GimiS0YY9DoP9ip7dWFBILpp/7VKNLu1
Ynr6gZNcvvfImREbXxv155kXEVtmI6kvP3jx77X09BVPiVqZOLKX4HwLdAKkxwNIU3VP+kt1gGYP
TJUdldWdDYPSeBddW/VFqCoGAB1rP02bkiFu7iALA2Gx0N9ODEfCk2RrlCRo2tWfvyu/9SDr8VEH
sAZLZpkAtzDdqxRNFiFRlTgF/n2wQ5Tw2r6pfpJACF9miV/tdZsrzMWsy3hiwSs/rHUG5Nzw48Q7
th9IKZm5VWcYS1ofaHJZdGeUKzXhSJZccvSLBXKhaQLvvv7L0ZPIO2Xb5Uu/6RaSY1OPlmftVBBb
dDdPt7qAjfLUKttMsRIJ5nr8ehAchGkVfFg+6mqQ0YInibz7BbvXVsOwNgx2GUbiXrPQuEsme8b5
d/Js9Z4xLcF4f/slAo1o3RwMhbcWXvtNGZQEVpWjUwZSUlb53WfN7YBinHhixSfdQ1r9dihVLWmb
jsjemvwRWWis5NswWT1pjqWxsos8TSUbGZx6TIdr1QydeJBLm3agZxLU5ipFj0kGkluLFjzY44/C
okx/9ZXhUNsbJw0fpF57SVfvr3eZlAGv+TQemKI9WG+UKGb94dFLKQSJimrH3BrBqvYysiZtlUlh
+CXWm/QqQD2B665HBHBkC+96VeDn6r/0fJcunasSyjZpNmM7XXtltR2sct7EWWezP+RzW/LK95oM
tmCICZDCpEXI2hJIlQTBKq9x2Vtv2wOySqVxt2Cf/XpVk4qF5ump6aoXRgnnAsEzKz3n5sEgIxhr
GbBHWpB1tuMf7uJJ/2bLe7ehAPl9S1UbSZQcL9fPIEx3o1LN3m9jkWQx/0jNmtD2NHAf0WicKG20
wER8kUF96kh7zyIiv75h38BWLrNouoNypLUq6tQNyx7gd8yntfs9ANa1WyYsEktWy+XDw9OQUMGk
ud3DirdJCnXn/aIrFRQRoLBDJjwSwCCaxpjTulT92hQvM7G6orAZXg/i2pgx93KhyPggmysYPAgL
42Wm7x5GMiSNcuvPWD6F5dmQP0WfqA2VCCZdMBIV9zriUtSpJ7pEWp4lUipQfOmmRnPBy3HI/iBZ
BArTrNKJ4DppJc8KD7CRdYKY+H38Ls/0r983Sv/wZSXI3WnJZczH0VpL0cmbE5T+rXl2h6GHO9Wq
9F+GfrNmuMMx0J1PfveJjvvO5uDoxCEXMavqrtkGJU002fVTVsI46sNkTZ8CXyV8CFBm8uKAPMXn
zrECzbCGvBe9jw++8xtjQcLb8CmLXvnyRx+i1mSBW7VVbEkfaf7uGwCKVtDigF//PN7LCuVaNUiQ
DQ/7YLzNcRvGyqtRPlz0bwtfzCP7soO0cR2hJLfvloIPtL2GjPCTuT7ngNUHaTBEC8/UurD4dlLI
2SHCivcKYlfXi/m+uVkij/H16xXluZU3nKzjL1qDqUp2qdXT0+QXvwf8979uCO2GZ/MumXwcsuYc
Ysm/LCn+Mn8+mVd82W8ExXcaICsdy6ap7QBIqggw8nliLS2o3ppx7XzXCi/J/lrZYtWh45zCnIKQ
MlE7oM6/1mofRTl3pw2xh8H+BCwjKU+fCVbH2jSDEo3TRGL1lnL0GzTDDxe6DsSupWBm9kvmZQT/
+4Q3tCIwMGukqglfALU/SMGyTlP1NLYWsJhO9ZS6JlYoRv/tdcgZSjEPqAJmW+r5PwO/9OV1+Ytu
hyO8Yq+uS1sZH/d+yUH29Yh0tU4/+3iRpnK5NYAAuLKGBWbHG0ZyX24uRQIYSDBej6yDePYhPQbl
SbvsDmKkEwf6o7lzbQTAQxPR0VApfhEHTs8SDJWGebvcLdKjbt5GWPiyiKtHSuMBA+ztPQcKYZcK
jUBsxeUuYVqCgmwYkDIXDJ0y6x0/1Lr0VJAEiAMdlEtX9+tgSp4ckJXMBhCkroRweGzPuhbFVUDW
Vf3rAWNJDjNUnQENnjy+VOTcs/oAvTe1EKH6U3aJtBCVKEwA9U6Lg0LEejxJ9MXiydigFTyi71X/
FL6Hnjy8PGTkTjedzqmOQoukXnEUAorSIYa903n+MEyDazKbEYqoUpiqDeQSDwryAWIcC5s+nebJ
NS1kusZV3D2BT/DMej5iaggOoncTcRH66/4ZyrpPSdnLkDkCM9nFiU3ePywnT1agp2cNC3dCL9QS
49zjKTFvGuMrNRz03ZMiDCZ6afX1JAfRqoGSVu4CA/hdIUkUqMORbdHHYhM+4enfc74jXrj9QCwv
kDiDG/CUbXS1i6JQnK8ukKzm1QEXBnHKqjxMhn3C0ypvSM3PN3eY1pDVuGvFYVWpIpV0IGHQAhlg
whq4ydg4IhOOBVIHS0AzjCdVO7d9EFYeUWWiOLITEvIt4yDn1vwa85HudMjKTCCN73I5OvEWKNHf
KA0VPW/CyCFolOskRyumeF/LOtCS9UguJP0v21IXcBSZe2MW6dOduEWtcbr3nkik25BRWkoY/N/t
whBq7k3aK+PpR4hyBcc9AaeCQBe9IFwybMcRE3+g3gw15JkH07H9CXyDAv1qgKK1zK5X80MLrYuZ
BFEhe9okg+J4r0LY1UGIqnHVFM2hOZVJaODkI2BsTHam5Q/0yHuudG4WXc3YUAnLhsjnZuPzT5eg
TH7ttH6raqr56xEBJ+cu0OBDX5YeqHPYqVd2xJCY7d6RbwBna8YLrzU1mHm/ZDc1XunJik4DldZ4
3IjHi7su7iYUOEUVirSwkFlVFib3385UMH69HRdJ0Q7tqAIVnSSueZ2UfA2k8wqo9Yo9oRrXUzv3
kU+2QNpbYqv7K8BRBYHEBKb1BRAbL9KTW4a0/jsHjU13jsHxBVQdpBq89tfg9eV70k/2J6sz7x7C
XlAqfAirEana5dey0gzAHl2FAlON3rfzT64VdUmxOONbH3IjHzfF8mVu61rLFYjsHKSoRTtOuxJX
wocqzlOi2ELNi8F2uewmdwraE1n8tMNCDwrUh6mae8LxWjvIA6CEfaAuuO4x10ajV520IimCT4gI
M+0/bi2Y16uqD4CspoM0xFGX0HZw7AvPx3WRZImqia0KZ9nDRc73KVFig5T378/AVTCQ/Ie5zvz6
e04KrweGjA82/0Nq8tWxV2uWsGtcaEPVUO+9HQqungco5jgboBjn4G0mTybtBHorajCWunPmX8tP
bE7FqPpglTA3FBiTRRmXfUFJrT0wsLvxMP4w6zGoL7Yxr2acshDT7AoYwimRKmZ+/UVNljftA+k2
AfnjpXWL+QIvrVaSeWQEjbhPtaSgpCVxVupVyf7tAMQidX7MrtK5KuQLxIIZbiNW1vQS7pphFpuF
IHwwRwDNYtFDCSexknkXLzradPlkWngXtOXjpQdpnTu19R/8nq/ZLd+r9TKgpZjGZaGZCXDrm4t7
e7Hu5iOl5iHt7fj4/CiATXbSZOXwpdPkH4ZMOHvQb6rc131HKh6bdBTTH+sjkVbliVU1cjHxQviO
XCz+9UvRtq2HNl4AQ2MoX/f28eEqM0F11Uwcf55zGpppli9OUq3RB3RxrCno5JlJVsO/jnlJSj4T
5B2ofdmIL4yo3WXb05ce5QzVYh4JazdSV7xQB9RF1kLzZM6hHUWfDni0R+/SFsz/VGQCSM0mbhyM
UzWd+PiB+36BvCSZPQ1vXdT2AcsnHrQ9vkym1z0R14rpFvq9oEcCrd0o6pp1dRAGLGY4wT/M0/Wq
skQjaAbAQ8PYfNy02qv6/8+AWZTdzXCIK6kS/ms6M1DymyB9BCjKVvVL8ArtjalCUdbEx3c9+UfZ
sOgb6l7WSBbc/rrAa0OZGbT7ecch4Y2My6ri/mX/jDPKOlAFdOWanDvEDx+h6Gnw8WIuzIvdyzJC
YB2G4jvlrf5AlDi6wPJZT7cSu7uHQpwmh7IGVcpST7rK1ZWQtCoDE7u7736/qnrfIB9NB9PEKoxb
WKDKV4M3uUv/SeuOW1pMGJcxv+6GIIqeuGvALiEXr8x9y+dHRt3S1qV/F2UWrnozia+1/Zj+OlBW
5UsfwY4X8CRq2lyntcvQmk8DLZNYkarK6bhHPL4fnjr0VrAEbfF7t/4aBJxLilvSCOt8NN3oTvqL
R+TfM7uP7zOkoTD/SEIzrlGxOhEOD11T/WN21h30iV+3uYSV7q/ys3LDthwia4S3nrMZvu8eabEl
X4oamQ0atGgW00Xvm5cVbzogep7ULeWlY+Xrg/z8yONL+ky4I6FLNXES+53PzI35IrcypZrNbrP/
/4yPXIRLUdVW8XzbBnFOyMF8+Ghaq0SpZksJ0spNNCotKGOcD2MuoRpSVT3oCB+0veaQM9NWDvg/
/Y7rEmKQRVJ6PnQx2I424ocFDO0kx4beE2Z1kTnudmKWaylSi1kPnxPeUhF/zYPn1+VkLSiKinN/
Vn8mxdwZkA0DbZQ8X2OeOWGpNJjmHkiVV7SWHpXEjfC4ezd92P8G5JJOeROTu9B3Oc2C3T2Yxvxe
5VndQjHYjg2kIwFh48o5e6wTBTaKUrPm5Y/aWhEAs5J8M7qyo3VJE4i+guzcq3OXbk6Ta0rNeNYa
zugCdNvB+fnVEl9cank1t+NnO6qWLD1U9SNp8xV7IE4nDNCaYT3T00WeDkUjKggQzzvOpYZ22a4H
BQ0QjfnED/tUuSk5RjPWBySIE2zT+EKPVeBAwhPGon4m8RfBSM2Cp0xNQ9UuL2EB030/YTXAfcTY
mj9tw7P7DHX2qEW7NFhz6gd4cUtGDLHCEWrKn1I50hZPd+nis3ZNG7BFzamvoxsQ9TD39vNR1baP
ZDQZ7CREv4z/Q+ootXJvFUcmJ9Wa2vx/aFy/XnEfT4ewqgdoCA/gMsyCePcmsMXfUHVmVa9efA6X
tRRqolSuBBl+oSe8lDkMllPHltDnl4jGhg6l+KYI2efslY+Di5i9p8qFP0fFuB+YMX8F68MF05QO
0SNPixtpLR20kmFbOMhdZtJf9VvSruPy9CmTLajBWZZEym5nM0jNfeorBtpsZKswQQ+D13U/qCKX
kYpwnjscOWGYGIbeBK+a6GrTR62/b6QHKk+1Dz5g22CHW5fyaXcs1vbIbYiSICLRl2EVE91nOQkc
yfgHEuC+B6xMBrF2yPvTb0WeRdkhfN73Y0dvY+hLbMKd6W0djCIvZ0SvI04MQYnwhbTDt2XFX7LD
0XFLrSRJls9t3ghi5gAAf+3G25CWUxeKvYc8KAVTi4q9MRyv1mKZYlIWQl1b8As860Mdxuw/jKtW
5iY9iQ/wPnYS/Vvb4xEDHQlJI/GopjDKzn1Ctom7Tx3ERcSogf0mEakUU+axmLnA4oxdARJkTCA5
Z0orQjwMald4WKzZO8NwOCSgT/P6eep4dzNEebU+YLcKVEhOjvnATRr13d0JTNJ+6pVn5herv6Ln
Ywv0IqLuiiohug5Dx0WdE6VRBDRInhw5bMlcysBe1aKz7xlaHSamKaXPHx7GeaJ7idpzpMJceqiG
ljgkQcn3l4CbJZ8vfbToK8Coppg09jiWvireC2GP+Fagw1wMR5yrcTsgXZe8Y09KpCIRu6xVQXyo
7hBUzAb3+SfhhkYZXDT7btxWet71jVCXlW3n0fxJG9oX46DjGchvMPYgxT7u4PV7z5oBB2dee9BX
TpSsZkhuBbswQj7Ot3BtZYRT9pTqiZZE8bQLa0DFu41y2sQ2ZjuvG203wckUKrBV7uZDJx77Ji43
Wwq68D/BTxr3vSTXSj0tw+07rxpRv/Z0iGqAsn8J4vJD5xshidqEZgJq+Ze5ZhTLAivcjU4FoyqK
7viqvmsdS2i9PT171Ku5VWLcLiYRvr6Z+n5vaGiga4lxgh1aPjuVDcQ/JrUjflhakJljvihlLJ//
B7s6xnU67H6pkT3uxzPNgsjQNmnpkyDctmayvH7aehLBKVHCcvB/TuEKVNnu+8mGzRKFvJReIOlG
nVzVXo7adK2FK2b1K4PMPICi8BKmbT7yvU2TpSzcP8vY8+LZiZiCQGInAd2v+GjRCRLj7Z66Rk89
Eqpo8q8WHVPBLU7aNCYSHoXk/yffE8sjsX5qLcdVG1BGYGCAhu3069lmrAGB+5J3YJtqTIqfnbcc
T7FBNxpeicqb0YrcIghPxpiOQUh9Fw9CCayCn7XrOQidwPb266zt8+1jvhp0dn1hPZ55+lzkNs9V
QlmPpkxMWIt84JW6do9DbQIGHVIJY9WYFDUUORC6nF4/DwZcHff14/LnZ8E7kC7WqlqeK9gu22fb
LWeTWTQ8qb7TcnKGEmUjBM4YWWFHlz6pe6si8MWZOcc9yr4H/X6dN/4a6aafMEOsT8SAD9m3n1YC
33an/ukHUP904ualsA/yG+Q7bSUe35RH1SpvwT89DBvC7IEcujjLsU30EdNjkEJW8emCh9HS/JB3
dmw9MoN5UdksDeXnHfochOuLVZt2wdOHhtYaqAk2USebrU1v+kHHmHKg9av5unD/DrcDxZXUgD1e
oZ5Zm5xyq79b1HIlDPqw4eoFWzqNS+LI2RmgmMsMcATKqggbkANfnPNPAlfj++SgOXe84+3KC0gz
HXh8oNXWbcK0+OWiLgKumI+mg2YVUZSAHxbSH09l8dr8pOftMdHVLXoxDsekMuIzRO6wveluUwMd
73pQM67pj5vB4QsJzuclb8ZHGjYlAY1XCymxdrCu4AzjovLWjBlAH/0VKSc/9okaAnG7KZceq/2E
OdRSt5hG5iuXk2vwPu1Dp+BtmT0wfsEAlU3IXBNtc//0hneDzdoGBhk3cLceCK3ae4pM81B8owQK
uZZ2+Rgg/g73qp6LUM90IRTAET7fsYHqK6MXX4anHCPIdh/Sh+8E4NnNXYfa24AYO/M4Aw55XNZa
W/8TJm1BY9vjaOwR6EBpl0iD2Qhr/xdx/0n4uzthQTfzDPanNIYmg8/tfFK6bPCc+pxBB1qK+2tB
0slBD7ehbZzoZxmEEsWVGJz24I+wwzraG5Ys4x2q331jhBVk6Z4x9U8OvrQA1O7yDM4uPQe8HqKB
BRjiDlQ+C2WeXOO56mfEBXA8Z2w7onDj5aAkTzEB90ltRcxfNS0VYPmdbFZrTiVoMVmf0vfA/B4x
mu8hpYTDPJGYQoCFEqxumA522CleNghUQDdtKRG1tpks1qWHz72aQIiJ+KSykzyr90hsIRhPXMFs
ExR5/SJYNrgS9uP2yh34e5oqUBU33iftNScaj1KuxsmWkmax6YabY3EXe5NKe8pllGc8amcOo3F5
s6Fgh+rn+0wcO8HBa1ARlLBZDPnZ9o/37EOooVHJMOPuQURTVrSp/UBObnaY3DknaSw4J1bOagQE
oEnKjjm6ntpE0pbNurveNEoKVCIXr/YNm4ythesnMsQOqrYczAqruneD+tKyv+/VqIMG2GqVzoap
Dz6OHKb/MX+nzXzkV5sHevAk/OgSctdirvErkxLmJru98kRJJqVpKu+Zv90p3IDjDxVn05HYMZWb
0Hh116mB1Pf0kUiOcdRe/qhJ5bxC6zXZ3l0aNLDabUOhOj0dNNFriJ7pLajWeZWDPJDREbXcVoz8
MAOCgaxKYQaRX4NJTXTx8wrjYG7vf4LEF+o7bejg0ERSRzN+NFu9ZYZgU1E4SgnHKbmueCo5mXEh
WHnB8jMpOWI9amiihWntaXymub0zW3aVrsEtwutBLvOu+PYMziTYgVtnY/dR7Iu8ODld25hp5ZFx
h3WCLStaPi9gH7o6EkyWMAe6I5EhHrnn06Gq3JVJWKq+u669HVUJiSOS6OwxUlltVNmYQc+DAF3t
p4p+EV4y0g3AAxY96GK06ROES0Bbp7P8Q9VKTdOPn3IjT/WsLMu3KvSsu9YIAzw80QzH7gIsCbMM
Oz+4pZ7FlzUvpK+To3T6zgDQ49vcXXzkiXlJTJbWE4DwhGD4LmJtUa0Eh4gSXtivnQnxxQ+w7kOC
M3cTp9D1iKYHtG5fchMWBEk//E0EzN+zYCyiF9BzhXR/EbLg+1dCoc0LNXnp9+rHb0r1Sno/Bs1I
LMybVrSCR16XC9b3tSr3oH0xTwgPd30xpkeb/p1fhHFgpt53WerQmNsnnmeJ+3GuaNl+n+WIRfST
fifK32/02LgOT/tOBmfQDjC0t4+VRDnx7lttwIdEnkGMDbPlnIJh6mFwioX8YFeEj4ZIbR63VdUC
xQNUWZZPJoRii2tobCKPA0ErlPgZDyLkiStb0P7H3iVljPBZmsjef2yZ6jbXyrz+i+CpQ7KxNo0W
27XcZNmsnPpR2HhXYX6g68h5N3Z/57Qo9x+bN5wZzfCZ48ZFbP8TN1IBoLnnntpc3FJPViK+MGy3
Vq7y3iRWyfwNmxnrCF5LqibpzdCT3aDsMyEcYeiC3GMiX3MhiMBo1fT8ST+7pVJetv7FWrIT1vzk
Mi2haE8IZjnsFZqeaXd8r3rVipx8+hh85RkQ+LExnq259iXJ/68QUelxCfD8BvBo0QZxY3yLCDag
mSxry5j3/3sEgS6Cy6hXKu+84lyZNLLeP55PWR2uyAYmSazyzixuZ3/lqsQHYuZF9UVGMdONodQm
Ky1Jp09UdS2b96PEGLJhCYTiu27hl1vbT+91E6T5OJthGdkT8P0kVYTLK6/AJzmpczuP+jK4kRN0
5ceAh7gK2nN0FC4+LFA6RbnHDm7ozmoM2u+TXCrZnFysbHy8HstDrRFV/imIHnanrGjH+85R8DmQ
uQY5z1VeIU30sT1QTW0cHiNbHCdJb8L/hJYXPv2AlMQXu3aNKkqlSko6i5tnbUGzWFJ3UWPXniyl
Qa4sx2wiMBdG1Erpj1n7mtd+qakooAj/Us2TqgDTSXZwy9FNMcVKwvZl1F07JvUk7XzXdbdYH4Aj
qlS83WSNpilaxb1CqiiMIHEVD0RpAGGFd65uSCN2Zt1VfWbCq/0zsFm58HgHeWDqJeTGPhsaZ1GA
WjR2YfDRpnEWbQvfO/WJiGiTdkZBLmWmcXbtu3X+VqNCpl107T/gXOb1f7vLqnczhMnAhqnfQ6VA
PHOH/mMXs+oZ5LhRV17g/mdnlowk6M8P/C0JRN/SGlJWu8IUvGhQDJ0WUREozY6dg3plELSKnKxJ
p7lpYhUcfh9ALEZIGek8bGc7h3YsnZ+QLaye9Imt/tGR/+YIkFdaT5XKx4JNIY+jOt878p1WwJdG
RPNeqtDu3m8N7sKik3aHGAJa2bgwIkds5pxByhP9QT5KbY4tFSZj8nHRPzTZn2rgnt0nVsAtwKzu
BIZavtDG74pluuXU1E7tOoU3vx+g87xPLxWA1ehghYfxXXfe2pjfUTGvtNooqVZoIwqmzwRLzRPi
qN+ANLMI8xtuH++AxK2BXMZYk2/vke/2kSn1J/wQihVxtEm/373LGIY4oKI1JaAmJ7mO2BErsEib
by1NJyxRAc76n41qPaGCzkTZDBMjPfyv/apsrAAYz2bo/vf4z87Fq5fZWAZI3QWW96YMNdnYBkgC
kxqQ2Xkb+X2h7k++6bvrgXrfpk34whyXsgjJ7Tix0XsM4gcSG62bIWMoZikmT28DJkGZD71DY0W6
gPSlLJKhG9jiEF6i2Sp3LTu7UjAk9/fZIJMMh93KYpd5gQ7RkEjrq72tjf7rEmUX09wwM8kE1c5P
OCfoNhGkSAGWWXpkPeF46dE5WyW1vUixWV6RNTkDTmE8mPpmmX4Zrh4U+mw/DcM0mVf9HGkzwnjy
/vRnPmJMR6Tt/mukWarDN+1qZyzGXA8Nrx+K4HhYBZ+lsV5z5ET081NTHxZNgvTjLBM5h29mHCKN
Il9nmsj8FwKtYy6z3bs3vQ5XYuxlxCL55GSs7Tp2AGyzsYbG91pOeBq/b2Onj6tgNHDHjr7ioFpS
2dCBOqocfqd7tGvylL/nxJRxlSnCU6aqtvmYATKPjYiIwGXjb7qKj8wensTspsps6pU22XbDlsH+
XKQNbAqtkFEvYS74tqQqh7skZqLBtWoPeKaBegMWk9Esokqb01XPnFX1FkETqS96ZwCfmQ2LKmfQ
aY4EqZ+sDhDRGUXHuacpbJv/OpbSa3GBGMOTT5U8A9awDq/D5m3Xmi11Nao1o5sdnLA6DrmCvjoX
Vsnrd/LrprbvdsUPP7T7PqUi7Alz8zLbkFSlGnuLsZOVJwcSf+WFn98Kh6SzorHgt7I/ix5D3irO
7bDf6HIu6mMcuOp6u6+d9siAWtf1+WSSAWCVCdhEmrpQhPJeEs8eeLiAVNaLj+ee+lqcgVSzXi3F
9naPCDlChDf16hCc9bHh8HKNixBCzny744ZoIsiAsXoD3TZzA/7wr91liMqhxkN8xaHeq7oi+i91
IYaT/xYoFnKJLXTV26S5TQo8d4kaUeAn15mDjDray5GkelRQpNSaVwpIXVs9/YB+fGxnVrqa3sNT
OCW0yvXAQbUrWHFXToJLf+nSxsmsQFLGf9FqD7N2M71n2UvM0YfdcPqzisGEkx/eXZZCjJSOKHx9
WBKXm7JWFSAoebxLfxemvgGMUkfmtAoUo27idYkQt5u4dLrxxM8DeG2XY5iCPbamLvxnwQxS8iOE
TfzEDdjonhi7A1YilBo04mHPB95m1fMBqujiSzwxu1ZPJKoFJiKcVPNMzfQww9zb8P5wg5qAxox1
kbVNssauE+CMD4B4CvwdVNDnZa4S8MV3hKBMS+qeSVPCIvVLn+mq1v5eXE2QeW8faDUiUHVLkh2H
iAzzGWW8FwRusO1UHy4ZT5PONBYBQz5h+ePGqTyJAbhy/qf6MRUFbYKGD+i6DhL+hqg2Kg3znHZF
0qhZ7LfZESeU5oYw34At0K7ocVjah92kKVbR4eu52J0PJ2TuxzYRIMNwMtaRByxTou8yyNbMbgJV
9q0LkeG/03n/kgf9pyShcQOx/TIvCZNEi27YIFpb9Z9f4zo0k7yVCxwvvmAFiUSOCOMLZxC9eR3K
/KHK5bebH8+M6oqiipzskoVDaE9GQFFVvMvzkXbEZw7647ibikfI6HK04a5RxGLzZbv5N2r3xxqV
zYfaD5+s6AHF0suy8q8lFqa+9rFkcI0FK5r4YIA90rYLfcb8Y7Z0RAWOidtzPhmz+L1g9OIu+9Ob
Bj7F76WKqIjIxpSotHHQsUReHcfNJ1jWYe5VXOtlmfAMzAo94fDHGkqfyj1GYxCh+eN0RiDED9tu
VXCItx75RLJJfzb6Cug6jTLtaXM1ZSjddZ3iT4NSdFHc4oWsJd1mQeipXBdW9zB1Q0TKpkkvmXf8
TltnyRH4H5l8H2D7Nx/LCa614S/WaaWZTEFrNO4lzDwF1vEQgmF2GQecc/q/P8Hng7EbTzSsXVIP
Da34rMnRANYF2t3mO7bJsRA1IhQ+VdeO02VDuqTCc2bt0ir501jt0SL0x4D7HaCYz32lEdEl39qb
w7brsLojiPjWCTuw5NMEWsPxAp4Jpa4vOujPFzCY3wZYnz6OmIErihXlwq4FQEcQaj+H/Bm1gZbm
BywQ6Zo8iZ8d8kb29OKGO/Zc8OdccIJZpi6RnDeke7Fbfl4PRAJpSak3lIEr3p14yVIzzyOtB/CL
Nj6W1uYQSKe5nDpP7FZNjUZjagyssGuINikR++amqmbtNLXtGtwfhiO2qam1eRwvVr0koipdxLId
hyMYChj+2N5NfGYcbYTjI2WLiciBwNbGM8GF4LvYruP8mgdh8Tbl4FaR2mgnRAjxH9pZ3djsGhAs
prQMqJKy0AgOelMdmqEOsNk+IxxuATo9UifWKCXC/guz0ZxLGq2NW+8IHveLyrgyCgYNHFL+s/vG
80CdiaLquqd6NuYr6hPBiO5yhSHrmqUa5oCxSKlKMbhD/48l2Bsd6r3ZRd5J+Z00OWiamfePyGUl
JBE3ZEXYeQ/viCVble8DzDO8k5/f3M38ITywnRDdGn+81Ij2smPPV5gPrjI2DJPJ840cRfh/UeI+
S/xxNp4OeWLh0SGSMi+Eloo3+XCLySyMmJ4vxMRwwqOKlhh3H4C9/HJ+evHvnYf/J1oS59427e8z
hOOpR3eDsq55SfeCiQ+b8dhMBBak1FB7zHv4AoC8GuQ1IvFSH+mHrh5b7GXVwN0/euQmH8M/hANU
2LQvbH4ujZ9t3aci+A5CKsK9K35j8VtuXxVdZxKqcGaOKZjZlO2fW0rB+WW44r+YG2VxWD+Gz4y1
OQ8N9N3M78uh0Q4ob2C9cl9qdifrN8wrmDwWdmDJ0eqLrr7eGeFjZOZM25DVyrxcJpbrFGgbLf32
uZ0dM0sGEwh8qCUvLQnqO3SErTtzOvZ9j4UbHpN68ijbHz9B558iAItQw4L9/XmGNvlimcHp3v+g
l5f8XOVSNoUrp6YBsy7UGsFLy09ABj2R6gpeKK/eGiUuPd47c5NUOY8NjBKn3CXBxaW9Xs3TgCwT
HrOB1JoU7OBTys4xebhxafnu01Nr/1RNiIJtTmbIx7r0Fd5RjX4NQCLfzVfE733zCD+iwhMKAo/9
2F+QLBi9h7skfLME0A2hdnJYbNJvyoVTqFmWmjVE/Rev1s6oHL+EFLPpx+9H31jW79xIhdDmH+Gb
vwv1C76rzToF+16XkKtm1omGqh00WQ3CT/DK6FQv019F+03A+jFF4Cy6DODNLY1xM7cEbuUdr74M
r6Hx6T0GQ0acHXpYngYGudhd8maNNd2bh74eUzU6VtEx8qZRiBYaqmeums6SYiHqihuKrtF2BKjW
CuzYzhX2V7IqRdSN4NcKwmdk/yEmOo7RHSTOzdbt+7mgkKSqrxMXeflXn6OEOqCGk3J3UYj+w89T
L0g/QQOcgml3wFoSCvbBheFChhTjaCmXXRaN0qguTq1EecE8qRF9sZGfyCpGeE7nIJuNkqvh4poo
jIWL77v3F5O479uyoik9IrKmGOAlPtKArVM4W5XktMEyy3c5SNCS+bNonFQQgsqmGzTqHcLUyr6R
0PTLT7hGDrVAjRjD4YKFH1ZH7+s4jcGdX+IC7zo9VSRtbTzmeQwOX1wM1jlpcreZi1K4ileQug0d
m2DfOxDK9kxipEewt5VewFgWT+TbaUiLGRugAw3t+kUfeY6/AnSPgUECJeGjpvQstv4B6TnJ4kxK
H63HF+oBNGogcTbY6lPB1ePaygky8xOWyYbIGBB5nWwDzdqEUNe1roqhWr9aZX5Ut4Bcy/nTOq4G
rioEfq2X5J6fzLZN6w1e/kbPaHHkoXwrxzSfYuqm0u35T7ieXnTPqKEuGfoLMeON4a96yJyzA/2f
MHCyxaFouJhpysbCHB/P0IsEPvKCVomBp1zxw5l5mSWE1gUiXiDAVascK89LzZS9jBbqeWmEcZzL
su8Rp6HTbFPB/GYzjQIeuSea63NaTnGXfLBNihJ1lhXUjwdmio1jshjG6Y1zdyZOQoRFxCZRLQrc
2Lzhax2mNuw4YgXpULJ9HkOcnYcRyVkDGesRA73+FbqZm4NZG0dFOLQQbAucd6u/PZcLlgEzJVQp
XCixawQGQy8G/61uxhainDhH1NyEUEwxfiSnNtfsfxb1/TdG1SrUqP/gLoNx8LTJmenNg/DzD/wK
1ezOZQ6X71mHFh/TEyBhRFR7jVHHMxfLh5aBNpcl/9VahCJ89a2DdNIbU3TV8+X2ksI/3ANLtjsi
Tt48aoylLkM6Lbg6hrLbwlfhLfxgFPZAVALZhj/sOh7eBCUX8MFiS8JiPeBIMzCU4tA+5pWyIN2n
rQhhRFEoai5YuDMpGVsRGEOC82HhIrzdeXc+VuLHHejExAJwj1m7L3RyGGvdJRoYUU6uT+q6+zAu
QrrrZBKX4nOQ2UcqA3T33jkVkrsRdcZI6QLxAC+LIyxcP51Hss4+ktf9zf6389cLW7FPHj0L4EdR
19jxhgjVqnqZTLWuXgwcymr0eZZFJybrLRxNCOyYQa5J/PPK11aYa3YU4rDcZXvE30eEby7jMRep
IxKJjp9vGu8rtxkNFlD02fY54DQkmWDwfzEatU+z/U8zlNHL+x0y7z/BzRzvvIczR+CbZRuwUhc1
GIPIQsiTM6DrGeo1LApYQpqXIv1SH7kOSCx32HrjyBa2h7qU01j1OTa3lEjYiGeO45YBlzWJQD4n
/dQk1U5JBFP77N/c56eqX5jS9Qv+/Bh0xVAQd51obs3jbTsrAZv+uEtPvweFDExl5t072MP2gOTV
ZkxdxtdkToXpBYamJtHWPMu7eEUFscfs6KFifbpM5X+FecR231xxdXNKDMYeUsjQXpYrtEzuQMwo
5hP/L1PpQh0/jLtxz3Z0mJD1vS4HJ0X1ycebhYdWbQBZC7jzHslTOOPx6JetMhLeA0WumMnAgfaO
F8prF9QEuH0tPSq1dtMfnFbuUj4ABHWh98/GAOIp+BihZAUpWxsYkZjWKQMlr+J6bJX3EqOGXJW9
Kh5WYkGCHKuj8FvT5xnljy7i56MDSQO7Rw1O4Nz3mXlIjNnQiUch3n+G7aR0X2Y+fS76UE0li7l7
piBW4zMbEHq6HQYBda17raleBTlkX0L9n5oaTP5NMXbcVZsrZr9YTv0jNZsZ4a8UptbFfPMaY0xE
LFTGH7/2qhI0kqlyA/tB08h3suxTdW1WfpzzKddhu8qEjW9xvtyAxpWWn3skkNa5j1j1uZbvVDWr
W5DASd2G4viCtSApFbw34v8Z1npLzXEtiPhAMhpimqUSaqBDBKdovVmbaibyNd9obyg85Ccxlg6V
PkMu0DQAJhFlz+IU24HP9Rmb1guU/IYCjjdV86pNM24dhFsi+VTnzw3CiHsTBj3mQdWf2FIeA2tL
Pq2mOSL86G4qOPYXykfRf+fQLCSEoreY8tMqfBGEe/0d+vCDVNrz1kueSa4AliuQXUUBuRpS/aBb
dqY5rbXre79uNF1DvwmwTOqqQgVI9euIyyDYpSLcpUBx/UZvG511k47t/L8sqavpItWZlV/NKw2p
ovs4xjtZYki8Kv+TKVzU9LcX5X/fKiuRFQNkDE+ss1ysyr7FbMx7lN2OCWCEarrFxQk54eMFQ4lO
0MI1png5XyCuw2oqu/YEZZbPhjE4Wu0QVsWZRK6GewTPMbI+fPhjQWt0AtWht2k0djQ2RRnWyGHu
EknAACZyHlnd+PlcEbXzpo/WWBqh2kueVkWbIQ5ZfOI/3HZDNN6Dfuu86hFilSuqFwudJq8FmSZR
JiRc92dPNSejtFFttUjNHSR24ZQEdfnfWBQV0KU8Zmj45nQxuy2devIRqZchFghPYTvHP0YSWpc4
Z3Xo+ar/kB1SYxVHkS6WAfu/QayBAXSONLQ55QfXuwAevM8TfuLBw8vkgH1X+sDn+JHvkPF8QW0E
/sj/RhYKKlDncGpjghz7yPoSiT+wRBny98yrzu/IHu8RUxyfif356+uaDBFykbAP2gNtf8mPWO3i
brbVd9IT+RrfstoKrhO/gW6uz8LQ6ZB1CZHN/O55MAFSLGY2gEaeFzYGnZTPVyCvZIYsXjbKWSnt
8nTFUMyOgFuNM+kymE0vrbbrQXuAXFILQQkqViba+RJXpteTmAwd8rZP1UGZrSPPybFOVAl/6Qil
MYiiKIiAaOP3NPI4ClBDV/IsfvB7Q+gU2kduHEFMy3/Vo8nKwkmOOj80gJcSl7BTDHchdPBaqMSP
p0kFwsh4KAnhg46PM7l+Ed3bWKLZtIAKXGUIricXTY+soN3Lgplcg3PTpQD0PFQ8WryOS6y2TSbF
OB83SXQQd4RY39cw6pcjuIqyCdJX3rN6jNBjE6HhGsuhSevymJg4C15rXnDS+i6FlbG1a0qWxEzu
HsZoXDX42CUML8K4haZeJhUC7YN00fkEvuF0XT53PwUzgBpcKlv59iru/QEX0VCwg2ptEq5AVqZY
E6FN1z0FSiuSCSDGCg3LKFursNR8mSX4BSt1+DoRLGXQTRs3LLKQinALuaFHcV8d7ekw7Y0dJIWq
yV2cKMTImorU9sREbCrjFZt/7sSwyk+F4WSrPusejcmun5Z+7NSAVKw4R7/NXxRNT6e+92nyscdI
a00XyPPot6AuX6Whj8oJvXfzzr8e2U9+PHAAG75WRxV18U+9c7y34abnth9/094CVQmw201YFlDT
MDwG/OHi74tAPbQvSPb64pszmAy6oZM+TofEjIrf/vfp7TtBn1C0SdEIo+DC1kpbVgRYEAgWPIgE
JtLJuaaAlDkgHp5YxLcd7/3oERHgyxR6Ld5zw1TjJCXzVA37MwsgzoznaYtIvrAiUpt6LQdU2kOh
Tx1GuZWo9nfiwLNZgNwnWvMi6X1F+YO8kmBU20WOlO4rtPMTAw0QxtWUUq1eeL+dEQdGJtavxCaN
Z5tOv4ORKP88ziSIrMr7WzbzpLMk01pha8saVqM66Q9nxVsO8/WQIlUIWDNmZLT6gl/9h4HMSWcM
37dxSJZIH+Je2gsEJnSPNyRQWvtKFP+54dU3JS7RurHb8fZBPuPpDV2VvQeWHxVCqKz/jalGEz6c
VOFpimothkA5g+yAdnh9gN58umjPABdbONwJhsL7GlqmleBuxVkgvmF2A/2zm6aHl4eucaFLIZ+H
qoOzjHC/mrPV9S0Y2fYorUGONFhkUJgMKMtfNKHzZQYa43ihXN1frgi6L6Ogul4WlGlwzSZGzLMF
xaACRrCSKG05uBKdjxHNQzt4VA6ggd5jPkCIt7MVkHIhi81MOyX6hfvh5zTDorKpPXQVvQ07Ibt8
n1RUkQVKCeJR3DnTGJt3Y83nsv8UdhnwF3llNhiOrPlO9v7/ctjSCtICaK++ClY+tQg/eRdchm8Z
t2oeDyDmhrHwvoVVQnpAlq+3z+6k109AGhNQ9ci7n8vDSFM4kKG/FCrCx1zGZ/iRE0ul6ARVdTxt
rhnjWHaE/vOcihC7Tb2fpG+Y8na4CZnRlRoVHFmWyf2G4J/4eNaQDcddEmm70+mL+jiOodcti3Xm
04zrZWXZlmfjTVWKcyDuxbsO5vKHkB1MRfpaQy0zDGevJq7vJbh3J72/tyyOHEbGapmmsevYwXeH
aTOuaN9QbDh7yit/Os3aLFrnqfmwgjPIsUbf55z9TWnVqpkn3/26a85KbMHww1I8R6nDWQmMPlmr
mAL+yEC3PLCIQFDiubhMYLhjzTL5Oh1Z7a7B3JfJ4swtt1PpgP6b9LXcHkwQx/Kt8aYdKczSSP+w
81/CspiGBkb+maTd8Dmfa3rRT2igH/EYaUwth8PDMuBoLvD5Zvofy/5ks28Lj0TLLrrNsG81J6TW
v9u6lKEs+6R6oWfo93UWstoGM4eTtPnq4ai7dqReSziiTRP9He6mTkvqWGvcVSRHgwhWi5ZESHOt
gELrxS3g6RIinFbA7U9eJ7vLqsOK5hxkQs0c5O6CNzoNVX6Mx1Ap2Ad2xyxfD+YMXs5xS5jqjZJz
Dx6Cp7I+vGUL/m5CRppbYOvX6XaqfWsbqD2+au5JDvBmduiZtwW/cMoo2bh1zS8TgjfeIBFOKbM0
IzfVHlPhFfPv5g4Xx07SoOFCjS4amYulY025dkktP4QDR+ykbdV+HITKUOd5SQvGRyiC13WSvJX8
5mOq9neLOF38QyKqBAg4+jqxQJ3ey4HJj0Wdudap9JmBZrL7cfeXvXMIWJRd7XVOTIY6h892ZGGk
XBco5DnwouTMrPSssbrK9LrgWR6TuPKSoeDBVumyDQmBZ1d8eqr2+q2ws3K202oDA30E1NzOJ3rE
gtafXW5uC3qqtx0+L8lP+DvHA9oED6EFOy1mbr3oxTQfL8o00ERF8nLpqkh23tyVpAoxOR2drHgF
Riq03xOgpEuTDNSFgBB89edZagsHvtEniC68WOoh8+jzf6TR50cqFbG1qveJBCdSoUSCEMFuyGOP
DIVMi6SJ+z5sUklIkYfgA1JjFYE7zauThdwwcx4ieyPK7v8Bm4G8nq3IIf5dzr2XAyjfzmnTaWci
iaWwb3FfFilMTso9UL8RzJw42qA+VxTxM7Lj/K2Z3eJ2rzsYhNori7HVx+jdQKYxbUVm2YK89Su8
Y0TKJSMA+6ccNk7Iw81Dp3cgCnm7r9sq4AZAvZ8R0zn6T4pq2BeUynXR6DMWM8zdGFpcmXQJWV17
HAR4Uio4iUaeD3McMwN/Ug3xTayY8ZJe3CGUtAYTruPIWmdvJE5W7bxLgjQW4PDziAz5QQqQZPcr
QLmuL5pK8vgcedos7jIeq6JinxVRMJ+MVbWGUNUzx0lwyV0P62t2HCk1C8IUl7t8sKxImq24gMOf
gesonI0lp2IIfxDD79UCSNDmvGO4PJpkT70RPBaM0M+T96tGx61HsGCPaVNN/grLHRogqFue08sj
P3UwpgFEbHBdIso87XnrjcvLbxDDHC0pXXqdJtGeX3ZsY2h6nELHFYmzNHstMSml7qIFcTE1i80h
r657NKsy1ktKdrS8OKA/nzcnAtpWRjUpnWw0oMnjkLgcx3wBu6HJqblc3dm9hLj/7JmEtByk6MMY
bOg4OI3idVza0YqeOKWDg9o+KrLh1B5Y//QrtyjqOoUZYjQpM681cpQVUQPdPbpE9rIRfj6uM0Rl
llpmi6XakJNZteUTTkNa0UCVroiM6fbPTO+ajbKU2q9qJagbgUQ3XPFXrlwp+E+v5Kurl4O4yM7T
X4h+hRLd+bK5iivH+X7SSOhdhpJVhI66gQoBWmaU502NaUcj15HGzwz96m73r91aHn3SsC72SUrX
gMY0rVy5Df+B0+v2/uMCb4EBoiyEFUoot+mYSSH7aBQjqrpZwXvUCoGeYmt49607bEAKqdVDFIXm
mNX8/POnkpPLMvnx6f0JmQdsYSkrrj4oLFHvMLQYOYOv9JeBI2LzVTuLrpMMqmyaPBRnxUTAVyf2
Wb/NjY6qqbWzUP478+RH19O2AtXqhGU+4enJYa+fyTzOC4kAe32gTkt8Hj+xxqGULxRgPkwnP9C+
GGNQHfuiP9CkHSY2hBwCt4xic2xfxbgDq0CGTza9Rox7ElqzGvaaYfXYtxBduiudRJGNO1oZ3nVG
elcX2godilASRQvT3GSK0hXbbb041md0Mz7OXcqHAjFiva7nsYgFxeDWszUy1Uaw2cUkMDopDDBV
SNwtA5vdqhqDXOM4E/hDGTcFQl4CimFOiWrpepAALHGJCZBX9PVK4pKsyXfE7O7bGUYaabVYboaR
yyvmXvOJhyQGk5FozYwtAvIyE8lagY7F3ikp6bWyZsc/VBD+jUJlRvvISG+879zJ2oD4qERd3S3h
U5j80HE4t8CGZFs+EVplHOZh2xfWAqw0GFJlbX7oXMj+a29UK5gzZA+yAIQkj/rWFjs0WGU9LlGj
vS1Of51vIr0xup19f13WDrS3PGSJ1Fy3epcSP3PtqrwyID+RVPl2coexHhcrkSHuy32INxmEhyn5
p7nviz0EWOEfgqdodw2NuTBQ3SyoMbsrRZgoHJd/Lz4X5P1TqyEMpcsh//yIFAB7Vx5wO2VI4R/a
N9os/hdmfdSF7iOUZEaYFlP/utfVWBG01BqlEDe7mQ5mHx8TDxuvrNskA4WjHtKxYvIKpISqgZla
LRj7KFSicafXmx3B1kvl1UKhZoQoSlL5kH7m6P4DaTLO1LMSlHxQspxgSywUwZUXQ4ccrzsAEHFN
YDH07LAhcX6mwq/kOorA5vXdaN5kEJoUxOaWuiIRNtK+l5kuQXJ5/+O5uO3VXvV7FDP4A2Gjg6GC
Nwa9RVUCXcdcqLYHMezg8uQGzfgX8vWsMjQH9Wq3I+PlPHVLlCA7M7dYyClviqu1HJooY8PKQgEq
xVkx7fCutymBcHbZorIk3WzM0v1kxpT8rZAjaCQ6SIiP6pHXTOlaaoSFhRWj5dzYpeo8vEksOlKP
cM/XwWwf0pjPYKucSIaeCBaouRdAbDh7mbGNjIpm9RiRBRU3mrQaJHyGbipU4blJzVidIbmd7/OO
UXRtP6oQsPytnfyiA21bxInGhkfHxyb7ST5WmoHaBu+TkXvTMuMpnjka6cmO+ZIX3NKigOkGdbP7
P3B5ZVDibimLgCqXxcVWEfTv8xeQZsJd074VnumIMPQsyl41/YZwBrPkozf7GW8RoP/5BVomMxny
RiKsaA9CjyE9nQaFriyjUKHuALu6xdeAjKsl9rb5tTQUqK2hd7KM1EEkBjdTXz8/hCJCrTfZ4AfN
bipFt5iDx9CIwS5dpTU0g9+zROw+r2FbESmqLgNLU6GdBe3Pq3QNbPfsFn35EaW1C3x89FW8T5+F
Eua6kLYQvUM5zL3RWnlNqWtGyIi16xeahyEBrZaixpPoQD5UIrHIDzfPjH9rSkAmUYDciO/US/PV
/O8gazJ4kZO2Vz4SD960B8wtHijgtFjsIusQP24MBtPd//omp93bvTGU3Dpu/xViAH8m2dkmoEYj
PfCBa5SXDaEgYxA2gHM25FY4yJp8I1CF8SQVbIpEfNT3CCUZSx4My30boBNcyJ1qVCD7zJM3zZuf
zSZsn6HV43zsp5DeyWOJwsVfJLt94ocM+YlvooE5DmulwagtuzgH4HQp7YHHST1wPiFbzWZJqYEp
GcqoVfqNgHe6q7rhHVrfIF0nec+kD1e4ebOSSWQHPbbtQSTYlXRwaAit6hofdaW0BdEBAa3KeNFv
oRrYnERIX1QSJ3q4Iq9cfAtWgf0ot02hCxv3OLCeEthTBQy1lEV82egYfEHa3yUn95q4X3hMNocQ
RrnFw7+cIft/3VjkZs/8HuOpwfLTRPBr7LjJn7uYFYw5if5QQx727yb0goDtCP9EDshlJx21dRa3
rEbEHpJcJGPG05ffKXfvdHcTvHVc+9W6WDWc4XxI0ls0vYI4E6vKTyB3DBJlgC3kNvnjaK7cHfh8
w9N4jvdl4nO/y2qUZBcRIavuhoes2Cuseb2cEs3HmfwaT56sC34XlOrcR27aZ1eDZGYe7jYob2Yq
DR3kYuw7GIF9WjPaXHNRpHaWFj2R8yWxbnjQUjgmYmn4EAjEN8OMeB0VqBuXcLbcNmFUKLDnTIRs
Dj6eN8EEKal0C+EqVdw32nd+smNwFAxlIipgpA9KoLC+1MLCXQJszYzEOsFrjqQbXZUlPfRptLyo
4kAjlge+AvVYznbSUZNaRt2W8YXflG9bSjkiAb3SR9kKtzY8/l9vWBd55UotbmK9kDj2FOoJXN+1
tK4aNr05tZWrOP9rKsIShNY72Bcuka8CZvdia6fe/Iy/s5COzEYbaQFuvxHPd0z5JCz9DjFVBFoI
TOXm5a3Un7o8ZDbyXIsZdqF37GofOh52M7LZ/Ui/H41izsgwVEnBqr5/pcXGJtQ5PHoeEqCXi8Yh
WnhGbQuNbc2HzX5T/feftQ4fqoXBFUhiHGJyoy9wcMtXxBlQPVzCcGo7/2ZwP6pdS8NT/ZmSgeVP
1luotgQV+zWCMHKhHM6DdvxAgEDKwPX5HGmo2gMQdmyDZ9h0PbJ5vID0x+R5BCy7MmmtSMt37LL9
NiJyVkz4jtNzwXlAkszz8q53GGo0tqmX3hzvE48JHgh5ZJik5nA+FUs2GIUu2xsD0tG6Zp3uXiJm
q5bB2O/26UkLI7vqShjvbLKVyHGtQJU16NgCLtZZM6CC/PY33ahAQz8bm/YgQLyUNXJ/kDhL7h37
UDPnoaVProytqYvDg0HGnRks3+6D2U0F0hkF2p30lwFb2DJrSUfL2Wcdb/BAm1snNOzLSUlxXH61
axjsJKCId3RvhP7pV05iOyMh8PTppurwG6o0kAO+gtF2yaUbpEKbFtUX9O876vlyUsWVAFMrcAa0
pVSAT3Zx0VERPSEoGaUXpE2B17/ER1zrb1OImwwMZzCJOkIha5+HF860TAIO7vPWGSj2Pvs2Bc+9
+YMhfVvSrZqgk169GfIANjsmtfRxnKvPekVevHfCVXIn5mjYWStXw2FnLE6ew3jkpxMJFXxgaWAO
5ll3eAVVneImb+cMsHKzSb37PzmDHMR+MapgeycyOhdZrQcUNPY+wk1jSBgmffL/FJiwNiu7hRGW
Ti+QtQSfwrZgMx4xu91joDS99++2tXK8Ia9/WZXA7K0dquh6vbd9fVJ8FTD0antrygTQMqv4pGFy
Y2s6rG2NdnNxrIEAvIkU7K0DxrRNXxF2SM705NuNfZk8hisLhYdqcyx0VMY1O4FA1JfyC8/Gg+aZ
VVTQI1ynI4IIJoovEJBUyD9gDO7U8s2YXqOyAhaouzF9VxEgGEQXANdEhiYxXrhIjo6m6zfvp8Jp
eW/ptzq6G+2sey0JVt9mMPlAqS7VLdTyCAsw5+2tOMb6jAlpm1Xu0C4Xg/js/YRqQF3hJVTBVZBs
I6uKkrwukjWPgZthuIueojJ9NFiks/cpVA2R+gmRKW5Hw05UWGuZgLv/YMgoLhghraW8T64mGSaS
sMRdn56T5tC7+30N8niSinJXeK2fgYWpKcMzqnzRU9ebKXW8EXyw5KQB5+A3aeRtpldH6AzGbIFI
BQ59D67V5KUZ+a+wJOLU7JDgQZU9y6i9AvbtlDl5+L+xzwDfvx1ktZ0qHCpJdyX6w9f3OabUXYnG
8yz6LtQ6U89LxbubRCEq9xLeYjv5tfYjcNPXeqAOy+tsPNpqx66IPABVDujsVsfxIDvxjN/z91ol
u4F/njZgNYnOBvh4z1usxxgkcNNjy6Vh0rBBznwGWCFPWI3fb9SOXtmSjz0h7HmPeelJ8u/CiNWh
IdFRKZr4OB8afAsMr+o6mnwoDHxecru/XAjXhSWbAc42OrVhcBynwXbDcrIN9oyn9Y7Eyn0TCZDq
nimU5NVP43n98gs2pShngpBJqokY401IjrChR13fRTi6MQZCma6VApdYBOFZQJNRVqpH8jjSIhIv
C5AHN7/r4mcBgxBfFcjjOyLj12JdV3ywDYCZG7kCOQEjZXwjXHWo0cWo6VVj2St6/vo2EkCJ74Hg
QaPvE7yQHfgsQE1Fn8qa5ZCYPXstsVwoJm7iCmJv7U55Z+WivSTxZsY6GbfNA7OcESjwQ/6Srv/l
rWgLglpIgaeBpKXLUesL2o1OVxs+zMKwUR+UohTVO3fNNJR+xQjSnejXHd8zggn7DLAfxqWb0oiD
LuJKa97T4pKe6coixStyejH45fIdp3WivtZr8VZHnyXRiiPMy4IuuiNAZACekMgiyUwXkZXTq2pF
V0s7x7qNBE5iMMNCnYwwI9sOhu4ycqDbszwtDskJOFN1UafRYy50NHKDJCsLqJMEZ01lTS6L1Ye2
NJQGpGUpBFHZ2oiOUMPDqXOj7+vQkHQ+RVBQfFmozHvES/IdYvNn7rgVkY+SqPaSO2GDqJbL01MR
ZkLLUg/4FF5diJPYBTYYNyFDV381DoIa316Vb57tNc/VkGgwuCkEelLrUQ5trmc+Fspzthz+86oQ
MzBZ9SnO5QjjbPAIO58O4N6AFIpnKq5snDN+Lz72X1UFBdcN+u9zqxPq3nHdzjUA1Z/iZq7AZNG/
+6ilNCpPbisxlkUoAbPgVcikfzSyz2cwlN/aKQY7B5e/Y/IdfwBLaH540K2KfoxKQl5QPsLYBYXQ
TrmRxLn+gYjz8NvbUrmv8vhcXNletYHhHXdsmiXO73/w7kdqQY6wvuVHF4PpPAkljuSP9+jZYib9
r/tl75boj1JjMy8bfQQgkLJMuxDAXqBOAaWLEUwMyWszK7s/AkY4iN0dUsgFy3j7x1jji69+ovli
TRcJ87F6okj/1aEJ8svDXeAKujtP6NBhtUpIwybqWtUaacnBdYEKBHjdePUMoMkpAkE0kEaaWNy1
dW6V26EmVa2omf9jmnwGhvnYoLCqKvvxGhSi0v9VXVKAWvO5mfXZU9uYRYcnSl3Pya8T63g+zLBm
/oj2CPmArsBndubP4VEYL6dE8bDu4jEAFXE5iVSq+kIk2vdrilmzRxIUsXmFAgbGiZ/9vPC80ThO
ZUdOMWQTRzYX+/ytKSSxcEBb7NBUhbQRrmf4lKuNgexS9TQem6Hl9sy7fHLDeeBN878ds/WmCkCE
Io+nkZ9tCLVAlslMUeA0uvwGgHDDiQA5xSRThp6hxk/wZDky65TRlbgAaPASRxI+i+ngGeRuivCS
ZsAZjfgoF93Lw7ZUA6FV1hmXZXwQjgqCaWjcDdNFgBlwOvgbcDUUTkc8bQkO0AVTYlhx2JubM27I
pJctjOlFnywh6PZ4lv7DiqQitoHmDk/hOx2b34OFG7eQjxBzznxMtfVtpk/mmfvi3SExDhQV5YP8
EO8Cll732Tgii5THG05B/X+xNdenimuKN3/mD5V6tRrYzZIENzZru/qF0lOMAYoP5dNhnQw6Yxb7
DwvKLMJDoLtzPfHGz9h8vMgLAc+gYyARF42FdD3SZwbdJ5T5yeRa9+QvhXICNsI7w08iZmIHndpY
HcfRBgUn4eiiaelaM1OXODWRLU6rXuS7tebth9/IDzXqmCmyFiZGdNoISgRI9LMy0B+63cR25Gmd
VUc5+9Lk5Pga2WS/if2QH5kxTkXTI58AGDhNJF7p8nQk76pq7CCVWdSyVcIo5HmhYKYoKDycySZE
T69vhZ5WwaHgnQ4IEz7xwBjzTwuBEN0pKVXByu4iFgGGUK4roCwlBKt8dq/mtNVmgTu74MV7uzQD
bKV6KkwxYWGulo9UPlAG6/5F69N2dUvlLkKjpf3eXKxUfkxBQZ8pJpnoCaIwj2/gqSnneZpFEyaa
vFCi/51NAb0ZmqSgV9TTuWsTDTFJkh8pSwndLVHIlsdKsoURzBX59NlFRcUnR99kjLJ5kKXXhr8d
I3i9rG60PGddK5D66oLewjasORNTy4VZB/90NWgO9Fn1+9Oz8dSAntu19ixUAUoqYE4fHGO75/gY
ZJGt/pYeqf2FBJCyMnjUaKqN029ipqbPxr5MIm9AS8D/Uo1dqIkRMlBv7l87qbMBGepH+0RCwe6e
JAAfTPEoq4S38Em75SvTUvfR1tdReKz73aTkuKzYy3V+8Ukt1fRbJUXI73HZeRV3SmK/JJycMhdF
pZm1UnM/JAyLpHf1Sj2+uWVjQQMVcmy2FVAiL0lTUdLC2eLgxavJLQ0I++cvJRCutHEPwnEmkSl9
ew8smP2qH4aJgKgCUB0bQKrhYLDHuwUIHetu/tnzPSveWceBjxweJhtl3cX88uL3S8vmSuDhpyCu
IftmqNu6GxFB1vScE0Rkf72p5CjQJDyexxIJH38Fz3v7wOBkG8JR5r8DFYIlFot5yzb2AJrclUzN
05yKaARrd/V173eqGaEEgtD3dd4xppBqb27Vqv82t/tIQV8WqzfXeCvhHjEHT9BMk+Wp+dh8H9ad
TQowUv26xlzwhjY0fUuG8t4cu+i1nvrotF55ymOD05CYylphIS5FZQJZs5YEUCGm5axcgEtMTpl2
lwXv90jtpO7vENvvCSpRd///K+pLMYhqHCY88i2s6tE7pqyrK26fSEvmcMm2zysCBXRGKuudg5IK
3Zu7y4ym7oHALH7vFQfQZEuRLaPyMT0xgK4o/uDiyOAZB/Ru0BJExmYTKOh4QMK+lQFk9p+fbcho
0r31mkLXB8Bh/FlhXXjDuPK4k8fQCzZW3O6J8dYq1YHyRLakBHoq32cjPNR7C7Gdu39/fGh5/yHp
bl4u4Ev2gy6E9M9ANQSTSakqeZA/0xgp947QwPE3sctyrEoicDIkW+Uc4xex61uf4mO/K9yrS3RH
bYHh8oKU6DG2SRG1NaHX4r+3domubpxb4Mp+cIuA7HUD6aid+6vPIcs1MwMkBmqePbZda6z6oOrq
8rKK3bgRMi278IDpytCcGiOM0uUiXUm2yzglAFm6x5yNfAGA81tN3flB9n7Qy91TyVNDFjiSlacD
BCCx8TMGMd59pRxjM2qFDmrY1rM8igVHCjNmj0ZlFrANYeWmSH+seByelS+5MOz1knibD4oGI1nk
fMuaR+ml4lP4K16nSS4W19CzkhFNQfqsTC+1+m2LkrKFn6zI3p/mAG4VuRv6ptxeeVu3TZ5TnJ8B
X0dLuhlohDc+TMnCzjGeAwsSt5eMiubcQHoaEtU+sTCxR34SfKZnxQELWEQ8O2oI0CxPgCy7s1X1
ZlIzECFTHwXvoHGJSe0G8MRcjzlne4yBukRwWf7ilE9mAME3z+t0imiireZ0VOmGN/xhcwMklkNc
T+r/soxQl9pu6ramGXqh1BS3aedxIkGsDKEls/z+hOeHiEPWOgoOLRi1eu1QsB8BYnapW2QWl6wU
6HapEeb17F158W+Ib3Ys8q4fU2VXNxYWQ6Ixvhn8sk7L3cGheY0Mi42XVsAwpUzZ+uz1VSOOVX7q
lTzleX4MMHDBjj3PmKoKCHMWRKlL57GwXIXvY9F1cyygt5ch5owBH8tBSbxUVB3vo+hKK6OFNyeq
trupJW/Xhd87ROMlZrTb8/0LX8eIHpIW4PUrz799LbCs5/sKLkKtLmIEC9ch3NHbJ9leBmg3LLtl
OOP2xLaTP+I9Oo5MQ6x4WQhn3fJUM5HV5PDLiO6Zt5s/VA7+pcT90bLIAmpMcVPWNFfiDmdzzzPR
0Y1wX0lWzR0pu143uDKpJMzaYaPNdbUtoW4h74Nj9Sn2GQ7shz5xoOObXuH9BIyV2xvy7fbUKsM4
pkcK9pui5Ba+71cur/u/NG69psyF/TxWbxpw3XRg6FcsVWMsV6ujfj2OdTkQblIIwh8HeR1GLpVE
r18HT+S1oNY8riWfowymp6MYrktmbnvQwTJuW/cpPNXBm8cXMIXsjJOB7jyNGOE5hmkNg9B14YD8
BFJox+9crPb+7ywUlHvN0EIPMwxD1UKgPLdN+AnD/EbgKlSNW2aLCvxhrXLKHZ2VSooUEx+aXaLT
oUxiqv5OtkF2zWV6bM9QISRO443QX26x17vcSBbdJ8hqL0sMbngHMPgTeDMNy637aFwjFt+fGSTB
ztT9vMuyssIBrxWIYsSWKP6Q9DI3KNw41EqjfBQOpj4PoUkliCS0qViXr59EsC7NVrohbeDzuncE
r8SWD0Nm2a93XFEp4edAjtVrNY2aEzkxnWcdDiFvh9+aSfXX4YDaLA5xIrUIVc1J59FsB2RXMR8z
iBMeyCNAbHQYsdWjNvB/l5SNcZGwt5KDjsyUVUM4AJ+sIfIQsKwViqIQUUm5w3DQhb025Oy344hi
QHT4anLWTKauUK5mBxCtNEywcQdRRxQGgH7ZoMTFWRp1I9ggFcJzMLfo0btrmGxrgJBwH4W84yrI
8tXUzpkq5Ic+nliKyCbAsy/1NtwBNXu63X/Zt49OUDHM6Z8OSLF/0Lzd8rAK4QPpZ2rEkpEOg245
3IQp8zR3i8pVX0noNbwcgEUId0heufUwfZWqQaXEUjVqGxAAg5zSKYFY1iw/qm4tuU5CtaFNhy8d
IIu2ulx9JKo44CYi2Fw3ePEqfXwcSKakxQWHKB3Bi5tjsRzZpD1mqLycgZKR/XyCt17uJv1Sc6Ak
7wee6IvZHDjnWGUVsNExQdDR257sP/+mWeMkSo9UiPyZxW7Z4u7XS2GsXxatr+b1WQOn2AazIfBb
GoCiQLjdDcHKX1RklsJZot+fDBz9nvnz056P+JhS7yOO+TYEPxsyuY/z1zuiWCPBoFf3+NVAoUsz
chgySdggnQ4X36gQT3VBOxODd6h89/2a9I9drxxkXqyp132KijpQbI6lHz/x5Z+o8AdqZBvPoKmx
HKsZYmAExmXmTWCKR88J8+R77ZuyvO7ZM02ZZsjNmWPv4F4AYD7OcQNiPZbu8LhZvqeKA7Zy2LJA
FI7X2sJtPNZFRSwLaioK1be+bwsdmsGgyVZw5lZSIw5u6GG+KCtQgZqUE9npt8CGZxzZ5EgG7yp9
0RR0w0I9Uaxij422YArwETcKPKwptojlv5UdQvy3VqsyDVm4tH3GTNkatvkKa0o3zvf0YnAF5DvA
9QA+u7dOlSAadGLoZikm7bIyVl5dpg2STEghQfx5/UOJmcmdpctd8wJs4f4758XDly2iijTLIONz
BNkyOlKfCILHfmHO3+ZYwTDbSk/bI0BZYjyaA+0rWySQ6QDYA62MEJMDfOlIBDg3YkCeYUnKmrQA
fYa0owD6TQMmES6vylTYPKzKmibTpkiyr65eKMv2iO+S5VO6OEgo0GTffmAC7K4feABvFsjTq2qD
ksjyzepGjjpg9H8elMNjegRXMdLvt3iZ1A+q62zmeen4as2Y+k112M8bdrcOKeueyNpt7NgA+iCj
VxLGkSZhpBuMF8dE6kd4xD9CawYVbXQmzAIQ9/iB6Aayc3jmvP+F6wCJo0WgbHuMfNN1PTfXYNZu
v457byCF27usu5WWmwjx6fLFWh3GBzz7fDAoW1JIYdKhnCSNct3/XlGfUqcLdPLBEAr+UkhvCYaq
LsnYMkd+qFj/oE7XIa6nBsuSnRRoEMZPa7vQ/LeH8nptvXxoOlqwNMasgZ+N33w129sHVhX8VACe
x7yNcJ7HgncdqQ5bYeS7ZQDFU9v4/mqraeVIh4mNSpSidWSIMac0TMz73P2B0DIyjG7hWI93hUBx
cPpFQfIXsv2olsE0B+ktzq6k+W/bwgdwUBQxV939NPXK0KVLLze1vdBqPdqmIFG6e+muUkl1x/kF
vVzdiEaYb6CFIk9gnUTrQCOoQBo6OQbelwOQbf0ZIp2/FpuuPLzVxLhzzTCCg2CpXLsQJl7FyloZ
bdI0cpqYmj/OKCWWffBBOR3Ocjc8gmgnknHoyS9AmXKj6vXuSEwRECFC5S0ajTsr3BqUaMDzjS8L
+OUSNW6+awW8qn/NE6WwOo3KQvJcaHPQ7VBVOok29oypXawC7vUac5ayY9OKZD281jn+nUx4pouw
A8KI7VR9chCjynq9RK3vRnHgcOztyiZQtLTj4U/V9pRtGu1At9n920WjYO1oxwxDU1oIWf0h0PsG
wxPJHmaZWot5u+LnwX02RX0dqEwKJ0qNVUDuiDpZzEMhD0Ny9nkJiil1DlwVH8PYQmwKJg16rT/5
2SXH203TT0PDIRITmpR3IDtk3/xXWRkEh5y1fJn9cVwTUaR/wM1dUfRT6JVlvK4rAadRCFqp4iNH
2Gw+G/kU8Zz3KrC7aerNPODqSeTgeG5IfiZZgLQsezAKCPLa2loPcPL9KpGXUNcK6VjljTYb5jJq
fdNgPcbxlPU4o9HERk8eEnj2qImhb0yzM+un1Z5N4mg8vENuYgPZZaSkozBVOrADq8FWMiwWUBFc
IHUenpj4kHB+QyKVFKnlwubzk/eNlQx242rKOXuG0AIK7rnz99kCoQcgneWqHd9CO/D2timhUJiL
MO6NWdIKt200nsO9jXJ5W/6jsH3y2Pw9VnJkopuMHt2KjTGRKOE9+x/7v0HcmHkCDAKQrqW3uBCu
RJO8h4WtcPS48jM2d9ap92ySTCAVojQG88e/W0KTJRJ4WMWS3C1CiTqjbjTGLmqgOUff0Qe2fJXV
qfsudvJL6nnVaB4cIq0+YlUJ6qkyQfNM9urS+bmLaHpkwcrqeSWbH+9pCYCTMG0WrR34CCGPOhgT
xv94mc7Egax0ICaTIshz7TDvu9FRTdZuKHN+zYcKFYGebyQWqerY+5xwePk51tpaJzD5CftwFAeX
unCmzNNfPzg3/TM0+6J6Fi4erpOTS1j0AFq6vN9ejtELERO9Q+14fW5mgIaHZiQEkzwksqswbBX6
uzS3wEJTwuKPSVkDcytcvmehUZZ9KlSLqr0Fg5diU7uu6kaFakesEyoijKFg7Q+GrsvXsO6zgprl
G4drw3x11t6tHcGkJhklNAMhf35Dtu9mm1IHGGFM0tInsFX6ucCE5quytQiDZw2GQ++LKVeDoDgi
8SzHjhnzTHNoj/0krLlHAddDPwrog+9+YPJQIWufLd0Q4dVCNwN/cNZCTkyvwOSnKumdUDipItXL
7bTvH7DFrDh3Yu0Ukt4ZutTZOoNgd1gW9WxrGDdHFpd9ENbk5sFnb5N7Du2S56fQyKgEuiuSxiyC
VFqbj6zDLyGiAbLuPDhbCI66wWUuu8YwmJiAihArKAiFEaIi+nnoKQPTLtQtCIPGrfJ1UICNgNeI
I/pOWmrjW7DZyMMWUM+vkXykelxOn2GFgx9wn2D/zXyhy4Yof5cZ8zrJ98L82VsVz/UgO7IBQ2rF
rb7GGtVI1CRiLWU/rQyE+Q42NIgZDhO4zbA2FJDD3EJuGxVhpabkQw4d7Pmf2zJvyjK3c3iuISnZ
eIHhadCaBQpuRuPhW7eZqrqmSGDrxSsj60AdKKy9HAxB6DxXHVXiirKLHxtIJeMRRXQDxbzwXRLx
sLe4JX6vUqWQGbN4ve6Aw62p2hFaW4pf0xHp68lro6YkivLubap5aEZba1OADzTm/WRdOzUSddwB
v5M+4/T6TwTQqAPzmnSNGa3PDiAzfeVLQuwOvHWzlsqOXKyRJLlXQg+6Zy58U0HP51bWE/by7JOu
SBa6iBa0sCm4iundELx0FuSpEH0BlAea/e3V57KCyFdrzDQGGckxtMqnWdEpgupcyRnuyX5/g9bZ
hOiCt1kV1P3guOhFKbhfl6aVERo7hVTUemSXEJ5k4azVq2h15bAGxNn6ToG+NBcEEMY1WJfEYA9n
OdwAxH2rPCvgKyRoEubZ0p2V6pkEBXylyiCdkpBQ9gxUZxfPhmylMk4KSNArGFGYQHz7twlb2hnw
Ry7BPKG/RDPXzzPnEyzJktntVv586g//bbLtFGfHNs5UAfX8s9ep798yEFHwVU4Dv8iVUUZzlCGx
7as0CgmP6oDczbVCe4ustOlbDeqFgHn+cBFuYa9pjUivC8My17joMPKUSN3b7mO+SL9gkbMS2IKb
wE8Z3tgbbFBbCw+BPL5qxdlPXUVeU1um7lp9c1aMHjJ7J5Ha7ub2cWerhwFJhucWVDss/0Zg05Os
8VxJcSzTP0HNe9uGO9LRr5gdaI7QndnfFHHOpt2GsK5olL8xhPkAj9jFMChlp3asmNM66dT6KPrA
xbYCIUO9ObQvQsi9Dr6KlBeltVk0M+1GrUh3vKqPvY+oGRKP7VALWnTBChAKD0//8nxCZlx/acq9
As/6OLZ9WjhZGhT4Dldv6bVpvQPz/EdWarXB6Xx6RAEhsSG3IkVaCIxF+NBzEm0QYS9Ags/UZ7BP
SEf6zWKQiUO+NKgy3Qi+e6TGuV7vP7JgAZPnOjCImxQHyCidRxbX+zB+BnJc2oUYl2lgCJjLkUFD
mBuzD1sVGoBBwKuMh4JbOkdiZXkloR5d5yZyHzOXfCEjwDBx/28Vs510C6KNwTHfX9dyW60rH0h2
gxtJDlenk5kase3CZTdT134onuzkz+5hYEDGLTg5pVUVPb1NBi+XYP+jl51CNw6h7DYdw8Sm5cz9
gZh//MMYXH0VFq6WgFD2yAagPSDhDGKy36V8gkpoCEZqegJ6F/j8i2AsZwAy68lTIy+Rjn/8TAtM
2i3G+AsFGZr6R00GaajX4WeKozKqtQXaonRJldsRrzV0O5gsTPACi2km7wkvxAoMhTtmQiJ1UkJL
6HNLlFixYNexj5aa3Bdn0oLci/Ro3IPOf5vYERPFvaEd8BkN9QacFKXSE/eK9/+kgs2hNOmvkQLI
dW/zyFxkcDt8NWl1TnDcqVbhYP6Irgv8PPMWkj4mANhTRBTrau6gu0SDNTC/9nSKhFiJkIMozmOI
WTuHLxi/iTdfbiOPU27m+D9Tiwe8igP3PynTxCB+i9YUczckT6kQq42GSrq//mYnt391HNiExH1K
e8RgU7TymtkcXzDUzzcLwzR6q2bNzCXx1vEvY1+Fd6lH2Rx+XOBYas/mFibZY/9UqsfNi+ICnrDU
PvwQbgQJ8VYp6OQvL02wmx0FLJozM57lC7MxfyqFnjxxDuy5sJUbFr4GqwupprKR8v3r6B2j6xXN
KzuxY0GyjwPFSVkyfNMQLQJay2EqMPCRQXmeFxCFZvgsl4jrd2iS+/X8fanUmeyZRxnwQ8i4SgMj
D4pSWP3Bqt7Ukl8+ZoLmCSXGZrtO9XnWuFf4747uiV+RI2eyAXkVtDHMY8reWh3WtViTx84RKLOD
Q31X32BHS+fgOjLAEX9TvRMly5z1l3dPLtat3PWBQkvc4kftZAtS5jvUi1MGyi5Sb7RFU8XHXKlV
+lDGQC55LSyUFd6QiTX2PWq4VcfPxllOQWhqWjI040HdvkxHkONwnjmwQihRIljtM5SgV3nkYKQl
gVE1BjcQOOqqLPpCfmPdgCTeKBTyEPsQeGd+sxRiatS4FYndlzvcSyYPej6xQGJBVaD1pSGFp5O7
sqW2K8yQRanEmVJEO3qPWxgyz3OwpBZF2D9YUaC2SoCFOrsIt71inUM3aynbkXlyTBkXa2esq1RW
L+EiAOghR78bubJWBifzdJhaewXTpZ+/uf+erUoA/USB2U9zAaKxzvzhCoswEaOU60/HwIQCZA2A
wcjwstASwI9na9VNy7je5/YBVTpSJLe4Oq7vF3ODrTQKVb5wkOyof4TRPRlJVSjsdNUwdNryT973
l6ieJAPikExnj75bdnEw5BFQxHASiwj5xOEtjdyTvXB9p1VERSoUNUXrYyxdjXhKcCGDGqkoGmJA
N/EZvafDbA6huH408ciVuloFe0Bt4FEXyDuHqhpCKm5gKncGhKnFDy4n7FiI53a1uqya+Mg2lY1v
gj4adyjJvcRelm+zMXSKyFfIDGmeRCx49e2gDcYHQ2sBMOgooNtJ5iFYksEL3QrjEYo1ki54WQ1A
r0jEKTWpy2yTjGSWvla4lY+SJs5RJKJ1Tfm+TWD58a+Jgrwa1XIrlWELQzuRR2wrgd1YFgWIyTZr
gMDyNslosIfDXNuy++l9A9M2NPPxSgWXazQxTwERlM9SMDOOa+anHW9gg0LCaX3J1YHjvIfxaFl0
JcODsxB+uCbtZJrgmq1FYonL1NRvPeDekVJXBt+V00b3YI6fqjr0Miq6qdca0nLt5xgzO3rXm6bD
QpbGUr4fwOeereEU6ic74kLx5HBvx8r1tvNt+G9dhiMyO3oBlqNj3djLRBLaVKQzb0Pn5SaM9H28
N2RYSUV94BIVMS9IqrAD4yhiVJOLNXn9BRkmFsdO028+YbpuA0mYtlnQSdqftXfSTW0oNfDhq/LM
ljGzTgxGtGj1MPQSuV1NBIY4DfGWMDQfw9gf+6OVyWNIySGMtteTIi+bvx71mr/sdM77r+qbwhl1
byXYoBC0WBLkwBeK2IPj1ZvDzKY2KUrAb57MhVp86XPeEZ6Zx6RZqOhsMwnsIWUEP5eM5MMZzMN4
huK37uKb2r8sWbHIsmlA693SCBhD7hnbTHNscYlpRg19DPLV09PUKhv3D2T978H2TQ1Kc6LonuHc
VocxRxD8w2PMDVGs2WQLu3dZcdyLDdsLAMfzhN/j4idEa2yPV+ooU68ldCnbbjnusl4dHQeXapV7
HpW3mE9rpQsMzw0boIcXEoQAvGO8ht/6MVq4RCxk+MlsARdVJSoNP008OxKLG+VLf/DbDw/CSLOV
jo+wfnrce7BJnu0OdAAntcFKkGYp6HEQJ6ZucNjL8112FFOACW7tA7v/8Sss4pCI6psmnVcp0QU+
yl8RIWpp/Vx0MYiVz+L9hFsedAbRGC9fULJMuw1UUL1sl5740UQIKJjuDmae4qbMhWwYmtjHGWxH
BmMm+upahoREUYZOmx1L4XEK0wcdhRBKah65dFKHrOHoElENJ+mtDoG5uYuyZ8lWEZ7nIcBEGXOv
ZA8TtS/BJ7p5jxJd+Sxe+nqdKhQtIYPY+nvL84hmLo+w4d6DFoeOxDooWts+zs9h/wJle83GPTHl
VUrqqpTbpq1DuOQ/J/f/ldrGBgJK68y62iV3W8GGr8OVfSEXkHa2BcdZYkM13prPwFagzH9NPKWF
aj670AjmIEtgwhn2WiFxMn7iuyjmH7N35n8djZJdHWklAQF+nNRMb+g1rqCVApf4QlG2T0ujZy5+
kI49ZnvUzMyJfjtq8CNVOsZzz9n/87HoVAXPtOQ/o7RAZdwGJ+gSx/dRlDa/DvFiTS/43DPRfd/I
eqP6QCsky5NdaszvWCxqz7hGHhmCSeSE6Mqn3GeG9CHlg7QAemJGxY/6k/941vpmdyZt8FtMo5r9
OPjesR5rry6xsnbMRbuYCTHwX0pqMYYgDnVe4QGONogmTEbhH8dEcADc1gQH2yEpgWwLBFBHtyco
MTUw/Kb8QkklbVXYrwumVJMbIbLZajLVfNu8AnyrVft0DFDG08TSJ53F4juzvxSByUbsw1zLSIR4
bNlPc41e9Dth667ToplSlzcnZYDJDRBhtZ7cmzOJAZOTWuPPwXXzI6fBHBKzi4aYVBochioc1eML
j7RSJWi/hQ66ulvoBVpQWt7siUF0PcOW1FTWJMR8LseRgGd+v2RoJzt05L+v718luWRasfjwNjf/
MXU5kpgJxFKKL5fspyDzt7saWALgkNaaDss9vu+FDjVx3opysgmz/DLtZJnPBjo2WMj40slm0Xf5
Ne9XTvQcfqiCUkt5jLOqK0rdsyyoJrMYat6CQUkrFzGgkz72P5AvVwOdGHIp0uZVzUDlXLf8ZyZJ
B46mSnG/dZuDvLWY+PDLoLzsCszkd8yjxffGcMEcrmiDQVYXVPZLMlHWvrt4U83t89MwAW0MdHxL
zIXx8coPugmn8k1TNOwZkf/l0SeOOUcI86fsBeBk8QwYIv+VN31EKaYB6JqCwzhgHlDb+2bsoRxq
vWQItVtffa/U+U29E9OudvBxrYNofFDEwf4dC78mfxUohX9dkj2+jUVTxtocp9zU9theaPgVhfU7
4/A3Ocmnezj/Trq7bXRIvkz9H71sDnkMDtBhkOIiLdXLkwHARElKTXOVLalDJlcZNyEBbwK4pUeD
3TD2obJXzDyHNeEpbdQOzOhVGZD7bND+QNscKx3/bq6EKielkpJKYFq7DM3Le1kXFT3sjat8ON3l
NYbFk7OfY25Qvhwu0vqLNC2sQB5CjZ0V+lBsA+3C3Gm4isUKm4b7QAEG88eESEvbs0QeDZKRStDR
MbLZRKtd1d0fH7TFs6Ql9HPTf8CR2sS2wSiN+4KM1Rxo0a23w9/91xoSJLEQcKy0VfgWofze6DOM
w0Xtljn4r26ENhc5tHDMN3xldjGsfpX4M50HD+OM4x704DgTzlZYH33+8i8yB7a8JnBPxcj2hNCp
S6SQwspFVbq+ELBC8GsltLkTYA2c0QmVpwa2uKr6SIkebW8FL+PWus3f25u54ydegsf8FtOMmJrz
Dhk/84NTE0HPWCXwz69sE9kTOQEB/06SM0Pl4zdKx5Rlram4TDR+eVRgfw93QVE066cGxxxx7DWQ
UE/DzPTFZFPeLLI6efum2B66Ji4Chn4O0+eFRmwWANojDB4+0LCMWEqJpbE/c/Mk+nuxG2j8tHij
I374+fVyiaXS5kvbnERQfaUmLmx9HaZiIAMHpc8+V6q+o4ksGTHZF0gZsOvMYZ2eERK5oNyCyMkt
GBA3/sdtoa271E9aJx5ddh2z2EosUTgQSSBin4+ZTIKJB1KJwXQBKKqA09oraRfBjJdtJfPZ9MXt
q1HjfoeXci5MUmekSZjgx6Wx7stNZr+etRZeN+Nf98bbv2snNUBV7pzNlR0u/jy2suphB5Bn1XY/
ExOBCx+knD/K+LcoHfwMz+wyZ7DmsOvu388Zcir32fBScDPNhETddW+uG4VgXv9086UG9Vm2XeN2
ePZemjSskBxH9tQZUIum8Kd7ax1cFfwEiQIOCKPzZ0tkVLxJjG+9gjDOqFUQAT/WwkVpnZNZkHAB
zNOv4qTEpN1x0INKr6rqhUHJFISLlX2YMQYfroe/8rae2dx9s4yuk0ymdE2ofRXF6D0kBmkuQPX4
V5XUqZlx0C4lbafLvdwXiBw2wBdSGSq3jAwZr0CCmeUvQDMEtey6UDnPpmcw6zQ52SX7fAOSSSUo
hXjRGLMWXcumBssW8j4tDSk1X243RDTWtsFo5J911f2+tyC7GLEwYQzOERNtxqK7LdBrTITLgRDk
H9JFyeEteycHn9mEBbWTnsTE1kOeO6ehWzNmrq+deAYKenXWL6n4daHaaCW5LgYufBcSRvkRKRYB
zDXXADf8dpxr8PnNSZycNgyKUkwalKDNVbPiIL/rz6gnVudFuUC5W0SFR9Gyso+DCqhSWrSuWa8J
6JgtE/Pw9x77uEKYkB5Zo/6J32jw/OHqjp+gbqS6GwQH17duSw4CZ0uU7nfqsOOP4WoO8r0qBQQY
4OAfRbKsHs/NCXnpUhe6S6PykQihbTLK+pxh9p8D1jwtMwZekZ1hCXQsjdlAWPk/ZSCOxgUBwqyq
ku2bSU7XiQkuPlnW9g5IAGdCeSzKC7rzv7qbDDmp2yMxnITX+aY/Qf3nL450UN3PJluvUAY1Xh2K
rKASAn968yNp33jYfX0U65P7k1qcJTHKhuztvrF7Wpcpf3CCQeJFKdNnKv6aQIIoSY7XCLxYeqhN
w4zJZXTR5jsWG5DdeUIzf+tc2Ld6FaBgJFfGABFZQ68V0cyC+vQ03WTTeKNC1emFkJOC/W9WBPmM
l/RyoS9by9RqQKtYF7ZRzcxx1x1x4VZhZtpP4YZJg3XnUJPHkExrCSE+8wp38F2s3rHvuH3oD7eS
ey5/7GF1L+QcsFkh1lzBPOmC0Q9P47bZkzHc5fCJxLwc7BYx9WCKVwJwDjRhWFXONml+traE166N
B6jRkNfzra+q3n9OHPqeY0noWfYRlpc6/ErNkKuqea/sc0bpjgLOs6yufNEVLBGiHvBUCWG3T/ye
veH3sgfkWT2CI52Ufp8t9E4iUmSAvqFYFKkS0TEVm6Zl4NBXoYW9huqr6ubo5ElhdLEdEJFQQNoB
dm1XyarznmF+XAYZV6rLcI/ukfk+2cQ5T9XIZ+T3XfdzNw71x1ODLNEbSbtwgPbzZIQ1IoPBxht0
zLCoaETJGsGu4q3+9b1YOPAaaVQZSspLoEzQmlWMZ4Z0BJ+Gdllzb8tXnFwJWch86I/EV47VmOX3
73ul8rdYVxU6WiDeX8bmZuL9NzCj6I9cZmJajuL18eEOhAskVCfRdmmVRFQzmlIesKphaYycMCwk
gg8KfiC9oySY2ES4prxs1oKpCksa+d+/mQa5hXenFmzVns9JY83572l+gQs2ZKBet1eqlTDJmgfu
v4g916GEtYz2F6I4qWn6oVAPRq5MzR4qaoPn3Y39PRfP0wb8AiwMT7i3mN0cBn/MSHVhKRIAxEmm
o7BkkznahXPNnkRXvmt0fbYq5mnEU0odKAVNqLN0RXBpkn+4v2TNRAaDeP6cCL+V4L08PaNsVxGp
lRgfWfDNUk587M508gFP6y0Pk7GqDemg0md0++j3oRoRqUuevbByPak5qGTDj8djRbWH02Em7rBf
mQZAvhNCmqKvzg9BDIGTP0vxXX80e/FGiCWvVmcbzAkYgPV00dZncIa6AVsyMBuwnXyHKNsm9Wap
d1Hk9JsGMllLsA7ZMGPKDJf8m4U1zyJRyR6OWTJHJz2ywdn1lfGvGxp3N5Qk/MhSGco5Nddn9yJH
+vpxpYyjV+IGh9ViwxGupkpk4+yDFCHdnTMvRKb68F52jRCtEB0LfAB3DBUC9nOF+iJ+OWVfMncs
gU5F8aGZdw7hZygQMHDCscpmx7Gl+9SznfqTY4xVAaBR/LmMp6e8pqK26SbjyEGsfJ7bQH+vjRiA
kyMgMdNIlG4dpxi2hOSX603a2gI72+O3PgS+/oek/qDQqfJqO1wU9JX80xI7uIdVbKYRN4fQf284
S1TvhfvDW8+SVytxqmFVv/7xPyJYNYwZ4c86BvB7gJtfuxehpGAv191uLXxsqJJBrgE5JkRw6Jti
VgO6qWHzaXtmNeqo8EQwkBa2m3fO6rHRjQpFFU+67tfgqmhmKKCE3nztdiyBDMVI02dZ64powtM6
W7T23kyvIGV1wDgYQJjlQ3Yyjy+Bh7JzeyROA0w6r0bRuIFqrfvyiDjTeSkl+thPEXhtGCd3fkRg
It1unBEBXaRqSV6VR5RtuT9magCfu3AosA7pephoukeQJo5XbZaD+pcSE7aXifOCWDHAZ45qGt16
anTBLFOu1dUNPCt9spxpj3SbX5wzZEyPXaFe+LmLdJew7GWhnRrnMnpyYf9X4fcTT+b9UVF6F1iy
1erHhkgbZg55Cpnni7OJmczXN5JSTFVx349ptsV0rxC9hLkWVZ4hoavc9D/YCTt8F9StOTMYPMJ1
whNMHIh8kju78afGRrN6GIsGHYtMxn2crewjobB9rp6QRFL9kIB1utRCYCWNcACSu5f1ke8bjPen
oA9uOoXquaWqFb83YiLi0uSY0rIjU6nGmDuE0RvWFeUiOoXO6XP7uWeIOYqzCoCQTq2nwwBA8nnb
k47B7l9AaEKX6ro/3OL+CXEU+1th86jFQjy1ZTAC/cBlg4FWs6N/RUHl6aAiEwAXXYvB/g6iZYEp
LlcIT8jS3u6B58l/yntbUqG+uahPATDimW6b8T+SQb0uOLB5u5UH1okoCQ29mQO69qoL4rvBEyU2
mQqwxMAmAG8/c8tdP4i1Cd/Co1576lccR37BTMMEH2q8cPLS0uf2FnnGSfv7VVAEdZ3B9a1xjeUL
a2EbAJrJqzYgSa4iupsCcRJ+cWgL1BEozLauZnB6mZZXUb4EQl3ephPEvJXgJSqrzhrHtrDg7QJo
oQMfwjXLfTLPYg/UJtVgtFQs0f1tg1T2RALbfdB4PB4EdQgYxU3HBO1ygSRMo8cT1oGEi9ORfGhb
f9EbFdetmZ1m7fMw14TMMru2cd56s2mIqfUNMVOTR748a7x23q4KUV5552iSRjxMTTApZ3ZM8TEG
dMMpW6F0u5vX0qwcfo04MNOm7zrjO5frJXjIXTe4n0mV0VAim/1FsFuVyQmyiGUJ+EGwFlL7Jy1k
/kjZMcSwehipwO1PpHyr7cr8COEYiYE7R0Ju45YcuUjoPXcSUVLBraDcR5F6j6dBWjSKAvJ13vKf
c2j1mAZMnEeKRUwKiYxwXgjxpVnXdHPOk2x+hsvGRDQ+SLnEbRhtFO9namBj95OFRKxWm+ZhgjGc
3MgcX/Ycqa9W4B1G/Ji658Cr7+iCXQgk79fce76+6Y4masMVoZA3ov07ghHpZ/PH+ukITuSxW7cs
MGLnoeEIj7aNmJKItFoIAJ0ETmoDDcK+RtV2M4qpUYLcbc2AKgdGRz8gNatd2L+1tJ49ICQUNGk0
gA40RJMrSbuvH58qrW+ZHnWtXnJ8DBTHeqWO77Quaqf7/RM+V1rDvNw+IQHN2ozlLAA2xAxe1Orz
LS05+A4te0utS69iek3eUc3A5nf7WcT7OCOZPS529E57E7IjbEJpXEV4SYjgIDNqqjMJPemqDdK1
IcFtXtRNdNOkNbjMi4eYyS7F2rQkF9V/0mFJ9xDMGspVyV3EiG04Ax2kT+tfBwURfikujOFRyNv4
xqScY0S4fGO3DcDNNFt6/0MhHI5WIc6x5cx1eeDIEc0qgJKnFB9D1C1ZhXwYZ5I3aijKhw9PWYPO
FV6FihuNhvlMcz9Id1w0nNZf4zb3JRLpApWbRZ+5ejJHmj0bvDA7pvFI0H8DmlyyORYMxiR9H9M/
yZ+cfQmLm8zr//5UazdIwqsWS44ibkTEOcrnddAJpturb81aITKm2F+fAZGaYfzbc2yjS/3cJWYS
bYLCl3xRnT19WeBGTYbziKHRXDoGLiL2J4+o1oFJXX+g6u4pBrGRWiiijFYL1MJoPH6OGvcDsIbK
wykDsWFibC7LIh+yT/q7fse2XgZ9LnpJvLC0j6fyUJmOdMe+B6wS7shsQv0IUBnWVa4QYBdIRs/W
MJ637Zhlx/QopDQ8+QDLYJQUHSGtr+PrKo69FJqyPyzsQzmRtQbV8FLZC5ssvpNNxj2Ou2IiQ+oa
J06+dCO0NJTfXdlsswQKle5MQfoI92FFqnS97QQMoQriD666iqkR3BwKYq4vEJHvhrQ02Y0HdHE4
Ho2lhHi6E4VIT6XYW8gksk4JrmrJ4Qre5zc2ZkySbOZRfMIBmwPi6rM+oMwA6lEZIfq1M9vvQWCN
eSoJfnxdMBmP1MMy+fEVXwwt7jZzkaAGYUFKmJhNA/2bf78UMSqpFnkBr3ZyDzpaBfOiS65OmjM4
qKWzNPTIrYTv70zu9WwuisPhotof4kSg7B1GRjUkI5ggoIm0sRSSN8rvg/uPJmDP0TtO6tlfsd6I
CXNOE7Rohq120lTz2WriMY78vd6AjrWpTlOvN9RgCBzvssgn8LQWZ+7VgBViR4gVbDqoQVSdkljG
ktphFZzbqgjnhAiuhXzYPo+g3LiBC6vz52jD0O4dCxbS2yAg9b6y4n3NVH5gElQ/BTa1LjN85XQH
WSf4SAE9z5Q2BtcGrwyC5j+XxgxO8vpY6WIUiKey5TwID/Wj1fbeTuz7qOUUKtDRxHl3aP9QEVmC
WxAMNkrvta2AretSswMeIRmATk6g2ypFNibzQC2Rnxw17RCImDTWQD4CUo+YPe3Xb0IVkkXjZ4vs
ZWvd8LmTfOQX9W8QQOYt1XhzcyjhRFPSLmW31v9f4P2COI938vY1yyK1bFPEHQjGKJidIKCBLxfV
WafVENo1vy9cVMTIwWCzUiIW7Wp1x6eoWd+zjZfcW+BPnY1SWir9IpGtnVVHq8VBdJbOgaX9ENOV
Xh2TCOv6vKJO56Sdv1lL0pZW4DN+Yi6fjwXLI4JPRulxRqdnXw6+u8NF40GcLSp5pm57IhWtpreb
2bLpxbdJshZDFGHaBkgb2IZSQCy6t3H1Fz8v7+ZkOiI9ufsGhlSrRuyVQ7KttXA7FPkXKqwbfboU
oSL32zhBPUA/buy5ZHlj7QBJXvjvsLmBDIy6cnqzZU0WcqqH4z8YolVEntV28IjW1NkwDShYqh7H
fPg+o6/p/kYHoJfUsIArMGQSRt/5xTkYjBI86l5LHwv/NLZv7b2qgW/2ynDquocvpAYHGhL7RLSj
JZzkFNPvrwBvu/vItuXLtcEpvoUSq7/1bbMWb7vYRT85e3XneR9PFIZgL+a/A1hrSk+RcerN8fod
fp+RCd/CzOrInPNqa9pD5KfCLTi++CzOoWYfcabbqY2DnSOIqZxpsZyhv5fn1cZXL2+4KmdcoTUD
y+oRA+bX7ooT6Pb8CwIFHsX5efKCTmsgbb0lENDUASp6140ZvyVDELH43S0IY/4/UuXH6rT3mXEL
DzOobjdozWqh5kBI8uzgf12dYSxdgDTPg1SuliVn5/uJ87Xj26b50iMS2LyN3jEW2lVR21QENnM4
egaUOzNCpSb5KYwPTHF23N8KoCrF71w5nEfpJpTwGTfCCdLEJyrvkCKGGT35Z5Y35F437n+GwwJ1
5M/yV2W1OU2XuFNS0Xo/h189JSgX71f1OnFRu+nrUCyhY4tEHeEzitsg9xjOTJLF3PY/Sm0h9gdW
xoT9kZEWVqNZcoc/3L3GzmfUAA/LC+jqlMZV9ycU1ujoeo4LAwV2Bdm2ZyOSoMh09YzYr4WqobMj
6D40D3qNAiA0gCRxnwn6k+k4C7CfFvf0iI/7oDqNZzZPtU6Z3mpBH84BeMxs1Pnx9oVcEQjRj+CO
exr0A00BycpmdGdmXF3BhRIf8R3sS2pAxZYteShVdNBFxFgc+ZhR+kkbOIkTq6QoKTWvIU8Ab+50
0oSTu74R/X/12tjPnUdzLZMRl4yuHmtyBoKWvOIb0wPcxykpn+sRtDNFwQobUCa/bqrVrAcr53s7
OCRwLjb3d6/RVMaSzZLCWS8uDTNtOiMj+P3W7n6GANpXunhPL1t4r2end95gbnRWcWk/oDqvEqup
mwKhHChhFmp4v1sVBBXsNnUlDkALASkh97lNCqZ7lj839cVlTbw7xoU95VizBJR9LiP4NuNjUjdg
ycWoMFoIPjfr1yn4dQSFL6XjQFnud0TbkoHICj+Y6/S/qjOEnMKeuASwpThxQWYMJiluqnSa6W2L
ZxEo7pKREAXjOnmZQUav0u1tK2M+fALBtNDjjRqxQg+U0/to+Hz4xvLvcZMviV6G7Aov/VR3kLBj
mPi3CH+8cSesl+KG6EdnMLMMaP5QKu+Wsfh/cg3mdwF4FMTzTzMoTnSkg9+jN4Mja4FqEzq+6ZLK
p63UMG1k3xfR4UAe/Sko5r6pvfJqFgLN4N2xCwa5azKlgafPelb5eMvrUtetvABKI9yOgIhD+PM7
Er58vpcxFSoot/BT2qEHO+aoe3DL/BV36Ab0PniblPMQgWCzXUv4GDabUP0YSMWKPs4rl/XsOGou
hCrQRzY5gIs7DVp31YY05PeEKD6eSSjjeGqbNpYE8E7XokHeCd8ztTNp++P4G0/y3Sq2zEZe8jGU
TV9UKLy3ioNfzsHouzI6EKx8wDwk/8Y0arZfmFJkons4ou+4T0jMF1uqBt6telnDTRVXA+nHWc12
SVfoJqtcg5BcO74ifNyBPnTZw8RC5XvciDgK1PHmlPw9yGYjaDEo37KaMeiuJ6m3b6vdX17ejL2o
GfI1cnOshNfdMZx30fs1TQya2Z2ptCdE6xTqBBvXZlJQKzwGzMQAVpDNlFYVE6bJkJgRQKzssSFK
qx+JVvsWfKoQN+j6XI2ZqQRAtgNN/QmgTJc5bVWT/6LKpDV8MAswJcOMC3dqnpXpSh1SyZ69UFoP
bAlAxYOceUcf1cPJ9q3cvawANNbK/SQLbOUcistlH8b7WzJDfyYLIH3E1q+dl7qz8gEf4dkWScJn
u8ZiJOUPXBl0oRpN9ug51cQ4y6ZXL9pm1rIA+ONQaaQBs2DrajP10iNCLfa+LikSy1ibfc9e4pu7
c2HW+wNQhDk1R4iAY1kDuJM03l+WUR1TpkGRemGzVD2iIUphf4raEEPz4gcaJpUKfqi0miQ658Jl
67HMLpWwT7eHfpVrh+bZEIw01KvQjyn5rWqGxzmt/iG/pKiS0BYp5D/61645evnDpE7uvgTOGPZL
q5MAIbF+vs/PgwhsZeDp76c3BYaozx/fGOGoAUdRv9KnE8HaoJnvp1DMy5f/tLu7WCff+SoPJHjg
SAXPzgqhxU4D9noN/Ur+p+xk6WOLQLS9E0euhSjoMzBJU3XNVnUK9Ifa82lkG2gpUVppee2ErVz9
mHv1sclZlNnaFrpqEOyTJgu72Nc9DhKbnedh8uO3diWdozAOPdmh7Xk84wnEwHlehaI0ikDFYYqi
kloRlXYxekIOuksWkbAznbLWsDSyfAmDAXRNX+qQYbKM9kmCd6HZ/aPNqKZXV8C5b/lp9RFnZa4C
NDmUXeYnz/8v4ZbHLP41ULRbPXSX+D66plc20xbEk3+Ndy9UQDGk7HHUKf/S32g80y0TlI6O8kTv
K/6UmevnIbd+qEKKRoXHFttxHFMkXpsi206JO3wJzGut2137SRDhzNh4G4IquFAxUM0FmNvbI7Ni
tm2EQlessn1svzpeLN+VxnXOZZN45kU72Yu2r7CuuQ1iMjWNX6+f98+fzciqfvUtTrDYT7qBadUu
REUWP7xPFTno8LUKQVBLGbD9eeBmM4f7x9PrET0KTxbjNbQqiGIWqSNFmzmGkTdQ/6UfEZsmsG9C
n5ytr+H6bc1JzQi5SP2G0uRGjLUaAv1NEoSmroDys/rhwrJ+sVNVT2gqi5xf9oyzQsxRVwLXXXjL
25bX4Gxuhc77ftPJ/t5xTP2vc+AyOOlaKdVGFm9dF5HYUWY5rIoRU5G4bOx+Y2zUZiyenDYQxefE
ZOUTv2XZCgOzyw5zNO/FaoyWoHo0znAMBWundzQDXedgrt8swMk9PzLVvODZAZwQMcyzouk95haq
u49zdwHS8xcDr3OFJCs0qSf+3VjFKz9cTTSkr1oaunVI6Wht0D6Yn2uG0N4dHOfwM9ojnapPN9c1
U7N8cxUE7WG4ZNe8xzz7M3hmkci9uQM2Srr/Cpl7ZpjdbEskw5vjbSS/9AVvlHs92/wo/nXKYz/G
PuX9uUAR42zUEXVrBEgAC0wNmKszaAuCgBYrk2a/GHOGQQEg0bn6BR2CAo3LMuvPuTv5ly95m4lm
ZL7sEVXA7EDo1f/TnG/u6GG3BGKk1RBrXvpbcnA52t8D3GWFAn0YrxLVPR/lnJ44o62c848LFYKS
Fwuvm3/3rO5uJfwHB86dqwZlFLEes3EbglQvI+kC4kCOtMDjHx1WY4kGSigx0I5vMoCJoMKjAWSR
y9uCY9ye4mLSAUmSlE5MubTau95O3ZxkOdbZ02zQuLDoRwYa1LeczXVXvsdhTF3fGDPsvN7ls/Dh
WO6F6C+Rt8mBD+EeKTkWLz/HbSwd8b1/wpV6z5ACxiGpKK7UdftyTKgGYCCMH3lIjq7sY1+pGVOo
nzy0/9XSSXO1uDRbvMB6KGhiZ7+gIPMJHlQfovdmQTBio0oLJu69Nn4dMQgtBoBHxoKwfAA3DNkE
4ChqmH+FEIidutcM5lFDr8W1q+CYgfxgqbTfqe4ASYTSm2gqlxKbOAne2RA+NrIaYwlCw+HDYb2S
V/J+iJfjVaR0Fr7YyjlUxG6GtOTrlgzaBLQcUO2oBUFQL3NnAILosJwPzEHwVj8wFeNN1a0C70Ua
FIj1EqZ9E7e/b2XffHbkeAmExJzuunx0RiCoi3Esr9ZZv8c8/N/Svgn5EX96NOknMF98CVFXRvUu
LXiRyaIAFnltXg6uncJ3Q4T56oAAEa68vXXJeHHc0GtXVjJkswWKSrhPqzOxOMOsHms4bXISPyi6
9nAd/McjgegTNujunY5PMysubYgWlEwszv18/RlXJFqLu4L6rAljXf4zaA/CpMr55DWkR0lLvSV3
gl5HFuT5Pfl4qNSV183FrfGtBPCA/juBDkPKF+31CCkPx9j3zxDW4NGVyDj4iLY0+kiNH3Huy3en
fvh5tXrT0CMhVaFJJ1ZKwUEbe5Jzk0/voIYz7X9g0xaVrZRfdFMUobdQcZqSIda1+Luwd9/swFkM
n5PiK4fSTSQn6Y8XF70w9b084VNniFGF5GHYoRtgUos0uJ3nKIc3krZTnHNwtpm6zgklTw7kSiBd
odqWYSh1imVO/jY5txMBs30ZTEUqMkfeeS/A82gr2DqIXTVceawiSkPMQlgIiDxVplfTPx/5pSOp
m0SWdRGkzhKa6iBFvPx3cDu9CBQJhR5urtVyUvvNOeyRwbfNUwSFNhKN1TpnRa8jVLab5jsO9bLi
aJn2JssjLe/feWFXNNexuMZx7XbULK99/8gcEI8EA5Mvr2AqXpcXHBryRB8mNCw6kdxg3vJjBu+e
e+Oz/0mJiAxxh9p2sV2IGE/2y9Wdf7Bs/Hm/Nfx2M+a+90zbVl7lpAa57lki6hCpnqV6uehfREN2
c9B2FwLBa2iutlCtw5BLHAyoXDkuyTOeaiAa1setTxqk/8CtU3hC+LYFYAMUWLnrYM/utVCARnbY
3G7+dLUZ/ovqbDLHyipFeZUYUCzIYkyUdXRrDTi4nZ72BpBUlKOt/8u2DbET0yTcLsanjcjmkVpE
CowubTS430yPyuMhpwI6cYcqVqcRSBv0CeFR2kFMukrvzUVEYlPs1/HBRYmyBbI3dETPLnU+p9ER
uq/en6q55Lfe2h9bfrgzMQb53NEohv+6GJmf/6kzJXqTWSosI0dy/JZqMJxe7QF3x0Kfoa6uJ84b
ff3LaHf2H+LlFqJsDXQyfRe5b/OZQKma82MparynlDoN7ONbVCrpIqw1S+BRLxHJbABxsBkmK2gB
U2WfE+3pS4cDsOzDAYhmaQjspYTZJBe0IkkeAnxZblqAdnlxgRZPRYEn0GNzSTs+8ZAdWRvDPA2L
F1Xjs3WidGVCXlxZfAPGkLxL/Tk35NwuuB2JRoPiLoa3mFcaaanKBPids7H2A+1PKWQYwbmOL+/z
4zHPts7ZYUcrvzvQSEflMFAOifzg0v6StN1o3E3TtwPVh6zDul7eKCC0jYCdMLWd6LrgLET/XaPc
Ly3sR/JSw2sMQAMR8O5yKXA2ZOCeXxYk3MSeqhUfut08ZcJsmkMBoaLxIxlqGIAKPHmYoHE1d11l
xPjY6fy+PrYMhKkYH3e8IYRxq9SUJGOj8MtK9zCOq00qfNo4pbdsF5SLWHFu5dQnllAuZezloLxV
lDATmogHApvUW5uKX7eAszfKuydsk3muTki+bIImuYH4jy7GxZvuddrDgVnWlQdvAovmGdVFCWMv
tEm2BIB5aqiBVnQ9Z4y1M0pl/mSVa1XE+z9houy2phWYsaGKEc1Ehb60aDaIVMeTmsk4tvAwP0B2
1Ovu7pwEXHGfyGIL8HTIxE4E08IJ7PkZu96Mbh7UhW4Qeg/HGBgHbb6JaCPSqAT+ZB7x+SJvUpqw
43uwXX3DG3JP70/r0MUuvcAos83j+AAdIqfC/16adKVhP50F6omj1phuAE16258tFaFuBqNH61ja
vI2MysDHnQsAaCYLCbuBxO0A4FdbGVv5Izxi8dnyJ85JiAf04wnusecoeEazNA8GWoIPWH0ZehkE
aD0+vHQeUamQYOAVdvoeoHE1R4iJm6I/6kpJ3rhjXU3+weUIbpQsbn/RQ8x5vabYoe0nMUK4Tgnm
kbPDzDqQnjIbZntclpncaIIOmbrsKX1jigNEo3CAFqVIxc8xf4xiYRkumWF88mDvDJ5752sgN6+m
Jy2v4juzNF1aGSYJTP8Lkc95Q7PiGwEBTo9Ydi0tm6qTO8j9KtP5V96zDQLQmnJKCHm6+uro6XKk
6svaaWHIOoviTuREjHSXf5iAGyej5qn7Vt/d5Dt06C2WpbbtAQppDrIKATKHAjK00J62wm3Vtm0K
sv9aHGbtnm7i6G08ov6C5FV3eR1tA7YiWxu4yFkXNIC4s4Tl0H9Upf+huajoRxw43sGTP5IL71Zo
DF07oQUinLLeIIG4+AsqgSGQVB3ff6yqpcg9N8YVIUs/O9uDD0x75fyKFHQ+l3nGJVFa28otw4wq
+Kcru+O1iXcZ88TG7+u1dKBQODb3HiUUwr11ev12iwsq8ZlAfZ5x8QOkhM5HwvTMOlk5guZ+AuUD
W0ReK8owPFZAtWIk+mrnrtUcXgLitVMuqcf8XVi764f4MyvIOWxrjPpXYoDZ8xqe4gdDGoc4hvhW
NPFLr6tnvtn5KDyKC3UFEo2osu8i8Ac0S1TttzLpaeo4FbQtnW7kTNpgtnw/16Jfw3tBdkEUXVOs
NrXJxdLLpDsKCPCroAtV1iyAzlXJOeh1y+S1A7K1XK5UslRI+luvM64yVF3kjadP/kZinS0lry46
BIm1eZZ7A92SvtuUIFA6Grw7ujqzF4IByxTsh7voZUuFufcHfXUQ0f5FvBYln9NUupk5kf+JBXPC
on5unPB/7dt5iOS/D42a4S7q3ppJhSSF55/vlBHPGg7b1I7D9o1pwMwzPhEYg9ZZx4MvQgS7RWt5
JKOG/u9RLBDNCBWJoLtPsIGWCJLhsVY5aKxTGK0W3EKJGomcuDQtL8uTasHIYRU7eHPezx+tImOS
19uCupjP3V1dJ+icSVr4Cp0sUrm2fUuXdAXehIpx0ywvtGRraV9suCgsD1yJZM5gqsRJb2izwbWg
mro4gpPlm1h6Pt3wsgcB7XVLBXi4olq39UhFyAJtyCj91yOb7v+AmKDJ9tp7WzdKs4slIbU2Vj0t
SrQVlf0RCL1AP5+MUGvO+ptwIozOCfOnQHm4tzdIn5SrnDlPWoJst0mwWE6PDVDy6DfcDusWljpm
Gw7kNJIpDPXtgUcUgftcnr9FD7yv73h1fFheFf+Hiy4EG0abq0Ds121bdYWoyiQeqV2ksDY60CbU
0sCmXgd+ZeW2AOHFlAZ4tgqWsRhzI3VrIkOUnRJ0ZRuZKxrRYehqJV2lMPws5UFl7PSuwIq1d7w+
3GqYrANY81Sdh/+0xJ3rXqoUWlyPosuZT3DDlvQ6aVgJGIw0MfoqXhr/xE9PJTLtdWk0krNTtA+I
+1rIbYyuGmh4ckaPeqP/3mqWTNruKc7pxKbWQacBkCEWm1tddWqBUA2bZo0SSr02hVzWRx5C++4q
32dsISGe4vft2S5cvp561/lpLfAEGDhM+jwo3xt7aIcJ2FX0tj+AayiY1ogoShPzTqjLG7Npg32E
nB/yz/F95B86XID496AS1pHA8UCIWPeCCaOdsOFL6FNJoIMiDFwU/ypjNxbZJk/X+b99xTeJSgJD
XXJ/e0MH7iHiTqzdkSqKbFMcojv6VdYv/kx43mgEITo5uxoPY4GtKRjKjtcd6DhemXg7FmS34aWY
ivvwz+9Un2gZG2lc4Wuw8wUjAPvQV5OHOWvSQL1uYu407qOrsSACFNyERIGAd+hksVTsAANYlfgL
RMPjG7PU/tQujUGtJOydL1YR0EwcWXFHYuUc9iAerSx90bm2oMy3f223P/vC5+uOAhJ768DVFUF2
kQDQe2O4NazKzbd28zvIagocl2glu2fhUtYNELouawbN74CPsPNsOzEUgsg8EtaScEU+RtEkFWnX
mDpQg71UIB8AqGZj42phm2lYTYIGFDhGEMD9Gf9G1vKuY3KNexMZ48vee9qJNQ5g/jgkmnaj0dVO
a8O31yHh+UuOtEoohMhtosu3VbKSj3ODzzxIkMxjk0HvRJLfOylYy/7FkJVynFKKu3/j+Nv1eZCH
qPs3Cb8JPD9JwEAUt7Q+HJWYZLTzLXg6QV/jhilfFafUitKVe26lVHByT/q31cw2sSg2oEQDt8Q0
txqd/ApCa8Vydah3En+HdDgMcO9Cy/uyoID3YwXMca4aTchK/7V34Gi2W1vW12ObpIFqFqTDyzJ9
qc7yW2IjVR2GAXufyf+7jBmhFSI2hHZZXv6Oam34TFNiN5GS6SSJkg1n0fkH2P9kqfMJyITonELl
2RN4L507ExqVXhV9I63Nmfl7mFPT5gv+qHVAhUcG85dldbTPSPrXXyGNcYM0F2/ce5mOzbxVKXVS
F9FfSc/9gDZ9YXZJ395DkM8p4NVn3GIr6yUTTRl/DbBbUcqkA7KfK3uoEFBVKi5yc8qoZwvKq+mU
kaze0IdPZWQsGmrez91VtYFXCsXY3Av1yxlhZi12q8Ct1yTjE5sLmh8AP/hfwcs6re3GMLqCi3Z3
bnmYWIjgjYAHSsMmrRGtuQs+OCYqr8Bt4fva/yV//tM2pmRDYf8fprWHEsZfQ/dDfafWFmBuMRqn
vqNtzc89h8Sp9cAMlMTAyenI4PYsoLwpyRxQv5uAkgRkPrppg0Z+UR6B+tfZHsS4ObQY4QiC6yAA
+aJG5qK5SxB3pIjxQ2hLqGVHzL2zu6TM5nFB1Dz/wdc9/uo3lhcJmrGTTrd6J57VLxTm4lMigOK5
4q0Ux3aIiGGmZPlfnWSBec54QvTGOQTEUhGZCx/7nXsEvJOFSsuYtb1wnr0jX/AT31xNrp9jiCdJ
TxIFn02eL4RVVlme1Gc6sR6HFXNS81VTXyeHNvYchBOArAyw73OgYevaQpf93Q5v0mMDL/ufO9CR
PPutscSuSWCTPziGBzyaGm6HxNS0YCkBbcJRGYDyLqsjvg9OKu05Z4uhGgfV7EK4/EhxaonOsdpc
7TVfPcQrMfpLE1+FcdmYMsa38Us27DHnNHTdvi5OStnb7bal9uNVxuhuhpOuCHU6iyKMq8THSnLn
FuFc1iPZGrfJt46fEVoc+BcJTOUFKk/kng+WecMcN/EdweGgBSSrLudIkuNhZqJalhjcQkOR3a7j
aFNsLuChNdZZZMDocQR6SS6MTIHFLZr20amg6eRTlfVWarqXMEPC2q2X7NUGn9uABjaWIDc9NHuY
tVDIRAiiTdWdPFIlR2Q6n2VKCEoTK1ooK0iPhiysyYJ0vbk3gCsAUO4oOnsNU1c6ziRMP8UPLuOr
iIA9g3KWRkHKlM2IP/abP4QUh9IxHcGYOdZIitVjfoVMquzYZ0MP8Z28klYXDOZzfcmlOPyH/beX
NHCpFpXie1Z0KnUJ65bNawt2G5ekv2BNDfVKzNAFjss7tVnf172lv/w5VeBjzTDLF4R1SmvCC5nz
sV8qsdNkzwr/AEOLM+KqxwNHO2fANvC+2OcEzOBNVwWkN3rNXHF/l1SkoEVn4DUdzp7NwHSjkGHO
ohWrisE5MdFT7Y8DvRYzpRq/mHe3UmZTzeW1pgAbV7ayeiFauaUigubW3DFjkRVV7zF7LSAqaesv
3nJAG56J1GVJZYANmjEcJoGTztH4lH5g1bGVU166aRiWcVdrmxsHatmrbgOaVHaxMiqp9ZHPyl7z
RG5H2VluP5DGHHoB7sBgFIuIaMOP+4XH+D8qzOwqaHfeeewVpYnZMuwpbOVztZD5zNRLTC8VHmct
5ZAhf8BEDD/U21xsAblUO5Bp/kNMdeW5HGPcTvBnmH+F7cTz1bvVTfi3lwp+f/fxSF6ce2GPmanO
tVZZWGOBes89Dvmv/GfzoJL+WWTl1TSZsM9fAe/AZ7VbnceNofMSFikxn1/aHolU/F4z4iFUWUKG
KsuuQ+Ps7k15EjT9Hz9W7i+zcwJWSS4oPDZDBzXwLiY0LD1hCh0Uq7u4TSODHjaxzzs4LoV7pvOB
cExmBvo9lHgiVCmpgN5YuW6/zTcVvtXH27L00Nw9Q5UzPbuNV0HZ9TPWsB0ejyBr1noooUQV5XTK
czjPeSAKYyz9FvvtXBUK1IEBJxjcskQQTrr3bj1AsVTXQ0+LTfEAfNSEg4htjZGNh3iTLM4padet
es0XgdNwwnkQqFNEBekU1guw9i3poguKLodQA+SXC7vsw04AQHNBIysj0t9GEFQU6MbNAqzxHWBU
bbnz7vmUFXPoHsx1JXbX9kC4NmjpID25d13L47MG2ptUSGMDqSOOZl7UFtuvK4cW7lhwtOF4rz2q
rDSHMM24tYoeDa2ob5tsIEK+w/ZtAKS3OFpvHrKw5YvduknwkQXIQkeeFasYsqF9RjUc3wWlfJTL
auVzJCbQtgqXdVlTbJbZtWsb5rUe4ifGf/cHpO/oUCdGhKsMnVvZCS0yGrSfSw4GctVTgkZ4AmAS
5h7mzyMFgpbWqikjq+RleM+OKFQ6EqGLRTuNe2ATvypdw2MSJvVCiD28xvawHcvIgTT8AjGvNNNO
WZ109JICiRGvF1fPbydPNZFls5l7qi25p1Bvu+G1B19vbVarGoRjeUBE8sqQbB12ojNLqYaNLZee
kF0hhP4PysFtbv88lF8zgXahexwgDew8d+qyYSoW9x61dSGS03Ueu5YCCLK5eYYQOJZkD+aAf+M7
Q3shEofOCxF/ew5twVXmUepKH7KWPZsji/HNftzB0vImnvmM4XGgpsCjeuKxDBW1aGbtKdFJvfH4
NcSPNCTtdPbyCGCUHiPlFCuBSfTq/D1OO4TnVxlKYXiMpgq1QgHl18lc82gVKy86UGtRk9ZIkYtQ
Hco2zMug/2u3IGsSAvvy9bImX/zIpJ+88lh/Th5HeKLDOPy+CjxrYojGcOxTciKkjSbL8Gpzs+9y
59RWZRL4mpQzysvyTQ07v8C8FSqUcAPYQKqF4mMquIzlfZmGtHIlcw/xz68OFQAcxBXdeqzfZLFx
+eVGfzihgZ+m0HEOXeFVsXMz1bGcl20elxyti1XWHEr5uOzotkJZC9BfHcIWR4Q/0WOXAHUBlH1f
EQopd0hPcLDBwByym4iu/5Q2E42B/g/fBAqxB/uGKcXFEubMxi62LU3Zw5AYwTZA5ufZ7YkzpB5h
m+dmll2vPyWbsw2rq+97zm5mQz9nLQsrFr3YRn68SbkasQAkGiaQmJJ4V5MJy1ssFqCxhHTzIBvS
RstTYdOFdxf6oC4br68HBbSrTT30UIrmobTfhNbsrYtD8j7/qFNqBm1mIZSPM643J9VJFr5VyOV8
cR3CX5e7BzmL8b6+LNYVO+Pd9/4db9e22MbNo1jlKfDmCUUgj1joz7iNFojfv/ul5rrnI1iCoDsU
8gymFvv4tcjYP30GIGbqyt7fNqiZdIZn5sM/3/VEf5//Q/HCt42KC9o2VqKVpt4ZZvzCgH60gufo
yNOKGcmJ8NdBeqkZJ3M2V690d+FUfSllCIzoy1MR0Bd8x/UK0vzX4ls1K/13jqXhWk+gSYYJH4da
yjJcycvtjW0R1M2lJI3bj/nV4bRGn8I+xvHxixAFZJ6A3vvdjDdiG1Nygg9bzMGCYeOkPgK2enM0
EoX+F4r5EDQ4BTZwQu2Zt9cPtUm/gunrF2/8JF8ptkbW7aCeT+UrNMC3SJ2saEHkPC8nhA5ulSqG
1tLxCkJu+iZS6tzhamiivtxZbs56YpPctuw1zJZoyW4Daw6z5O4ROXZPbZJOOfmlvgnjp22M40xz
FvKqz1D+Kzvp7vkSPUhty0L7cGmb/dvBqwjXsdoGcdUZqQOR/Mhh5+Ir7iQbKcv0+XdX4QffQhGx
gSmVi0gbDShb1BYQLMq2KrHW+yAEPpm/zgcmcl5iX2gANEaUZbBkGlQ142x+YmkMF9bii5pF6/jY
AFo/W5fA0/CAirNm/aKK2pkLIktCW1ZN9xx4iNQSkJWEKNkw1e4vGJxhgW7hoMXzu9j9RZZF8cgC
mPXT2khpdj7APjDJbBcAH8RKjVsuefkUWnuLjMXBnQg70duYqq4N4/KprT4KiwrzF3TVCimdYDTp
H013N2p5g/ImhDSa2hA8uTzGXl/3ybD6oVQ9cBc/RXyD/cgYcJb5UWJyoYV5BRcvKRkByYuW8oxe
aRUArYBUo+9++9Uc/8+9ZlGOOAtxix2fm+rCNP1LbkW5TvSVerhgbduVQBF6bgSou4bstNccnfl1
VTjZW9e/iUMPU7N9mIWg6a8ys2b3kAdvhTOXSF2M0V8lbvHRz+p0L39qjZUmrxNNiDcL42LWqsFl
w7CnGd/WeMNpL65Buq/+AV22O5Dmx9pc2crrFj58//QJX6J+VmxA9SThP5YAI+jla1bADG/7xwZM
825J2gBl6LmLlBkz3B8blweceCZN7TwOAzSGTNPp5+xKedJTG6U+KfaOVzZHneNnkbs1jo1Rvz7U
LuuWxQizBz6AJjHN0ILAI+8X/4FVX3bV3N1nPrHw7S0NSyq/O7hY3teCuAoQAF875FzRVplDEUkz
KZ4r7Trna52N6H3pB1eSJhg7Vj5H7BFJ+sBmVypz7tZ5Iuw8CbuaBVhM929JdD7XAcM7pZPG7Qnb
LROAhEc8068PExZPO/m/FDReI9udovcpV1+KW/dAUCnQPbrzZyu0LujG0CFJESyKRNAlaZ5uY2fJ
E1OWycPoI4M8zfaIR6aFCv/GRgF4xNPZN4YUGxlBTsXkBJ8KEFdnpci+xD8GifB1rTKlH43hZdH3
OvhIGghm9Q75wOmKEGKKauaiUUq8WAmI5Hau7U2NBFWvlN+uULcJd4QCm9h/eh6fdFltKGsYKPA4
cgSg4SaKpAjPv4UkcQGW62nUkmbU+SB2OlsNiqzWAknCiq9BIqlACBUpZci2OGC1mHa5Mw9VifE/
GlR7caZbxdYxdK+1ttRMtA2HUu4vXDXCEng9pnTkYmYFjmoriNrSMytl6e6nzB1ymVrWN9KrXHcb
OEVd1QA11S8PcxBzz3/rJeXwz8y6jorTa3WNN4zrWe7ndbWic/azW2FWQjxxIXRV3neYP1267i4r
jeX7HDoiG3TwN3qBcz9+JH8SXWfBZ8WcpA4QYdp12ck3sTX8M+jXTfFX/kdtvhMFySMCdmIlvRb+
3iE/6nWprzjGAAJfSR0wOPOf9Ur3FSGKgz2aNdoMKfTHzG2B95zdyb8HO2mU1WYB81StESqSd+3u
u1OfQZHr05tcs3FDrTztjWqurqoXwkSvLAZH6LW0SnbwXz1KAyAkoTmqoAHkCOsaLymYydwRB4uj
Abh7jcZAK4hDBJdjJLuxAy+IKNt90hv7p8sl67R5OkcZQAXAj+W5Jkpc7nr8N3stqfDjgwTuuT0V
QCAYhnbDBUyZuVMU1ZNyzzCvpDqJl5a8/ybI2jbn2BIbPMo5+c2skBAjLfzxUrdpejScEkyw34Xe
q6rCFLBtJgJ0QvVP8NLUku7ywrBY9wpapJkK800iMOwrchaiTwa3KNsBCWE0/MJcSxfW9gecQfmE
qKYNd/7ZRZRlIk+lo8hcRNJ+ociJxgGkLYdqZo6faMFsLiy3hfNS6cL2L9v+uY0sFaJROhTuMjy/
+K6QxI2UBYotpAmmLUgajMAep3WbvCRJDuyfH4+QqddR+bzDYHGm1zYY6YS3S/Hkb4SoACcmkZlh
bzm4sBDao9Ou51jgVNPACyoYH+R3ja3hF4P2Ixznv4L3Y29DwUcyww9OFcD7th2dcMcerNzA+Q9k
0/u6dW7JIx8Tiar2DYtvKsJYSqH7NJxIFXOgx72m3F6VCH5H3BYzbTF5CgsSdj8FLmcvybAIQ959
tV8uRJuUGNj5m13GruGjgZV/h7yjJnSIWE9G7t/V/nxRH95WMJpvKHgEqKJSrlF2i2+1uI8yengo
2mI1r+PUpK3BTgBea0OWJl3kI5oCyS4aEGI/Wwt9xYMngOwQBVKeZPoeoDK5kC0CkEbtvOIUUdMQ
QPCl+T3TPP54bF01ZO+ooI7u8ZxROZK4ERoE8PpinkBJHf1u52cZsMPymdCxIDBZnX8GvkL1gRFE
YCQwnXKMC+XUe3ac1oEughU/0nCX1SzvLpeiWmpcjFx3h6cuaI+sm1iGsTWtXK2Xus+yjg1REpF/
G3bdRzGwslt93ZmXcS4JfStVpXio74EUgS4qdzLNU1L5kw/pHz9oy1L27E+qV2j5Uk/KNh3zjtYA
5H3SrHJqlK3/ho63FFqKNBlRe4vWk3e9KgUhUON2Cn8J6aFA8MdE5uva5hX0rJfR4UKURhUD8Nvt
yE4tNSUxgM7BwSiew0hXDmHbD9bVwlXdKBj8y8z+Re4VwF5IuUPuY2Cz3KV45/P0FJOnIY/GmGsY
vcewmPI3v/Lh2uKFrXugaiPSRtEES2zKTefAtienMgFvbL7dqJhXlA0QuW1ywC8jJ68SJRxfAlqC
fKN/zHLYtZQ7W4wpgsonJM5YGlN9cw9pIbOPoxKIKnELAjZsGeiZKGuwv56Ep6K/xLg7S2zao+E6
T/AAWXJLBk0zfKLHrwxf34H7gd8YrBKUzsjq0HVGujj/st/BndcgoZenRFmkeT04R+BiGSNzJIN3
JNueATkRR7Q6zibMQx/83eH2BrxujeG3pt96uP6yKBQFK50M8Fr8cYZKo6VkXpC46MyU4oyDdH2/
gqemR8J2XyzE0aTJ10Hit6IQCxZGg6M8+rpt9QEvgXlFZel1PwyCFXcuxA9vq2nK+ZChAAE+CDCA
l7UsKSoYu3BEg9A//TosTs4Tl8DDpk5wGvz8l/Xq4LLa7bi14Har/IxPZjDW7H+k8RMWb7Sib2e3
i7u7LFFKLlZusWkqJ+9kjOSFfWNXwQRkny8KcK/zVDHY0bvzBoafe/CfGUTB30SNBclZGCMmEaDv
rAUYtGwfyuM7fPhrbNcHqF8MliQ9kGy5me2Os6eC5c1L2+9ISLTRiXqgoFOy5qV7IQiMEYZPewiz
3gNcIWnpmmi5yEnV8/dLZxOBuku7ROpTa9dAc7BC6SMaxthBOhx52Dl2cRGil3X4VFJrY2VmVNGU
bbcCMRB0t7p/PP+eUvNZDsN3Lxi59YPIpFizdGLUgrIDPOIzmENLxKQ9hlrKLf90kJhfE8l85Gx0
URthmjEbXjc/IUbZ2V/2wkRId5nb18jzlcWSzzkNyzW7gnJt7VCGKEuYtNdH7wz9u9H6RjBix+ed
WgYon/r51mgPvAlfcK/8/Bhp9V36raz0lb6sEDf6DGQvmYgU76JnKuC9CSI2w3hggwJ2gNRkBzmt
DRUEF9Ia9MaG3iSbsb7V1LDqm5q9R8F4hrmYKqVKytIR7xOcR6fWPYPgtUU/B5MmAj7LRCjqXgQf
RPcfgBhuiTGkz+1PZNjnWfDQ4vR3HjpPw/9KplIZUwS3u9OYplLzfjUTOg/3SeAbtV2jFInP3HWr
AsyMx9kmw4jZvJZxesfOeZoTNsBMTTw/tSvWsCtBZs63u00NbbE/JX9EAcN4aGdZhAZE4q9KqR7f
j2UUeEL/OdQLMUtpJcEMpncFE1WjkJJfEOYiTm42uExxh+z2MwWUkfWYO55ICj5P14Dm4Mahp6Oz
tIQvDslTEhptrSIEDwwouVrk22W6fxESSOoME/iEdE4oDnk1/qtc1YqwiLRUtBZxvg1USt8Zh/54
V9ZddXl4HOhmWm5BuhHoTGbVGbP0BSUBlZ14TPO7g5dIVzszhYqJEc1q1GprcHqKyxlcxFSfNhSz
DV+YU/HIel9dNMSKEToH/Osa+lQXQ6LOmGghjhKHDbvf3CKoMVYKcFi2lBaZtK4KO/QAiahxHlwU
UCAt45OvfEUSKJMv9xdKU33E6VVy0ogwialJy4exFNG1MdKOCLMvbYwdJuMhNw+SA25qw+ErvRQK
jP0AkSSH33XGhkGzgrSH2xPvV7iZGOSDusLdrsLCysNZKjvtWG85TwyiLaL6GPb/AQS+9ePCOXNc
pF8stouBFVhxnvJvg6pXb3xrPzyEl6iCLUYTtBCRSii5M0BqT/ourhxgkWi7w0XpOleAh1vasy/O
su+CWgvP7EUb2kcTPjrksmRrUm7Aa+DVmqOEV5k1yWcmz0acfqcoyuqF388zCvAB+TCKPm+pCWka
ghIORwK3YS3KCg2Wg2IgqIAwTVJ0KealF45Vf8z/pHcgE/EQTOG9iq5zIxBuRgKnwpQLTGgLkncm
S1OvVQH0lymQJSPTJDv9tSCOFbnZVbDJh+m+F0h6/isdtLQZeYgkoZpBqmOJu1zEe6vAL//1c1ub
yp5bAUHVlZWVsqE+rxXm0sEdbjIGvBf+7ToH6DZs5QndSDZmGru4rlIHHOtJGsXQJbbhyhNG7vP3
u2ygUq0X1BGn3lnhIBLrEz6ksWjLvX1ByfDQttG1eYPfc8j+TFB+0bE7mQMrNy3E5aNjGtzahhCi
WMKq3nJhYui+Cg68R+2KsHp02ulzbuhvm4lN1lENAkMxpEUhWfr0eFK1BUY+KYX3YbGHgXVt84K9
XGmcCuuXJ4+BI2d1nVEkerYym7pTPlP8dhFtQm5iCBhA3C4+dUStNHgmDYvZkfEpjcWV+z3aHYj5
sBVxVPbGlD+bjYyNzOKJtPWlcf09wEvqgo4s5oZVEFd274C1qgIp3ntacVs19XnXWkxhupBX8sEP
qiBrklgnJ2hgMDwS93X21VyJUiDGdzpRxRD3FsrJv7cdrTkBDTLhsZtJc/BU0/Wsv6O19A16vwke
sZPqDZ6mzEY8ngJ3UiQGF7+ObU6RxB4R8SEX1kKobhlCjlC74fhsuHGcbd33QEOpVVopKvIxhIcF
XVRznjmRDKUgP6jLNKXCcLCZ30TQ0SPAhJ02rmo1HVbWiQFslgcJrDn2NAkwsWm8fNt/ZWwy+XSA
gxMw0vfN5vRT8/DIBO2aD6QrsHgZrzmsIOE4JPJByCTfi0FgimCSlTmCPmJYoir0iyG4lc/rw9sJ
kcVy/oqkEii8FUt6FBsKXdWN6zgb1OW4VfvDHOz+3vSqsx7Phd0aFsSyuoVpAqUZ+Jqb0jZXJb4z
h6oGt/l4NjX/SRttkAVimQGvz5dwtOZTmSf0wGk4jOtqQVLWEpFcda3uj7oOliQ2mGt0X8MaHWfa
X36eZshFN3KE86BsoOh6RRyP7ERGYYwxiA5QxPkfvZMKJEo7m0WUF91wQH+UVspGL+lUB0E/g+X3
yWi725E6RBVBx7wbxfC/1WqdhzlNZT5Ntl7x0MgNfgte48yei9vtiaj6AO8tr0iTNG3qUn5sKcXr
2XZMyvVogiqQhiUvW0x438BLDW9Q25s84Ob+e4TzEgKD43ZltsIOLSJwXxo6w5UarivkjjVt26Jo
R+iCSgUK+1V6+HUIYT+du4Jt/9Yh60uiAeDKKdwzQYD4MDdkD6IXMq1HUg3jSaN3bGvu0rKHYvcC
2N6nEopIH414V1EOUOvWI7ix5xRNJdPYr27vExSXSwvXuNbXDpZl4Vp2dxtjs5g4yt8wCDOKVElO
SuP8HOX3A5/wVZyIBfH6vFLC1GFt1fnk+X/JQroL6INtL0622JDTtK36ddRX0UJPEKG3S9wp6X4Q
CwL28E++yGUcZfx68sqOrodKkqOkza6wyj5wsK0aF5kBWbEyv465CS9w4q3cRN3BrqS/ZyEapb2I
iu85tfnow9UdH3aB+2n3LohhSp6UmGsjzaltJ5Iwg4lDUo2pX5kI3+Tq+tHLJEJw1jD4b5UQkgxU
R8WPUv5cvTXbLk2hO58aY1jVb5RNbz47FNJQhAU3DKNNIxRpCo/UtHh9Da5DLEv+jHcXltaAzJkg
v5Ocy1rboHX04Ui6PJ6o3JOH7D2y5uIwC8bDF1kpqqHRqvhgg29WSMHL0jBcQj6V2zb46/AHpcQr
dS/TN1rSgcR2ubBS0kZZv2dJmmCeRHYZy/VWjYfatkPsqJ5CYCYt4XUvnwbRRtnq1vlQIEzOIMFk
i0I6Vy07WofiOPiZYqAy7W3OjeV1bsip12OEfQAPx9OynMBCg8G2yFMGBsHF93P+eXJf5i9hyoBL
c4ds8P4IFT+2TqpNF5o7UsHLuorhhaJ79wMZZIATehy9jUyX0ZnP0cwcTlA2KywJ4BypB6ZcQsQL
14R7EQ8mB37c0moIrJt4sGMc5bQrovJQlJArv0gCDjbs2SmuR67yGeflAF9MFtp31sYtS30gx/zH
l3y0VJqMau2WNo98wfSDTW4+5R5rohoSE5DvUV1E1ApJaTyi438xupHWOaRe7w7iprkb39bhUpXx
FyA+/PBBEXLSl3/R9QhH8nstDXbmIJao6FuRYzBZLRp1WYkd+Z2GEYmViub355GdmjXOLQ1eeoc6
0KKMnHK3g6exwKADZZPTAs2FZH6x5SlELOyWpY/x2X1Q0hzKUnWI/YQOrHwxMOQ1YqzlOWc4fMeJ
KysB3Errmgr2P6IRBJ+x+BMEW8lQHu8lQTs5XWiiDA6LWtnFKcQee9h5sblD2aCyzFlIKqhPr6VK
HJOqieaGURt6oTZnOIIeyhvzXj9pboRNZavptyJeKsQfjbhGgYxkTzm4ATlcHM0R98DvGVo6xrIt
O48VU7FVN9ZvZ6GU0M/A4aFTIqv2hXXc9UmeMpzK9ttaS932GJOck9of2MDRcAMzOtN8bHpkjpEe
I/1EZW13sKUA7lDz56Gz32a/1tr8/7Fn5wJRubM6eMqfmRb6FtoN2BqWXIIjvyFtLT0C2q5NRsns
aHlwgboVPmYhYg6UUXIsP8YQzBbjAjSneEaArT1MevZNX+w1B82syv8txOylzlt8MhApER7MXRex
5XIfvz/v93n0f0Esku4v67VyXbN58EDA2Ll28xxLsHhwLABFjZwTY9WogB6WI6z3Pg32/h5uGtpd
IZXCvV58lBXxKE0iueec+kvpwwx5+g+p9sVmCNV2qPZUVwyx0n+Chf/fu6hVM6e8Lr0KOC97vwBY
k5CtDp6o7Z9BUhResAW98TlhwqzoxZh4xHc7k3MIMTEKcntUjsRbvDr8f7X9LQT4chIWMoxJNG1h
4Z/2L6FBEQrKRyNnGvxgsrqusNePSS8U2m8VFMtGJ/DtG12U+fQ5gpZSgR06NHqLpZ/bqK9G1V8A
JxZnplPTp1xtxrk/UER4t3kYLsjbjtMDer0RDBlMvd0vQrZDfkaqVdmpF5WB/c6QCTj3YYJ3pBkM
ciFLWVoIOq6xOjUWB1fg5QEsbXh32joqVKGLX/qDmsYlZqgz3rwsP3BoT+FCvJx6hl7lhTdz2Qig
84gSF3ZTnThT9tVfI7E2O/6IaNEtsPmc5TwKJ8D7GLenT9gyLoUm9StafQ6feG3k0jevnSXYkRGX
U6bhjIMfTitHax86hPDskrc3mLE/RyyCAZjBvbq/AQxQeQJImB/A0duLtnqz7nfOcnWn8G8GH7F6
/CIrFdEeR4Bbcpx8FTLue8E6PqAzfOGODDXrCvEWFWF/5mUKWZ9O//oAXkUYAjLEOYqnJlG+Z8Vw
ME18A7cVsdYoD4M208EmJZZSZpRVkMf9FUnP4E8Vn3pVHBO48fp8AXA8ZaI8DArmgHVIVtcel1sV
BHdnPp5M4nMdpNjObYA/G9dBEBjfyvLmCUXeUGoTvCMUfvKyNQ/3uB4TmSwP2ncyogNajRDAv4UN
eQLfigjAnoKtU6ejivJjVD5Gk2f8rv/q9rJfPcYzZHgTWc8z2ds8kYvKqVQKj6lqkIRBqUWRQuwr
CFbQKheUIqvx4TFdzpx41xACP3VuFKC3FzLbj+a0KDL1VbNCPaDbzvemgN4U35he74YA6J1HvOBv
dViSfJ365HfccB6AnvL/YCgafsVPgIMk6IsoDY+Gq02Ivj6KH3vTJTg7r0t/9xdX/rNZF3lhPn9G
f9WDCQIkYN114PfIQVf3iTuMOUO5xtzRRe5qr+7qQoBmFgxPQMaYux1z8MF0lZAYrpVZfkh8DzN7
26E2pDK6BogVaTP1FKDYi8mVfEe2vIt8g84sBVxOnmUeC/iCdHLEY2/V23KMs4ZoTmt1ksji8o0P
xojysJ+3fTw33Y/GZkgqyflZUj0dqrSkYqysRaTA0UpDfBpcsYvqNhN+IkVZDlYWKXJ8UMDZ8kHy
yEITqC3GSiXpecr9fHuz3BsI2bpvWdAbu8bZfwW/wzYzq26Ijv6/pOLGmcr0UqGd5v1e31R8ynbY
nk5jVBTSaabLRXP/ki2bYRidafwSMXijjHEPUjquYfRJY6Hb4v5XF8OnJvsbvanOKoS2hSumV+bm
OL8fPPcsHY1fNvm9UYCTym0RYanPbfQRbeoA9H2vzm1L0/tOF8BIbZdTKs+2snQy2G0X70lhwZTb
j8XMYJTP8E1IzznP05QKGuy5D9vjnfJ32gE0x8DgGDHBqGFOiMKJ0Z5YwQtTVdSp2zyHHjcEXe4c
F9REDowWx4hxMyW5Iunrh23gjAFCWTXCiQIoE3LXGeFL+NvfVr6pz08AQF9EgsL6+yT2g50BT1Um
1IZDii3M0FfMK9ksZ1qjmCC2gQkiwFQ7FaiT1fLAoU5gGZ+F5hnfQJZ1dXgysAzKgb49rqNo7hM1
GtzMzmu7Uo5H5UCVNmYxrIMwrOIYLikMCusbvm3w4inf13WtXBd2tNXWS6+L40VaW+UBDdhHDG2C
ll85XbzZDvNJ81sha0zlU+A+XwX0ZLmvq+xz9ih6lmQF+ndS20Bl57DnfQIWaO6eIU2b2kWDlNgc
x40xsIMxS/ZZN/9fiPiyO42zSZektauDNfY4Ttbc0ca4AfIibsHnooOyrn1yXZc3EZVVHNtrTJv1
ZiVNxjjeK0vQUjEuVbAyntw8EsvoCxE9kxKCV2QZ9UL/2UMNFgRDUOH+b/8BpWsiWmM5YcVPPHhF
VTpeEm3iNnOYNpLzCgFqRDFfuqUxbBlGF02dzzuMG3+XIfKpV16grEKo0nt9UuA/h7TiWXwql3lM
8X4udW5BXk02T6RWzI8GkNSUt2dfHejT6DCrbotjT+/ND6TZoXpfT3BLkZc+VCLlUl8tlc9Qjpgv
4lfEVufFlVATx3ecvbZyXh/flKMs/TFI3b6nINCFu5YtJ4qthnj7RwXX0ahTbU49gJR5vO8MKElD
QLhLtjIsSKTVlL2N6tuvrg3OpGS6HDbuEzCSPXC03Md7DRNJgp6wSCoq4pdX/t81j5Lo/PE8sMby
UXUfgKQnZP4yhwA/B5oy5cPzMzjbceM1elYw9tuh0K1c5p6wZ7BFgsbaieVizYRYeYaOINeNgj1i
vxDHkrivzEExR0A8IWxxDy4LC2aVDImdx8MOf+5E+qfe3kPmtNEsCNVdQVRfsPiGdq9hutzxQt1z
ue+KyZ4HJxqp4p4a6bQbNT6KKSLETG8h+vsJv1+pCzNS1uO5TXFbtHe+ZcPHxNcYJFseC71RQXHr
amDik1Fvbl6kJZ3+NUcxhKgZVEu8/HNQ7xXT3JPUqcGjZd9iywBltZ8hRTN5d4PX+k2L2Q3PPXjk
0MbHsIRI7h0v6Q7GoNfhMvoSxDVUA/FMDgnKbArSYMyuX4nZdNQNt0lmZNfC1y4/lGJLPq0xftc6
2MPCAHpii0kP7Vqs+liy9VMvF+JDGaboInTGNhyCVRvHkqSsO3khzVtMuzOMJJ+IWRMFbiqu+KAt
kj3BENN3DcKXO+UpDqnQRZjKIl5wnqoucWn/516Suf6feZllez9nmTPb6dRnr+Jsy514OGjks8K3
WH/VKBycs6vMjOhywBX31KALDeakvrlX8fD9K+vXHfU1KJ+CXJwteTm+R+5sj8BoPq54ZTwnZY2i
DimGZVumBacm2BMbIWLsfaxqf6WaJAiWm6igq/KUjr7ptqJnUts+K0gdn0KMLWEsF85UjE880FFf
GGpx/5QqvkyV7oNGAOXsIRXdj/oD9MA0zc09lxH8CXiyXFWCQDq+pMHpkeM6u+vxufbncCOZ9uCZ
JkUFMBgTGDGXyOQcnSkbFq1GO7zEbYJjnHVcqtTxGABZgzlgR/cinn7Cl3HsT5SI8rOBE7wxi+LQ
7dYlBCCDP6lZtakHdEdHRPLYeXMdt0KELGuDKAXxiWNt6lBPqNniiuDc02MHmY9Msbizg1IcULpB
MGUIaNGag9br1zlQ0b/NZg4QyQ/w50iXiQK47ZyNeR33Eb95Q5pshWg6HjUa3wgyD1rkhHI4hNB8
5LZKIWXQ1ra/wx5ZpOZtKKxKziRLg8w2QUptkKxZCudN58IujTAPPl/kCyLmDGNNkNXOZ84lELPE
kTiEX2zkrBuiDOT4vLGG/WXKduDNhjOl3Cj2aPuYGRQCpoSWGHc92K8w2DFvlbvpfNPXtB5l2H+3
9vSygwgyVIi/2gQBeOIucrO6DBHldh3+HfwDfWIGYpdhHAFuFwKtf5HctqOtRVhEU9sMC4ak73C7
NYpxqwCnkjNL0w9jv0Ssc3Uvk0W49+RULdUbdNh0K258N/TgHoumxde5vgFmAjI3Pq9JUgYBDN24
9gM2xBvEHT/GfE7obbp7ObQHa3zZNVwVtjWIVuJYaZmhvOathXz7+oACCmqjFUirKujNFjmKq0cT
ScBKd/ZxIWXfx/EW6BKG/qzxvho50DZlvHqtqle2BjpdCbfk6Tj3pYRi2Ud0+paJDJsJllO/9lOv
AMvPwwFs3md18qo6UXV8OjCNyZoWkpnjsmbeLMGVXFG1e5PPVb9bzZMyUeDYgIJfKyjiMJrv6i+e
j1t0pjy5MHWKR08ot2PdIjCqwwwLnIcieGFrIOMQRl8dGsTw3LZeHCJWtpeJJG4/tohG+fnQiW8P
2y2Eg+pbNznJujl6Du44jSp4IB+FdHzSm/HGe+geWn3x19qMSXJxX3EPsuglvzT3eP/8rdJ1RUcY
ccuQuVZuszboxJj+3n3TUe6sEY22kl84inRQluk6aEPcagtDBYPx1Lbp2HRYErp0s9fZQ2WepWFC
dAQ3Og7VpJ7Sro4Hgzej7hd+GjhmOqTbaxp/SiKrhO+FWFGpTqaaRcvscLTOAn6PPs250rGzJH0P
2GHbeKCmCk3wR27oUR1iyh/vkLnMUiNL3YgqdFUKWt4eiwNuqn7PQCNnXZXLKm7hQQjp0EZLiw7Y
uGzvWSmWk687XDOeTy/kXcYygC5bIL0JcE2KP1OKrNjk6O99/xDZZvISvtzWpPtOgCXTYILyFIxw
KInItFaxPkhT72vvoRM30erAO3sBHyu2stpZiwjW+DrOHHYDA9UP7JTZAgXxNSsuqthEd2Lo4ETY
vVetKP2Ddxocw1nmYWD2vYOnXbbeTFCHvF0ZaJhX591EFrtuG+ojRRIwyluzD4tWHgRjF1eU1JAe
oKFtb+iQ1W35rAv7DX2dgXeZpQpzfQz3SPVL8/nI7PRfJDo6rdY5XpYSn9MbZC30Ny9gBrlu2PkF
csj194YOInNkBxVrzRhCVOvxWyQ2L2DwHVszrUjPIuXRRdId9T81k2FYQTSVl6CMhrgxRw3gEEEJ
vM+Il5En2sqP5try9cWUoIqGZL+nqjrDgBi884PeVsONwrRJStox175xgUv9hncVgRO6ElAYZsfD
1pPKP8GVRVPCGFZAV4Iy3BKQ8gPxEWsVmG/NsbsmUUwKZzB+JBw92U6FUzAIdCFamCp8N7MedgEl
ZKp4BO073vcbq+KJ/rHVMiXtvXEGp9ApuENMQcxQTr41qoglm8nx8JAk4AbxAFozdAk7SmrVpisc
jTZyHRr1AAk+Irb/N5XeBb1IM1M3qgV7YbcHY571LhXnLYiZ/A6Qsw/FQn1jVoMg3nJ5QGiH9k97
Dds8G97O+eIS436aIOTPwg4Oe3KovvjAKTAWTOCDnLJajHTzh8/04WsjVN8MHZR39YR82glLLdLR
Ez8X+DKlA7CPwHMU/77tHn65ahhfhzd0iYLrFR6JoBsJvZoTTMx6HJldaNRf8TOezBZFO7zp1ezj
glOSIwigGzQiJ9N+YNA+BZvU/rFLhWhC/xcdHmTufs+XqdfJm2ZI1k7BWfNuzG1dYCRXr8hRXL7t
gDUWeuLWe8l4i5lw1WukoRWKA4dVdzuEzL+sKGEY/aT71HAnacfZeOw5nN1bJSkt4vi5bK68LJrM
/p3/49gWEV5XSxridPfQSW/6t98cz7luZ14I1HqYAhrn565jrva352abmmLw5FmpjpGap7ms4EtY
pYTzRvoMOWokhuiePJqG7u8KcOYkj7i7rVrSGYsr5ywVewNKqYf2Kbnp/6zrng0iIcLcDc9wApbD
ZcmnuH8wEvNuh3tYRSY4FlHpLJlIWXE+2RGco7+ejdKApaPRIXr0u2Cfjbdu5Rbia2HYhcJ5C/4z
ogEoRUukt4hFg8NaHWGhdRF3YRBrBNO7T+LdA1QmjDMxjE6T3iiDUcImDrktYSjuzbAziOn55x/n
XXff3uWcPiYUo5/c1v2tknvLIPeqY+MJDq8ZHD82UZwjWzcQnfeaDysZp5l9l0xI0V9ixKmv6jp2
nNK7gwOPZ69yuXFgvgkk+CfvttnDwECGSAoiwD0gGG5CRP/OSAPwxh2zHGdGLUbj6haKL+dBaUSc
nGAhJQ6szXS242DZ43iQkAXtVIhjE+2ytwhxWS7133kfEgWvQHV29sjQTMRNtvjP18uGX4HJreh/
hPUz/8MxAoJU8O0pPm8gS7kPDhPx4UeYHMBX3+9gfYYDQMLVZvDsMgSu+tFqzezDvVV9M+DppSNb
HZANEDkI8SpbRK+CrZs+k7D+9rOgQW10GX6TaUBqa0JPp3X9h9PasWGTIwfVBM0kjwQvuoR+n74O
hKCmzd2ZgK7aMnUxxJzKyip/oQeU6smtwoxxkn0duDvjs/mjU3PXXuw8F+hkgLyBO3e8AscM5zUS
0tYQVmdybVqQxLPKlgrorL0qeXecT2FQkxh32DcwQ0AHhwoTPFAzNpu1r+dFzfq2SPdzDaoUuCpj
O2wnephLV4vOrI6j0qH8y80YG4ubYnVZfaz85REhvUQLaEVK4UOIJR1c6sNXLifsE45rzgwwxjJu
V2C7c9zEYdgA9tptiHYBFTOmFfEFRaOuhvDVj32moC6xZWeU62yewfyVLIUW7CFeZdshkTe/uCrj
es/yx8CKbu6Hh/8au1JxSIg6OJpWXq1D+IGvjgFy1ytWbEVnXWIxjAjSD4DDMgeSJiw50Gg/JrFT
QURDa20+dY0DUEtNrBvfDFVLE1Q3EKxGr1Jo0jk62n4AOCHT7lNnI+cvboBdscGMZ6SNLOoQ/1Ik
fSe2fXakO9zPCzCgn6sxuVoWAI8+p/UGDzRhb+mvoYzSOHjGqbduSe2u8rc4/ymKEFYZG1rKQWvn
1SBgrU0lHyx21EmkoXax4mqM5lwdJsb9MxfWyBXvOV5/NFFh+rTPI0NZAI7XNbzu9iu2Iz+1mfgt
XHW+8G4yhLHnUb0n6iC+UMHgZaYwGUA33gqYygaeABdYH8Dtgm6v9X3mgx0SOUZnKpR9rK2Du1ni
hGpXl3OG5pY7XAmQU/pvjlLTaLBNFcQrjBVcG4+tIuKuLDq4aDT2GMY9yQbFNJoHb9koV3MyGznP
lsU565+yNv28l/IwhE50JcLH0erzPItkFMCx4ulrD5KGLAf7gfpArxrGN/ybPCDPEtsyPHsLUz5B
Id1FDyNyYrN6o6MCXmRc66BZAoQkld9cOcyEnC9haVNwjsxFSWLtWFUovEHVCDocs5T7zXKPsnjA
10URVycJqjpOAtXUkjIvqwTyCzVYxgJmZwx+u2v9kOHruqLtR2BMYqsTQ7xnpw/lZBmWahVQxT0+
NPzgQjbYWoNrjechqmAsznI4HQPz0djX0imCBiwSZbUFtG3LQ0rOq0Yz9qzc1+cnaWHiPTAE/iRO
hZ//UO49FsAgp5G8IAvjr4bNgErIyaSPyqgZmouWZvOA1Z0P5pPteyPDL+2+5pJd7NS2x+RB7+E3
jhYeQbAde64wF0l6658DxenUSjs7b71b7STozIoNle0zA7C/ALspeJmv9QWYf1PhgLYL3wj6v8AJ
bfR08d9V5ITbuM3GGWMIa/PNvshkcUPc47sFnYm1m8y8mCMN+2vobd0vvlBTIQwyV39gXV9OrtXD
WvESLF5+HZ688bsLA3GlhVsf0Srwq4wtGZwbxynsa2uFmy12QHsQctvxCrkJpK4nobBGmAvDvl0t
gY/Z2IW7sJJuJuoKRE/vQDTHyaUsyhtAibTef0ZRGx3jDvy6SVLEAz0gHVdd/AG0RIsf5/fjeIOF
8zSC2hRvVNAsOlULY+qwJy97q82G7DUi1PBMfGEflaH6/QXb7T7nkusvCygXYUQxbM6VoLMJx44t
I5bJlIC2XXnHHxsvAK0qVUS6WlSX1mrhusFN7td/bE8hsj3S90g3OA3PlBOwxTVwrwHS/QUHKvJ8
tlSjh/OVrM9cAQpZdviPlVQXLnvo84Ok1rDNahsokm9kkEBh7B9fxaRBJ1vF3x1CoOs9fsl6Akg5
zZv10NWtVFzFE5sDe14CDy2H7VNBzYIS5qf0p7ciKg3UWvdudooOUHb/5YK0PVE1nCnaUtk3oG77
FJAY3Z3ZnceyO6Qalu9hPfTE9E1zk0V9ylhMvtQ+OGIRYfB5ksdSQEkwz6OtCrqXamVmIawlfRXp
yg3wIxPJ/sy6ATdbCD2SDFzJwLktAn6yPMW7QFv9YH20AzjvXVc7ZJx+pwzpbNiVlBLEZwNafsMp
hD+/SuubnqweSe1yLh5N5LDkkOorPnHIifXTj6uByyz5U4g/nbaIU+R4GkS9PP8zASYuyjaDJpUV
LSsRum68o0Yp41xrD3ALV00SV+1ydCaQ34spbvFpSe7ig+bDjlqMrNhF831MYF3Quz86EHlF+Fhp
vGcdWxPr8fIQqfewQRxSVYUmauM3GZKHKTNW2X3xmdJf42+Oc87r4ZjVX505sbWcYT8XBIDsr4yz
gU7TsRoufSuPD0X8247PIBwRlMxVzkU87a1yjvTwZvDo3DalSJ8g83S/ItmP99IzyjTaShwTNJJe
HwYNz8vvwvbmMjR6LjtaI112S+CdDKYYSNVcCZWimATeSsM/D75riXBAgxLWFMoMp5yCelv1e8MV
kFanqbdC8YBEsuc/svELMOn+jexouiV3RxIHlFkiVgLsuPP5oWzN92XUNga0mw36Cm3QY9yrHjxV
kMtdFm9hOPrpFwODCocTUnINM96IOEzjYt9hNF136Iw/kPa7k9CYd0aPOMWJQtYhXSgUsHcmHE3S
SfUd++YIDaJeyy5+W+RWqo6dxgon4N5gvlz55tKSZpysNSJuOqHzj5BhCT/72vfjgOJh3qqZ1X5e
6luiQlXLI4VvlLxF59ZcCXe0zaMqACbHuWYJCme73nxHm7K9gl8QpXXRzAgRIdmbPKrt+UzxHX0G
jKhtEa9LWizlZn/Sier7ZZ6QvdT/nNI6qPyqRfHZMmYK8jQ3OUWQJPd0jE03TXFEkac2Tporem+G
Iyihlsy/oM/MuOWDSto1qMY5KQmDoccutPrqgC13xr9xnjBj1q8IrtDBY3MJYWAAppQAxQax0wic
OTqf4WNZ/cUTkfLjEPJ9yPKNDqG/W/mo5bOaUj/e8Cf1ntzVA4k0l19B2x1Ph5IS2J2x5AfBjMYc
9vVzIkf7qb3ZBb+CwXJEUhVszymoQax5DZsAz3hWCwWcY1VV3BiY8GVlw0/KwF34CoX8TD0cwvZR
z7mgb0eKJgXsMsgo+jB/fw2/OqWZZpzI9DKMCP+JGOZvo7s3vvE49f1nBZxnYwkycfUCYzJqBG0L
Unkhht8irf0zag/2nupmpVMmB2j11udBE6B+ybSltuYXL6NTttCTnRrPpPkkjiNRZI+VkOOYt+2W
sJHCYr29XF8uBIMk7oJd8E3Dd4KdLyMYEYLqc586BUBNSU4QsbA3opD3nXsMSfaSH9xrT/aZi+TK
GLUJzthoYQummxd1J3ID8L/4jVMFOSxXIV0SxPBGcWTGV/dqw+c9IeTPZFvCeEsEQeZXRFOgVj+8
/kpPfYJIPqCv4xI7il0z4tjuaEKJtRAaHhyC5PmUbfKgkz3T9hD1GxIN7qKxfDUi4TZa3OTSeLvm
iyRQW+DpsM60fqYwsZm/CUrDFriqA6rlVGqyj1oAWhzfLa6SM6NAzvJnZvUHYE84EXDOqdwlTFC6
cchFofhiiDfNdbRmcnwZvQd5onAWDnwRTpkjpJ+rUrBDb2skYHqTPxXBwUzPLYP0eJJZUbVpAR2r
pa5xFhD+ND1v0y061qKi/MU7TPTrV4DZMwgdMZgKyMUFOuClZnsYPnYwDZdMdC/y3BZzZ6f15p37
opAkm88CwcH8lI7fBMV7t7oQF8NZZvmRZ1DaZciJgP0u5fQxBuPvKOOmV1PB6teHXCog6NnBKEP3
0c4xncb0xYiLg6vCjJb0sKBfZnA8mYDO8GuKt+bRyVtb8uCzO6SSRu/s1fHQEPZUePDY2yfpN4UT
WjJ0q41Sijr6yIg4sqsTi3FDkMbbsBUX14wSli28rwibgrFBnONW91CfkgFBeCNUIwep0ldd+Vw6
dn91vEPPuuVc77nE7MRJOXzREU+DL0SqzEHYgcm68zNLsHm5LfRKHZOVs5lmpSXAs3w2RyMym8tB
ahdVw9bcTVSQHFo12MEgvx94EhNPe2gwpWi/OI6v9raDi5IIxE42cbobz60wsGZK8pb/Pxl49RZ7
tptwRn8TX7Rz7oqdqLAHXk09ooFcdtGWfxU9fU1zMJ9Vo6CWTFuwM6DPsu+4X8Fkp28wMKoIZEdN
yZPQUA4zw0cLgYXMs9ByfwyiAka9b6Js25EXClveyyTR92KA2PSTCTmbHuNPkP42x7DuKk6hMAux
kwCslZKIl2O2u61bCZDoJFDrVceaPP0iCyIfsexD6OdD4UxLGuYwsPtzkf+CUZ8B0EIZ3Tk7Y293
vbrq/XSraZP+G0AlFojEv1xHxgx3h2sdHhyZLWwFDfC0flhm4OcQrPY0mlWb4qAODagl2cSCrern
ZLiX3M+oQNcvujpKbsxeU6k+H+k3j7vX734T3KQaCUhdsrIKyb30FHJJuRE3WgPKpfPhmDidavkz
1jF7NZFvdb6/iBjR1nYa47uICJ2Tc+8keA45LdJ0QgI4oYEpexHhofdtUoYDp/fB2CG292r8jzoA
mC2+vnz46nTuaGUgevz2WRHcQYrZoLhrPWpLZl1atVgnlZqWs17Pxe1ocElGyQGL2EwYs9aP7Z06
buuGkmlPTzhxSpfK5ePwYAWEAYAG5zbvrb1+b5E4hb/75OGlzZHxiX9ZSpbf3lX8b5CnccUCKtaY
txCKjlAXXl8xwHSw+EEYBSJOD8dOqF3EJ4YATSAhXk5uD0xCdY4AwIOlUE35R12droa8JV97LYYu
6mKKvadlng9PjJ4J+9UL82onpXy6OGnM9wKAnMzFEg6YseVrnz3JB8AjqUsfX+gnkrVqDoQ5wgsB
E2OwD+21jGf+A4DIZ8SbTE9V/AKDj3haPlkIxO9YLtc2FQkGmQA0ySrrn+VSuFCecotXMXWKw9V7
oIO94JpFatesDYcS4QIrQmO2SyLGg639ZKONiNaDgs9HN2ZKvGPDDZwvsZ2MZyGfRSsIGFUuPraW
8drYtlRoN8HYjktxLRq8+s5fzjnj02wKzCvfpdM8ZYZdmIgNvsjq1uaFuFvvcKe5XB0wbeIYYO9c
uUe9In+0yCiLsh4bI49R+vuq3tL96SulhhNPw9MkEixhXiIgjoHIUOUfecg6M7kju6IoiioF0ysZ
SWmzWkX6nhY1vqwzz8fLMo/HgCz5lA2483tQTM/msF5+xAVr8e0abhkPZzkSj3wEgIQ4aVvkVEiY
mafhTLwEa2vrSAZ6es+VgEJsZN6CNi3MLpmJiy79NPg1ExAGJug7LL9I0jExeMhU1ER6T43dPbDT
lI1fKX/D/c6Uo5uTO8mxVzUroNVUebUcBWc9z9Od68IPNolOllQfCLHL+9iqA3+v0/MkWbqrEeBE
ep0dlIPiLvE7TBYfMXgERagsWW2tw8HRWlypB9iWNaWcfwHCC1Q0vxg0iWYsl+sFnb03kmXHzVZB
C/idtKmPOXAIrLivXlIbSBOynEOdWMl9eoE6dczwvMyqqqUWJrlbnQYedp3EaeUBjbvAS3Rf9paQ
CdB1hUtgypNpGbM0h4oaOeevQlOhg7VSRxIUR1ZEHcLnovittnxYyAHPCLmMH0J59vM2w/1dLHGQ
OepjDifABA1IJOJJwZ5YNSOWDfH4tEWG26N01LzAB7qCUTGW9O//4vvhDJBSybWmSu2AUfNteeYb
2LTt8bYighGi72T7yCqNjdOOIs9L/Ju4yMex4l/MKXBuQZIBtenCjFqfQV9P2TZDNP0FOvtgsQ9l
mMSrjiw926AIyhBKb4+UW+sOwDZAYMp6yoW0Hi1cF+2i6Mx2NxZvu7oLYLhmY2NhRtxh8i+ZtTdc
C1TQ2nnBxgwzAEu1PSpdmxrjcb25qMF/NOp9prZjSOM8Dl6rMtUY818TsMMb7UETf/ng7N/kQqga
sZaer/0i2lSF8H38x5DqNg54jpIkU+K+BXlkygI0qLzRRu6ZuVWKsWLznJsTdHrj45wr7GykTLtU
exB9KDPMA/CREAVfT9LdabFMq4XAlRXkIvTgSSACK+OuT2N4ZC0wibUuOm9BZNuc2MHI4k+h8Dip
Aj0uXC20JpXQdOSbWlp0n7VeE6QtvCZOcjDeUng+0IpS8EjnGVko3qpqPQSNWQ/O+Sv8N08Haerk
bpU1vwu1+Cuooy6fHc39+1PpfF3gdSKvX10ATqXSa7W0pL9JOB8vySFl3D0LtNHpBpxJs8BMeUru
YdTdIZ5n5PWl0V4/ZZ1vpfHdPDMLPs4IvkkPnwtIZxDfhlz6/t27TvMMqUTJYQwrqeNVfx7ek85F
ABvj7fBDQY+8NNCDgau4dm9+jsgyDKWSKSnmR2Hur3/VJUTLjBju72mHLWE/JLpbP1fj0IopeDEU
9cg1Dkk1C03/QRm0Gg7AAKwa4m6e/ngx+aDtKOlGOigxJCM6dvDb1v2dZLPYDVqbqaU3F1hStcMq
PoMx2IrhdA6t+YnPvxKGeKu5PPlNffru2SKEPjbIic9asEtgf69UZixyeci0VUjbEqX7hdZMdVTe
tVNFjfQews+8e25Eyf0H7NMQixwhnxSJB8DKQVbAMXMEg8tAA8vzL5I/3x8VZr71NfOIXOSnI1gO
PSrBjyTrP1oCE+eodJhdxcJfvoPqzeX3psrR3B/89yaNzIlAxWmJF2PX1wfjRbrbd3/bEHXt5SR/
VsQ7ifTWY6b4TyNJkoM+RLhR+lvI6fBC0IFR8Gev38jVmha5D6yVCCLZp8TrS0O3CXTRonqmFaGl
NOOU3lZIJUpMjEqyIuxlUC4Gp8+bSxUAm9HyHCwlXcbn2SM4rIn5q/s5/qtuRIHYemNSsSH6vHKb
QOedQIZqiLvJEtz0Ktt5rluAeVe+TD35Y03YgmKJ7S8HqRd0Z0NIzePvrokYRjewuvhQM3owwkbf
9rxwanVzSP2S71CmnMvhVib0kkNH3Zg93Z4uaUYkCCHwOK/A+gpyutyLQN9HASGXN1wATznjxQag
ZqPs5VW/H9iu0AB0wF1u1+P5g9tngrpWjka2k43vPKJPAurBA/krlpsTR4n/A+3IVTUy2DxjSIB0
8VS2GJWn7vhEalQdCtYWL50CCL/0JGSt1OJk0eR8sY4OXchn/V2PBOUNTV2BnHnuwuMxKdyFJnfw
R5+rjDCKGv1EWUFeqljUsYxfSaRhbYkHdXjPDV/GrT3SyPVpUYU14e4QedqG4bp/dji8//IKke+6
/XFKolwJiNKid5hSv3tlU5SuwgIR9mwjkp6OcNkK887IlftznFswkTtw/pjvMaJ1zIRdxOE/6yZD
iV0ffNhpUEBvhqRKa18t8sRHQ+mP/w2Rrf120SVNxa26NhYwP6Y88WyEvK9K1mHwXTeQewKyLYNa
6tqW8lKpNsEAHH6KHoJpTWu2o3E0dlfCp1K/OJjujpL+JK4YHiGMnBy1c+NHkVV2+NtUYNlgE7Wn
y13yMoMsA4fmmW6cZHCzurHO3s8tVfdf4qh29AzidWG3aJbtDSABJq5MtOCuutd9rBYoTA3CL9vq
EXKGvKoRRsBfX7grN8IjWBxJzYYlDDXw2Z4HfC6yhz19FBXdI1zoQDXRshf2Um2DSAG1A4FKVKCI
yae4llsTIfQ9rkZJVWilKZVMZIaYkfLtrzw1d9irhwjH7qH18Wl0RMO79OKNJ/mJcDy1XWoqinnP
5yyxtwTRHYCKUC6/xyD5bf2DP5/JBJhAoUz9H71np8tLAslEYDoJ/Qu0OOkNKE33DuJrjB+XLn/1
ynMuvQd/uTNPXHO9nOPlrOjrgDNqIgcrzXPm/1MrCs0gSsATSSOsdxvpYfcHnnUx5zzBzKGhZuNb
5qowS+e8Rd0A3ZKSWDKhKKiCCWKS7gL81S7tuDHl4TupBle+Vt5W5T72SNme109+BOnoxT3BvCX2
k0ROYW5LYiVPVe3e6pxNeb+I6Xf751buV+YmQIrPd14/QcpIPHIz1gPzH4M1KxOFfe27dsJ2lNko
v9rUYVFrYn1gRa7ciHWl1nd4rEkKXiZfqnwNRqgq93y9INLRah+1dsYt9BFzNFxwWAooIm9G6A/V
zHqLy2sEI4Wmva/tloKCRjphrQU6SCV/UXhgVxqbFgjgUhLvHaYXdvzpy47QoqCvNcKrUHb1wAXt
RCwgO/XGhfaCmpDDQx913DtDb8UWXtRtQ46DFrvHmEAQagfWev51hwcZ/0nehN1ospwn7qpUMMHg
e0gxeOwynaNk03PQ3ML74WH/fBxetgC6+t0/0xllneHUNsSubinU6WPuDghyBgA5P1TPZHx7T2fM
XUr1eCbCjmGssyHquTmptwWiMYywUJTNMgNb30HYGc0wc6E19TwszsdDOLChq8qydYLos3KyTc1R
gVhb+gg5n3uHOplbRbDwA57i0s6C7VrxCwBkTVX/1FqG3De/jHnpfzQ65/ghx+KBfqzHVtAxeE79
IDZteI+FtAB9S6zzw7mWvYaz7rMG/nxNIk/jkT7iS8DXvTOFzmHpnE9llanQtJzk+nT1/rEwvdla
+HV/PPv9OGcOu+wkUjpCnkFxclmHweFj1YzVwRjxAL4fGrmOI3+sWK8aHO6EhQ9sp+FEPPUhwnfi
H3xd5FLpPmB+THfbtOjSrj24ED7WubZo3ai2rqKBvRIafL1a6L4gVrgMo2C9ydEL4NTRRiY5R6cl
lXuYoHbbpWu92glQWWEqWTt6mV6hlhvPyfT4YjEih7fU6N435blcXrw3fLvqOyIHYAx0joq+zxop
m70Kja0WpJnUxGRFAHPwnBhulVv58lxSQGxVunUzFpfAjubDtzk2Bh9ItN00PBk5dT5PQmdhQ6Wu
Q4EHxCSNykXY+CWV2bxZS2fsPnWQiFfIAec0HjAZkYDRECxoUw5RfH1B9faCpxQ5H4DuuIrrF7Wk
fPH4IcY+4nACp2E3rGIv/D9Wg6ea7mmeMIt+mfLziDXeT9XTxGcs3Qxc26N9jhhajQoeplgY+p8j
xaPxquioOvUZZebC1wRtp36JA/XuCdDoE+hbyc84xPuTeEDxBh+FEs/rjGIeb+rctL4ZPXDuFDS4
PxGAYIVBTE9XuEKJXQqhpECmNhIzgxU8/gdTqlvWoeWxqx+EG7f+EJPqjAHrbbFyfTA3TbwgGhPj
lKEaOkDPhLxf3J+2drkURdFfE3GYq4CLq93BfLixT++nqT4qj65v8+/nwO3mmWD5D/Z0s+OjT/tu
XyOCFOowhqJCw4pT6TNeaZHWHolWLnw1mD9zhyusAw9g6128CRGcwVQw/BQXMnYhEOHLcbOtyx+U
44SifpIZjnHMpJeN+qDK0eZvRkJUqnYC5yOHwOiUgU3TlQUKUOLby5ucIEDL2mFUzgvRq+uKBPtX
NQPjJZOa5+wc1EGxFZcrKpUxziv8XJH5CJaxOwwK24yIQpwSW/kxOJWEm3SXJxCYGKIOqBEelaix
NbgeP5yMJM+SjX4t+1Sih8ty0HQ+u29XRrkklqs/h3Kvf4jTUKNu21GMjjLvv8h+MvQbTZbHGLF5
2b8Np4m18D6g+HypmxOwP7nHhoGNUFbTgFHkhC+NhEKh2fIvb+bkJ7sE5cEhxV4j5Wq3s70sORHe
wm7cd4OSLkQQol9RAtuAqPPKdxXm6rAS4fyHrp5Q5QurgF3zWu8FUmVo2x3ehjae3Pe9Wmy6dUO5
X2YXvVX14PbnsQ0QoP8kj+FkV4yFZAawDgUzlB5XrupTVKPeqEiBFhROpnWULTWbS/F8DixW1ksU
ceyBG1MbDFyeqTmpRwmr2OhZSUOJoMOcy9WR3NnN8wRLdnyLUzkgSzswZdVQmSXYSwq2KlApIyUW
HaDOLm7f3UuHUby/ADlAbokGYdkNLl5AKUTddHxi7Udxjnh9ABPJDnbuRkVys83+20+4Z8bPxDa9
JQMGIpCMzZX9AZpMDVIWXhEqgxW/MjokylaSjsUyKJj/e21EEDbmyeXc2xO61P6uBtw4Z8HiNLwa
jHhixpEyYk0O/+qhPwR5oFJVJ1RJ+QhvFyBtyr9Xf6pmMSfsbQfWaKB4xbqzG13iZj5t8pi7RBbp
70JwrSF25LuOPh2FGSPfSkTvoTG2P60UQrXx3MxsP/1aH281we7YavekukF9e0TF2cfdvRKxLVCb
Cs6ALQAUMYhCXyuiikK5U7V0HzJ6MOsYNtC4MMGcM3OlHm/FByePBl9NRpJBMB0Ig8EyYoM/2Hqb
2h8BArITHxpwaihCIB5vBORTd9Vn/V9CWu/Lw8diKrPY/TSrttpHMK8/BS8HADSpSVgcnY+82/n0
XkjHn/81DJ7hN30+Ym/W3zoV0wosjlhSkKrN5xXSvuNzruT7PN7Nsz55BxbaQFYLghPJIO9W/e8A
FAESl5rsd7KuhTJUuoWBUDKsUl9kSYxRdn1BOfeBryzxs7H+ja9MeJw6ozTi4spilFhw2wPntGfQ
ylY5kPwvflcUzpRRZOEdFkg+95TqWBK+aXxwq+NB6Y/EPqkWGZIMZoQTRY7833NcQZbM/YbiJUEB
0moeKI8ucEzJIIkLlo+DMTmE/7GvhqpO77ZgHyzvXmjEJAAGOfFmKb1lS7OmirehsHpmAeW96zvs
OQcbebcFU5PDB7yCLPxML+28/paGhakXBj74BYO/W4aZpV/i2uiCnHNwhGn84oBtKOUusRaQrR7G
CtRfDZtzL9SYagQUaK+BHq+HiRT+xVvXOzrqjdozighd986HIINbZzyy0ZGXXB89bh2tGgXTYTd1
OIlYa+vgJIPlhOFWmqtz0hvPKyO2663d5wayUxRLYWT2dpZSnD9InwuHSSyBu5lp7VPoPI7g3UwB
4SfzfDg0Wcq0ZHPZI4t9yGqhKNj8znKvZDp/Utg55u7A18g0fHf3qNK0ZRu5qZsqCcFY6M29x03g
GWSH/oCbZnCLc7DdXn2B3nYjVjKCld1a3VeOuW0aPoDNvy0GSrjk9YZ4ndjVi4Inn9DvnQfJxg5O
/lu2Sa0tT5NwsradSIGODASrQlxen5VoXu8cZYxaQf54+pxK5Hu2v0k4eCnzDuRdJ+vsmgxMjazj
8KQehSLJMB1fxSLly8FtkG34rIkkPGGiR95mIIZG65VKuujjw2aipAqyKy+Xvs2r6UxVWIe6RsAH
1cA7CRiXb6Zk1G6wb4/R+QD/tbPU89ubmtwpvtHYp53HDCHQqULOlvuRWSHetiLyjUrR+8/W3cxU
S9C1GpDVFOE6nZi6zJ6kD1pP5YhptiU3MnDGRdkx6bXZz+1Or04nhAigLjYrh85M8MMMc/RG+k2l
ka15l9uVZasGSHLIRcGm/0p2iVBfZqTw/V5p1+K5m2dBWboNTnOjZUF/g5TwDa/Ev79btNMZquJl
k2Ukem1f8aH5pkyNghP3z+r25Bxo1xzE1mpePiP3GRxMbZb/qzi2Bokmz1sXLkXvblE0uUS27iO3
QYdaNcbYI24I58KCVlGpZHJ5qfZkZNFVXxkHQBRzcHlRimdQza6bdh/zQXCojI6Lg3Bk5I0Sty3s
kiWtBo3uJMFl1ktQpFxdL0uA8Ztlayeu2XJ8fsTVvsyP1Cse/EgaXsR3s3g/fU2SZQOQIgZPN1Pa
/A865Nrgsr25EnPSZCCtKXDG84q7iM0MLTDM8kr0pLgV1ZfdmGYTbaTPGsx1v/ejDfwSy4BXhGR4
uHY9ynE7FhJPeyvNQPmhGYKFbFc88EVjE572cpf4enamZ7DWRnhRu6oOtOIWJ/CotW1ok0uTurXX
tLsdv9dgkBk8/7yo40a8bocx8lPz2ZQlzl67mKJl/lGglwfY40GGyfmMvzs5uDn+UuCB0up1v5aW
KcQiXEH86iXflizcAwYBBSBIUBbyQuD5u84+WD5QuPJtfCv837lUFE6yBaCDnNaGTaXzVDTIwdMH
1cHHJykQs3+zQkkOtu9gns4yuy098y2lQ5yllyn66Uq61hbbnukS4pOj1XwZeHNsA0DSbQf1Kbvp
OwfW6QfWJSvD3NKl5wzfi1PLg3eNpOpIKxRfrSoMf0FGxetYJLaiCVpGHmp9/TMqUoN5ivmRXXCb
o8Y+fAhZ8DCCbSxm/a5VQ6A74w3JZliFxQ3PaG7oiwTw6Hhymsv61O4NmzW/miaPFcOX3/b5LN2w
bjvkN6Dp0k8WLgcMT2Y9dasxcfGIDmyNjdukZ2jFVwLYYyhzLZq+GZVkg2iO8e4Caoc6SEusLxiG
uOs8FeKdW+QpQGsxS5l6TgQNw5pSeivt5y1h2HhHiLCaVsj5eXG9cEXsQkcrcmk5KlXyg+/9ZqhS
wXFeW6l5DSgV+vRR/jmFTWymQTtH2Cm+CL/f6AcAdXhb4Y0vY8GXoV3SOiEXDezEs/J2iZJhKFYX
870AyMbZFp+G9lu1rh4O9rmryc0WjVrwJxlKTH11GRX3sqIM6A4+2hbYsRkIjUIMWH/N1pTSgsb8
7S34OcJfDiTL4pE38ey19gnlOE6SLZXFd+nfoeyaAWIOMboPrFprvhNvmJR2gAiwi2qyCWd1zxqh
kfFTzFSoPuvazXLWPYRKTAZWjSrOoKccBLIUtwrQB8G1HZU1WsYBWWOnXzQsqaahVDgEgsmr6Kuv
Fp5HR+2UEbQskAZkoVei2gGq7kktLnnEhRStadPVci8WWsh0kurDzZ5J6ccFqfJFXLpGMfSt4/ZO
5YnEfi8IBeytjMe5zhssKFyDGM2JsGJ1lGSTgZ1LGcq0vvY8AoELOyAO2Cpkb0dsRcnjujaGkh83
6hw2gLCcltm0khdPkAvY5dFO2SSvaeXZ66xcxZx2LQsnvbIwlo9rxNl9w8RcXgmYs2zHgJI/IqBo
haMmAlhhjIyEgpkqsPNyMTv932cz98UecFpP3y9VfeJQTugLro7qQVK61y+cvOrB4wzm9Sk4LgQd
nyiaIuolVo6VNNdhBDjjkkHlaCkVPrUX7CS1mEmpG7e8u0KGjSj17h23c7cyawmxKMhKCsXGDpZe
dvrfBXzNh4PodW09IDQCnExgZ8oQWL8iRevPeVY5qiYBDZDAUnVYe8614/ONgHsRFvDnl107N5ll
j4EewsJ5c1anRFyJFX6N/BUwrLbooBFMY6m70g9YhurM7usrT3ssYp577uSS2R8Z9OT4hZABiaY0
mjDo6iLd1skg5z/1es24NngrFV20t4BkXTb3pNQ38NmmJ+X67YgMGha3a6eFJah0bwWh1OX1rMUQ
5SoN929SBxkQ4ZQPoZAXQd+njT+mPiIEdCZuVrremq05zCPNYVSO9+HyZr9QFRhz7HxThvLmwk/x
vnz+LrTwjiPJZFMGWJaGFisn1hYK9tofrgNaT6aOWTGwhNY0gv8hZ7eOLfomKfQQXvv96+d+J1E/
002bF2xoYvb5qLtyWy+GUN1DjWpzK6cxGLY4EMbAgYccOLB0+XuKPKIkZzBdsAzGWZzuJlmaCh6i
k28xnqn4vtSLqWgHJTRniyk4r3w6dD5YlUw/2hDqzL+3ycV9vo3U0sT8mBz8mH1+WAnr6T/LYcXV
LrwvUk5pBxe1SKpM5ewJi40VpEl2LAwPrGIb0pvG2ryq+eTqwtxqbWRCTNDEeYk31pkDYmjEdHJN
kQRGPC39EOVaHFX3rc4Z8Z/cykMk5gGLMwLxIQkpk0JkL4trRQmHUkgafkicFUpzinQk4FuUgna8
La7PcqY6X49sJDo6uQQBvgJG9RJHvjK5+f/9vXMkbBIMNihPaUzfQ8wqUektt4MzZausBmAYjGxl
I7Gv6WZekH+uzKOrtxrYvhdKuILvWSXwdG4pQCSQ0u92xCMEJlhKJWxkCg7a4GS029R18iUG9dew
J3SSdzMCe6y+QAMGQ2TbGbQcbho+vgINhwtZVdTXtDnzXbUNahQbfcsfAJ8izb6VDmIwmN3N6IFw
s+zbN1zvwGLm7wOXXJwIOh+I8hNCt2lmIhB+mlk6AvzjA2XkLKHuY4tAnlojEY4R+lfCQEhkpy9w
O02WxDOFeFG+yyDOCnKPHgSwVyVf34o6X+gXMqzd7EchihcAeVzAFTb620YR4+UMRgfmiDSWwJM6
Hnn0T4LC8Opp0yWZ//R/tlIKpTfzwKrgSSeVpU0cZsAFC/ZMwhwDyFglMCIhzGMYQggw6uZO2DyP
n3npX/aAfWggSdeSI+cbHT9uU9pey7zhE0yt1hDqmAg8KFid1OahbpOz3xDPNva8Xa74Ecj7ARmX
3RpETxQwix2/ckvPdZlreDCYFkP93LFsIjOnROUbtzBMFbofPqApQjwamAU4HgxKGsQcuCGk1nFR
UZUVUVu+OaUrUjQwPa9boXzUVd2PNDgYURcNrTLAQPXRV5/iHLQYLNzKFnYp31A/9+uL6C3cabXo
h+Oqt9RNOtJbkKxk5G+gU7q1Aw9do8rzVE5YGn2qdDu7EkQdz947ts+Fqtp9Y3dRaNXbc8Er+cLs
QcRw0my4jRKauCKWeRwg6f8FI5IJuzsfFMBq8Dxe6499OOgWMqt1liU2I+/hfl5rGQquqxrpbivM
RVCZG3hozF0XOGjOTtBuYiYN/tKPjIZaeoPZ5o/QO7lqgLIsELOtp7eUnsjTED+8HVVuinJeO6ln
uuNn9AQwwslUQtWY6mbifbYT0elDIBkR10xMmhgYXn4hYX3Y9X1FKQjP6anAZHB/ziwn/O2mYiVs
R2RZGfxXA8n/DXQF2ZzZacWwLBDQsqKpBBUH+0rJ9ZbiWoitolBG+GCKer7wUd7ZlnQzfEGkDiH3
LSxpDcH61gqth/r+Pviih3b/YLKZGaS2Ek1z2i0AkYFN2pYD4m9RJXoKdVemJ3UAOhUEG9Y5Xfkl
XOVTd/2BdcPPT1FmQwQYkJBMUHeHDKSnK9k/yxKauqyEwSicMj6xqhzyzKH53fa6ZT2gJsIHdgyF
RV7CxDxBuvb4nn7Mty0NRFBikK4rMtUxw1G9AiA+rqb0yAk3/ZuwdCRVqmHExqQsohNjl3MO+khI
v4aIOZEzlGWaIalccC9/UEU5rcJJrW3G2Dh3FNPsPwO1sM4p0fefNtmDP4RnG6uXDqECb3nUaJFC
R3gB3uRAaTrQu2yK5GZnu3/TRGlDf+9ylVC2neme4S9MuuEORmP3iNHfcLQv2aKxytVgCAtE8UOK
NB/2AmPZcJME0zIupBNcMp8BLXYbQ5K2m4xCIJcgEReCAxwsJu/fENFjCtAtUjT7HYlEI8A3B/fN
r0+LWSkL+jBwmod1MMbI/HW8zQPOL0ZZTr39dpL/LfXfBokwGHGMf6lelQenTKTvpTv4As2vR1Il
/q1b2LPZ+ZQM+txYJP1cLzLGXv58e1QN3thmfGmbYJKO4awPykpUKrV6PoDvflpSU0LAiOaNk86t
KlCj9aUb4heduIborGEXQIXN3hIhIUbW51miPvmTiaxZXyJgunLAgHeQBaS4uxomfSzbLgaAXy3A
CINb7EVUnpC7Pjtulj5WXTjLwQhHz7bBQDRHdAmTHRn+R+flOO7iX3nCoEOvQnW+qWbhyDICzgbL
vmTD8DDgD7hnRmQABxQjdJOpSvXndwCzBgu5BIVoVP0wF3VNNs1aWS1PtoXj00WRgXMLwhANXfit
TBVM2DF0My9Ke4n5NQIucWqJW5BW9evW/EoUMWqTsP7hchna63+vAjnME9VcXbj3RYE/Z71I+gMZ
lSn5GTOasywz4ne9x+XwuxZTwxDLXVgMxSI4rjYUpXg5stYZXzp7cUNwePBBy1GJYS4B44ouMqYf
6V3ERh2p0ytmnh0clLxz3WT73reFR2aqK+MLPMMflfzTvv6zr1f0OZGJpBXY0E4kPpH0OThJ62yq
JymPiTxjt0oIUX9+D60WCyBg5dO7afdKIeb7byqqi7407lKuHnB/oHXPU1X+m/Yj+RZzvKs4dQRf
1hFdcJg6A+JPjVOphtBiyjru+ImvkpLGuAiRPoKGxLuzLwtLOLSiWPbgL6BeaLVo3rCex9pkiRnq
UBQSkPrRWkONnFjhtMd39ipup6X9BIulBPKZ38gPaxC4tRGpfDzgg3pJ4pFARcUK0vZxjoznIXbe
9LuWlzvrXxkVbvlVC43Cyon2G8IkYnBIYF5kcX/mVG3Uc5KgjeSvbPFM8Cmmes4oLUCeEqmrsMN6
jC3wPh1uaNhZDuoS19B2ry2Vudn4+ZfegKD0caTrTo6GATis08cBAjdSpa6LpIqKLkvGmcnQvDEH
qWLTmwhAsZig2wfiBF1Vg6W2ZDoHCXXvyM3HgOwJgDcFC5fxCq7peXPlBOvwNxgUoZVlGjuTAtE/
474bEiNr/c73fkJB/WyBXWV4qERD+69u4/1vSc5LqIJeRSgg7fcOEN7jcv3o787u/4yaBxXlWVSZ
3wvUZu78o8IkDxpP4eopQTKSidBgQ1VW0ZtFo7xB9LQR+wnA6hL/Mw2chEXckI2YZnsVmCXUhyYx
sItillNdI8QwXYrIACR8Dgk5jtjT9rKaKA1lpG+jd7sKD88QxB5PVFKIcXVByf33yGxiT1RE90M+
WpD6b7nZhFOHEpkbeZdvMS6zjcUF1XlBNCiEfPXl7uySf9hmtT7zDSWbYjd7JYUnJvqBwCoD7OZ/
AfagODKGSikKeH3IkqLDbvnMDxOpHSv0DaoqAuQo0mW7GmclQSKoQBdCrab8Ir6wUEv1YtByjhIf
WDpo4cz9pWlUXroUDXtCBzy08PhLT914iqlDyACYAexRJoTOtE3aXkMjbMgwo5gsYm6LXYIIbO8l
HPq+lAkQSNCjK4gXu6qz9mY6xwFEt7d6i8XyuGQcP1JitbVONuzvKC0wUDtNS6BpjbVr5nJjNz0U
grdHDiO5mf65Dmy3WJXc+niD7VGbE4wQb7W/p8XneDGJ9r/sYw+I+5MeQ6gQwTZBIRwPX9YCaa46
iWdmCLv6NGDzvJ2VrgfVzbAYdtjzD02sx1CjRW8cPQaU+JiJHjMGmIjbn/3i6fhKyzL8r0LbmOXv
wlc6HVASh1hOAr18t8h9kXaH8MWN5sKzi5s/XFDba81pAs07wA8QARj2c6f+QdMnNJLTMKuH/3JE
2nz1gnzGhSFaz7SMwI7giadUiO8MnlbaZtNnjf8FMINBoqOK4S0DzhvwFV+k6S7H9UYKZyqt0nqG
KEJ0FxHvw5aVgjAzYUOr/OkRsXtHEZ2esxm6fTdcouB5ve26FvmfaX2DfbQH8/AwVQ5NPdxb1eCm
r+QKbRSZs7ocVzRJjkVtycIAwXjvbag23hu8bLo0Z1J/NAf80n9V80O3WmuBnupu2XnCSaDukgpa
YFCMue9msf9J46Ma9lS4KPr7yxSkcSVqAbwzeUOumYsZlwBkXbD95YQh7N6Ag3cvothLBjC6co+G
9LpI+TQi45C02oAyidiQ6wwP4NFFY2H9KUFsdcc0VbbpkbM+42YWuHikP7/2YoUmJ8v1nfuJ0J7j
C9FJwoUIKYoxTBSJzm8jWOY3JE/gmu/B28u3WtJ1CQjnGXM5uTBcoE0oluomTChtAy1gzKCM65F1
C6Rn6ow5mxkX37L3Ik9zasBM34nxzU9v4Q/Hgi7NPFBDfG0+2yVvKTtpDeJQtP/yK1aDsJYLNzUv
JEZCpRT9BFLuUwIdZlkXWw9NzMfD5lyqAwVILG8cSv43id9MZCZeuuWqUczwdv/6HWMkBTptFuh2
qfDeVH8GomCRs7Ajfln4t3RV+49C24PFowRoRlpsPTXgw9xdUDEVEp9O/E3Lw0wH1EaJVzD9VnBe
9eQ/o2/46gVe8meUfmTbpUqk1o5v9JxA6NquYaRVw7QmbuGnUiwjTwdpDRRBqRRvjaKak26r4wQO
qSayrnSIddBHdP09zoPsYrzo0dTxsuFHQahIV/x5nBd0s/9tq9vifPey5lexz9Nq7MEwqC1YTrfy
ncMWzCG48Y4Gu8TMcWMoj1XtqZlRwMwW/80YTjzBNEWCACNekjeGoQXvD9dc/3ETMEvcJTkId5/d
wiTfXj6AhEslkAu1S9WL7NR4WQSWqoQX/R2tRb9KPOJzxBXqaAL1rOBpbbPl/N0NoaJxT6nP3aXW
2JW83LAg/yaCM0VHH1OOhTtqaRRvcooO2Sv9wNvTT2K42mN9nmovnwB0Mt8BHQQ73SDVlx1NQg2n
2igPkVIQ6DGZRrnAtIoUm1Ij3nxEFmuNNvf4JLbsJmpi1cfNwAlmy3avgHYrrogm9fFT2LmpofQ6
0F9YqTPmXjaHYyQGfziapsaWYCdbq7Y2iyHMDWOGSrdSml/Ll+jwfHM7Y7ma29KlJPEOcI9TLrtA
hfaK1kf/fFd6GSlkaHqWHdyrPLTOwLDsvMdfBlcv6LYgw0vM2IQZebvVn+YIL9+VGCbowu429dCB
5TE3lXAolLZRf47M2qYkgpi6K/YaaZT3WqHeGLMfoHrsLkFtnXosss3HFvoNXNCsk0lzj4RloQx/
0VvKuu9fgiSZlUTLlAFX5kdrx8D9dPuEuUe7P1N+6oRJVNMhrzWv/wdESS5ji5yWmY+AFnmz86TP
6JLK/ed7LeRNOLz+zhkdsR+i1DrMrrtT5mSvR3U6HRfW0jNpDWDeqNTH5CelBzpPEG4E/Q1+Puoh
L/LgGt0tkH9iYQLkLJUGN5Z9jL2AAtqpBSv2Yrb4om3/mHBsaShT/gUdfsFo/TeYz0F0yBiddJcH
zC1HNaistF4xxzD0Uoj8Aunt5jyKsQlpnp2C3Ei8QsTlj0IJ1OXnzB/j2yR5rH4+UMKupxx1t0A8
tIiiAqpxdXGOt9ONKQGqjqN4Poj3xl8OqA9Hb6d3f0woYpJzPir7QoMPP204E3Wn1vd0cqcsgCf1
Nb2YE/TC4t4zcGtfUBmagYJkISIO/LiU84Dbe5lEVgvvxomfTSjPL/ZFfHIAMXNxBpELp1VtqQhf
Ec7if8lu9GLYoskYFxbb5HWzfbh0G3TV/fYyWQ/1vqv0GXisiHqgiiWEzOsLT/ymRemDL3egsgss
mPagJeMe16zbpk8PLbvJ+La9Z95D2Qnk6sURhUr2MFmWJZtxiYHas1CXOsT5xxs6gBM7is0FSNLl
P9pknMdHNWjG5DuTk+0hkr3li0q2O254Ai8jk05lofeSWvKPqxl08Yw7JtbcfqN90zAlfIhdIdBY
KvZ1p+woNSP2aW2aql6nfHho/fVmb94mwjlBAHwOY9Lg6FTPwB0zr6b7Uf6wh+4dfOX52iFiByTc
5NJ9g1/uHgukUGXdCAruW0hcayoyFf9RY7DhBt9PAFSrAXRu8c5+Dra/T5ikiJyvcQqFcojHV/Xp
wmHF/GduRE+3Vvk8I5aR2MI35MigLSDxoW70BrfviYKj6zO20ClVMw0ciI2/5KLUFQPcQcPnKGAN
9+gp1jCVrqwzCp4/YYWgmcYT4b+XtFvIAGBqH4P2C05BTFOU+97GFnJ8g8RU0dN1u9poOuld/TpS
xUJnTIzRLVhLIXZYvHIMSVlzcLOpjh+w+kNotavS8xURvf8almMuwLZJsQUw+P0gyJPVHOi5Cy9d
v3qwDQSfkCNE2K66F3eLSdRzYNdlIEVt1zayIeCZeLNrPhM6teL8quMTzIiv0pkL4nwlu81mxfY8
Lu/1jVkmhgLmrJ1ZsfZNl0fwvPr/08qkeuRReXzd2wvy6PLkVfhNlbk9ttK4PQsGPH6hu51wb/Ze
tr4ad2Ci92ybyLpImfFzaqjT9h99DdAZ3W58d7hJ3GfYfSMOm9egGuuiL/hglTxLhnxABR7g0nW6
URM+OjlCp4Ge5HLaSeR2Q08rqwEccZn5TR5hfUn9swbBd0TIdcecAcx2ZeRvyfnEWXy3bCsw/qbr
prvNKaD/dP4gPylLgCHfdnr8rcR0ZTcXv1ugDwl9zpZsauo7IRRXyaC4Dx39bYnCUFCfJ0TOaJWQ
p0+E+2P+eXrgBu9wcF9OnranS2XirnINlGpRuX1+FkKrGUtCmyin329R9tHhyJz0P+YMYmo9uCMh
xGceESNMSwcBfuM0Z75ITgRQVezoyWcshQIqedTPO4XQtws/SPX+KtZO768V8PC7SztZlQOQSCWd
qZMaqzdb7p6XK8XOP0OUMq/lmOfHi9iCMA/1nsHTMWPqoH9lEtuDtnOUgl5hPMeFKqkqqJguCVxj
D06mnWkNnIDLY2Q1yi+E2CRNhMjr328N7oR7S5LC9cstxaaEcHdll4w++RHhbx3NsyuYGpKAaoYu
7aJStD4hFQhN1RXK1y4GOfUM67J4PZNQpErt1lPZkMfrzQvoZCcGYRnUc8nnqvOsSQ/IW9TRbwTJ
rF+cO0YSJF+iLCslHNQPFEgkypyIUlyajAjE6GdiqrTLnNq/SJJkllUlqBCDARUF8/vMPoG8SJBN
0gVh+4kcOg/O1TCvPJct+b4KP/JflBkBJ8URwmNb3y0+jzHOwW20IkGtVsnKlJNELHzu+UZv5825
QVXMXrhYmagmz2Lbkk+wut+ekMmIMH7yJQ9IYb19OG7mvmDYcRpDdbCLGONhYKm4BRJrvP5Ib/DD
D0iblzlIax1xMuDWT1ZSEpzPHZ3vjDYxjJ3ky+7FGrPYKO75UPc4cOW7GkgIKvsPvvIkAtDqG+Bx
RpfPf48/4b17Ye6Lb+3SUTO5ra5LNW4+AU+yR3u/RwWhYEGTXsbvXRmG2smqFYuAyJAUipGm75Oh
n8uIjSuwe05n1DWbNz/mKB0gBaxpgrK7JeDNZFMi8QkVtEDXo76K1ySfda8PClc0xfTNONwXxIse
8oLGrsY98gQYILcHOxjff+Q9LR6QkeYF6qlWFsfYvpF8KaPBk2jik6turm2QOrWzR+w3thk+ObjD
/BcWbncNylV0f+Jy5r2Yz2xioIm0avoesdza/N47tOKqC5Hsgfpos/XZyn2yyHU2pYASKQHtEawz
YOBM4PZ7SmEfFCSQnenIhF7a4wvUPJa3Ad+8Yqrpm3yC4Zzkp4UIULJNh9XE4YrIWdciI9qoD53r
Derxco9LYc86ZzZLSWvXvCuNtLQj5JBXvn4E1gXUvSRXpIOexNlnV0OELExhmrEeUbjs0lzBJWkU
vIC//gcRz/vmhW7VjEvp8P9wfmbh46ZenUi6Cuq/gskQfYGyzCKxz6P87c3IUP1dXFdUnOOFZgm4
7Y2nl765CrqSq56Y4fhiAVHMvekSu7tkkhmK7D4QE+qyYtm2l3tNoqOHZFhpiC50vZD+CYlVgUmQ
DNJSjuOuxgP1wNoDdUEH0qhbIZ53mW7KmYsS1YVH66JFh/s36WrZsOdfNfht0IWq4ZDJIeYr7mks
GHnbPpxEtTcZZtaxGCWT3zzvyTtbmM52db00Yl86vjBqiddb49BiA8AVAxcSOgKKKkCtBc7y0lBP
xuvn+ThTX52q3CAgfxEByPgnK1YG59Lq6f4mWMC/tx3Y5UPK3ydD9NUOLkcetZv9nz/0gEyAsoov
xlaP+fGXZ8iyGRK4pL5ryHt+C5OZe9xrUyZe8oQGLwHf3ReVxt9qc1UUdmlX7MOignPyJ6Hw55xQ
w3HRm+ShM3n5kx7eBDtuzn3Jr5Q37m+WhF9sCxgvNNsoLJKOA8OW4FEmIW71p9gTfCDYAYP/dCyO
6YCV0gfomgZRMP1Fky+hmFYvabAzRyfq0CWVSQ1bKTV4OHoYjh4lLOgVRGHi7AaoVaitpdIhTGDv
JDDdSrNe2uZVpKlDwaamxKaM8piXvI21H8v806ZmizIbZMy+9q6yFMC+1ILhKETnzAqas6//8LvO
3663GQdhr33QZzCP7e1aw0UatSrofbm/iBuIeWJTXPUBlgyPKxKKIjhnbT7ldTQnbS2qN50RztRO
hr7nlfAA21Pul39Ki+hBhOCyfIcKRnlFx9W1w46nA23XVr+ZqIy3PjfejoyKe2FFFxXUUYvE1WJn
Q4dknmmcqfElVf+qq7CE6g3H7XuAzm7pw+lfGlIhy0zajygx3TB7eCNzpeLcS974FuX9xKqjS59v
I3jShYJDlaJlnBYAJT2gWnlrcfk/Dw0coiLl8TITEwYBTRBn1As6CUAcuGZKQK0b2H9o6sUUVLsc
EjAb2ubWP4WNTtbVmUWWBYA9Rb8ep34b63vD3NJ28OKSfuHyKGC7/u00cf0POn3pLWRXfJmyqNsu
D8BUmZyUTC7YM1524Guqe8UmWpmNCSZN03Qf0HnZ637clhUP72K1ad9XoxyIk43106kwlW1aa63+
+CISPIfwGvqJWIeVc98ZwE7bk2I0jEmVjbU2mbduq+NnHGSI0Cf1t3nQfKxhCuxOA1ohIVrze8yo
XgEYycVnGFiyQjlCdLYMLOzARHHbRWh7Pb6GV1h9x5Vb2cec8ewbO/F6ioaZknJGpFvTjfsjLTkR
eORB42mRmSqWYAzTNyXVB338vg4Y6ULfFIWegpkVxL3BMEi1MtCRfINxIDv9+2xAKVRR1cw1SBic
GISFOu8qhmkgqC5IR9Nzc7tz6VtCQToTpk5EYpPyyailB5jpHgGJVW+tNcUsATZJ3FgM/KojsHMG
yFLq+pJWpiOMGyDUn2m5ubGF0AA6B5ygnI/gh66xHXIsVLJqPrdDP2CJ6ELXDFyp6XoI2IDjLg8V
4k8vI9v7l6SRGYLY+MeWPEMcHwWIL+CWZFoOZwLcsOw10gGMbWvo1HuRMNJkJMThxC90df20s3rV
+vnr34CiBvUDDO+sWcmREPU8gpPipGWrsHNh5LqJqpfI7I6Ik+qQtEIJZU5hvYt4pAqzQofWDcD5
Ol4hW6ZQXJem+kiNipPO8SgtTz9bp1ZBAIw6eun+SDl2uLxlPGZEt+k2mrJXdmSO82ek8ImCSJZF
A71Lt0KKb519hTaPR0SvKljD+GbN7HzYVQyk5yXCpRVDB7Wn6nhtIIwHLQ43EjsINVd13hmabwDI
MW2UPV1N2Mkl8ZSPNGi7b3VEeHGm0L+7U6+FtQX4ssatf7T6bsGEaAHVc6OoLLN91DxWvVhUtkdm
iJ6Mdjkz/r7w4LtBk1o++ytpIsjL2maClXpdfFNG+KCLkVfQvBZQP7yeHt745vMc7a6LOqMSfgPs
K6PB8GWgaTOvFLHaFbGYsU6nFsL95B2dzqgxtVEC/WnGi/RvbPp9/P+efgcOHv+RGqDFcHSmo8n5
CAAIFpiiqDD8Tp9Ft9ESXze0FvdoA7Sk2qhvpdSG101s17MG3x1JlkoiXtJghw1FBzrryVrLRtjO
7nSf1/02EopLnfGAFDM/WnC3cIJ/m9UMnWmqWO4g1HjRfQaRgTnuFKX0C/0gxMYfwXtVJWxHkyLh
8OfYffRbe/e9qns3ktSyoSVvshqkdDCMAWiqAh9v/V4oM84V2cf4mPLih/LJFKEzVLHm8QvGYwcC
RmO1pPe241W+bMWORERV0l11uVkIHnzdbeA8L7CbFYHEF6IJZZfDQ1k4sPiHfAax+o86P8QkfDA4
fpoLqdXN6mpWfcmDRbGzzloDPVh0wLVFp5GwaJYL+dt5IcjfqEpKvtODQsFG6ubfZqrqJkNt+wth
3WiqZLYlBk3Ldn/gRuMi+aRa6xKswL2ZbGA2HDuEuAc4zcI4MC1wnlfK9Z+BHAHGVBfVC2rZN0uD
8/zpK/j8+3hTUKD55qoTqPyohN+VdKca97hAPogxH+C0L8L4dskWCJL8fU9d/wMxv8kA1BJ4QkwB
vSVOUWRTxoLZEzgkoPfEngRTXbIZBllTlGyuzin4FFUgizkBhbQOhVYIDHJNjcAnhCFbe6zQ1hWF
A88BB9mrldoEC6iOTpuQF2cYcKSGD82FYjuwjvQ28BLJGlW3k9X1SN0/SiCl3GXKAKWsY4vbU7Hc
0HZzZj95XDalrUVaaDty4Q+2OuhxGLgux/ovkdW3+T0S7M6BFpKUj2Ud9JUP2j4eKZi//lTmX0gK
smunO/lEZbX4gkSEhxyUiNnv53SfXV3oUwLkfgvZNqryuemHvOxXX3BdvjcORO7U+IupqA0oslB+
6HQRXOeo8NFPZVoGS6/df248lZTXba6cuws5GGEPgY4KoF4Jyv0r2XnTmFd0e6G9HKP/6yJNxEWp
AQEG2djEOn9ZR/rA783TB8W8W7o4btz8nZwR4tgWKqMskBWwOL2z9cKjVbaJewEZr8Lmqs/vlIOP
HsRZCbmX4BUl3J7SKCfZV9rM+bPPbopKj6qnVbWZAKQiz/Fp0JBJq1DEEpdtMaDyqClqQ7t1zf/N
BrQr1E2jZb4y6BBI1bPheovj4sK2eL7qPkz+LEDJZRZpquE1reL9vaoN04LQi5Tb9yPKeEkbXM60
rCcGPWE4l5qd7ePnyDLsCRnXdzN+EUkxdk6kCxhfxj0kIiTVGzbF5tyNoThTmIHQ7uXJJroqJqw4
iA2a3XW6TfSTs+dA+hrn99Pt4/U4Gz+34yd/cWfLGkyL8GE4kdO58Z38W0NhwpWE3tv1RjkjgbXB
7TCOtDwH7CFhaZ83QQ9/aUxy2sF/QdlTAnB1T3GxjWUXKnqUnV+IHvTyL6UbN5G1q4uEDcaZT3cu
QW5X3gc6SD3lezUWsI/Ory/YYEGcow5+6Moa8O/HU+UquOrYt1armeDXrGLN862y5eHFgilcX9gh
JNx8olWOzgsB6UWc/iuGRIDJoqiNAV+pwdz5ks7fUGZRGLkUkUSIk9k55wok6dRt+wSonLLexi0w
iJoa6dxCLt2Lpj/AC24NTMBuAOrGUIVj9Q+XQqHbhTCXlpsu+eHatL8I0GJo3wbwwRUzBfU+857S
a+FWsLydST7YkLHJ/L3s9LK2kfMLtuYYXyK3P8ZvIJw01ZhLmZi60Q3OX/NMazayMzHyp6IFkKtB
NTn/2T6H7+zQl0G8kG4YyczFEWxtbRTUmqTQO3bc07phhKVsucPPZUOcfzuERPD4EmNyEBIj2Qy6
Ci4fWY/Wy7a/X5d9BzYJ8nIK/SARMmgPZU/PYpjQtGNr+V8iog8i0naCFvqvRKGCsFlij2823BKJ
sUbi4avBwz5+Xs+SNer8EMlSUHBF82nTmeZqc7ZG87PQbROIUBu8ALxBq5fZMEFN1X6ycFiA1O86
u4K/Kvh7CDDV1+4tA8/9kzsETQXXcTtGn3Stkznx+tXeGFWqYdzmZp5Xl0am9MUTSivDq3wSvX+7
VAKkV+4AiHHyBIOID80yoluGHdYoaKqZnZw+5MUZiX6FZUCON/9I30zX0hsCqaTIP3bkLvBSMrKn
IIFMNUHIQdRzLdrTF0Rsdo5ggaBVlIGf0rN51Kvh6dvU7z83wu5dAWh+RMdUYQsVI3RpMzQ/XNeK
WfPRO08A25+2Owgccj1n0jzSrGHXsqN/8Oz7X6dKDWOr73crDjsxSYry4kOD3SWz3RjKzifr6QF8
DkB5fehj6JfyuPqNAX+KaT9gSUGjznROqhD4mSw9nKEyDQxfkpdSMYjrDMQZztXk+qjDT3UIY5UC
3C4bH4R3/FBkLOHCigBwWOsJLZ4nEfa5OH1ItLsedrmQKGgac1WSoq4UjUy93WnAq0VkGqlE9rEV
E8gBwLnNjwJS7D8gGYzXUxAEhR8oPfxsY3c3oTemEWDy7foToL4elii3o1w+Pjn7CE7Wr5i2UUbQ
2MYBG1l+pJ5CNUK67H1Mw1hprLZbkkpJmHTTtPtSfZhMG2E8rD40FikLo4qY7Naxeh+gGP+r9n84
aqNg5qraEq+upXSYr2/RR0gbq7v0xPJgtCcDB1As1yzn4WmDED6yBiwecJawNDcmT/s1eGYGnfGP
x05/0HOYyp3NH/1AZBKJCCYv6lHcXVqLs805wAPdPRJgmyLihY43RyybZ4EMtGzr6umkkxUZTe8V
+jSDl7tNOH6P1UUzDaQR0ZmxDr3SXFLK2B9btgYUfWAkxMsnWBMmIxYdR59aYQihxncaIhmw9hyy
dkYrH9em36Wzvm2aUN4GBPa5KAKq8okmdAviKn3gb+T/otz13GP261vSoPPeiOmFPz5QC+h4icp2
R1TI6rUV8Nzknf7ZjaQwrcYZtAhv31lMxGwQQGoMnuO7f1MZzZYICrw7Frit1zL9t5xeP6aHeSpG
RYQQ64WDlv7jd6HuC7Iz1yqij6hNj1GK4HRu3Y1kAJwOnEmV4KEmFTdsnBGteSP4TMj39R2KJ9Ip
JRe2EL1y7ZDD3pFuCHexpK+a1xaoK78JUbQ2IGeQWU5r6++5mliJDhMz7UWISL2RXzUQdWp6WrXP
Z3ZRznPYKnx4c0WforKsJnR/6dnOAaphhKMBIXARNCW9rewlBlrDS5D8vQq1rKEC7LSMlv+6vrbQ
8W11vxOcyMMZWMdvGxKLsHOgt94lQyVd0AL6oi6iLMDRv5eWb/f7R9HO0GRHoVyZh3oZWbjM4Cz3
JjfOk4bR8FMJhL6gjVvG8IoDoh4pD2DpEEhls85wNQ0Tjw/SPbWbdInLW8suR6rTGolA1o8ufibO
/7DI2XWwaiK2TMx5ZkCvUDCacXf4XFeZEyfaZrFdayhu8//6iJknMfrdfi0ASujlpoMf0UMwKoya
QaBMFPews4y42sTytO0vFq+YdC03Zz8O5Pm9gQT6BP438ys6CpjkbmH3acUYsQwWreW3dkZ0UCoH
2CVNe1YYoWcsvOs+Fzx4UuMqJZBPM4VmE45Ecfp9Z/niwHxYeTG4aPDsnb+h3pJ+m9OGFkbja7sH
8xcrpXmlsxgxT0iP58zQ5tzt+xqM2nkE0xHvsct3K5RTdeKvtU/hevdvRM42gGuJFW0gIfx3wmyI
iw7uzsRB7ibjiKTVlg0cN4GVAPcB3dHvwHnBCaPd4bgRdM04JPmes3Z6K3o5yXyL4TXdy9viXChw
6HIM8JWRHcwEd4xYXZO5HHgIu4XnYq4j9X9uYocxxyK9cN1tH3np8TOXCYYdzIAe2+NSVY7UpeG1
sztoFz9W5IqWbPeiitooLd5Y449pHHSQmWPx8W5HpOawtsmQOuFov2+qMfDLjJrlDl2Q/IkkN9SH
BTO+GVl0eGIY2IXR2e5H6Ea0O1Qkp38wD6hvIG1YfQH9+TIn8xlurx6rDUFbFkLLpuxtgnmMyyrs
7Zo4PuO4uS7zXI0+wbRCRfW+HOfdpiZ9LsDgCFYRtHj5NqZJtyqyg3EfE8w5KCAxYh5wZpHK9DLl
zFrU9WUWxPvz3XKeCbQgcFSLWyfjjNqdu8m67nI3VbIpUMyoki5muWIbSvLExgOUeFCbywnWND9s
OV3PNexbrh+guUQUeZuknipZlNVQ6fiEu3oLe5xwT1dcd7wBNyV/h37bSMwRBM0fBlG/iUZFv9G/
Q/brmSqET+D2MVELiClAJD+8jjLzXkUZeV6ejj7zlLCJQNBvq7ZPvMW+BR0fcXuM6COjhznfLskd
A3ijZgNiJj5bxkSRsIXixhEaoCNCiIjVEWYAZuveFoSCLXEcf1GHrklllV4J3ULBv+fSmS9GQlez
1i8v80Uub2YZt0/S8ObSzJ5V/jTZWPP79kVOpLcS+ZpPFzK4KmXkUwFQi+JHxb2SVvGiYqy0JL7j
zngbB6e9RQxTsu/5g7vP1YN6wlBDiS22MTCp0BGetdfV/JjpwyaK01ia4mB8i53xb9GytK/GNvij
TItPWlXUefHBe0khKWsysLgkNQDGnNmuhpZzmjEeBKXGUrnkEvEH2PDRntDDxEfYw8wyy7lhNuiW
GIL/be9rWjDx1yDWWV41nYxBebumGX418u60M4WM8lNkWEsKXYm2isIOJ52NT6dS1ZZWacFp66hg
urJIXnO5tMN9+dKL7+jJdRBg3mUS4xkTjYxlJmZRLoGWyyKO1k9qn20iWqu56r0ojNKaUhK9WGOl
9wUmXDQ0+z5n3FNHalA2P2PXwSu2Oy/TyYdLr/0a7AbhGvnlXhiDSi7xhBcpBTr1MvR/U4bWsc+g
8LyZLle+2YDhyee8hhgjOFEV2g/CClcF4p/OOn+iV8wO/9/wbfK2IilYXoPp3/DLSXbYtLfaHoc6
I4DQb1lCBR2FuKCUO9m5ZcCueoTW+zTlUFXT/wOaR7xqiBr9jKjv/60TNH5/bsfkui9hopUN7dG7
J2bkZqirhV85p8Zh7bQMWrZ4DwBEZbbOJPtHDVYuWP4F6bi5p13AyAyAZ3UQkhzZBz6u6+q21j2N
di10OBXBlTC9XFJmXP5ZK0GLmp6Ze+34X89DeOeYQkH2SeS/cm/7YdJ7R0VoiOHO6SUqBlJTJGVh
dN/j8LLB2UhpCUjMgZM3NX8/q8n8kGTiLzMltr2Tiya8rR+S8x2E+rdsy1wxP6OGenU6sDIFs6+o
Jgqyzkc/57BKfyqGIuFT8/jcjchlOLoiq8R4ezEywFzYRDM0Xj+thbq3aY2s60dsoF0iYqJus1vk
6Rjk8cMspFdBMeftfMxz6le/SNRz2IsY3zrlVC3kRffk1XeLxFkjBwq/lJsVsAgtoXqDteO91D/E
BJkQtdHxg4Rk5wn3zBSDSjv7rBenXxvhhJIanRup0Ypnat1d3WtWGIQQU7IAH2dr7VQfJjoKsySM
oji3H+CpKAPRdgmQZnZ5N2DBjHHt1DwlDautvoEBcQasZ91o/6isfJbBw7dzYfe2MQvqKLVnqvUP
6F1brtxNaaOoeJyKyo5fkR8B6H9PrYQdaM49AvS/nzx/+1nmarLPF6oYA9UYr/igZXlWRx2QnLsW
Odz50kiSjHWd1NrhFCp1HMY7Ut1vVqD762EkKB0wApXJKqcVJ9o11QO7z5TZrKrvkOG+pTlZnDCw
gUz+zR5BvrvOiJ46R+KXEMO4jsmQ1S9ujkvsbLkbL3ACFKqeQCBjsBBxx0kLZ0u/D+hss9oV6vxk
BWSzFNW4IPv0Qm8fofPAqAPmuyQ7V+/BtCUjqZPZ7nZrVYiF1RLoD+JQ5t2oEsi6483JC7eVIe/n
JbEQFEQrI83uDlTyyWUJD9RTkuBXg6SxF7svSz0LUHjERM9fyhV09ix2WowAlHFNn3IK42ieE0FG
tRjtk3LPS+Ci7mBEHMPauhfUL6DcvUKFwjUNE+62XddO1d5B3Fd61CeT/3bEt8lIKtIa/AvHmPmt
13bUQUPtre9EoHWArQyJuOUQhzdsElJR0MEvdCZQr2hCCUZSsutGo2LXhrdIl7rz1mDXiEMU0PWQ
JbRCPa/3rrTNy7jT0bi5QqY1YfCZMCx9jI43xguvFzWz1lZ0dqJw4NKvv0xujsWXGJhGykfkCdU+
73IJZQzbkry5w9q0Q9gjuM4JBZVD/7HHJokFNUInieCcuhu+KfhJyHKc9ijcu1gz6TMkHiz7oH7p
FkjAcSWFtcVKG1JIK1Ph/auxAbXAklqlqo0V2d1jenRBBtXRpXPgTMhz5Mc883ml8F/4C8eJmE+R
OKBSxhkgamzOzxe4YOEDoLJb6Tby+jUROYwG8lsf/xZCL1tRDc7iZIz/jwVulsJIpk12pTnQ4dyP
3Lm3Pjasy8lpJX5WoBisa5qfJTYu0RQUipZLhHvXU1HldzqLoYRjlsQoRiQlSk/kSly5eqgNFdJk
4DJvrmyoa0WPsLKVw9PlEA+xH7ywJSuvln2YsM1kO5JcAzWcVR70k7byehUxDRRLuYuu5bpjctDz
8WP52oK/SBtv/NmnaNBJi2eZb2hCWTVEdepXy8YZ2r7FExnRbW8KjH3sXz+0UWGJNtAJEEyxBrLl
Mxl/l3PTkYyF5pk9781wCvcrN1mBg31nQQO7mR11fDKMNmdP0ku/uA2oh47M3odGfVZoEH4zxIkt
0b9fK1kV/p4OtxPKhdYAomwB/u08VvzbeNwqeW7HDv8t/pz/8gFXuSHvu9Ff8QqpjiNNxR8TEHCv
wpd1My2LgZkmP+qaJYXqpt4Ch26DqPTjtvMaPvm3vtlmfhyX13QXzsVIDMz7YQBQt8fC/YYGXJpF
EQwKY3Gq1sK2z8OHNde5zplW12uejnXs+c/h+EA3DDqE1NV4l+MGCMBSYs0j1K86KT+4NRq6o/Ap
XlCe7QmiGh6l7cYPUgyouxjRAOETPLRWyOUVrJDpkWdmriCNJVFRJOC6wDsBQyccSEKGFvJ5P79/
e6FO09m0H3FZUJ2DCcxcpCcxcRtgIviRXgHyFv9nqcktT4LDP2aJlP/i/B884JRjk2TH/QlUo6Pu
rbs9s2KHh4SdI9yM8y7hBHoPKy31YnZc2lRGq7gpG/gFBC8hFU5hyh626IjbeDfRCiogEan0f+1A
M6bxVoEG+U+u2PcTqPGavZ5c+ZzuJ0A2Onq8cAIDGifqyONn2EGZO+dLBBTe26sG8uq/Hm4VbOUo
QsibSzot8nhaIp5eKDaTeu9Zj4wEgTqMbgC22QxbvkJMFtbFtTVuQU0sQnbCVKq9nJ9qJ5nBEbsC
g/F53oCT33ru9v0goUvML8ouDtiRvVw9/6QweWYfYOTBMbNoLFkHKQ9mEqysbIucOwviTFjM2GZJ
/hnep2otqjLldePCxdgVJhsUTntdKD2h3gniKfMfOjsxuQnrXPzf/XBia94Mqv5xaRAt4MWBZo7Q
TxSQyHbW7HgeAIWk06GgoZxgpwSkJkkydRWL1WTOrNznUzSjxIU30ZYAMp41E8S1g77KXXp86F24
jnZevdw0oK8K4u53Vgi5LOC4PV/xSt4LK3iFoxuXGZL6uHV0tqAopBQzPvpJ6X2fifnPONEOsF6G
Kld846G2r53MkmTduVBZjbpj7ViRtqtp0+iS+VCwJwCOXOx2cxqs4+F8iGSMnu4dXnoP86yAUw2g
ViLpmz9dDv+A1v60fFShE3IVTy7/2cOgUhfhvUD117cZxYKHC8TX77mlaO9tVzCCRQR1xI85j3qc
T26toq3iZuItLuG9/ZjgkjvXpYm6fTw6315xWVFd79y8t+MPai0kTDC29vN+vUZRUDllscKpg7d+
nSjTE8KOs9IadZFuhNT2UcvOMWW23aK6swN1u1EvE4pC+fOAXJfzZFln4GTMvfc1VfqCGir7Vgvv
XyGx98RDBgaTHuXEn08pAsMAa/+yDUrQEPaeKh/OjdobpPomACcJaN0PhUIe7WCz/yvOYNQ0fMLJ
AdfkcUF6vhFhM2vw7iQzSgueP0wFNpYHjeJqgxDjlIW7P4XjLnSp10BoKNxD+XcnqQ4YtxH/vRaO
Lj6DeTll7MhqThUqHg8OxRrD4+HFHTYjgTw+e4AC4VqUXIv4dzMga7EExucDrMq49LfAopdyf/9Q
UVSTPEV2OKvNU17/VNQfC1Ox+sqhzcDmsOfBrQVeDg1sxxMNUQPCYk0edOwb+hu5U7t5Ko8vwvFv
a3vN0tP08mYoNcCJXylG4we9wk30s02vsrBs8Q3AGOVNf4yNqmG3WrlZ2k6lGpQfDCprmPY+Ay4D
IYO0RXGEJwWizIZ0HqfivDP+wQ8T4u8ME0+sbv4nwemJkc4vVab4aeP3ogWZxNwK8iio20s82JNi
ZSr0dzSM9gKsmXnzIKFYiChgF1ORFrRy8j46EQJTXo9aO8HIJlNGI7+tEqXYkAoCkJvIrNGG1P7F
wkI1NMd+Nwg1lFV4ZqQv/u3KBofAO43fGq2HUXQYLhA4HaMOqERP870UcWNaW9u8rLLNdfejqKAC
LWtp31Vs1xWEBYxiR9j0ILRQurzvF+YMotg/yCXfbvHrhaF2/piFbdXm7V/uVLlI1xEySt2AxI7T
OHgLqH2yXXff0zBpf6yFOTOWxRU11nUmFDRh7zq1tGJI7PLknr8XbRGpR0/jH0kavcFoKwBZyf+M
c6PePQxJTuYiVZdulcThXdhq3JYV148dohJVrJTpxnr/RZV+PSTeEWnebxBjxqzcu7OUo65CH2ae
kxSLo2IgpbEZGIuRgaZYo76c0zw5T8CK2WrhP0pE7tTfxwDTEOsZ3Ox5tLIhbYMbxaIILe3SVaj4
8bQLFRW2KglJ5YuFoYwr1p/v6H2jzx2wi7/lzWvFPXDPfh5juzuPgyjMVOCAWKemSv4nPjLx3zX4
NOKQam4otg0Jz9dfgitUNCKc9lwM+ip8AS1gW3R5dYza0vbLcjPsk5Vi7thJw5v0117BRQu4LkCu
5exCyypr+Xy9x583Wsav4sg7nalH2DrE296621IeTfqy4o9AOoq2Nhz2SDJaYGCrvTzGZqkk2zo0
8RY37VSklJ/pr/NoYJG598yRfQTZMfYHwtLPU48Yyz0Vnp9rbS78Vr+iNGmkMXJgEnng1Ow3xAhq
8paUHO3DLmyOGjI9LytTVCQ6CQniyQ1eZ5mgpkurh8chQdQBPehwprzaJJuYAdZuAxftVoibfKEX
3h4Ud5pSwp8gZl1MU0fT0Scqyp8Ui/jogOJhr5ZgoXoSxYl+Cr6aVg9gMzifeimwL8rRPyfn6qZz
f53tN1GjnLao9BTzdcu3EBH8+DJ1sXIWyGU4crj5Xe7DPYJp/Su5iNwuUhLF9l52w2Ym/f+1uR4D
Rt/3IlzGXAyvMjxS+7PP6E98OVRTzFiucigUhzkud3vLbrlKsCM0YgOXxUlj/M0OB5PrjOwRWw8V
6gMPWxi/RFioI9G0hIjzOXN0EXtE5M3PxobxsDtkyG9jYzU2TYM8BVQcXYCH3y43Z3GsYgN95mcX
Yah7uIu+ThrHP6KXr1/NTxt6ehIBb2b4ZAEue4FoaIqZb/45brBV/XaMomyeYfxlnM7gGTn9ouzh
1OtR17jLqpTZyci7dwA5Ro89Lkw989try5tQGmeHUXoKYb5ppLjRdA6f7lu6NAaWyyo6cMUtq+EG
kRW4RIb++sEZG9oLxZkmUF5aCxkI+2jjXA8lrotyaP2uGWgfj74/aDU3DP5NE5Gcq6ZyItfSkROU
jOyh3C7wWoeLgL90eEpVFQXy3iXj8FdEghmeL/O1zk5Ahd8Tu/MV7VrRlR3u6w1nnFsovnUbyBD1
3hU3q4jkRvkeoiAxf68Pu0rt8Uok/vgdXkasWRVKSg+UCpeEtpIZerG6V/8r6SKGX+BCEjozN+B0
ZkXbFWuhKB1Q2jITdBYtn4zQ4k03PQmdMhuif0M4f30mXW3DizVjG1PG1xDpKoNN3eXyQ53TJx1Q
jYWLkNEzK2M7UrQVIqhoN6VM6UKyvAcJALBsTXOaijso0TwozzIO5N7HXT1AYWUuXCrMdlaWesQC
uEB+B/kgzhOHirtzXb+REm9KS6kNpIH6keDYTcnHnHW6zFh9I8PRCkycFEL2ScVeKaVP409w37Sl
ncd8j7BGlxDs6IpIFKKQ13hsDHtADcY3H9smiJxru8Y8q7bYRHSOe3tsXdGb4oOG4TdPjtv6Px5l
7vnCvwqh5hWHgT8Do/bbGAfaT0CeZKiOZuXFZ5SmuwNm+wQa40KLA+crShYxB8e9Qif1etQN6MHu
I11ftXhsYU7nDglipx+CeiPIs67rD5x9ZGF+EIkXgRvc8Q9Nt4PHdO/IFRlLrn3FOKLmLRqoBb+B
pBEGr10IULwfucAjx8IYe3pnI7/b/1Z6nCBD4Hn603hTubFyWjtzUwa0Ys+nGNu8CexJGXE7HnyY
+BnDZGgIn+yGi3mSylmIkfNHc2EaOx0mWc0ZyBxy9+Vudl4Ucaybnk7loaYVHg3f/PVadc6O43bb
TUdvVXXvpbuvU3hWel9uFSMjdyhQzdPrdSLLDvVRoG/lsTrFvCgmgQZ1L1VKYiPpuugfzcfGe2tc
5WZGy4un64u6vr/sRJTV9uLCNP4QBD5ScGk+WuxNUDTf4Tz59wvK9J1VreDaNqFNGZxXPg4YOfSh
tVpKnIB7CAPZOL2zr4lDJNAVR2XlXZAOh4LOrcYqViDErPIpKPvNwfkBCzLZCw89Pv7wm1X0Hzrs
565/sT0i+JbftIZXuwZqMmL8WtlUaQnxIu4BtTJ2DfmUPYOvzexRFiEVRX00SNcnCaLQZ/xCwy1v
LaOPUms2dLpr9TI0R/uJ+SN4z1CdfROssuhEZG9N19DfbWjrmDwN6Mjesp/z7/nzdlXasVBPGmic
6T6y6ur7Jep7BaSGeI7XUWuXqtVl+MSA7QZ8ZfCKIC0CWII1u8APoAnJ7mgJsLjuazw1UNqFAQVX
ctSRUvniDaHLKJV9COnbgySOJ5T/gzvgSjzayv/GsjkizfP0fnM4H1tsjaQgMYQK8MoHfCDOUlMp
wXFr8hDRqjKHpDpIeAOs4zCl6VYik4dzqfpaw0c0+j2WL5dwnqc97BmgvxKpovJio5/nE7jjhELp
wLcKx/J8qMtSKxZaBV2t7NixYMZu6ppl+jRCdAufwRCL0HEZfia/QsotAEXZ+bnL5HPvEO9mc+Tw
g/JLRecxH87oMnNExKUWAItEDXuI9aexD6Tw1FCeLWwGV+QAURngahIkuOIjTUbAlvKCUvdaJPQh
RjqJO0jXyveZsNrnMdIgQw6yJU6W5Z5MKZ1SzH9ark3tVI1pZpl6EVyx4paTnFAD65iWC2/PAq4n
unUDLSKR3awpz6DiEGeWVYu8onWzCWYF7/tjLhfThj+NwTkQWSVk3Vb4bI5hUmqmEx9gz9BGVfqA
7zMRwYWtnqrTy7VGCoPd8c7UvUaJe36pFgxXOOR2QGdTwqUqU8+BAHgeOgiWwk+BHTWvJCQEsYdw
atzuVWYly3E8qHwl00x9zXygcshyTif24AKKDTJYml0q04pe8DYluRbAzyE4HK8TNiA0u/JTkA+Z
mLBb49284xvCKjZsmyoFZMFBEbafVPCUVQC5V+a/avNixv53Jh/5va6XJ4/m/r9ktWsM+IIhqfU8
A3INVDP8iIWXS+0VlERIifSLLK6OzLNo6iF9mBIWmybBQgfCwEBf9NnJXygoxmXop+JYXEab+NSZ
/K4rlLD8LnQ8TK74RaOmTCfD+op1HaaPT8cgMhgWs4WG7QT4kCPg9fvZCjhnsvneJRMWCv8WpnJW
LM2dbytYoYaGI6aYzYYxL2y8sWu9/OnCVGFtY7x6+gRqy8lGPqRqf9iKzg+xGbE6N1k4ooFH9Nuk
iPzyHthctKtA+LsLA3haVJCOBeECDBDukmfWNAP+w+p+foql6pEfpYpHbp0vd7igGS+nVp+zQfCC
Y3U+UGRTjitZ38yitMem4tm4M6YVSn2gnuC5GcuPPpF5SETHlht9urxvXU7UFmH1KyJMNNLoTyoF
3yhvclX9RQHFajdJcaKTFW5h2EjLMyt2ARRPMnSfdN1M2ab6oTFnlsdhfVGTPvb2q27a1BakUuYl
8vqTTiBNBE5TXi3rwnaF6gYYf3UYlWOrugROKr1zBdiF5webf4esAz8/3V4oy4gCnDvXC5f2dxcC
smGD5gt+72i7wnPpFo655S9LG9KaQVoA9Jk1ilTm3rDSQHpZ7jGUeHiobFGIyFDhfV1ZtNMMt0eo
SHtJx6g3IXKTWWf0sAwLk2EVz+tw7zUUbG+x7YvpkWHfwwtSBgYRLjdKFBzjj8tmA/HJYqkG6u69
t2QSKYjtyJdX5D3r2gjw+t2fZVov3rE9ocQsnPBZNAclCmM1Mjf/Uup3UtAvqSNv5pbErj34OkQP
Qkp/r1WHh/izRnMz4WoeqAuCRVhLlf07VJi03flHVnuYL//5N7iqrxb3uZmJv3xVxvNeJJO3JzLP
swdkR3aL5L3ibvZtaqxrQqI3rBlWucRX8MzO5azXtMB6QexqJv4PjeuoZKL5SpBiBphDqhik4HTB
efGzx0OZp8oDr/069Tb3andwOy1RFjLiHoBQc0J4VFLWyxKrd4NXjq4PKO3axtMQrrBih8KDSZgN
RC8SdMy75aJpdDb+Jk2vjsrSr/4YhmnkSMddf/vY5XZ/kxjjGy1Br/d0TC9OQVopptaL68lWHnZy
Q/s8GWyhQbAqUg57LJog1mplHko/jJv3QGSbL9UQr3V4KwPWHFfJD2jjUECt4uQfaoZsQrSpg/4r
aDbJvB0IHftWKy1yb4iZd5LxGj0yNy3Mr0R/vbmiGgy8RzijhksPYoBWTrVDXTVmzfcKW0qFg0Uj
nNnUc8HQ+WWhcoil8UqUPXrUNGjCctGrdyPfPQz5r+0V/YvPI1P13MGScctkxSWj60DLBeYUZSMF
gKFUWb8asjpx17xMo06Qc1yIMHjCEqo481u1DadNdvFFj0kMbrRlgMKxYyEzedF3QBuDbOMFU8Ol
GUxWbl8tHr2ArNASDlVCiTKKdLZIpaWBv3Gv5nO+hw5x7ysX4CgbvvwMoVc5SbfrglvOGD9DZ9jS
4PO13JZ449Ge1dKJuxg5RwWodKHlENtSvi2H0YrMyJXa908RNuVLTZnOUUa9x2nWhao0mPg1t+Rk
CXVThrE3VgknIB5B1ES6+X3tA2EoL8uU+tjHNJptFUNOxhEVLSc5LXMy+Cbm9UonFEpprU6fa3yC
8nBB04HFG0XNyS+19Oi8IQNptzUwEAm41/gcZyYAl+jt3Vce9asAGjPGWcrG6AnnMd/kAW+UC9Dx
Z2V36ocgVUzsrWj09yrX4kozbf49CRZuLMKNVaQgGyXv5Tk7FegP/xX1vHNFqkRD50qGa29VviKK
rqRuZTosa5kJbzHwgt63kG7WLcZN9d7bfFYkSkBVl8FtDf9sDLjqFPnsB8iWKp9pZequxTIsQhKY
MEBldZzcCqXo0bfB6bJoskmczy/HNsjZM5GSPcmCHicxMbLZI1PeU6oShVV+PcX0LkdFIK835rsa
TEq5nFepced8uqpx9wlHObXY+yZR/NCpYyifC1HeWziqq0sOgtdIebnQqXEKZwuEVOVP82eE1HGM
9ZrZilrSmgH7AXKCLgsqtoUl87pOn7GDLEwWfRM/MLfq51FODDAiY0qBsyHJwAuUsISSD0avP/xw
8IMDJPxzSIdJzTfrDhDHewTz5AJT1RwWWQlAcswSDOQy3xJl0lv/4sCUI6rwdwEQGKLWSUtqmYGC
7hRHtkyIVTd1yK4f9oqWbrOwZ6LpJ8gaof5tedn6WSLhB6XAeimNpuzJkGcNe9PNvWsIvX7eBry4
0pPiA23oAifb50PbVnNUQP5H5zSdRzbHupqwGSJbO5v9XFHas/gRFUKuN/B3n2rFJHms/5h0HuHt
xm3UWELilTipL/x+epYYdOuhmba6g5cPnM1icU7klnI0j//2RpmG7Wizp6WDiVOeZiXiXGAoVdRN
x4nfGw/5Hvgf6VDN4POLVj4gqH9ux3N30HErjmpjF2yWSNmH6nnOFwvVaouNwYpfdzoR5dsAtM36
dgnZdBaE1+QvIm22hNP8TXgmHLj15vMZXHeIkhAd5LRRvpG9ARP8y5vF8OlK+gG8ECAc5NTidw67
0BHyUe/HlJdlQNbWfpVwEDkrMhey/ZyTxMk27ifaKHGGp1CBchxgSDPsz4QEpasgldx9Fl/fv0UW
NE3vNxoSJ7JdmtacPHHg1hAJkQZ3G/2vqlCtdkC/cB7us1pHi9uigWBLSbhLTdrMP9z0luIWSGwR
83qeI3sRUnF73kD3KznuG3MvOvlcIPMYMe4nGQszOoS913eTck1ApaMUL0LFPjczqxxhql/RThLV
J2nFc36j8Drcsxxk0ih4e3e6Z5/p7mMlBdv3Z9LL3Ra7rvHBpW1W59l2kpBESYofgp9wBnLYhhLV
yHDr9Idz3Db1iLMJPpAk/kj+voI1JA+VG4Y0pBpCEx5TmC9/bFnZSlUef1Sc1wAA7s0XOOqVn4t/
IfoyusRd2QmcTMgcQMTUtRHygds6ziaAfnoAmu0YPqQQRsb+eVOYoDXfdDy1hHcKH63nUEACxULq
e5Es9t8/LvGubYZPXB9CqTflcgkQIP20gR2MPiCiPdflNC7ZczFwFAtwlIEK7XokS5JR6YFHv2Ua
bmSqmx3gO8slUgQIC79zoUVj+dirM2xG/PBjk+BPDPH13bGx2EQFSjZB8zhFnPToKblGu6I07xNs
JY6f4cOfQ8oqxKzEgIwbeJvwxVuThqMFqFyJjjUcSpwx9LoOiaENp62eXONy0KuXgq3HiW/BfjHN
oRuH7/ZXeS+H4IgEKt+Z9sboQjt/WLDGibvQIAfR4pcGHUAbb8kJmhBjlOB4TSZZh6Q8saXv17xf
KH2GXpxmRgffkXLL/AYRllx5l0Zqg1kk9dr6+1qeQOhRuR/pG8Wreqp4/o7gJxO7JyLXHu/6tlME
Pco/hlpt/5gVvtMrJmHBG5pKH6vKGTMmA5gB0xxjMC4o1qLa4d5LRhetUurDu6wDsZpZ5KHP3UZw
408lZbwXYMPRR61SyhGe8/O8+cTiUU1nFf6iCkAAJNW36bukATTb3UPBw0tJ+J2jwpavyMiE0bfx
VnrM174OeANo16MbCUQe5YqIEJocZCXX3vgRnwWahaqn54WF3hVfHRXRmebdpRdZjQy7asg7raH9
CS22E/hy6YyXc4Nyc0R6REkcY3Z2Ovn69p2sv+0Ite7iMm6GFqsINWjTkwtO3p/Qr20bUCBgZFFt
/pZkOTjTWyKtp7+t6oURv8RW0TbCfV1Kv9abmdDsA09y+LvMJFOCygIv51i/8rT0x5l8zkWsOME0
BTNK7Ym7pCorhCYAKwBzE4TgMACdKsoAnjdRitbnHnnuRYRkjlyKD0cAmBMC/6LUNaghQwliRRcb
0HRbHz9bzmIgI7HCChWz/dCp+WtxE0/h8WYee+5/4XBSegwbUAHdwDpoeE/y/2WWp0s4t92/zpqD
7f5vxwnd2sB+1je9cEu+UBrrm/Av729Fu/4/Yc8gUL6IL2ri6r+01IXPR2cc94wQt5kmqyqVGo+H
axM9jqTyoTkvNUHlr68Tq8zTK9W1ahQWYt9oQ/xS9Xh4q+pXtOIdvqIMJrH0oAU80nkJA5VdKAn3
jjQL3csTXC3kztBBin+7WnQ8RWvhDfTxwHgERuY1Awczp8Oci4ttaNL5F6uiFqfAmFlf0X5Ati4j
ogQ71YYg/o/kJEwf2xc2Gc7OLO+/yB2YJXvSdicN4qVRpGaAj/ViZTT1UG5yHI6eeP2X4P2ZiFzE
HVMIJul1F9zDvJVj3RoA17pN2ZYyja8FuxZTNCU8wGrKGsD9WIJSDOqve3NCErvvJqGedBhvMAA5
ICIDwlOJ0yBO2itzoLzJRPWb48XL3ZFYGK37gWji5ccScjk1VqInebM0WAH5/HHc5fBt/cfSdsKE
4or87SU0KPo2+5z7PYtQT5lg1cNX8Mzw1gHPFSZymMQtXRc5yYpbXkGlRkfy1i2PEzmxPtOhh3Oj
Z7ntk+x4Y0+vHlDKzSZxx9xZwm9CiXVPnrSx/wSIG7+Igi06NvcekS5cOghItaB14jB4Pn1FCLsD
yrs13xcDalQNQJytaBdrdOONjqIQbKu9vrWRqXSjV4vNxe2TEV/2L97/CP5VhTLBJxUElBEcBv+z
33ZHp1gliS29QXKHnPAnnf9QGRGgQRbm2MTwes6aDfnK1h/A53GdAZY/L3cnsdLenGf0pmGl2T46
h4UFx8voUq/U7/FFLZ7NparapQ0pjYUjiIpcU8L7S4oGBLq8cdyeK2BJoTSBAKNZ3kRm9+JRcEZo
eAEtiBiPzP5O2uYU6psVsxAbuvNZbZRk3mszG2KwRJycRqjJ0j9pLU6TR5TI6Qkv5dnvkb1UL2LH
7+yMdGA6ttvTBTM98dji3ay5J/cqeowrSke06jyC5FWnGP794Qkop6KoR3eLcdlqM4Fdv5G+JuOT
TuZCK3LvPbFzqoFnuTQaNPP6msvqkyEER6e2ickg685G1obrJys/KbNyjdRyiQbxJ+/dtuo3DKmG
ytxL7WBk3xh4HFvgxr+MQAA4Sc/NYZxX8c9hHfznl5czSYFJJhpbR2Hb+mT06ZLFh1TFLRpkpqcj
b+7H5wsXfUTyLxMij+YuHrfit48plxMJLAJ8U8YXVQ/SMWmn24SzOl7r6Dl1Ygcfci6w1JlDdtcW
aJlL7Te7RImRiHZ/2Vs/JpIclYXwmWWWUm3pMCM955ClOeFBAd9cj6yqmYNgljDdPsNOgE7A16tS
KwlkDnJJomCuFoXoV5U+8WRKEwP9IsAAVzssXq6/rlX2asINMshFxpk4r7R+NiC+5156zzQFCRFK
7DkALzvAPi6ascTEiBYpQ6Ti6wbgp4CkAEmuMJdqeUdl1i2YEYro0UXoKt49vOjxMVJXzMnDMAYK
oeicHHgNBcO9Rrncf4/bE9Vyk57nWYgGfmqqYt4pz7HgREPCO/ZN2X1eGn2iIq9KLTHozQvqJbTx
28BV74qBGThx61PHblKA/7cOCE0hY2RtO/TsXX3AADVlfC/1FagCklgnuNW3ZLNlCR2cEo4X7Y8d
djyqCZhtR3N90wX3jh+jCzYd/Q4lD0DHaZHb8SDFDaoHntr53cf3OB8B5g7a0jaa/lryl6hzPRsI
98Th1K1HrqYaNbiRVxbKD/AX5M6JU2puEqnEx8f9+9xT7r3GHWvDsYlrewEs9nt213rUFL6sIgTV
Ea8xwGToZefnuyPS5weeKELjuyhXURUHc2iD+wX7olvfhI3y/DPmG6WetK4tzR92/hHBkKKk0QPJ
QWJaNMUcc09dKAO5bCea+lUDL/WeSwTq6/gfxQpiHLGy04Ie6Z1inU6mQaqqlCOhAjnIoEmz+efb
OOMCFQyrheKzMhwadEBH/CuHuu9xrZD4Px8T1gKUKeLOt4xdjlqrjjyoRi2GA6ZbELG6SrWANUM+
yQt7IbLrTjNviPVrk4Vi32HcMVhYuwnUASiHe3KALFwr6akjZrYksm/A8aQwXLbw7yqRh/hqlTJ7
TDs09Z598F7nCugOu7OpivcgZntUYlxWTqH0ns05dONR3eGx+Dld6Jtw14MeH78rJ+niI7wsqt/5
NM8kL+GsZy4OimWxl0yqcr1RkSZR/gaYHvgkFBg5PXDDVMh/I1Fw4gUiw5Z1ZMr/2vM4BkMs/PI/
nzPQr+B/L2k+clDLtFWmcVAtGdoswI63I39v2HUzMcefOp0QupIby2ZBJM8c2glkNlsyzft3+pJ8
FjhXolbQUAaV442bI48m27Q46F1dztCk2Tn//epOrXeqs5lgYG7MZdTuuiVsvBEeVug6/TTjjpdF
ERtLTEUwfvXEeGgkEvRDMEC/jP4hoXDOPE09q9DDi3TAQNatXUKljCHU+Y/tDup+wMde4+AsMTkB
KFYbVWd+tQ7YlHrLPxCFvyOC0VCzuiojiEzUWLVicM1U+InLb6Y75d6c8LkZ7x2ep7dS5y5h1ZFa
+2H7UWC/Uicn3QjqvApj4KQzNxmcwBS6GyEMKuc7s3kZXRQDwlDSDckguc+2KkUtDO6fBa222rft
QI7fnME1GVCT0dmnMTxyuKB5ynweorCwnXavxOnLOyV2zeaGRlOXfmo2kAcBtF+vl2Pj9nhLfyzy
qdtycQymNl4GoAoXkvzkk9yU+6xxnmwStiLyn7lbtj+av4Vu1GCSkG3AGkEWPxgP7m7tzJk607Hd
30s+52FhXa/70kebh16F0bt9BrwpW+fQiIh87qrt7OvpjY9mPlblV5rLl8T4iKhvPpSlv5UHrKxh
d0feCKPjH6VKjrlW/pBzREoH0rDoSva4YdhSnrFavpe5Fl2rCJ5qJ7DdRwrg1QTop1p5+Bn4ikxP
U9rpt6saFiC7mNJ11ZpT6U8yzIfcg/+ElMI5DXo7fKD4Qas3xiY0wkuvY+LSGN8cQ0OKGMZz4ju/
GEPrFYQcVTDrRI9cfLmbFW2gRbQXI4281YR+rF8wRCb0wDJj53hFA4W7UEBk1yXiXlXyPBzGBf1l
jL0x6g9CRnljA75cXhFhuzCV3/hm7O0qsQeMGxYJJizGU8ZnKFFtrl6JOHX0vZPf3DhYLvh8yOWO
0Fs+MQ1d4kQYCK2OZ2+HTW8fOyXmo2zzX/JJU3h6XpOmpFgkmzq+nrQxqfFmZibu8O4fTks6uCdT
JPiTKXjEnDKFKG772n2CWD9Zyw6dEDJhkOufUkttNqt9wefwQCCuX/8VGbSbviw2s8BAmmfXDncZ
by0tHNFfSO8ulRSHUMUxfgpORz2Gtym9eImIUVoilxqTHe2e0gVvBdMr2sh5fMnKky7M7t7gOSHL
xQdVt/9pt0ybhHg1/4lrywkGfwNZKaTG+LiZoJtOX0W9ES0iYfVWmvwAwiuB2dA9EcBnhBWZ3pv8
qKr1MzhcHHCtaEK+ksGcG9JULKs6JaWbD7+iin7pYvVaHSCBXzXYf0iWiLhaQAtEtZXsKe3MjXcb
DBTuaWOF0dTJOBIMznEUwFSgQwRvtY4RGLNkdLdzkg6mC2p/tJ3MmnR+x6axIBb7+nEqKRr9+KlM
Waw35+K8UWNzV8Ku0avhVcwdGyScwLHijyS6NmSX4315WR3vYjHJu1vQtBOBcCNFan5SC7VV62i/
PUWcFKIHv12Tutg8xXAbQurGLMsByIQ6IxRyUg35zI/cTxLRUe4leHhdkYawb6izU/0QQ8NNMgMu
/3TvVp+JrgiWR5uV4R9Tfaba1S+0ntUEZnILyGwB1NZWHhv+HtRmUxj1Z15s4cEBctg+WjgzwRnV
9Bu/oOdfuoihNolvzKPfjpzCaTq+Pu2/j7YKqHvc0Q0mhPFQ7HRwnE4C64BzW4hvG49K1WZAuKPf
9goPKCt4BREgbufiTvUJWevvQyXvGM2tPg0509qPnxz0PvDUw+j1/PcJxw5ulVuL8JV9VGSZhFQu
uEXKA5uj00vJlWqJZ2j9g8/d6rns7SY6OGj3lC2MlnnF8CoE1JvRIzBTapL9GqCyZk2uW5Sj7PIa
djZAAECHQqs18f9WUgb6Av1xTOWbpRDV1r1DYgW5ptbZGDoTsgxMby1aKOYn5+XIv5od2n18bAbm
CdtBE3qGZZ43kkyUAePTcukBmF/kvO6IUz+KDaVejs+tE21+6GFW9emdXU2+OeV5SpunN4B6Pnbh
59vIhWQM0DNiJj+9vzgE1nEFmLE8N6vSh6++osCHOOEqlmH78CZ+pIisruj2ckRKFa0EwuS8w/91
3elEgUc++pinVl+IfFW1r2liz69H7RkRhCcn9T+PQAAIYegjo0kGPpT5X9eosAj3UPBMPa0SXm4c
s0rNt96Hj/kKaZpaWPoUNCFLc1vUz2O++8zzPkiEOU+/NtFNXTmCo3l6V6oayPIR0K7Ls0apRPTt
kwM3BhTLOpbLtpDu0kxAH+2fxZmNQEKcyO7wex/P1+FNJLau5lyTDil/3ZtlTsVRN17KdyFr+mab
tDZ0win8og/WEogUFOynzb7cVSpclzVsHR68G7iZE7MHA2MinQiBEd6OM/pqQI3T+PHZyYyxE10i
VeaNdCfNeRoQBHmA0bwth4AyanoB2nB94KhxgKOZnCDfeXjKnR1jGigiqYmtlqHq0pLcKxSWD0Cx
LHgswgQO8fqkCgowq32hpDC/HdYlC3dX/8Im1N1AfhEzrCGwf2Sas+fbKPcGOSLWov/Hl/5Nbczj
xyxhJxFvwk8PU7fvHvr9HgRVQZsQZSISNk/sW1TEGjgiNLC6AsePK6cnG6cF329z3EJchuq8Lvyo
0bnwU+02wJjxogdQNufBwlNR4zf++M4z+CwnC1YU7igdUG8ZwPSigSxhfJ/uNz8KTiy9pkc8Y4OA
m5Mhg9Uwek0p6/udeM9EMATD/jzPZ2jt+5yMryrHdOHiSVYItXBVcOO858HSSo3Pwq6iMeJZdc8G
nohauH+N8LJBSkIlJ0rIOM2GdHTHwCof8UXrobCepGt4BtSlmNpRjiSjK3IiVGPkM58FnaiL7Iv4
uL2VmtsFhNhvldcN4cjQ+XOb0K0slBbgK81jP/hflfZtjil19v5hup0oJNv54RCScONvlzJNRua5
Fd7DIDZBPW4dZ1Dph8WiqkeL40sXWDg3HTOlQ+NRhhKAlOm/jaXffIUTFUUcPlaSPoF26GBZScUd
XmfGN3Udo97kRhKiICTjDRooiDZmH41jqK/abPwQzomobRMbOWKaWumbvlUPSM3e7LXbtkA8E4OI
l33UYBHcBZaUYSvllO/6vPLG2NQHDBOco/YndWck68B9aHMNTren2hBT3w0KNPRAj1JBc/j8KHq2
Q61DwyfWz9lwhSKrjHtY2jYqpaIJ9b505L5bl5u78Pmr96lRX6g3qYkjC5I6ZupRdBMDDv3O3q5z
qegxH25gERSJ7OykOYtbHZ/kEWhDsqjaE9Mx9vn59CQ4NQ4PABHUyI1YGMTPq04zWLDNyb3GgBYk
k9LG5JwfCM/rJCpLN8DOp5v7xOjW/K7EPpTn0aEaoItRNLmKEoNEQ2cT79I8I9o5Fvou3+1O7Dyw
PQjKs2H+aKt7OAt4tyfFWzp6Ju2nbqgRWHsIaolMmCfGPEeNx3MuWcG3zcdw+WQTQ4movMYzCUoV
IckCeO+rqEFC0KEajDA9JnW7vM/YcGWbNsy4Jd50tw06CLVzp9VQYHoZwwvfKn3UDsBbOZoJDoAt
yXc+YW6J+Cm192VQ+JYcGTCWURei++hEbLabIdef4rpPcdM3d1vxLaul3Dls1KxdwtYlG8TGjNh4
hYF5yfVRodnLv47GYaonckOeBkdYFfj+QqxtMwKDsPdDwV8kUaa2tJHv9YBUewuWWSy9ZI1R1r0c
vwaljmfzMYAgBPEtbxwGSthJVJ0TQLC1n45rU/b8LUQk+LGWBGqK73M3xVcPYhXjgUubu+b0kvXd
ZC0J5MYFOXPXJdJ9bjN+QmdyqzLxBrCDH7Ms0V8LevCBRWEomzCYamTSB0bzUlDcH1erlsFFKqN8
/60v0rdMfntDnoYZSgwwSrQMHKlpcUDdbJZ8CXYyOpwB4JwxVlpICUa77t7tD10hUcibWWJs7F4w
AeHqoTxOCK238+HdIhqk5nQZh1YJfZA2CqAnujKEemGvoUQkkzIvxZPgtzvHo9ho0+BaQzjYuSeu
puOufuzV9XQUvMpiPj+RBgH66+WUgMZKvWZQUDxnJw/Svdf9SH0v9BlOJxft2NQCUUjdZAH/eIU5
FYQbfXMGQaep+CTel2K3GcHyiw75UjjzK/Knm5CUGPTWxQ+2QuMgW8N0NMCNS/6Fwad3obm7p5Zs
LzTOEJApIgIlG+mQW+hZJp1XXl59+1uauxdn6Lekro3lNyMxzTV8qWrngpMcrmGnv4C22WVrx+OT
SdxRScTjimYlrm4ag/SFkqA3eni9Ex+yqgNXEsi+iraCAaNdGKw3uYDvwXSJqiLrOk1iX8C8MS88
yjwgXAL0zDRpcWzjxfjOwIBfvvQ9AOoYW8epG4roSS4qS1pjpdoq6HItuo8EQCn6Md0iH5YNzjiM
npx2uSmJkH7ZIDDbDjOfaa57WVrkJ+eKfroxJq7VVd0WPTYisYAt3wa4VYYTPK+tHHsxNmRITkQl
wkSTDHPyomirLJQrRE223328lmhaEDMRSf6tKhmPwNMWhnqyl8TTjYqkEG54uccSl26Ag4m+3WQv
syi1Tjzlwx71RvNBFC41WgjHSPV3X1SJK1CbvBl/VP8TzWnJUjVyTK4PEyWNNXveTHLrD3zLrKXH
rF9ueCye5tp/Vw/hu8TiMbHTEF0rWk1+wLkWCIA0bt08Hn9G4h7dDPnlYdfKWvCRZ7G+c7XfnIqq
1JwjcVMLiBb8vJmWR/rWqG50isVnMfrfs8R9VgDj2ntioNo8J/+UyMPMLm+4hGeryWPHln7KI6A4
Q6BLElrKeKifdOXckDs24n8pHXhlaqhGcFi4zqgWdDPgFi/kqV0aRbDkJ1PGKOytYsUo4TtATsD3
UY9xoAPTdbMfU5I40GGBAttW18+ydCH0HIeCrc9iIKWTtjTvIm5oJJ4PEYb1NxUf9kU2Dvu9oRS8
WSQ3RT/D0Mo8kyokoe+V5wzHvxpZRsn8Sjilyx+IiRqslnrZivBUEFn0bETt64saE5JYbnEbXE7W
h1J7bgMAuXkRExsgD+5IL7IYjGiEk2ckHA4OEC4NVruWC+2UzV55qiJxYRdxY5ZhB7CmHvBvJFi3
pQVLELfc7/FnuYCB2K4RxiMx91y85WFku+9ymfp9OSCNfgJ/GK+iWwQDci1Yo9xI53Cb0Fc1wat8
XNEDHmbpgqVsV7qChcDlb2vGTq5A+vH8iqM/xH5jqy4uBwWw9lDM1i2XNVtIjrBGWPLtvqzU2B89
4QqpiUUPHDVJsUODIxzDy+/8yYp1xUc3mXdEEpffQa5HQqg8rSPYg/rICxRqF/uqSk8SrumftKDG
RUx35qSrrI83a7dKXNG0sMkBit8XOCplWttQ+BowUnhFxNII/fCOBomOgBNGTZ09ecbtBQDQSYgw
kS31nnWk/MU6/ex0nKqWHbRMoUMxDMsh+XEgZv7fZQh31xJC+fu8/6ClcZlJOnP3ui8GyuRr92i5
ewPItaJKCw3o0PN19FSgsBzPM7/fI/pBSyjRGp4IMqCM44zIopeSipSRNXdF1DdF11/zlejmjWg0
1j4q85A7A/+DsMt9peo34ljea9HABFpZYlcngbd87XIL8n0MWTLUdSVqoaHTzkpC/JBtiPHOmLq1
Z6qZ4mhiAsYKf1nq8PDUtO+ryp9Q99Hc4ul0q4YQPKgFxJMJ1GzdNBo5pqXcgcz/kQjc0SU7HRYX
Hroq8lxNoiu4jGhUaUErUh/6FT4VeDNRSC19+zTm8CBmvILBgD8ghGVK9g/XJoO26VrsZBYsHuHx
nBmdt4zo04KhJqFFJ2Kxqx/t91u3k4N+8BZttk2QZnVmnaGRHjlrpmtDbyJcowqhkDQu+D2cVcIh
0uc18ocr6GqrJmO1e1IqbLFDl5S/AyS8OOC+lCR8Vaajtlad2kpVPJqCx/LJzNcloe/xxwR+Skwo
Y8X9IT5QPIB14vNnnMAD2U2oIkehrayFuRxycXZTJaPN9ta8SvFq0AGJ53vHhqP0/wgtgxDpfKq4
0jhl4/8/zCoNc2z6a+LMOFPFeUjruAe35Pbpjr2/DCYUB0HBZ/RBdvKESRl+AYrvQ7QUY2lPWxWt
SZ2KD7e0bx5DHJFqeyqYnz8pMxwmkue5prpN7I4M4GrerMm+L2q1AD6DVsksJMKvIYU8EXKdsVfN
4/2aXr+FLR0pDTK3vyErBOh9MEdPcJlUJgIUtrTpc55/62yp3dy41BsygUEBUJ1XpGVLY0dEp+OF
d4sVsJSKEMSxRNGwYJEmqXcVZ7fK8S/g4WqwXFv12qSwq90Gh0Uc9450JWP11u6io1znca/copZu
byQ6wkMimZfM5qhn81EttmdzEbTZn2GWPDCAo3CCiSwRfPGLWYQIH/j5LL9f3ZJ4B7qT1y9CoYLG
qzuoWgWTJDY5rszbQAZAyLFIbIGIMdiSBT8wZ/4bQyJCHgo9anUTaSsgEQzc4HDbHuix7/Dw3X/3
nfoN5R3wu1FWcCa9F4i9ki0S1qziimCUc3v1lVR1Z5YSSPwxTdtFBANyuvplz/ar2c0DJgd/sv31
+EqCdvzt+TQ//zbzu76nk+0D2UyNuDyKv2l0BHfl4B7AtRW9Cy+XAJYsSZTu3MoO5Esx06E/Y5AT
WtL11JoIdBPwlRd5dA3ZRm6d5bzYG6TPCUSMOtUQAVOZgh8sHfpBYfESxjEODPQ+zW9oqwLPPqub
alWFnnsoP82j4Ex9Ycx4zfUR8q/PK2ANSktUSw9/Vwx2Ha6iKMRhOwPpbhOuYnRwTpmvaRIzgOn+
DF8BeivCekJO62LoMzLrN8SbhGzbGhHZhvVkp0B4ivsPmFXtc0mkT/xY7pin0WmWg1nuDlKfrW/H
gfLBjaxHlCfMf6rVp7R3V8N5e/ymr7qZjL0JLoz8jzgw0du6UhNcHz850ZBl08CS3bCTzazfwSPm
72BaHqxk98UnqSQKahTb37x+wX+IHBuiSwTsFgzvUZRcG4kMEIGAaOajeU8FXqw0hg06LBR35KYb
oRdmUZxS+dZ8DUre55WxHLMdJBCnkxMnsM0gQD+qZub3+RYK46Y84pinddY/0fu91RgrqP2J8gZZ
iOLqtUiCNt8q3IIaoh/BZwkNnX+KKIFbEwSocfq0tkTV73iaaDaso67WayuimPp2w/bl3bCRKACm
HS0yYo2yul2YHI0t8iMewJFrHINhV/D/jUUGoW9hgLQ0s+QcKO4yVh9S2mllzlYj6eYXFAysYhc/
XRG/MNn3DR9cpLUKPzgPQ1Uej1FYkzksnbmDnHX63TL42wDY1s3bORENBb5m9xt3yQwjLU7SqIns
vGg+e6cnwtZ1lT1VGkgeDqjOcXrfnGQsEj1OxP8VHsab0nzaFYzySzoeZoSb61AKJQ09WQgLlb9Z
UYrAo7Pr+2ay3EyVct50Q6Ycadg0J9RE1t/t9+keV01Hk9eOK7RAlfQYNZ+a2msPcuekpCldJgle
c9LKA9KLCglsOn5DtkvsTiDU/6t2r85/kGFAKY/YguZhPQSMgdEsyYo53hea/7u9Lg/Vr/kbDMeQ
8Js17Mkg676vYC/DbfRTkdpWt0IX5ozWDdemdueE7HqpGIDKXJEsx7Qj2OcOdtmnKs/OLIxdARKv
GCTpKk9i8Nhv+ZG6VLOw7qzphsfu40slPVgBPoYCBRteJjQuRDaW3Aiq/9aCOs4Lf9SRrYPharGP
Rc2JpDjVEKJKpoyYTzomJvvjmyiOGQLpvHsr1JXLp7xplH4XHprHlimPgWBIkuiGRmfiJoowdeKd
8FfxmdoluRK5CNaEM2SrDewdCeC4wVxSJ6q1pk5rQ3doc6C11EAa4AuBvuKbkacyMvXQW/s+Ml1L
XhNc0Q0PtQ7WM07nBusNOFQYSdXUA+0RyhIAStj30ce3VtWkPrun6gGiSJp49ZddDx//x4f9Vwrm
nw0fpSIGNP3u2QkDxnU+mrtQ6gDDwgl/rEUp5QeopSxtHOQC5569X8iTaZPWWgkSwlE9HEnjAsx7
eefTFb9g7oTSxZXFD3M2vbVMteNpzQaLDL1FdZGuNp8DNndH786x0gL/7EZr9K7NXsjcEQSTpJQQ
DhB0vhq/Z32zBwSri9Wgu/KqkIrPgVmDIYGtdL9rthMpW08pJSZ23lZ3CltjLgM6YloR3RyKiGxY
FHqQYcArQ14NxkVakjbYaizSVmsFPSYdruo8Q2wgroFhVnFzR+8BPNbbiS2nJZ2cLsPvbEbvhQm6
1V4uNkDcemN15+xlgRbzigeaqy8bjWU6KkYBcUjEy3Z8P10bzL9xVmW9OXr2OAgTVzMEFkytiK8m
ahM7X47ud60S6KgR2NSz2R8X30WsQUWF9Hewh4QJ/ADo9/8sIq7MHYK5ztpODzjB8WIjtaMFcsIJ
sRRhFQU0w7eWaX2bLmoWeRVCnPa2+NK8vaR51K0yOehdhS1zJfclsmICFlcP8X38wIX9gpjM/LPz
08mUss7qrv0ZDG9BgIl9kmDXrodqscweq6E3wklyo/D/tb1pjPQzVGxKH6OtJyOKn3+/OY2mgOR9
tuvGebCqHhz5gv8oU0zN/2c0BzHsYHSNebPJR0N7itleOAXMPpygiLPccWL4L8LnTwmM13r+UUNA
OK/APd7MKwWYAck4XTuLZZTZtvuKTwf3CPgPHFwT2pZHNaLk+DvUAeQJkwycgOUZjGggSJdSgQQC
M2X1jpjycj7Rbant58vu7lx4DThfcp2pU+G/VG0pxaWsSzOMdWTiV95Xy8RiDitPNh8+RTUaHKDe
FYIGJCOCP9u74Hv8HMnfuNbcMm5d2ULkF+Xv2EzUgT25tI0Zch7icyNlIlwZCG5CQ9Ua2V4tM1+M
bgJdJJJctADiszTLecQtQgnFX5jvo5kabybv6ECHpKG6I7KTe1sH74xD8FbFYk0+UGtuayqNRO3x
fkw5G5DUsc8jflneQ/mfJWcfy/Ucsc+gmoDn/2tYgjgiNHTfaAgqdKDh3MhUyPxTwjeTQ1RPN9dB
FYo5x8djZJCEWY/EogevKnK0Fgx4utAXlyIzrm1woDh637O27RDJcMJqmbG68XfDOVgnGYkfANOi
F+zzjuMeU4UPzThESyaC/nLlbhgac2BQFe3PEjFazcuYV9abhdl66p88ltH8OJ3WX2oLxqqO95dL
TuAiSuMppEscQIYYFSmpY5m7YJayirtKWq03IJosridkpNm92tBpAtgAvML6JJhoQ8TcnLYPaLzW
UiygqGfugQTh8wk+8CgarILZVQZsOJfGor8fu6yAR7BCoRS8aAqzXs7U9aNfb8fdzjEfn0S9xVBI
PVJaqRO9OC0yfPYAXZrxF3EsE53zvFZsDtvwAKDcZ0pJMdws69PZhNMPZvyE20HeDWNfWlDGrn8Q
NDeiPt6YBVxDSKK2RRiOfn2pJK4aURz+GrAJTL8eE+/5wLXRQm/0PVyaRbaF+15GD3MnnRoDPjE7
q4vFSFA9O8aNGB9ZVvoPE6dsBKXAihsyzPLW1bZzfmmk4bVukvkD0z0GqgKxTpHh3oL8Bu56ZPtr
g7B98qBYOCJ2xgtUXW3rsx5WoUbGK2L+cBA6CKylIrqum2uhxDbc//oBuAAwX/DYNOix6G9skXNk
/aIofAlEwYzwOwUpWBdXn0d0SGkODbNsqAC69/qsA29fkPvIIyfZKQTmaEkHi8a55MtdNXNueDvs
X230ubg/J/ko/NnFTVe1ZLkajl7P5d98UHY19FMyI2dcUeQKl+v6YcnxvluJ5MMms0uv1Wp1/n4/
Iz+dNj0w2TSyHwRKLkZKj6voYkXuudVovJ/wHnNHnzeTYZN4vtt5rgKESNJwR+ZR7E6oCtoUIVoW
GD8lUuzgc0pBvIn8sbz2yPRq4g3wn3ZNNX+NYQw9WD8nEhAZ7tP+1vAtVndXfMTxFVP7EKojBALO
17JZplOkM8usIcJyjlVOfXC9yk991Z13+lVZ9lQQFzz1DULOCjVyF2hThypPX7PSKAtsPMKs72/G
Ksiw1oLhGZJiYUMtIUwFyCfFzEobWRuAVluuuJB2xxpLZfMHFNtzdbuK8j8DPtAqTR8s+78BnDQH
gO675xoNeTxANPVAMX3+K4N517k5Kps7JJVqzIoy1GXSbJoiEyFKg3WZ0DuqmorzyUdGTqa/AsXc
it4KK7V5hSKava6vp4pL8eF+3S9npwJBz4tJe3m5ajlwc1X3iSceUSC8tlktA5dNL1LuLM/rEZ8W
hOwS50j/HGqGrD1ghOQ1r4bF39UpiePjjmG6iF0See81YEuKYGhSQi0pSlNOQ0VaJrPCybzpaYfZ
rlvLnjHBrb+bgj9STXhB4oXK+CcolmK2sG8EpL+qg8oZCr0MLZNwlB7qltxOgm/sanS4DM4Cqan0
8ceMjgX2E/3kz79T0CIw1FoPT2yKrZ9QtBIUYgD1bHPda9KjEww1iAuZOxtAVwOsyiez17YUVMf+
pATHSHpxf/zXcZcEoCbHt2zLOboQ+GmYFXxKxqumBhMBzLY2QW9cEf8d/gAqv4of11PRqrxMmfDQ
IbMsNQJMMyqWOmo5jLMlIb1xppWvcDOOQJbecyJM18cs2ogVujXVy1lm7/lC1eZGtV7bZhuVWYdz
YK7nPClKlITSXrbNTVL/H3QEMVGcjlSZHdr4fZ3BdhWk36A7ENz2vMQqK3BpyagVUVk7ndPpFtWA
4lE1IDSLAK3ZJ5FUr/5c3pQH6m/HST8ul61R2LiIQjysjMqnZQPx8i7Wv7z78FgCvdlKRBh/vGIL
YOHWPYtUJaIQNPfo2y4ie59cQCG+wqPmuZ++cyRbxpDxAxPCVHWjF7NGN7qgxZMRxS9ZJalLr+jB
8/KLDCsIBvfhIlwevp5nrMslcg2NTNA00dANf4yfg9V37Mb0Pa/1xqFRt5H8F/vP3WWMyOQnVvvE
cqny/2Ngx6iPXe0vkHwxW04mB7CAQknPQJl5BfS4uMrEla1IW6bYXKsWSbUKX25S537evjLT2ZnD
XjazQiV8oBkb80RL09bzsNWndoCeUt1BFRmVXC63TjwXhbN/bMI489e26Hhe8cxVSHERfNUlvzdq
NBudzFtf3Fa4ZAmswHrDsvNGnTmc5IHaCdmr5a+8tVsclPNAwufZ1uzWpc6UEUZZWHT+KFIZTlDY
4V6Ly83RmjN5l8Z2Ce+S+qMtdP5UZS9WhYgyBEpZnxm9ZAJ5AF8xr8jPvCQ2rs9osnoBnQ/pKdFq
jrdYz97VbbppJaz25RTXLtPUFgmWDb68zsCaC1tmG984dYNPHFCmX9bcRWmvBqcNxSBSqcpi+z4O
JU4RtTAnizCAGveLUBVD7Y0lxSC3nurgWhxWtIzOdxLR4/6AKoWTtSHRI8xpaSeEb1oNbT5Ck/Q/
izuOdM9o1HmkL2wMTUXkM00tuXD/XrUI+655moK6GtXDHG0Y3dNuIrmYM9nFxQMZ95/QXJ6D/JNg
h8ZWrhXgjoiu6E97qc/VADKhOBNJg5kpC+vndS7gEy57IAiTIpT+/THUfjBkPhRsQEoFGqbI+ZyX
GlgomJU7ggtJt1yFWscqWS8DQcvH0zHTqzv/7baVLTvf0euljfkgJblIwJn1iH6ilufnIyMQdD+6
jBaPvxchhBuHGeukqFEs2pcgEQZ5mUPdkhxQATce2e1pXpCEKB4G5/OFejGieDsFFapEcH4ExEC1
kBUvWJE7pZPPUwcd97D766e0jedzEVvtGsPQciUzDtSRbUxnVU0BWVwj8Mw95J2j3IcmUBd+Uig7
pNyy0ng1/CrEg1j7oee2/68Ccwt2Mtn9iT9QEVGvUDmpibuctjpK4EuiQ/UVdDUCF+4Jk7RfpB5E
J5EcwZ/ApgnJvIDkMd8eA7sedJMC2OTKZxC6rgKkK32vWt4UMKRDVk6ve714/+NZxT33ZQNUIFk2
pbwBY8kXUh0IBiUw9QJoGhOGxjOR+uSkgz2q9Uhor49Am+jD2GLuSSCBxGQuWYtWZAC8G8WlpENU
M/U6+qloi7hjzkOGh4pFOzWRF+zzTCem3bTav+1GqdKJkkzdIzB4attGbfkYPpX7yK/WdnoRZxHh
8ftCGR9GPFRN+IJkbAiREynv1/43dn6ho5JGIrfshu5zhi78wbdqpg0XYPfuZXNqtoBtC6pvZfm2
ngzB661XR9KQDPOlLs3JNixpcdO5vP/CIrbTKAGwa1JTAsQkHG5YKS3tpRo6u3eKvl0WWDum1Z/H
L4y4mE2bRpL5xRHSRL7skfQyaiz2qQEjpbfeFyRLngIJc3Px1zQIFmqqAZTp2cl97YOCTLygSyMU
TiIR7h0cC+QR+oD/YA8Bil0nvQxvp2KglpXXjwDZk5fXu4wSIf8UX5a9vEGE/BhGg8JxoGFd5PVd
5d8f6gUhmGI47NwegcOFNmTZCeoTzLqSptoxLTmln+AcivOEp/dTCMtvgv8AuAPjbdjgWrcyaWS3
nyIoLbdZVy+8miod0h/K+FnAaYQaXcvLeAKbJXJiAA7tktumIg8ABT4PXIUuT1LGd/EZ45IJK0FU
SJYCM8GajcIkRse7CI7JQDSDX3odQTlnnDFYoLyGT3xDMHvnIPHBgiQ0LmMJzl30RGA9OF2r8ZgZ
EBLGd6OrNjAHa0ZsLTGjBcLpv50KqtK+glxuXxDabUXi9lGjcGMrwvqtIruik9UDOmD4VWxIvNaL
JbX9lnS0xiQdKbX2GMD387Ka0r6GXGfcCZcDpIO5Bkw6mATUu7gKbG4M5hUCqV5bogtcxhniUQLH
ol/Gw3xuWVYHQMG8xUDjIX11yLhk/7lREhkB/+xQNpf+s+/I/46UfVf3Es4lGavxldQOBUcZK8J8
6jFLTICNcuxu4hMt8CidK8FDplPDQ1hC4wFVs0B/vcNE+Htuh2PdDPbvLLQYqZplFW6rAK5hYPDs
TjhXWCMflBV8paMs/4ggYDoHBbz3uPl6wBNOD6aq/kwbb1DPZRAHAJnpcWjxVwsqiv3jx98uiYK8
McshwrzgBrHVPD9LAAPTWmiYHU+dOeFXFEqIXPYN1wHEOAj3PBzi9diOMr4o8i8tdN8gzomteFLo
tP9C5vC+RFDFL2f9ADiQrCpNvjiph9m+gGIlFuBojG4YlndNQsZkA7ZJhHi2WVdG+2lpXQLgK5Af
ubJbFb+X6MTZHb4ASuEzXQkeRRLcydnWuy7qYcVw5P2hJbyvGFUVtQhWjaE0J7GpsZOrUGCsSaIa
B5Hn2OwV5qCyADVt8L+KyAhpp5wPdhSNHH4H82oKRxOvG2zIDCZO0WSKm1MewiD3t0qGbSzy+In/
py11r+cRgcYEuzy7xHwB1qHAQiHwHxsABTOmnZGDCXsxQpbSm1BBKHeJ8d1KsE+z52n1OqRwwInd
bmAS50wA+sz6k+4E5YaPqTIXtTMt5Tsw5VJDURGMu0t75Y0ewLLHreSuX7vjIsv2IGGGI3ZCb80k
LgB6q1O/oXwtVOfyaSJ2DKj4LAKzFbXp9yw+uAHvS9MlBtnjk4xuoEcjpaz5WHzs1fJFfeChI+q8
iDpxh1U6vPpJGpIKLO4DoY4iKlriWCX1Zah1CM6bfxdNgdYkBRwDBrD+yKReDmGhV5qVB5bY9pSD
LrvgiDia12Ds9mmq92cWiBXxjboaADfNTwjMes+dSn1YbKzXWpoJHV9ofjXEv7HOMwwY9Hn1sIPG
G3emzkQDQE7meDBvki4ClEnvU/ef9/DD8PA1xY30ErLAwaJKa9OM0/d7aLR2GDDqjtDJBEyGPSCk
omxkRvpweeWSBshqPjFZTIDYeea/85OuNkvQQGeSydVbFymVP6PN4AyLmTq8bm+iTnLkS3WRKSne
i50FV3YyzCaDRLLTQj1FnyymynkiZba3E3TqnWGGPHvseAe9vHjiBLyF5s7GpTz23iaqDQzc+LIw
jx6628FqFMw979GnOGTzc0KbM0USWLA0iN+w+URj0C8/a4MkiPG9h/1htUvq72TQ7F2FHJEMvL+Y
KeqMst6Pv8qqyOooRV4UGaqvCLSwO/ZHhrwZeL+YsBSPXGWTLt6oDt5HiyrzAY1wwhZP4WosSKtt
XwVP8qAZSb1ZeN91vKb9ZoGnoFeRf+IgSlFW3n2hpVFJwtjS7+rSV4z/UrlZTPFN20us+zH0V+K2
J29WzHPOrhN0cNvpr6DL3AhgeaV8oRd/XPFX+KEIZBvPFKO0Rpqo70PUt6AXeoan6foW9dwmoJxA
Z0HKj40dF0zVZURJZL+8AeoYuXVFtl+1hHAkoeAuTMbk/qqnuikgDcCT+Ub2xZZaoJnJWOMIohCU
RUUQA8k72v2gzMCsSpWHCTD7Rqisg26oBRr+l+kyCPl+9UMTk79zIcIegGdXgCJdwamnruc8RDV7
Yr/oEVuqDC2KXybjlYdbzl85iF6WIsTYLTVlaVvOzXEKZIanhJEz9PWYFHeyv5TfQAxg4YfG34BB
q4JeFyFfDuuSe1F0JK9zQKHfEN4UmCf7MXzRvZLO8xtJHwyi8h1G20meEdSMQ5tiB6PecMnETXuj
vIgiUtJ/2oZ4UiFbJ+uW8utX8KN7YhG4KcBO1B3yH67jQOpA/EzK5oKAaoUJExYQj5wLoF+nIoxH
IrJPxGz7gVg0kedzTCitaPc4hiAQwgdKwz2utmm0HAgB1t3W0pIL7RFegUyJBJ76Af4F3abO6uVx
9kIiqtVkx8b+zwXQnkTugR3uzu1aKXC3P45hu3qrRS+0W44G+EfVbdvGU4AJ9WVcqifIgr77+NQu
4+CZwFzN0OG+gJ2mCxfoxSrGArqGbmz2Y8o7LE6i7e/ES0Ac96F/kX+/ReOI0q/r68voixy8Ebmc
yl7flvSxdlJgarLBzff+EE1tKgLUM7aqEDs3BBGjY9sgSroIllwAt/ov/ujQFWHaJrdycWXorAPx
Yb51XGYB6qxnGZNT9sceR2qHj3F6rWdD4BX6r0/ZwSYclXxsfN/beAmA//YSuklnoooUmCV6r1G5
ImI2Rtt7yeA/CZyz8S/NqWLV2m+xB6J2i2QrrI9FYYzdjyrxvkgPLdGOKn8aQcA4AT8iX9RQOxXg
W4IxqBosNzrU26A1vuzABOSd1ZJpbFVIY25kDgVQdJTTajClHUTTNr1Hr+ULzxIM98AbXVIYsm2F
AoFa1+9AvjTn5KVF4gKXyJClSY1+XRFyqGf1t+20V0UmMuYIxOpCOs6yBGSE/ULrfxZGIGQSeor1
leuMs1Z6A/yOBDMjod98vfEpzy3a7FlUROuzFPcCy99VT92xoub91pkbNYVTPvSkx+0XJ3724Juh
gqb9ozN1pCeFXfc1jZjmBIwPLBrWver0nbUexK89fV77qs99/aMq1Lc94A+VhF0Jpx7yegvVoLmn
kX1oOOP9zYIG/L5ZBCdu3Hit0V/qeyvKEsy957MEtCugM7n5N5VKbcfQd0zzmfZzjHNxaV4ZwnRS
YS9xTVSE0Ej+9bYO73YcXobtwFvEdvzyl4ydTOXTPadIYzv3SeAbB9Mbh45vLFuEx1NZthA996UK
TbRoIknEISA9Y4sHL+TLO//hx6Rg9BICHMV0TeqG5u8hJthTjWUOWzBVrM0OK+NhSZKYcMnRrC76
zdp/7ni6xEgHQ3aN5cvXKSkp7CTGsjkWwye9XJ6OeKEQLLUbIu4ubOzITSOABZUmiTbLfaexu6k3
sOcJB8M4nMth4V+QPAvsWnnWuNwge/FbDfY1n9Cxi75WWdBZ9V8H9EDwttZBv8SEV5j0uN9rrG33
LEdBOwRRBWSqXSg4ryyRI3q8DaJbT6UiwjTCHFr2VnkmG3nNyjQTN+w6zr62V6nU20sGAyUwmoph
aMGQtz7z3NFCXvsS57TXQZY5Lslf9AZKdbMUAalOiduNc1YWsR+laFN9RvOuqsb9xKu3ntyUckUz
FKl1v8848cPC0+GrI4uIwv+8tuWkj8lTt9AZ1dKuacMTxoQE3bhd/9bA47MAhXx4nxNMvaWr9FgQ
mSsjv+WgrL4npUWg82OGi4fZuGJVt8xymXviCUvEaLyPNi6VYNa5zj5JgUhyB9k3cG8oBzyw+3EZ
SB5RFGDGr9vmyY7PFlGZKrp5gmIun7pZTYNPXV3JTRxBlRrLvVJqzjXWHcxnBW5l5fV0IoTGp9JQ
hmDm1HSoRvho09v26Q87AQDRF9Isi/Hb7/H0k/K6fTgZ1JnlyJeS2UHYpYH8mGAzk9KJen+Mamze
AhXfBjIQoJKrhc4clbR7NI3OYzxGLL2i8drLmuW9M2RRRtOnyzlAwBP7BhnuFGhiFiFuDkc0iqwE
T98i+yHWwoLIhn/Hz6OGpUvoBtDxFUel9vygXBh8QewvpBSLIwZga4qfooIosS+E5Yfr97OkTi0s
ILDTV9t5VdjDf7XByTv1Ks9rrNTSzGH8V+df0gv9oIcnHk5+2KrHE1OqP7/ejZPoOWdw+o2KCsV2
TfQz/zY38k8Rwl+F+31j3F8gOELc4Z8Y5AEKZ6M/1uwRd8u13pIsqXeFzP24QFow612/XppeiUYa
LRdkBY9EefZC9hbLkT/vkzdHCtrANWgQ7ga1sJb1NfJofwZGp6O6Rktbzs/WVFv5or5lLSUiIrKr
UerEt+6q95KPk7n8WTraTkHhh+ggXK5KXo8wMwFCvpyWZlD1lsF/6/IfPB41sTJepkGz0RAnkJO0
A0hdVW1t+7WtISeF3qc7fyAz0Ud6O0GCp/nCtOXU0XYCPRKWGevE94lVdg5eY3vsFgdPb0q1a9Hr
K9klrLSKorCnHUBlxKqVnHFxrfcfJyBou6PxSfV9El63Rvq+Y1bmzfWK3PzDY6Urq04lw3XaHCAy
1YDrB5wJ1oB4GCmEEqo3Kj5XrebktCqjKBy9iu7SLaTE4hAybp6nQWUiHty7voNecEgQmpQ7Yyx7
VMYXIz3qSiyi0IecL1GFE5b+7LT+8OoIFmEw2wpqREEQkQKKVUPSyvZvQndzhh3t//ZkRSNxrV3b
zik2mmDpvyxhfDwkptZiA5zUm+hXBAv7WdelxjBWyVo0iPZf8bB1Ugx6tQSaH/PJ/2pKVi+85fVQ
kY+5T0Zpa+LzpD9d8vn/b4vdU1beMAAhalyR1rMGoaK0BMC5AxiQG0WhFI7K6F2zbRQ6LF9vMTSR
RoLGLfv1FwIrc+XlmAVeWd4FjrNSc3bvBioy6kXfOjDc579FI6H4iqIVBAfeswX/gzvqvH9AC+fu
RGxTzjt/roYqtseT+tR8qGtTl+lZzSyt3y9jROPewqWB0LpCRLtc+jbNU1VhzyhHFP7nLn1aemjd
AVG2bz6eWlkfgQAOyB+0q/Rst8H9RTxhe9sK0Vre3vBWBYX1qieFMx7w6BIqYJy7HXCZnCnuFqgk
+/Vu8lEqxnCuz5xa/6Qp/L8053l2gV2Yvbv1wVhDaewtkYtwgGd2JlkpPZscdzo0/XjubAcUQ9/d
bX1Z0GPOuMcd2/1ZqY/9G3RHab9D1A0C/RlkoY/NQJicwG9oLZbnyFaWrpClzxOphtADqkJjq6Me
1s2zPCSBIj5zSX7ESqZ8Zo4OdKGVEsfLmZuoW6hGk8+AQzVxfWb+Hvf2T05EOQXA8rLB+ImLaG/A
QC6ZXoAIQLv6WkjojcUkqDWLnjorJlsYz5CgIJndq9M23Iq8uujkG3c8OnjSX/X2LOwDagEdXvQL
zpcKCkqr0YjKIeYx7LdaY37mddZ+eJP3ebR1e87bd36zLi1HzxR2iqQQvmkWpjsgP1pwuPsLTArN
ulei69WTePzwbw4RnmZGYY6psa426mGjBVlgvxRJZbCTj1Pn8koBBE03v+/zPNKeMy7iZkshAmri
jXgb54+2uI9TwHFfGZED9VF8l0Y/Z/dU3JNRGlMnUDrfIAOBrsE0Zo6NPjrDiKmJ0WvRQkZ8pNYJ
4y12UJM9gmCShW+9PyaRn2gpmEusZ9vgc3qC6RyEgglkx00W8mWhIT03J/Wj3L4tCIuJUjwnmj+a
ljfte+SAjQW1WO75ZLojuTmmmu0NWDiQQfJ7lBEE6xyXn5GIw4LFawoMxtmNap2zsdYvduI0i2Do
pupCj9pbs/UK0MTGpQCOtuie43ZsM7N/zqDSP5yHPrIA7GJefRPOLjjGZPoNazcWXuJm1Kn+dQFk
H27x6+xg1qcA+yrgnycCtC9Uh1cnlYYnN6/uh8vMUVu7tLjDEtOl9ee/WMF3CjJZ70OXfsXsHTz5
6Na8gLYdcklTchFARBNKGBRuFK2BbAcPKLmyJBxrcig0JFe+bYi/pxrWhp54xG2NK0VZBeOroPrb
H/A3O/HhoA7b6l4Ad4ByFG4p2gw9lHa0fsUA/FnSw6cDY3Nf5gLEMP4r13FPK7QcycpkXpVIT25c
B+UDotukExKpYQ60o1KlUzMfWRLPMJoKxyhFVY7rme7qfsHv6rWwnVzYibZeNIe9kw85fQ/HF+bK
H6fPMVUEJ//WDHfU612o7hpLdhkC0JG1mKjaGxzxVPgrQKJFybOSyaD2vZD1svo/4ZF/Zyts3SCU
LP8CDBf8Fm6xUs0vuckKfs3DfrRFvvBvYpeDGR74xVF/SUHZBygb7nCFP0onTjc+sI4gRYT5kYw8
9g8GZ5L17otvyOr9g1s+NcOYJwY7KjR0NWZ/0ibnFQaXGI8kllzUSUBid7UJ2Vik2rTzb8pOTN8D
fte2MKQNEt/m8JDbltxxuy+aZA4QP4mB/JQEHMWaWvYWeJz0n3HnSsaEjXPTE5Jd47SxrdJjL/d1
LybZRl88QfXjbg/LylSE4FcZ+ICi/ttaq/CeFCLNd1eVax3CJhvjs0n8a3kAKN/AG6OS3GPlTO1r
gU5FeXpFu17/LUDeNfwk9iElzQfyd2IcxtIxHbOpYq9twwHqLy0zlOuA44rwzm2yGcKOEJdmgxGB
cacqMDLcLuUgKWoR+Z8LDotsZP6YfjSdrrNUdXwNXQdyoz8F3Yxavn7FA06/jQGj9MsxlpCy5HVa
YJ3GR0/kohMYwd7eGL+BCKCaEcoZiHs0eyNe7i8yOfj/iNFAUr0IiqKM1lL+egv36gXXawBObQTI
lBU8EStNiBbTV+lVcprXTbDvp5oMJd9etcbUPJIBfr6b3KUsTAQsGGfDvcfKa3vQ0xUA6GwJ6fBV
nUNYZKkDsUkbdEclni973qjCLk4d3nZZOmpfhW4ZlTSiBwl46pDUOQvPnmlvyx55y9mJdCW9+ojN
Fv1HOfBtLRq5BfIjsclos3uVByglze8jNmX/q9H0HRS+CpOrQpjx+s3wlnVetV3Cf8XTgKMkrWeI
CdrqLNXcY8/rAwz0SC7oXi7PeKN/AjB6KsMEfxifY+VLJpaPlowNwBgOHWbP+HNMwmEnuzLXLTZs
PXwicBW/GZa/H5MPyY3txQBACwVTCWve2LQpGbjdpSYWoxTGG/wbWQqlv33Ccbs+Yp7nV2O/SbWt
gPm8sC33iWSbAOEtATSAjJ9qQD06Optd4ALuQMqvsQgxmC15HszFRs3j9VafcsbRy67zq/eop0jE
/oStTMKQvsHqIqlbhDLH6oUH/vVXQ43vZ3rZBAw/sCzOjDmplxCB/9AsokF8ZM0Hi+4dy88/S6QF
MRRzRr94J4kbZK7noAceg6WAoPzaJ0MMl/hZlXjtO+TrlUugrvl/IkIYI4A4QKmoTtxSiUSdMrcr
remcBpRxxsTaKGPn3/DwzrLB3zBO02SubsMba0B0ivYXmBV/ZAlyHhVAfeQZQjICqyyV3M9vScP3
Ad1l++huupgJXIPYrpZEqxLJaUYgHy9fk83zCBj7sDRlOu5KM2O0tP+gXoWDm59HB0xxRf69uk7k
j7cZSenrBA6fnQBjcssh5O25aMODrnGd5O0vUIS+VVb/TYDy+QNGXX8WxSWdTb3sWTOiN7mSqTjM
i2fwU4CM1TT0X7wUPArE/A0sSO/6VdpTNRquYyMZb4FqybX7hTHKi1fCxV0NLKMkV7ujzHowuLRe
hRInTivLVC6H6ArdiY2Tig5DtPoKPbHaslbTHV8MQ3Vj0vt9qUoae4li6Brao5Uh2/ROSZ3h4KBN
NJNyiBPohzUEizrDrj2orNwd47w26bw2pmZKQW58t+ZVbHHr+0bXBSFza9Mlzw5vLFPFhSuIaPiG
owzn8zzsOeRBZ6kVHybFe2Y+nWeMFsTjW29uaOfyY3dcMimEZ9scsdM8kbmgg3jL/YunrzQpcXju
1YsXK4eHmfOomtnNnV8WBBjAKjycFyJWGdcqJMKXBFj3+7kUz0MA22m5O+N353CgYdBoG22w5nuc
8VilnmEi5EUFvK4oj+2opiLaCOi/2Ow//xFIHEJLZMdO18Fxd0JuUVe2sZ+YMpVGrLEIaGoss/0c
VHlz4H9YJCAHUwmhrsJF6ul5tMi4+kLImF+Xlvs0YrAIFog6CadSaI9Y7xaRZt4uywSZ3SSfdqJ7
g+XzivOq50Sz1fZcrzaoYqpozHEN7crfE9fRFnu6SGluCgozLX7+759oKP1V2sdFGzOBzP4S49AE
jSyYegNuS2tCTPF0ALo4XfoJ0oDzJ/uJogLilcC6BANePG/Lc80VIZlmohNFxpDUNlwgFTDKrD5Q
xJv6d0mhwc7qBsFjXdrbG8/Y0CJiM710QivigyL0phB9KOZ0ulajxUWK7jBtBie3YWecMh3uTm96
mLncChjV1jEPfbEgk2JyU+HIpuGq8IiSBpvTvPcxnOCtweQjkfOn58kUnJWYjx//GLTjk3m5b1Cx
8tANR78ydrq1+dON1kbqlruJ3UA8lYj01E+Iql18DY0aVQnUnPsYdWVUwmdP7fyeC1t+cfHzb8Jj
ap/O583itaEyO+qdm77cvZ+tisWzrK9blv6HHPyE8PQH4wToLwhhKYAnwsjtE6ryhcjgP1XEwgAx
ASpKjnff7oZbO9PJUvofamAf7xZINQeiYjOUkUZ6r70bBnRee9uow7wPeSgQeTuyAGWbTN1sdKP3
qYBaG9PrR8cXfwsHC9xaj67j6UPBwZIpVa0n5AmM8BzwEemVlluWHU0VBGkYGjn+Z5pD+4KBQ65e
IM5itycEOpg2DN1n0U8h+m9qdLjlqj7uIOoyx2UP1e0iovZUpHMLXY01OcyuN07eiw1h+5ZEWc6C
oxRja/h7f3LV2AFgMqRO9axJskbmj8/UWFhR4FIJpGPfDU5WOKvTvMJxzvk7ZR9CDbcSq2zz40qg
G3qQOFEWRfUtc889NHIvQVjjg6TwrKUTABWbLKPddvfCYSFFOQacWJMXIz6wBYbDDzi538X501rm
GAJv8VzsJFNuJPviLFlV/+bRdSuAywQkCz0vmEk/4o5z6fU7hPqd4HIbyue3lPSGWnu417mc9Ktu
U8kgaYNDF4pOwDDNotDcAWEthjlkacsmdY9ZpBIMpS+xiTXMJ8lqdpmIb/Ph9O4j3g3yenTqMxjb
2HgtYRql/QCN3Yg9iRJJB+FSlzuqHsHPsdkSnPiuq+R5TagsMOHL3EvqIbqMpWKMUk7HkamJ58qZ
XmGno3wAWt//xKyMbfuFvO60TDsHct/CN9A/geubPCs0Sh3oPJU6m1ipkpkGdFW2Qh71rirZK9s0
ZUnP+ZHnS+1fJXyAVJYpExZsYgaCS30Ug5l7Z19ROozar1dIs5CYpZo7pKDQ6+pwh5FrbdewVl+C
RTuM21eWiHzccPzKGxnSbFu8b/AJk6/zizm2n1h3XqoE5hRd6FGD1PqgeI88cvQYhdCEcPjiEJBU
XCkZKGLXI7hQM5tfigK6rMUJc6od1pF5YuA4dW2lk0aNqxEwUd/osRwdcpAoOddPY8yr+5m6B0z+
6Xg98OqDkyOaE4PmRHtnIV297avMOhkBwgSJ2l4lQz12MWqatV2wCJgbYsblFPunDhpsBdwhA7Ch
zcWdbJFYknNFy0wDeH040S3uQXE0gAq4Zso2Kjh2HXSkX84TiZGwKOV/FwEYb4OELcoKYQCqf3hF
UlO8HHWUJJPS71Qvx6FwgYvNjiWkGXv5GITidNHt6LFULzh5qrMmH98buOY0AmjhR7HQo1EBd97q
SCB8RVMNYVn+uhGJEP1hGEiGhPhIA5UIpy6Fj7Kj9FZ+mq4xM9l35Qva8ymYG3H/rnSLnlipCykS
SdJoGcHYk+10i8obE2wFPQnVa72w1AkBUhhdqA6YAq0xuz7PFgCLDylyV4IVjOl+Vm89mx8VJQfi
IXU8ll7d0ZBmXQ0kYpye/2iAa1cdLCJpMbuCrzrOyyvw/ursVMTm1Ao59ZQE87jOITPj2KdJq7DQ
dpyxf7jKIPXgmfhdk1Ze8yCnTU51/jPIt+4Gbqh7EUSfEOu97p9BZPf2uJYhTXRoepe8JReyncuG
9Aac44gz+YnacXQw0m4OsIt9cSVXx+JA57kZ8sOK7A5Y8NUUJuyriAGmpIIeq0SNS6cXgPY9VtsP
MliRuFrryMiKkjuPpx05uSlns9QE5zemLj9gkonhe41F7pROnvuE9YSSUL+t3PTJZkcz1WqMqzIm
8KbFq4gYxUMey1zUMfLD97q1UZG4yOsA0unwMa3kGdtEeTibd3OPlwW1whE0fDeaWMulF0gsSyJe
uV4Dtg7JP2gjgzlltKkFSI/d2QRcI8VHLo3VZrn/TIX3hxxjKXSbhXZQnJTIpSDL6jMdw5nBjOCs
zrAvcIaoYnmliQffbPyrW03Py7YiAEKL+M2KORRHL/Wj/EuVnmk5Xou6fCfK/981B7m0BV/UdZRQ
Y72asFbulj3RnfVlhbWqFpzl4VdFJ9Wk0S1Aq2djoTjknDO+gnkcIVmmOxcVZqvcIpPCDuK3hYNO
uHHHRGNOf58XiT1rGQxjUt48VSfcTuN8V989eq4aImKWCICsyzbR2rAhHGLpRa6o2HKQe/kjDAfS
BlB/2cILyEfbaq4R4V3aqWdFCigvXx85i9LQhuakpHo2s+bzOAncVYBAcomu/WizUtld9uJ11ah7
W5AHfo3xzfxwmxDy3pd8lkD6PAxQKQtt93PYR0wsZ6zyrMZYP3n5Y/YI9+fd+w5nmdF01ce45ptC
uFtkNPExMNEFRJrhMfI8WJSqKA4BYJDPYZ50GdoJbLpJEyzESveHUdu/MnAPEQcG5rm2d4plRDJo
fUZiwrS0r61qbb4Ckogal9RLrR80+cwc6MUl6ry/UdCBKVRYQvNyhjEHiI3kWRiVPYKkGBNXDoIg
2/eg3u7pMOLLx19cHgC9wKHsu5QROaWIYWVgzAetu/M/34CWyrFyAcprp5pDiH5tbZpZPKL4bQfy
fFqISnyXaDE/pL4DQYKiekYV1h+u0cciz4Mua8Kt4zhvxMoNIoZ7sGBTtGD5p1xKFR2rU743IDgf
LOVveTgzK17hu7hL0/Wbi9Oz6HUY/eb+SyiVBdrzNQWy7q9wW9fX069f+l/H5eQKUm+dG2c4lVKx
EJtn47hlU2aONV4LSkyJj3t4gR+Ax1FZy7+wsuuaYnSDEOsy7F5i+KQb8YK3d6ZqNEK9EqE3AUSG
ggPZAP1gHHJVTHKqDe1dJceY8D/ReqS3W90/zLIA8fnPn1l7SiaNyDlYJPNXuehy4ZHrUsFtt4tJ
fjzzClMYjhTmjwjYs55OpigWdxPUgiEoHfRlNTjX0ltfqMPK4TzRTpnSxzkw/X3DWAwGEpkFPpgL
wKUpov5RGzkbUAShWQMr9bW/9c9B+BGqOS/7BEa5EwqBLKR72YzNtXkJSwDqDZpN5JB7YS4huWgZ
eWyNCpRLFCbmNuReLNPG+dobm6OhozEu5GtMqfVNZ3Oa5F8Bw4MQ3/pvFr8fRWSN1M8Y9C/87BCP
ye25YWQpbKZOftNOKMRoZYdjlKAdd+OkVr+S8RwWnta7s3iuCKnVAsbgY8dW2+UBdkaG5yYbk68j
PEU0Hwv5jg05qa6bwV3MWrARzFLMb8SoKUhGSv1L1/wLnZRq/jsb9uG9O5kUGHiDK5FLfJTiNUSN
5C0luIJ+vJKYdcFGAXCXfAMymkNuDvuKkhWL60IlC8ue1vhcdBUdPuuGh0NmbZli7EQiH58pTyeb
Hed8vA6VDDqTUcf2HkEmxA8ilJbFDSuTf1m6dvFSG1F9/tfJHj/eLCAbKMuNaifUTJGuuqQLNxIu
vW/GVikNwQTSJqGkjtmx3buiO/TbbV2Uv+0FD493VE/ID9NGl6Bn4awDX9SSpKwjyK0uQMCMMU9l
pFGNC34RxfkZWoagkvAsgLI24GA/QI/JXuIs01u4zIpFD2qcj8Gro+mV9QH2Khhnj6ntG4x08CIa
YlGEUucG3rx/dWEkPTU7xkZILZIs46Nocj1WcFdwpfMshXgBls6e4NAmq+ApRGVKBKGMdzIn1h4u
vQ6fcolxnYLbLnY6x5H4K/JkxU0cXxK8BxiKz5G+jZZjjNfYZKfP2ZQTaMUe4R/Q8NqMe2nGj+wf
oC2FNU8JGpICXiJrlP8Kd4iOkJYt1OPKi/1plQBAqllEFqIrkvR2nWsmu2q9AEkO4muSXsZpJ62w
8Nas+LlGrYCUBd+T5CbOv7W18+sa2lBQwqlmfMGRsk9VONgOmRl/nSG2/zuDV+jA9ce4QnQhjLIq
EFehp3aWxTJ0bAMEHY8odJ46o4eJ6M6vRHyZN1RGcz8ZLSCW6ml3xFoc/T3hi+ZV0cg3zDXLz43s
oYQkoy7224UfTJQw+vvnErEKcRi/5AK8O0SCGxhPPi0tlvasy07m1CCfCs/pAYLZL7xhH+1IR1aV
b/p8IL6Mu3UcP1NUViVcXOkG1O30Tz2huYLAO2hIgzcRnop98ERLUc496x9RWvrWfKTS0RbMwOCe
q8fAJ7YrcfvU1WeoV0A37mCCnH1o5/HNi0Qt4Mrfh/cA1ymc6LcpCciav9s/LAgfKYUH4j3AyJE4
OKM4/UR3kdJqpuwwOfnbEEk5Js7HPjvMKzWr3LSZOBpJj2hqtciTGJTmrL4Nd0LqZXXrswYGj9aw
TG1sUdyU9Aid4Ba9xQQO+5NEm1H/5y8IhZcSZrNjItq8ZWkchRxmBiPQbNrJ5pjUWpXYKbC7vE8u
OofrPaye75wyZuwUyAZFAAxSQOdfj4e6+YogwqnshXh1+t2VklWm3RxaCYcm6jas0ivhqG3YR8gD
VutIxhGS62Q8E2WV3y1Jca5S4jr+4lZZ/T2/jbj52likv7G3sUUQchGQv7pOYAoTt8hd+0QVKj9U
wx7iiZafCw1sZPdV34/xkfjr99s+2Q397c/mpqmRy2XxqNXNbG0+K+HxZn1Pv2ZGwOMyX31FNm+8
gt1vGzaO9JdVvbFVOcPIeXycdxDO9KS4wDLOonHl+XyPKc4vvhZaqlmhrlIxwkrkFEVqrlNY+wrA
m/1rpPguz8c93+zE0VJDEAv61g1hvVFq3M7M/ZqK9JHri++SDmKfRSCDvfCyA3CEYk7/wCukOyHv
YMpbDREd7F57CcuQ3wTeBMFCroFnL9m8uFq1IGI8cfQX75HLb1WdZt9NJa2tkFBn1UZDn821JKy5
K6uq/xpftoXLfcfObXrtzfKsW4k92KPrmFtM8gyEKI6MmmmWyKAhbDpiwFNCs9YG1bnyWxwsD4er
dEovK/yVzS5CBnwP9rK/NfjNp2U6fmMAcPx6PUx6SayI5/V9V7jdhyJsLPFpevIPXcIBh8boSy6m
ty/SaWZspqBz3nsyO6ug6uoX6h31WAVImSfbEjEnHjDzcijtF421IwkCN9Rv9eXYeGYm0zv3AM4d
52dfIm7TxCRWRa1VmnRj/g+BLGRbRd2XYVaZHGihKrpK5oMcYIjujt/S2xwZdsNSv0COVuNhUw4+
fRxpbj13wsp9F7Z/kAtB2gcpoTaFExsfDkgJMCchf7HliaW4142pg8lMQgFP3GrC4sOirUM1SXBF
4QBi/v6T+PQXqcR6HggK2eY7QN5fuXCUjnDorvlo7aL9Zd1CkuH3UW7lu8Enm6o4pbBhPFIiaySx
n24R5WMBL5c8H8l4jhMrLghbKDleewFNt8v6zuICbIvnfs6XcsStDLyaFrVTo8q1QOpJdJKwhRe8
bElYKpstChCqgQZ1gI4VDsSKasKMQP+tDy7+nMGXHF/kFaySilSZ+uRxz9+g8/Cv+biC8KsKBlqw
dICkRiV1sI//2UHr5XHaq3nrAzfLSrbmkAIJ7BEPNxvYCeqMtjiivT5dnnSkgZFt2/MzKgbc0Ykk
IKr3pMJkW/QfE2CrhackrLM5fNC9LlTVGLIYXGZ+D7jlFTPuNJt62hMLd6PaHAFSBHqdpw5srM7c
kHg8vLUsxaE4bR+8HafRiS/dOhQodBm3uzez2Bg9jB4bs/SkG+g7+wvxzNKvmqG5VnpaEUDo5CnQ
m1/F/1beE4tNm3brgT3yPCjy902t4ZO+ZhYwhQEm+x8+3KHUh3pwcKJ1O9oFElGNanc4DIgfmli0
zNalGmeWWo3IypWpCeOZJNYBLtDFQITsujOj75GUV4pc9ne54YQKSfYPNtu9fTKb1lal1/idac5j
jRfWvedoPi6nEozGEeaQElwtdab/AGFJB6N9EH+WG3j8I3BpJiT784S/vxIWdVMzWrlcm0UG9jo2
c2VH4L6AANVBNEX9UXB11RsnKAAhF+JJjJjtxXzbjZ8OQZOK8IgQIDBoQpTh+IBTyg+2qbDQBDfe
1o1jf3vGhCc4Vy1nS1BZmNSe+COVZ3krRTT1s2X+VFCg1A2q8r7eFfdai445yLi1rwWK5Miz9CfT
DzQQjLOm4pmM1n83qTkHgebw0qPmZeIiIt2E41ayIuB91RGUxolUfJHapgCq4voIYs2OzrXmiw1o
yHmPl+F+JFYhs33LzWwzTOkIsCPVZQJXldSrrxRSA1GuYIrxdosQ6UB2M2zIeUl6PbpCaD4Xw9vJ
PK+o6UKZ6oQgNz1c9WErlye8I3roOKOce/MhNa1MN9NaOg9wYCGklE9wOBtcpmf3fYhyQ/+5zwQC
WzkidwL6T/U3BGfJ1WGkyc2kla1vJBokAIyPR7VzlsooukSIGaF6QAk4SJxHuPkk69I1f+SMH6yd
qJTs/v8l/zJGHZuJKsPG2oQ/fyw6bvsWhcDR4v1jvElJp7698sjfJLyBDDUsCKasUj99fdh2q0uj
hcTgkJ5hFG3XflRiG6qhXWcL0ROm6zs9xCTUEydA4pIcRFQJ160HqvSmVPuWBcjj8kRHmm5NH/ip
8X6ttVAp+5JE8+g8YFKrWlhImHdtTvrqvrNGPcSoVUGQE4VjOQYeaI62E8U1Mq6Xj2yYUxKha5y/
Gw5MchU6tUGvr9XNYTCXf6w8T0V3JKTieBvUpev4sCvcKU1yNPy4xwFHEzFpL68BF+4x548xNfds
PIssMgG0eoGFZtJ+vayVHAPB/SeER66iq4x9ruQzWMsnF9NXlGraLjFUhPv8AzkKtzuWxO9uToOF
iemu8FOObOFS28MjVBsxSY5M9QH0xGWkiquE3IFt030fLPoP/2eqG6lsPtWWcQ1HqxjrQ7woVg8K
xHhmNpI2CLdHZHcaAIT4qs0uTfEaZUbo0AcLmTnGJD1QOI873uJCnyp0ETd3LrSdBZ8NtY4xeBud
keui21x53HYLmh2D1xn9TAkHBgkdagfU/bCsHwJbTWphKT8IMxvulYjNh5VwgIubIjEqjztYnqcK
b8xpYTmEGhDC0fZKAIWh9oIVQgMzpfaIhk+9fuOhmlH+H1ZWgnQPDG8xzLoA8wF1sL6WuZ6fC2ES
IVGt4zr24PJQ4D1TPPrA0Ha4MzrtLYiSZEf8/aLSQTe6XivaAEyqaLwtHs7uAnZVtUqXRDpG2tlx
/uuvaiwxbe67OqJhxT52ij1iMV3rKT2YkAHLx7bS9lBzI9rvEb80nh0e4/pydqMDYjcTlcuJ0wLt
Je/6o59XnP6HPsWjHoI2DDsLIpticx2ZplW5PWJkQEM2D6/eqlgYWV06g/+IsG/A8qQ7J+3092kz
LnR09pkdLuNxHJaikmBjhawZA9xXSeGNo3f02EWy+4nunrHH1Crweb3WiJcEi+/3d/MGdqxxXMrv
lZrlRR+iauHanCyz5QAPUbbluPVyqrCXxh+go33euBh/W2yeYt93iKy5JAedUINcmF8uwcsXS8OT
WvNQSwprGTwTlKOnmYM5xJ1GK0kI1B+s/WLDorJHq31E06gXSgTbiLw5W/99rK4sYA+TO9ZHF4eP
0cdYBLjtfBLFQtcuzkHlw1dvLrlnfkQQXCEEtbWauzl4cFLVSF7BHOPVT5uIo0vAFWxixWP7RRCF
RA9kXnHH0Pr/ELhZiSr+BMWszfheJ+CxR8rndOdwi/8iM66H1M79o7GqQpevQi88J28EqNLE0ulY
l6NcX56nXoWmL9dNL2OheUVEGME1YVlWp4mu9l/lDXRto+YwxWr+9cTAMcYYXwQaEFoxIe2rf7AM
H0/b6cTgWvY+pkjDJAAJeMFVzQqM703r/vDzgobhYqv1tsLQvT5IeFVsa36QOBacR+OvZWKUNlXN
rrUiom488tHG60dSqJFrWZo7pbv21JOUMKUonBqgcCmR9tczy4yPc1qmnWnMRO1J+1r46e8RYUS+
W+DgQ6CS7EHMMKjgx/eXlZqv4CjHZHn93W3PIyfWPmTqltiJWZuE3ILXYR4HIXPx5VO+/pRLnMiB
y8XyUQX2gZ/Z+lY19FMr+Qvd4Z6ckmHQPpFw6x49vR4Vi0IkQ/+t3SojBEQegfhPkuPv92I/2GuA
oUWWXmRThWjo4uZra3u2Jeyn9q97oApXF8KOLhnGI9aaHROi/10HTMx38++jH4LIS5Ld5w5kP9Qn
EHnyDzHg5oJsXMOrEPRYmnPW+K0avGcztA/IqOUanFyRI3y9KL5GzP/VStwZFJYmIfKGD6k9C/bx
9kt1nbSJR4YPPKby0RVP9Qm3bBlZ4dpIe3nBHK7bJW+irttcsqj4aqkAntfg3UyOyPYXt1W8tjJy
U5CEiHh6nQ5ilD92wxY/zTzVmD4vLNxUYh6NjXbfS8dck4jyDPF3GCRCZ59GThVFro7b4uvC9ndT
N4t16Qn7j7JsBSMXwXjZyYJ/cPdpLeqLl7GOFtmKrun2h38DieDAk5p0C8mpooKEQiQypYpr8HSP
gNwICFZMOG8vtCr4Y3QW9I5wAqi1G0zy9CtbXooHS/9bt+XRTq+PW5A2ecKrEAk5ZCdFPpBsP442
NDpjfb1VXOWqDQkbBkw6nocQxdF5SMSvniCzxVJZQVnRmi/yd+7N+H7X5R6cunTihEI2dvn0ooX8
XOx1g+oAR/M/DGstzmrKtWyBHMC/0Tf9X325Mz8jVIRRlMgvF27k4WzU0aqZQ7wQPjYtslHJqZKS
LCPXg7sExwC/lL/cxxVtskDN06nUQa0eeS+uj5UTEl6GP+1c2VzH6YeIu52zL/AgazKdZdoPe6EZ
Vo797EKGidF2JmZVmVPjiDYUXAiDBe5UYQ1swVNa2Tpc2/NwgV1CmEpEqCTnVvQ7e2TWKq6Ixipd
lu3Fn+cFyv8vzWUBSo79pWszDp5CkW0ySLSLl9abbSI/uu6i03IvHSRM7fnYW2htBVvXjHZW91Yn
lMqHsJnvuf/8hSfCjnn+ja25nDE14m4WpAhpu0X9AYUSlSioYom0Oa5YTk2njvLB2ET9WcVg+Ftk
bcPR6sR8nQ7Z9gBjKABCSjf9+cd0g9fMx2Z9I2uy+1nhAkVVEP5zJFCG6wCpVJcs9q+w7eVqhLrD
wSh6oRJIaaczRHW7Io/ma1C1XIRZJzmOe2MwZzSuaaRN+N5F7UP5rg9v3oqAU/06T7UyYvdsnQ48
ZyMmHPTVRQQkZsF8DkZKgjD3It09XwZQdd2+hJ9t7mhu3OgH/zWtqe9SLCUfxsxxI+rwbd/FkHGl
77qnQMU3YZupLxTy61ZIYWBDZD0JJlQ/TH1MTTT/yWok2/GR85UsRNlz6xGjO0C9KKVDEipx4Jgh
s3OW/HEb+eKTZipp8mTMPt/kyQbeUxj73M5GVAWHR2OV0zXXOaHcxEmA/99WFpfwlI0v3o62JV99
AuXhfsAhABqfpIQ+2mu1gDcIERasBUOewWfs1fah1ZVl4gOhb93JgliMfOi8V+KWCFdR7n6H0ulh
pA1AN+SsL9JlunpymLRdVjlgO0QfgXqTYXbFpPbQHBNzDS8gnXKCMEPRPG701hiqGZ9+3qMV+/9o
W9A9eA1RRXgznuu1aX2tWYNTQqF75HuqSW2i/fzh7qIspahlb045NRahT5JW9A563QIujn4mVUNI
rgVYV+b15rtcup6vb2F7tXn92hkDYH8YbXXA9nS+plnjexfUq0nwAqJEAAmyA4DumTGZVqCSGEQ+
LntMy9dbE4WOAqD0+j6W1rfpWk3bz9snXqDnGInhvdpK0rMb4MLdb1oJP3PlLwSKJaFjjzm7fWTi
IL3TiY/iGTryypMVW8kuHRdKeOAtQzvKkNYzOWfr8RzURAyP75ls579fLWld7orpuPAL3QqDVdQb
lPg0aMAzjxn4zp1UrrR3Ei9fbUBxH3LlfyzJxCsfvjvG5Ti1LnK6PgnxLDIe8mqy0BVZ7YiCZSfc
lbMfTo1pgEvD0SFbeUTJo0xYJgQGKEC/tdQElRgvVfA5OA/e9O7Xwqm7zeLLhw1xBVFBn+PREv6Q
2RIle56OvkikYckzOZdoSVv4wpmHAPdY1B433wewDAta3EZ1Xz/PcPRTVlbF32xSnn2t3XEHUKri
0fIAUnNb9TMbMVp5sEsDu1rezeHXFwuQk/dRjfAKdzKosBX3CWpkze6w59iY12PmmEU9RrndSFmI
TPO9GYD//8/xlC77yD+m0Wsi8ABBcKyDEwVCEownr4nmm4YJoOMmshnKpIlIjgHXmqnt047J+Ih1
40vjoGT7SjbQ9UjgSCoYgNv/HBNd1HS0UZUOpi/9cOSC7UjJnwnH68ypcg5SAJtJnrYFwahie68N
CXm5Pzg6mlbTOSK29ZWYSABSawwKZKndS+Pwf+sJQLGQSqn2vpbikSsMMM+dbVQRaMnI7JZ6x+KM
d541QuoFAegTpnOfkk54nyxjpjAZ5G6LsXmNSVXakB6sJ9quE+gD0pVGNF4in1U5I5zLpkc1XnjB
0pHcUzF9YtIw8ITIG5QJ+5DQF0N/XE79rKsyHoYABlEVmhjeIe42+elEqkck0TaEE7qkECKF5xQk
bpJnxZ+iG+aFcjOe0UoLIupaUZFvYAI2yFLFxCEUIqaUOYPBc3X2uznpnheDyo5ZiHt79zSJoL7f
OGOgPAgpSSkBNSVereogqhfJmHHgTluwfM/FxeQVzXbELdzNONID4UGdxBNtmlRjIA0OufkrMcXl
1RTztC4n1WYMi/nlYo2ArVlpAyfE4qqyaccZTvNLm6ssluzVE1YOYwMCD5ENenIRL7xCC1gkQMB0
jwUuk/88LcH15Qp9iASnO74gT9WhKbwGA/+9xLEXVIc8W8LRzz52BpzukxCAIxyfZ2DQwU7byN0v
ZNJhszi400+UmJAn5Ig7t/B7zsiv8oOLGVs5QEVwOhLoONQ4X3+CvRbFHX5gnbGa1jePjf6DHh5L
Wggsx0Qxr9hHnkZVQQ/BBmbi2bkf9I9DTrhT974IdYNKfjul+W9fnrG1NBXpFwoGegRRYlxSvWg/
wSVK6ZhoLCt3K/04Y0ly9hwwb3zp4mcuNmLsfpMefCMGVpfVRJNn7Tr8FmRXsY5Vllp7gyR6f5tM
ZUtUWrUm/TZck0XhwNNlQ4Fe7gZdFe6Vc3ohT6tPZ+ByrAoouGmELa0GAU6UpUWp1q7CTFHjvSKH
nnCqnF/Zc+UOmcKH36O/ruh0Mn0opK29Sc8VMSlBqhF+6zXeuXJPse762Gx33koCNepc/cdP0DfE
ePiN70lGoa4IStj4EBI7c3fDWGyFUwwoBQxvelsoLYScSJq5yjsKU9lYN+i07i60ZjochE56ZThZ
qzdFubw/WUP/4hcTcQsleSLAgfoRX1cEQGyPolp1AWG+ZzFvxMhOVdwcdWN0VqeEbo6LCiqndmzt
xIz6z7hQCfgIciCd3w5QIqmT54d1AUiSUjUxKNGcfC+Yf5k7piVgZlHQe8S24BIVVhAVtFUo0e7S
3weNTaHGFb1zTdf2z28c/7pohCpcEvvrdYnujvRTweyNqxk6+uwjHGxi99IycgrKiyTx++XbL8Sw
mh+43hHWxwv3PMmLIixkEB3VdyVmWaS/zA+cWGOKUxzCSyFcBfCouQB7eOXIM5GV3opkLsy7yDWB
DUDt6XRg9EZV9JKcp6Ba4QwFK/KIIE0RV1nYHXBDqnGAKwLprrHKsebDca3K+UdLPqpwKfxbU3sU
qFNS0E+nIE8IP1+zNAWjmsOS0pNO+DPpDaT/Vb3wDH52iZpuBjxHJmxum9yFQujfwp1nm7ZM62m5
RD6DoCFF94dfradRXSmn0oX8zTTtIxcpn3jX4rkQB0bSgNVriWSemBD50MOAQv3+y83HH9CV9F0d
9PCDEm1piZGqdfoShT4Tx5iYHOD93j3A8yskJb4FUhGhsTyV/OCoeXxYlGIik9oU6JD38KYJWB+n
ZxR4GHKV+zJcz7XVjjfwO3ajoDVOYpCBDnLYeX/pDRH4B2XjrdK9WkXjfL/vD3ASc6lMWa59JpM8
I4heuhN7x0x8bNN2CNg1XqLY+Hih3fBjB9mU5Wc+tj7YCvo4uuWWSjj4/wHTaJLvA4wdua5tS6C0
OxMXkuWDAA9Ck5xBOBMeOpb4ncUm4lQop0SGEheDXQyEpGaQDAnnRpGmjSGGl0s1Y9M6wob4M7J9
NmMrRgor8ac1Xg5N79M3BnFjwcddOymdqSPRBxDMPk2+CM8AqPsjZRMjPx+FxybyKLdgystPxsVX
O/wzR5eRcAAROM/G2fyJoZzkB7jfVB0GSqHrpMuqsNj+lp6zdKNBUsKacqxDmzQ6RBmqqnTNfAB1
cO3Zo5QIwGv87TTLiDUe/yt26VawCmJt01vb8iUCsIW/ynOKB65YNMzwS+kiDOCXL/cULMUfWnTu
PAQKXctw+C4QkMczGWaDnsxBcCqd+rPVzYO7LozO8Lp1/xJC6aXe4Y+xEMmFGwF09YnXLqVnzmre
no/HND64C88gFitdIEBfwx4RLzrIpC9KsTtOAiLzcrV95Ayih2QzaI/16p+00zRoa44Rkb6WiAUQ
64TRSFk9+51VKgxiF7oYqdSz6Br32Syms0q2T1lltzdB7cLTtafKF68HLxjB8tnMcOEIZS3Keasm
C/eJ4UnJsWHZVjMUggbZB9TTNrfWBYFLvq0dm0VL8n61rW51fOtNS/2M/k5YiD0VsrwAih2AGWaZ
c1P5S2h00ralQ/Yi5vf3QbAXCzy2OLCSBKiAqaf5BYI9zlPkDCt8XzMIlKPE0zxuWkQ3uy93mVF8
DWnBmYWxe1Ea3XYJheEsMK3Rn18C9LRHmQ/dGKMGmYiiIinHwVE4CNauW0nvM+VCVVYOJMiVfi80
jeZ5RMJydyk5uxWtDNwVpA1CExdFk/t5EHRea9nbPknkzpPm3LU1+1Cf2hRGqESBSN8b6Gf8r717
tWNHlA24s6lVg4/ruxqRTUbFKC7eOZw2zHkR05zUqJiG2xC/9gFSlSz+UXD6fMTb+/ViDtgoODTx
G5MIUBaHbKpWRLwNMH10mVZpeE3pM0C6AIPlVRAQ85GoEB9dT0nA2XLx++2P3tHzywIqEoJX2MFk
vQtWT2USC6l5slyj1Fbe/6Y+H/LMnAnMo+sBks4xMRIqHmyZNW+Cx1sftt7qis08e9Hh+J0nug9T
4nqqDUTUxGDc4KAHsqz6T9HJmmHLZ1bd+RKXJLcrvMqrRq84rKy5plfSRPh0SaqFfkKlX8nBQyr4
nVZ+M3jb35cpL/hJwKVX+rIL4TaSUpo3BhwrkodgSUUnw7gASy6KBOP8p2m2Vx41ldFfOd+wnkvR
5bQDyjKKVFmluQIeFtgswCAFy83TVfzk1213rdJsGCCqm1lY5znGDxil13GDQ/lcVqRhTdV+jJQf
woa5+7s0lm371ZkJIFqmlMH3Fy8mhYLZKzcj8TbltraBCoPD35rLn9VJtDt9sbKYAjaM9rbYHtOO
Q5eQVsNgrGgvFNqG8reAnm88U+QZHU7OjcO6pZ+0MF1qVYoiVMa24DK5m53O+HgUDklSQbouy9FY
F9XqXPgBFSXhyL7T5tyrv3lDccuy04HcqGALfI4zQe212S6sUp+ZjRbq600P5owCw6ErsL/8la2Q
iF5FzyjFWIVsEW0JNz5jqL5W7u3df837+4RG1rRJC6IFdWl/DIgil62VlXAt513u7QSG3lI5BXGH
9G7UpbshsYSUNobI3y5P7O94u5cetAKJq3EiVLtlffCwjBkESrBnmH65yhX3I60qd02xRkDthcZK
jyOwD695e8bBAIyUU5+N8O4JEnddI1MSjgH/wTLh7C6AddTLtf0knghAONt9C0yVmPCZRyoxdJDi
Y6zL3/pqqEIlAPSummjPwPwB6iSCCO6BtO6fYZOSM+zGKXb1heOmSYFbCXu6+E4eeEUmWcGPDBOm
tWBPG3WYBp25biWvzmuRed5VAhK7Cpv1/HCc1vPVPIpElFQWyMcW2F5zYjLIyZz42iMm5JSq30oY
zXrhP3FjkIFrg/0sXDoaokdJV7xG0RX2VTzvh8zRI5iBkbKHqHivRP3dS3fvh4gzxIJvsmFq5xTd
f37vnILdAnCMvmV6ewGQKwsbbfUjkKHyDfyT1pQOakxK+QQyy+nSS+5DpcEw4Ckb1CchR4+RkahU
Dj6Ra+Guifrr/BzdrelINUxfKuS2bn8rcL45TCwsIE6efCPrmviq4LRWr4WjlP2kqlNcWf6gpTIS
dTmh5NEWZEefUPfTnpzYN+NOGJN5G9cFRxXAbuUeuDbemIs6uMGNYSC+xnTS8wpDP3lw6gR88Szr
gpK/178QFv9HBHU/B1G7YxTUo5cEG9cr5KFMUy5NM6HaDHFxoA9zz/gGWsJW+5m6NSj8xTJSMIK4
kO9yZ1UzsmC7cy3DeDsWR/SouEiJ9la0oMZcEqb5wL+kXKvkSaLpV4ESPfUCBYotItLbVcEmAI1k
oONv1TuL9SE7yfjA2FUUQ8e8HXrmTbUw6heQeuHWmByj+R0T/AjCZvXY0nQRWgx+ZXpTALeOnwQM
lGAHYXykV5Ap6qpVxE4kiuDzfIe9/C1ibGBb3+OV6Xwszs5W2zYftPArX1L07Htu9etVIGFpSZu/
chUm2BFN6snnJFxl3i61tj6duqDYylA7HzwIct19aj6lgEWfJCKYBNU4lT5bRFW3vGr7YabaPwpR
UL1oxk/W5buFBSLFVG0vZBvAPtuTwRqlG7JjDlZbe2Z1/5SP0AmvGiLK1DKmqBuOJjqFTtkdGh9W
G7rJ1YgS7PV8yCf20iwuRswyE/k9ESYZ/ozGhcOP1KtpgO5YHPltwcKWLZO7j31Vc4C/nV9wHBDT
0yrE1vlF67/5pwQTC7Sqh697jBNTwAcfjJs06+BBp8Z8V31ShbCGaldWCtm4KJZ93XzypY/gueCo
dtv9eXzZOXSVqOmd/HwJF5A5ox5cl9s+dB36m+1xB2VrXq7cie4IdJK0k8tlnUshEHWhfxVoYZg+
HbG0bn9fgooVcDyvYMcVCk+zujL8y7rPw4+UtR0dOh2t4ZbMQ6JfS7rHB0riDqeep/kdLpUdsqXs
+qz/AWrH4DGCUKWEW5oFtNfbHyTQMBAfp0TIbj+zU3o0D4BZPUoBlmOjhtN+x0ISwH0NRW2rzp+b
vZf2pD6zv08HLCSijIHvcACT4T4DM2C1rwODO8cocj/eyrcWSTnupuGA/wGoPAu6PesCF4F77wKZ
EJ0isrmkT8sEuM/WClqWozh0r7l24CYQ/+gl24Wp22R4jELSbzUJUe7FNM7FK50BQclQoadREGh0
jW7IRRZGrsgEluE0+HHwsVL7TCtIfTyxtIY6c8G62gh2NPFixyZFDRAriMJgd9SdGp9tJzkO25a9
sy+yRcB9EFQ85DA2lY9d1y3C/tp/FkhTO5ypylGz2mkM4T1qb47caC5WY+NTQnw18yD7udNSWlpy
LF6M6wG4J+nbHmcKypJRFbQj7ItEXhB+Y8zOJp/AG6CZHTdEE9RvCfSZQV6xxNaBOJJwSAkECnLd
zu+FKhn4B5Oc+Z2MxfKilSDPqiGdKBFRntrVYkyCfxDW03rAuTX28zDwWjkNZtNi4y4iWIZwWcOn
kUrsgHKF84NImLC/4fgdWqshDEsdA21840YhaojAJKQtuDcrTwAvOFIs3RtjrmrhrB4kf4GKrBgJ
/5NZ0tMi2lx9UtztuGeksETq3sshbbDA6qS8LHKT8ksL0qZjqKw7qM14huFcBN6JKJwP1Q3sOra1
KvS5pDqvCuivNGXYS/beYcEjetCHyt0rfGAvXU9IPrp4WMlHkk03fN+nKD3s71bC9FOcm7J42DIc
FRjJnINNtKIVqUyXQq5ubRS7GJN03rgtCRcIZy389c9vD6BIU8q4hqHCdswLVXNCmhxodX8hbOjw
xLDzz1ndks5Ew4gbjYcLihYQurpNf/T0i7D0/9WzzuDAVEUaZxBjjvwQaSoJwk4bJ2ApUcF0gqS1
s3JhI+J78JgzMTNF6Xi7+5KX2Uo8QJRaSsZkeb58QyC5C5kCFUVT1DUWuJpdtEpm6q/4WXxVBgcW
BCN9LV+DC/hexQuDiAJNE4rIQ7iL836t5fzPyN2sw8QcvGDIZ34Ip+cbJK39Sgpw5dyQsuKC3f/n
XkokciWn6qYYY7LEIzLB4IwJl3qYFROWR0BoLty1CSuMA+EzGblz4rmhUfYgN03bo5eOt+HdlKP0
XDFXpy2b97UBjJDup04NdiG3rEQWtiTzcRQsWsVeGCuJ9vC6IPPclMemNEIw4AD8HzSEtAEqpwDx
HIDiU2/F4Of1cKpBbYNSGKf1laXT7zqUTdX/YMKk3HkWOHF3UhMHChSngi54ghA5+lyJ4UjyLeRs
6ekWg3wwP26Irf3BXDPieodIenhT4A8suNzSR3FKHHhHdEVezFMNO9hp+T/F7paFuJNzS20/TSC1
rf718r5CY8IVwKaETl+7Sn6xU4w9c63cFNt65mjBv3+Ui00TxhhlI/O/N6ENoo73o91Xjl/v7ug8
cRVa/3+hjFRa+c6JetZokSm0rOGVUwvndUfWj23/Nu80HnDnSp5eqI4nLOf6GEswhWscMzrhLSGN
ZERJ/cLMuVFUynVYJ9zQLG7QH9X32VgRqK5Xkw0BM0mv7P+gBHa4OQG/TeEL8b8nk2IBnVUJBR+U
l57RCj+9CzZFPcLSXb/f/+Y3Tp/NCIL7guw168MWqvTET1YVO4UzliR8bZoYUaHSlqCDqF5aEYmz
j8UeWlA1tS8vycPn3BRM9II2rfcR19r/s2vDePf0ae9ExWI32/L7WukdbeVLuyLSsSVoVNuUxV6a
mHVg+IyYHi5N/XsM4NRggGZnkt61SVRXYDNZP2KqZBcYEOHGm5pKtflK33k5ml6jWPPLV8rZ2Od1
NYqx+5vnsNK+oE3oH/IaPDK6KizCTbBph6C5R1drTCDMaOvLvbLHHz3LQg9eEccTic3RMyaGqunc
MhgJKehRuj9BQBLpOR4Qw8O2nxJ4mzXEB7UyUVb5N3XFTfex5P5U5dvDBlErUhR9q/WGQ+DliSWS
nfnjCpyO8b23wjtl8ALAcTkNfJ6Zx5m506KXFFzg9lCd/cfpkOhwmIOCYTFxMHsq6HBxZDcd/ZQA
/d+v9bWU8bPJ6vrXRJkKUau5yajNrZACVvhnXqpon65ZdecncInLM02KHz7DUZFuh9ccknbiD6bX
Lygr/LDMVyrkTDnj+HvhqPci00u9RPV1FBYloVMmaKrjs6qOPdy8vWZ+4gvURyQ9d+Taw7S9DRro
Z+8riNVE9ZOxjuyloPFJp4cTsa9JVh/gz7g4Pwjgk0NA2gIVDT8PjJu3YP+JSRm0C3CbYT1QHuW/
12jlA7iR21V+C6hf3/KY3CJuotY1SsYfMLRnN2vg3PndkwvgwSF8uGMPTTlHpbrKPYbkmT1g+OLR
AUBFmUDieAlDB5d0k9sCXjaeusYKSeN6/7iaI0TFEciuZrpz21JQLnUNykm7hZRm2fjFkl+yr6Xm
eLrkU+BWne8k9xYsRqpjUTNAaAmkOCe4LGZXgJ3kE3lPUw5ImrENjN5UsFmtkDPnWD3iI5js+taP
xGjJO0ePYOaR/eVCQ6wyP5sXQv2SSX6IVTdtdvWHxmnNSst1Szfweq8pvu+VodLygsEh4A5mPLkW
hqWqhuEELdkqQsm3VXMM0KqtcxDC7hSm5LzX+c7aS1y5viWna1Io+4BvSpmfLenf04Ta/lnJL6XS
NyJkY3pxsjgFIcSJNt5hFOF481vtbC0zUrfh+Pm9cXASXCxg6O+O9XQcC1DReH0JPgfgmp7IoLr9
g63MO/JxpEgqDuP8yagkdhYAaV26ibPWkUwTfRAa7tJMWdXmgKxWz8RG58qTFHUeziPkUbcs4Hmw
QrT869dC7uJryho3jouRTyAnu1X9KdWjJl1yYSuvwrEnmAalXNteTUpEfG5+IbH3oC5S/pRDlJ8Y
Y/wJkx/QQiEkQ2WCvtQ/IBCoqiwU1vm9Ziw3iIKXuU98364aQVGw2OdxNC57Ipc2CGTpKWwAeAly
PKWSDtgd4Kp0TeexGZPxrkRAFaeE9zdx2TycPsiTOg0Av1s3AdOUsxOg2vRExjR//yDxzIDZrUVG
HNok4w2MVwW/IlEFnzxXGDShF99U8IUV2DSKFAaGkgeX3zOD29k/sJDPgS/UYScpl7sm4k7qYUWy
Q4R4cC+XvNkF0xaZD0LwoAefh8hvF1mqz0exGcl3j5EZE9c83reaDe4EC6DdHmHkXYBCq7NEUWhl
pQsdoYTXYcDhc8MY18sxGyorDNSzKf1O9vAORhSakUfPW0IJxBO3daJFOE59oKteustXH9WLABGy
mekOpqJ5yvdjUakxVom1PcobPtJb+ocjuTtgqYMq6Rro5yWLcXTK/fTM7Uo6/Bm2ud81kvkWJvi6
yGNv7Tev6S9vjmy/ETU8HSrw3sKmBmN+e85H0xKpwBMDQiD6RtEOgeHL93Tunv9ursFzCTo+LB91
/pNVFVfd9NaD5AVJu2OBKs5o3LJGusQKcx7GL7Zhucocki+a1uZBs1W7QAYhP/ycsoT8gawg1yfp
vE8t8KyQZg8fPUmXyZHHkIaoOV3R4kGiWDcXpL0C34pt+7HpK6f/8E+tJEL7bUsaQesXPwwl1DDV
CAHJRgPfxDGGJGcBnkc2ufRkIQtcDWCyQFqyIuN3lJkgW1tzbslck3s/jw0wJQYzYohdYfKiHdAC
hKD2YZ1JIkF067NrKtiEh55zjwVnweH3PDNeqyrkwxfrngFjPfclw0zEWKAtxIgPnxpeJ6euwAoW
JCscA5oYMvcvjcbj4H2GwUq4d15GYRK5YRX6Fri2CkRfUfoDpkacWVSEBaqldzn8TK1Km07VrMD2
+K7DfjWG3CjJGcnle0KNQaJUNWWWWZan+rUPQbWZB7pPM8YsQ0Y7wykB82cVsNGHOYr/j+Z4U/3a
dlqh4dDUGj9Jn8UYUBoWl5nxyHq2BAk22c06eP2U3pds2k5r6Yu3XTgdHHdf28iJTtSdDFmup1mT
T4dFapFb+hL2D8zPG/bRWTiIGB/X8cjwtllAUdoMHHhQg9B4QLeGSuJsSr+3Ow2wCESD6X0cgiMT
Ju/2+/QFVC7rWN5sFBuFTA/XGZ608F51k8LwyGsPBMA5gpRf+sulYTKhimxuLBtR+nujNLG8aWhP
WeMaTEwlhP47rMtmBLocmHihPtqpch4AS58OQUQDWqUtUBZw5RSb8aIg6NCF3mgC4aziG9RTM6+D
bsUH1VDpfsq2SZRC1IKi6ldhffU3aPRw8RJchA074cMKmdsvNHkWqXyHReehNb1kyuFs91U2VKJW
hxXZSJe/+zrt9+poaMp5zIdhb3f2VDXENb7elAluf3wgH6G1nL0vWM4C4Jr6k743MN+xOl77yurj
nbLAOK8wI6iJwCzlK3Xg9CruZ6EfIzrNsGa8cqe/kW42cMEV5VEAjQfE1qHesX9peI7LnDTn70r8
vTQJTOKclRFrrddawwBHLZ2/m7ziJlx0Bj2xjcP0CH0s1DWCh5pzHE7CuVnjTITJu+yZ285+yEOF
mq2CcvJwIv2t7WytJjxXHUZtn/DupurVZFUs0azGvrrS6RabUeh264BJAFvxNL3d4b9+emPboavm
8QADH632VedJoZTLdQjyDa0MpJUngvOwjQo6iHuBxiZDnfV8rw8o8SKw2HxdcOD+pPkOBqmXDLdO
49IqfAmjW3Vc1JaS4daalfZc21/dZOpBXXzMCaFN9w/MvAkxcVMjcEchmdWoqnltaE149BusgEwI
mutjxWXpLORyy/mIo7seqDnAtr4TyAvcbAIZHhIAn0MQRA7lkLv0hNJnXF3LPlzke7s84nLRa6DO
7Y7LaovbLrqaDjC0ifZpu/Pye3ADi5/n0pTQOJxyrS2wbNjxLNqAD6/oP0pVbBFK2/LeKNBBZ7fu
6O44tubGZ4ae5XS3d0Kia0Pkb7gN/cSupxHc8rzD5HuVLCBdbhUR1vWjcU7uAEiKlRqqgNC8kaAS
bWrgnIhCTJ17nHGbvHBRtb2CpTIqb5kC0k8FlvHT2aMFM/qgy6tcFxT0uZTZclt7Vupr2BD8imIe
iN5XxPx1XPM57jcFTmojxnlCxRg8C2AfSe/7B5jBLLgSCQ4PDdQwRRgHqnXN9kFNjogUuTs2T7Hz
mIEn3vJsA4L8l7TIThcwQiH2rWPto11QIOb0KnZbG0jOQF749YKGavblTIQJv4Y5yOlHuMCrbFxQ
Bo6JHuZrqWCqzV9/BhGlY3ihkkmSusKFZ5FlMawtyUVX27ekNjezvjVz/lPEmlcASYCDSTrCNZXn
DfOo4meJCQ09bxfo/I7celYq/NkevW25y9FqsP2/Brx2KLlurfDeCCO+cmFVs9SyMPpqiae2rKgu
noxythyoYkxzL8zjx9l1nB24aDUJt/1+DSjIVwLE1JU4u1cqdfc3q1Rxstkat33aFB0KjaSxXTLb
jrfaH0jN/+SoC01Rms9nfU9R2R6kraoW1R9JnKmaoiYry4jgOUE1hQmocUKqFJU2wIbR0q+qZ4u+
3tMcpRnwhh9Pz0GI974WqCcKw1JDLsbG5I4W8sIypFLtRKxwDYfJ/oK8MIJnQVduj81EiC7/QXHw
1TmS7jvpqF8VVWy4QChFnmycW10zrviF/6+ip2lBpcc8eQXq/ZxqR9n+IA+GXzx6CjBzbk0pbrE2
7RJIlGGClEb++UUcdzn8yRuhRH7fpT0QVVSVy08AWTM00mLVpQNhL8uzmZNjZsrFnMm4Zo+apWvg
GLsCT4S5yQ0jfQCn0wZwYDbXYtomu7/h/lmTrivjnS57BzWcaxBP8kpjboM9xDKN2DH842DYG9yV
vrlqPZwtL24sK1XZrAh7SZwDq8YWhQtutfiia8rjqE7aoS+//z+u9feXrEmJzlw4r0oW+9pN+at+
6jl5WdJoe0yWHpx5kFZtdr9y8oHBngLjjv9LJcpt2xpiukQwVMtE41hH4NR4pkc100ALtmDDy4B+
nNirUpQB9cDIbwwhRJzQy+xRR8zLfBvHnqOWTUAaZhtuYdOmoEibvKdBYK92SjEYl/z5F5bWUwYo
mtUCPzBjV7KF1mYEZ/SFn8r0JdA9mNln1u+1yzMGXReUIbxmpPSgPi/XH9FWppqwfRAfh2QbMhmB
B5Fj50ICblY5gEYelat8IJCLNXnWZ8T6COhLR7JLTqgTHii8Hqe3b3Z57YCG5/YfMucL/++ClybB
nz9otnp/AoGvidWxIedmlGw1DZSXFQQzKdRnp4bWkYyYAff/IcZo9j4XCs5PAztrGmx6ND8OWLOL
hj2OxbdTUcJHNeye/iecLwDzE1tjytcNk/slueHb1meQ6Z0APDdE5DrERwXryk9qP71f18JIM5Lx
2quc5RfpiUc6K0h3gaFbbV53YbYBX6okr2q0BS7fy7ru5ENNCgMNrFclxDOjVck2n+B24G5TX4tN
tSAQYsYXGPuDHD7ngfR1G1dkswzitqYRZKT3kSh8MyUCj3Eez1VwqSt81n1y6pIT7dE6341+mGXY
U7qmahfNlt11+s9zgt4S2Iayu8eTf1jdwKECkjWhIwuZs4nn4FqGzOAunmzNxt6qL50bP1tJKCmF
7OxIN3vhVU9dWy6xjxU2dkv+B7tpqb6xsO6rEPcuDHttyc/rb47jDRmWBm+BFj8rHqGI3W2xHUfR
Xns7VXO0gu+ZjumX/2VAnML5wh1HMbTN3Kr7+51clGHmLZKPDIG09/DCNyhqE7kEdVA3av1TUvrT
Mk2uiM4bwydlZO+Pb+vmY7H3oy6yuf+91gq/AUflTzek1DkXg2sG5+eZM1XJzKR00P1x0Up04b3F
oa+736suITcxYvQp5+0cN/asgHY5+WcxjNwBjYxy9EkLoK511F9VNfeqeP0gnq4H+xxICIYCb9fQ
/IxOKuFFnPPsofEPY4kBmj3Lw3wGzuybxAJP5XWz7o6hQP+b1iEN1ATQwcVa4r5nO9AsBr9IBRCa
+R+zYyj3xtaqRFClwe98EDza5CeIPaEKc5/zhejDubO88FYMe7fGcsUGMdSRWAOlcQCSleMsuHHp
bKah+W8kFzuRcEu6Ez/a581dqRVOfL59TpS8MbMVnhDECecdJvjAcwr7WUFnyPiTdPi0znxVq5L2
rpMUBdYU54mgmUg9VQWF76Mq5vywW7FWWxEoyeHDTa6m9RhcQHNwPtZDAiPpEaCOQkKIAj6X42+g
RvjpYjboU+CVZqiAH1rMtj73ieWm1DSFZpvb5OWKUDns89KFruYK7lBSgru7Xv5NMzdUzHh/saUI
RanTQxReM4Hm+Brj+H0NxaOaWdmSL74K+2umB4hQFBGgOWi+NEIejKj7kbHlr56QnsXGfCAjdFKC
bBd+PnFSSoF9cHm/YrI5vdeBTtIcR4668Iqsj1Wv93D+yPKuvTckiL771bNgYJH51nohgaVNtbgg
XGMrrq7Lv6EA4hexrKEGdGMeQNzfAiEm8kJYCUzwEeoCCJUC4Z5zJXdEPOagxdmrVdjs681oP9An
Ic2e+twHZ7PKttmhWSHgyude5GJRfmdiswk6jxcczYdZCQodGhI4q+oH3R9o+OyIvIJr1ct//Rml
b0nJ/O+Vv+rEkUX70QTN5MNDLNHwhwriZdx/SdhcLIrDaUDt6c0pYh4skjDNbPsxlp6YrFDPERb6
HvSJ00bhfKxA1C/tiG3IZPZOZR4gsvFuQRZXUPQr3I4s4+GqTUBKbGMS7jS6amF40byYWu0KCw9a
U5Kng86HV2IZPDC10w6dlGf+e/t0WOsLG2aGbbb036ldLJbnAclb9NOe/62C0EJPmMTwBNU/jFHp
UT8jAKtw7mzcjo4HoVQvagh+an7JCSXNCrs/uByUQ6XQj/2MgqNi/E+U8oTMmBfvitv7/3xfOsVg
4WiJf5noAhY9O2pLmRWAq2OiL6o0mpj/4f+HjzK4611hNYq/RQkf+k/BPx803+w8M0T1DogfvhXM
bn2qZGHpSmoVgislcYlo9WdUU9TKrNtTWSkk9cSjOoCO9FyCiYwLvdcSV4VP5/xOYvZmWEXjNnE1
w+dC31FgSHzlAzDGVfOar4Xf8j8two7xMyvXpjm941Hfh48tD7jwawAvTUhCRHLYKW0iseY4MUsr
BM0GK2/jHqG2XKzp8LsZKmmMXCFxqnJMGrSA0SWHUSvQIxgmcJJcsBAQeGh/4dDWDEhtOB9ixEO7
BVXaxppOOyG20iGiyTPq7JALwFGPi2oe/xGKEELbYry8yszZr+vajbxgFHCGnLyKWceSCWz37+2c
um2eDmgPTixIA8m5TBIrd0c7iYIZHGddA2rKW4pWlJjpFgmDBCqrRXEv3VPd5fyG+t8JsMiwHvq3
UXh615soR7MAphctMPQ0M5jmM7wMRitvrfFpUh2EE8eCGmicN1em5dILm7JXntbARg5ivdVzGyFZ
W7Qi1t3CLPdSBYz+FC0YDtH+b+lpaKYnUjy19ZSLA2m02ed1595OCwZ0Gkhgr7YUnd2+mpdiNvKs
5caz4wZRVXLdD1TIz4kPdh7H+NLUNdfdNVcQyU9OYINc2GqH62ngPb8r5tm9VUqA6d3XWNKhi46S
KqrgeuIcUAcxU9zi6eXynSdvTlava1G9r2nqU2yTwTrUWUhs1sRE78bkYxTQa/cTqlvHwNlXj4AN
DRfrNtWMuahHyelI8lsi+rzj5sf2fN6ssV7Hj0I/Pdg3SDj4Fa3MuIfEGXh/nNe/bUfjWWliqkVn
5KpkUQdCVdQg8kf9oQwhecXBjCqlHkWVjgwhrjvOwii2FkzAPctgCq+DvTZH064RiO0Po5k16KBI
MA4vsXYu/lDi6udt5N8c7A7rp0DGOBRKUa6Obw1qpwHsvHO7mmBn1+xSbTY83zWLJTApvZFS0flQ
tkbeyxmWQ4Gu0emYUcdtKMJHbBWvjDc3Nf+YHl4OnYrAlQrGbe00hmLePELR4WnLk26s1P5XROPi
IxLpaQKsUECDLHvsJHPxjbJ6cJE2AQ0sGF9ucxhyDtO73mwwpbKfKuWleT7SJQaXsL0uvODA+RT/
oqbZO5QWrcns3aIVqH6e1V1gOHTND6IEc4G/NZE19oPYCu+HNlOLgzcw2dX7hyRSlJDZYo/mQZrM
WlK5OsKp8/1bDogfUHJOO0pLGE9KIiYar2LcbYVHB+17o7gLtgKtNhAEOnxPHoiFBTD4dqaY5Uzc
5J3xEcuhtqlU/k7MORvKpQyAvFl07bpO6fRhvMB12j1A73pJVJTBtyLnmNSwMoKWFE1qEI1JqUMn
YGlNYXTm760e8AgtxcdTkwJNt3QuhxJCQ2ObhMdqeAeiADbJsj1jdin0jeqIqxg8KSTFfTomCBLh
XxhlJl36Cro31PmxaweppPVCIBRklDiKq773Mn0Gk0Zuq/FViW5/LnaeTJsq6vg71l32slnV777D
Ip2JD/CC89sZl0JuxOYVzfuQAg9wHcdcodBSb9QxhlrxnVkIy+JZMAZA1iMSvl/hBA2fPHTVuyAY
luJuo/wwu9Si4GSjoJLzOXl4hG4FjpqskOZhu22QS/8TmhbMTykMW4mVBj13PfNkhNDsVxOTHrR2
xrh4u8WuyKx9M1teFD5C3gyC+QOA7v9+qEviKNwdy1yPjPJDY30PHSrTKE9WJlpQrFra+eGA9aDG
83tGum4rkt4BKEv3dLpPA7HtxknPaMCDJ2uLvIMkXSXHVLfXDq/9A8v31TvFp5qaDSjHUE2yXfkf
5zXxjKTqbSnWeqT8CHfNgrCW2dugSzEvSbxtyRH2OqvLULvTWxM52JjsMv8Up2xmWOrkI1qp2d8O
USIAYqciVXrNiKYM7+cJILjNdoVtmnInqDNIkEWPj1CWx/UtjBoa/ldwB0N8/lWUdlY+CnnJOeBs
fDWcb3oDthiLrb7qvuNIfggwrF7CHsg2wNhH/W+IFxmd8/qC0IVT97Jly1h9pDtoq6Xg9C9Uf9qz
6Q92euiCWuWhxE5if5Oft29L5eayqt4J3V+a1gH8bMAfrIwBVThpIucgaYMJEe3wFmiZrfzdxBLR
e3X74biUGcBAHJU1/VCsYQybiwCLwueKLCN2qT4w7zPhYZSBowc/ob36512FcZlwWN1Z3X00WTFs
xljAwEB9l/p5m8SOWA93NQkp9IHOrDqyPcyvSEHCJekm1YX7njU6emDb1YnURUgUtBjEGzNUboWQ
aC3qsYYX2SI8ssHL6wnvwQ04We5AX7ZUvvu9fxjOyLxtBBokSAyQkIp28KwGE6Zxr4Zde+Kxscy1
c05vVi2KHjIxFcx2AI0JHP0Dh1ofrFppFb8S0/RScZGF7vyz6MJ0pEne/ooXVGRB/Qi6ESdKWZ+D
ihqFBEtACFrz1flaBADp46LEVAjy4x8Jluc5HUtW2xmQorUN2IbwG0OTaMMphzAUbnjly/zXYg6M
NbVbgCDQdVA9gJV4src1ZyPcW2b9eLD8vW2xgkIQRJf7fRQ+y6GoaHO3i4UTLFX57+aC3OLXhNy9
uwetH9H44IAtr8HWyy/Xo72CDR9tAVywMroAp7OtcOOJp/viLDBIrZF6oN0liUNGJ5FrJBgpwsUR
OgqyZDrQV8BQ9PxDIa3mB/fgawuQOuyZWSq/XADOsQ+mPSzWtU7T6K2StyYz72rkm5HhimirwGyU
26IEewfI+J+GEwU0DfZEd0zQrT3SlQcw+97uQPtcpvcwTeoRR6MlyTzhNf4jE+Jyx4Ye5ypBiLQP
Xqlv0UJFgnNsHYmhFFuMwBCXSjqg/uEX1qrSUmTI2L9aTFga/Y31XaF7bdVE2ZGY3q4QSwPCPsBz
ARsIacsBd1+MFrCXdk40GKrlN+KWqzQrGP5xjXJBvbq69v6WmdsrB/97VJAfx2mx57zFeY+Vi3mF
wzhfQj81IhR51eGEOu9NKA8i18MZ/7YT9U5FOarO2gjPVMPmc634scF9FvdPYS2w1Uw7Vxn1B7LM
bz3aMsMAjJzy5htkrFYYHdPfl7aikSwAdxWb73vgi9mzhO4mAGWELNgI8VJB5GCbCahfPXlex5jB
q4HbPh+m2u1SFN7RRLH/NIGM3JHTbPy6C8CsP7wZRv755LABq5WpRe7T0V0641K3MTkAF26mn+uP
/SMGXBS+U83cvphE/YhbB+JRGfeyzp+m5veooTKuOGUaE0Zxxe35ZDvX438mVBdwYphB8bSUOCDA
LPu49sdTcHFvYMcn8saBxr8CFWOD01y6Pvobjudacy68IxAlBlkOBse85BqGsezqJqB1/m8iCOIP
iAM7WeOOxOYIwPhEphe6yu4ocNcDWXrS4cQVu18tOo6qMPILf9Y6PIAZLHZ2mzSu15+CkqEljWF0
ZS7mU+nng+akNi8H42NJeO1U9IRekUGzNzqtYSOdhEvWLTPjO8XwNML+omcGJKijz7+YJeOuqap6
Ph4LsCeq1TeATZGmmkggNxx6dGwo66dZXwPYaRO5Z1itPU/lXmT2q8R3uqNU/nHiu1YU5O6407gY
gbjUERYq7cy66GKMwnjtGjx/TAEeGEomvYPmzCNayZxjVHHDtRON3PmUKdtNCA6aWscYjanssNJW
w7Shoug66zgyL4QKVHgh9daCCbS878dLI356quhFQh6UvtqXHbaJVvWpfdEktRHQeJlOfB1vfLFw
HCSgVJqcb72K7+Xw2ak4xsvIU8xvjWMZrvKK9wViMcucI+NbxyMTgkLIE5HLyn+kTuRK50YD+aFh
0RejjNgLuov3rg0WqTHR02Oo9v46UPITMWhZZmGr03HB5MdmCycjdD85EHAwKDHIW4nXAGPAkZzm
49c7QifvDuBevZv5ml0IMt3rh/wf29PMlCk0phdUKN3VIMX210HwuGcpUUvf0G3Bk4J6IWy5bD/W
d1O+EvnGA55IehsRnQAaFEENDPt0Ag0SnkLjW1UkIFU/g05NH6dMIgHaIoOAl/BTNnuyHWF9LyBn
Pd1JqVnh4vs9f5xiUKyU0AFyXCdcOBUpZU72FJLx+y770JieiCviD1DvjYfLTy82HKT8dQzxsGcA
PQ1jU/pLROWFo22V7hUno0ekjjRNrtvzFSKW7R/DPqYEeyTnjZLZdjy5qQZ3aEwA0c9XovfaPK+g
MtbviDV2sDncLrGfjnPvsAlAiE5+EPZyNF6eAOMbq1rD8lZh8IRVRNPe877s5ZlXWq3pdJwh03cm
BxgxJP2Ko6HeTSUDYhFx1yP22DZAFkAK7CCbjKD/I6ESsYtnF6IvePAV9IPMrx4+VXk8Y4f4emP8
FolGqqwWrj9sLcCn5+6tERpJgPcJvcsr5bqI5YmBVrf5gccw3q3vC4pV8XEq6ImeULKE2s1fTjBp
nrEkGhCXJJcjrlzky3I6S1bwGaoBOLwjrXeE0CFk4odee2gS1Ksyc7IBZovJw/+sF0nmvgI/I4LR
vtt0hEjGDSLLTlVWMP7a1obXRRVbYdHMlye2/T59MzvrBTyn09+S0kwWF2CHN7X2pg2rafAzOypN
5VMnHEThLmSLZlC62m79E92tcvbL4/9vYLLItfQInSM4mWpD4hMCAXd+UZlElbu1nNgIVXzcScBZ
BjbElPvvMdzeV9SW4g7z/Ba5DpMy6YKfyWOphLa4EWDwYcz05qtunDF7Ej5odHsXE3hUMQbBWd8p
xaMbFPrMw01F+Fu8wJuO8Pa/V3CX8PZsJjwnM+aOImFT/b23y4ZjqGcKnmrv1pwhvKLzUc+khBRY
ZKMn2Bmw7I/aeao3Rncw9TVFmisYpobDJ9q5/VXcJqW/GBN+dzrOehuJo+VOVfcMYWzrDN1tj88j
ySsuZsT8huLr2eN4KYnrmBfqXaE0TxlWOdCZj2T2CBjNI3LPAe8pObcdlcjTeXPcwGvshEaRC1zs
HZN2fEhJPmQkNRKk1WJWwbwf3HkWcmBFTW0MbH7MnZZOKQd0X29CcAFtDa1QEo0ZocvKUtjB8df6
8hPnAnj4b4UUI31OLFqvW47+ED2VV2etlXwABV1uoGAaLribooiYGJrluZNtoHLGBmx5mosF7jIV
UmYKFAY6hA7iFQW6d0bfsEk+zOGiBgZLOKN1t7jPOM7zAzPla5SHB/u6MIxoC3hMg92c3amgPeR4
AaWqlHzJbBpi1Jm6jJkl9YG9cr121oZStG18uPihPRYExJxXN4sXDSsXeXpvJGz0G9K6pohohm38
pZ71fo8ZrXKSRP3pwqH5ddvQpTDCa2CzlnV/e2rl/51TUc4AElJrJxvT/QhoCHpDy1M7pQFscxah
6uwZrvs5b5+nhYIaim2XV9maJ6X9U0ZJ6dj1xIeNDQHmYHIZ/BGF0Q4MdS965cY7bWP1C6sP/mVR
NmmqpJd0Hek/CJfnKE7jpeblcmag/yTQhqBxIyaVNnx+nEf8mZTcHC25j3Q/gzHNlycsZCRHSnkG
ir+qBHLT7YlBE3tsAkCTgAO0pbDi4hRPwoHpO6WUlrIpywA52zzuWf7qWjVTQpOLYg1Gx0tf4eEw
keg5O24LkPMLvEsIE7DpEIgiC2S+kkMpuhcgRSSnrlHld20+OMFn+O8YMWLK433Cm83VqwWfYrck
/vpjRbcX0kxuJISO+Ur5jxUb4FuI8plxSisCR6y20KdK5IHEkavAE9WemyxEGAYUQPxVy+SOoBSf
hljqdRZSQZQ2BhSrFgP0SkgH5qU1mXWNF2J2oaOwlC4MLXlpEn1KJI7TfLaJHPqZ54HQ/hwsEWkc
ViTftyFwS9KDDTIF3a+mNwA9Ue9wCOHypTK58qNT5KCKg6Om21nFQwh5ee29YVia7r8RGXLqxuGc
l74htcSPJoU0zow2DrM/LoYV1mqfZ6fCOdWISVtNgzX2S6yL3ebjj6EJY+QG/6fMZtM/IcCWqswG
SeDA6Ie5PTUvim6rDHRE8AK2OVKUrwriEh8eJr8lKCXJI2xgkUA36DQn01SAJ/hvurbKOUhr6YjQ
9XLDsNeqks0+BoRBQzlT2r5ENUyNN3tiN6bTQRHmLF2gL8/7/KSdzEsKH72Z4XXe99I3brI9bald
L2qKDaHW2rvvjl2KnCQm5CH3uGtiCdSUnT1d9KGrWq3hop7rQJ4EqPUd3EpxLPgN3BlgHIr381V9
kTJlP1tI0fERn0IDNhX7tLU0dPGyAlTsjPKQ8fuXMnha0ojFJ8wupBQ8YqsvnZaP9NtYwqPfn7+n
hjLRrqv2xlKGcnrIAbFVcLBInD3XovaDgZWKXzq42r+odE52gpEC3Kx80jCL3Q4danTmfql97jAN
c30r4M9OMbbbkZIXcZjOjM39IOFZsND1t0MVfDHxGfm1ZmYWI2KzkI6R40QmHQNVurSi81AYMp1d
luOIV6LJSAfbnfehVyxOjYdsG1OMM7nh/xJj8EtNoDs1tn4H9v8MD0b62fvnRHuC662uY00QoUHv
RFZapT+Q8OtXu9pZR733pFIn2ffFi4SRirj0WBIunNggb+SK92uFFP6DxsoRBpN4ZgOMblmsyVlP
k9CDQKki8FhoXWM6qhYVJJF93n+5l5kuWxecnIHRjxLoikRsmyNHaKhMzpEe+CmqNwLyxFPeaQL+
BUazVwiWr2GqH813ppv/x7TsqtV30Pc14ExJtyVCUp34jqYE/f5F7qNacQ7s0D6UsSCLvoxjxZf5
0VssLLZ/sPFDtn6fOUcSLL+EJ/Un3gYR2AfOs+IQwL2x2Bu3j7BUiRyM3RODUyhvogR78M/RkoGD
bOpCSrTR41xX8Uvui1GKe5iwABX+XFuXR5cf8Oa3V8X+dUmnlkGdVL3VUxVZi3/75Ob4FH4j1bS6
K6OOWD4ooFO0oKp7drWoURfpHVr1rPWazizzlHj7Gckd94cfrwDBqS6HMppI3uD8qcP3DjNJLoCs
zDDo6QiO4UtQJMBfm6kvLmgrQRXKweYSuYX8vAD+/Z/yaeLHKqeXudyHuwHN3fpDwcbVbkqsBFTg
GlFdh7UuIoOhjGdY9ueCAuit2syKu1jJDg28tKt9rSobY59pC7jjZoZBuiC8018JeReg5sPxAxfG
BxC0xSGM2hGLrFGtDKVcoyYOUHnThsw7ftLCXWq71YafM+3x0sCGsCjd8KxmpRnSLsRXqX4QLlds
LOlpSQUH6XcD8P4i4i0rxN2+nCwOl/9x5vZ9BZKlAB1VCtkASnFm+8KzCjWBLWyspvjGI3BwI2qB
HIjr7IPOOsrfYYJfa0CCrgh3L0t9hdU6Nei+UV0qDnGwISJIIlg4xJa8vzqn+wR1UOhoLmx6Fe27
RFWfrEuh5FgY7Hi7Vx1SSJcOonmajHMmZisRx+imPnzDcshwg6mWWFZSmVqK31tVrhHPc1KSRc/S
X8/+7BSxKc2R57P5DkoUB7rT0EM/eyCBKZeCuc96t8vam0FGjum+D4Au46H7FKfxDjNU+2NDniwo
ObvhP7gZ9Mh/GzKpj53HPJ9CKNuLgPRAPAifwNNYubUQ8dK8KwBmY5XJbwYP0CC4j8KGiStxV6H5
Xz6hiHzrR2TOyAwk1fhnFDS/pQq/SdYfutH3uEA47+XMEHvwDIzp3gZHQ2SGsYkUAU2BsX+vNqV2
dEhWz3dpCCGyisU51znHH5PbaYmJ5XBaHA6SAZxdsP6gNf0beSY7VY22oYH1gvuC3RXudGgl9yjO
DB5vK9rRkllgN2NPhvKow4cZzw/DtnHbL+qeW7mFUobSixKbegplWY+/kbdPxdhG8COIIHKStUD8
r6n1hgiQQGUO2BM2yToMHVWeY+LZvt8UIWgSd8f7ojpFmbrWI92YMAZQ+qY/BouZe5C6kbxeHASm
g3eLdaUnh1g/KXAi9ZAlUjfXCRq5WTWpQQoDR6UaN+ZzIYvvMErK8KEYSqnDRPgF9bZAzEeI3us7
Eu5D9tWsDO7/XXlSRfD8ruvAT9NkEbNB7h/cYdSlIEl8P1kb2TloF1u+lftD6Vt2SWqpAHZ2xk19
FeRnHZduluS4bOWnZM62Pb022s0eTZvv/FA7EazzLnls5wQ6wV39I4+dIgNTeeYEJIdxLg0rdudZ
AJfxvVTGJtjHdYfjzX3WZallWEh9AHmbBNW/x0PGgmplhPg8Ynwi+ryeVjHP+CYUX57UgBi26k30
+4R+R0rRyqxSeomt4OlpWIqbimfwua4tQtu/iQNCG8hU43r3KxmgO05lkxGeyAXOEi0KfvurWysN
B1GNl2ILSdTILXpYXXKawZVYsywKYAyh0oYWcilQpeAn64K5NJtyLyf3LqHU7Y7zjz37ttSvpJDo
FHHkfYnprB8hFDrla8wFu2sVZFjeOu9Fr2+toVX0W7XUHdwncx86rqmEDQFQAEpjCaH315MWb/xv
SSbbhJQNJLaLF4p3Z8SNTZnWHE2oJdRNRiXn5OPoq5qTMegub48LtcKni5Qerk19RzOoDP+Dn72a
6ejOcodXu0rTGrtD76usPD1WemINpckTC3pTeZkgbYZpADbSW1aWG+wUzQGYh41ODEmMw5ZVTezL
92hQ3LifGPuhCDDlPdkLsp1uJ1+8jgr8y3m9PS9nXlAYuK2CrkK2SM2RiFKTNvE0Ea+SQQnMxEch
phtPIBDc9JQF2VHiFlotysdg9uG9IJfCpWUrajEhdI/k64TmZIXxfjsyORJyR1RrknTMg3SJa8aY
UqLqVzJe4m2+o6lsxQ+0xf9Akp28BWnZJ/d/ViMDsIF4bONSdcpOENaK6KXbpbFzijPqSjDhgerF
f9BaF8xlWCvgt4ZmJCdxe72xVAyKjOcfls4f7oGSn+ouKsMxz1XRRX8Si173zTcnU7OEg6apSS9G
PkOw5EGIXcPaB0OL9D2dK5beOg7nBABNJxnBSjKRO4W3BOEIY6afnaMZfiTe7wGr1W83ctVMjr4D
X1ICdeSO35zYVAPJRpePCd01gkEwCJeQN6+mLHaEr0mncZ6fVPlEoLfmrQXf0sO5SmaNJaUPDYXO
vS6oWHQe5jQitqA5bmodsxSYNBzmlWRQAOZ8lVZ6zf+gC8u55k6wNgZlwPebmWGF9vdv6VIzpHBU
Wcbp+4PNXGGOf4bLhlcYBTYVwlV74H0fEH+os/uwr5uPxtA5Po+XGQatydLw+WfpnR70woV43bOf
tC6NcSZfgGMggdsi4HBNaowYRR/IEKb7aix85ODqkqWLMiHGborH7Rdci58KwBX+S28itzwwNDPb
RFa/iJO3MoRN+FScF974VaXpV7Do/lVPPLwbpbQJL+tWEXzeW4waRe0qnzhJ0r+JvSMPkGCAVucm
UhtHrWu857LDONDKflsSNcIjo+t9nAoAU1PhcRJWkjPH3ngMpKuypVZXIMI/mAISAlDDZp92/hu6
CG+oSj+f2cZAFda6LC4Eo/A2vNx+KALlRDw0jtheVG5FcHweY4CL/GNm41OZ6ESn8dhhnwL1J1n9
bMUo7RPqCPPcifyY5NLNcsQYRsuoYuqwDlMdkv/uSivN/DcmxQp4KMKSKmzYfQ2Bt89L63z/Ro0Y
Ua0MhQLbWx1u+XTe67WyWvKvD2IhlcSL100+9SUZbUPhzO7xta2Ryot3vsYM6i6JuP4haQep5fa9
bDemfdSJ6HWqRLKMJ2vcF+UlvRKipDdOS3h8kDbZSihR4huZnD0YKA6YGrPlXlflaplgGjY0l4WG
egAHIZXUzu1qRK7g3M9JNY/X6kSJbTRim1Tq2A9evZ/bYHgDxL+xsguxfkLRP+UAcO6cNy6Vf6Qj
qO5DMUuJYiSRSzHWaLaUvBxlI1YLY1FyFz7E0BKpt3mZD5dcBhnO430HrAr5dlMXOKYMlpKg1B5z
U56kKD5jGY3lZzXJVC2YCM6esuPHN/Z/mx5dBJh9iMg5r5cF/ZCnNxfYJCuih4jMIRgBG66FbmCs
ujz1OLWF/6XfrliveRCpITmuyS1ieLy03jRMdZKxBfX4V4bcuTUgTHIjE+JfxeameHWnQ/WGpFSY
fNMnpCh68xeirS+ozlV7WT2eQGcAJYdLwfKAis4N8Vl6dCprtPpfAdCh8nQ4QmJpCzCSzc5zenBg
ht64Qm0SJkyoLi5kER9rDGFkvd7J94wZnGNbuvBFAchMnUlQTpw9cYeKgpyHar8TtFmzqk2d4pHr
SGJUrw6N0yYO0Igv4Gy+/Nu+LdpBDEQrvVC7jSmbNooFFX61/S41icOPKLJSWFa3996dGc81XU2i
balV7xxe6zDybXexAK8N5fiYP7TnBSeK0voSwwJyk6vrp7s8kdSCz3+c0BPeOmQ9LH0njuxY7Xcj
ooifxS1wUEjm5DSe8zCux8pIlxhIbQjlmZ6HG/3Sp4qQ2PYl4hE6z+dIcZv5KvrfNjvxaRMQ9U0D
o3+AlgXkeFmEowBCtNGHXa/XgJ/wJ6ruSQY//eua/uoyIHQrks3Ivz03XSpxbzxucTXEpVTJkVll
8cItmYyYCGMdF6t2znjdTBSW2666GZCnG3D2Biq110F93y5mkKSKyyUr1f+y25Ha+TxI6yizBUNn
4Z2RpC/grjO8rMMnBbmrrbSog9lb3Cm7L5w6gN5KRfmO06ZqpXDpLAogh2uf2X2nLdo9bS0EoRIF
IetL31KbO90F/OIz8RJU3CAJnnYuUjfKFBQK3a5gLX4XXBslnP71d6W+o6RWcLCKek/qTDLuB33B
JmlcXc2G5Z6V3RNnD3OSNNqu4TQ0FqB9EcW3gbKlGRVMziLo9e0z5J0c7lTE5xtRXtQWwVqcQhPq
gajearTPVNcjwcAGus1/RNKUa3mx5K8yQ4+DiHPv4upMRfkc0c8Gcly3X0nxR4M2ZoKHhA1m4V7g
Xc6Ol1rs5V/oxYiybjvR3/2Fx/zc6NDctpkMrdo6g/cAdLqf43mFNZxbit249CMKIR4ph30zkJNt
Zah+n5LNvoE3rcaK/KL4Ls/bc7f35MfIR5cMxUhm84XBWL5lezi+1zMnRhKT+ytpWoGHUbHMOcow
3IcjWoKE1r3aipKoa5LPYrj+qEnXJVcd0HUBRmJ5txlWFPwe1QOZ5TR5fDx2WKkYkAMY8MYFWO5D
ZDYOIbXrKjdJHmWvPcC2WWbWcg8kMJpEvEKPf0J2vkwYzTiFCXTA/iIvLv+UwhtruE3Dw59dYXMn
8n7FZZeWykOM1oBlz3onqPvo0tqJpd83r/pb1qW2cf5nIrEBgTQfb0erC28uOWUGIV9Xjk1lQtUs
c+Ya1P7psVX1Od/HnkYQqO17SFNSjPsRdx1RboWSVEUwnHwlj5xdfOgTE0Cm8slqRj620ciKjc/w
p8p4Z0ty14mBow9b/9RMOiLx/jNjIBGs4hYVS1sIf91MWt6e3Kda30fu2ek6zeqZuQSzzABEzMKy
AGIkNEmbjOmQIj2CgOzHh3D7XxBqTlndbGsQYiJKrxeitG7NFqODf4IXxFQGZbfnqqiLd52vkugu
lWzoyELP7sN9ItT356CviJr1XNv8cDjEigoQWTdwUDMhjZoCEKkBzLvBnmPYJhPZEHMRp1jWj8Wp
3c/b4LRREdH7/hEX2+4GtxuqG8Zf7VgFImrIMhm4hvbPOtbnA3Ty4NwoNyhTqXCCcPb28Uo1PnuB
UPjL2Nm7k/CwV8bYszzIUGbVGHb1o44bZCGQrEjDqBceEW1unRM2vjGItjprzHx5Mw+WbDkLfTrd
rB34GpoFsqgmzGerMJzD81PR7e1KeghAVLq1sQnHyD/9/D6l6hHkttKL7fJgWhmzCBw8OP20htHl
U/3XGEWRSqy1mChcBv2Q+o68qiHL3h4e51lhxyGZF9IjfF3H5hWVxvi2LgmSpYflI+UzrQL/k2ZU
mgPVTsXLYEVmYUsInJ1OYvXgg1k6mwSbvNkh4S0CiNOjTJy6qzBRDjEFDanWepYV2Eoc9E4kKsxB
y4x/hmlgfHlHZ9S8pVqjiv9GRA5MPcEyaUzDvYvLevneQOKjOShmEXS6vgnp7fxJaYP1ZaZnQWmH
bMSnEequPkqSaT0X9wJl1WBIn6goUta4B7kr3HAkvY1DPzydnHaM+IzehSR2f6EG1IqzlAew2lro
7mLq6ELbQyBnwXk7YcLEMhDnuuZ4kCF8sMRUuMxL6r52HqrsoQm4lHBFoTV6j09cEVQtz4F+joKt
af5s50KNF+YR9xY/RqekSsUhZrm7uSr1sXYgMqiMnQUUj55MqrxjHgvQMjfF4EHzMSkoGdZ3opkX
V5PXEnzAPwGe1J/rmZ/Ri+kDY6d47bYxdqa/lB4l7lZiDC2i4T9bCM/q5lfqjQyx3c3vjfKUyora
vwSB+Ed6S3Q41ntGgASZy8CjwQO8cSxH74EBOCzo3fmJSrvMNwRMoio72ReTpkk9MYbsRQViqwBQ
0r+82v1UiRtd/rq1WH4rmGxWo4tJi6BmiXS/zkQA1P5IyNP1w520xNhfChrvDWDfae0XQ7KOhOAu
ETGQ8gSLKJWI706K/6tJET5ovR3vUfbIZ3sIvX4/L6NdGyMYX2TbTBhsyacz2PU9JHKlQED5Jr03
ct+EObOnUy0PvXE39RzH3YIF1gflsR4F9qNMFgGN6MECw6F4oyEchRTf9G86KtWhFQQ77kJZsSNM
bvCpklDK6EDbKKqvSFpiq2CUvX0C9G2pI7zWo5I4nJ2D7OojXs1LDqqEA4GKGrWSs84bDeSD7RLY
siAe1IVrEJBysWO6uizk1wRJDQ9HUVU5IFcf1EnOp0XQahxMkEkBkNdKT8Bez//u0B2yVqa4MGuu
OHv+kQB9Ca//aIlUMt5VUIw52m/kZYbEZmNyZsndw9WtBzIu+nIEBUNNtOUeiqvnhYE9B+D646jx
JpzHAiRQW3RLch5ViHNq2Z5mhXYv/TOscI1awcUyOhGY+DiUXCa9IHrlD4yXBWvd+MoRiKP+sVaR
iWlw6RbcXrvX7vLw+HV/4FXUAKxrsavwHQ1tuAHOjH5wWp/7FLwAPLUuqCQjESwLjd/tTFgKO+3H
9lcoFegSkZAj1dh9Svo732HISnUshESiq38prxBqHElQmYTcBXKQ4zzr+Hr9j60xGxNwagW8nE3l
C7HYml+4BkrrgaLgTxTDP8c9wWIEGUmxgottn/W4lM0Bktm/0c9ooYJv//s8o5JYDSlnYqvtI+nf
A+BTvZYtsLyZhRamJyYkhE2BzfhDU+6yZ+/21dXJih6KThdRjU/oToGLQy7pGJpV35sjbKihVxMA
2QbLECvOYuqK/aeExgfCTXpriIgQ3caf3nweFX5qlHILM5A38cVIgeFIt4mi6WneFiy0JCpN8XMk
7jRop6kvh6magtytREebQjFTZZqCfgKRRHgrwsLO6WZ0wNnBwXnNt885VPbZANT/Jz5IsfxX0XvQ
hQF690P3dDe+464cc6Pe29OnD6SIRaGS51ssB197UrQ5EE1GZuPcfBj9uYboI+mOqLMS74dy3/+8
Cb75R8gxGc6qRlGyrIQ+fZXF0brCJcPd7pbnalRgJhdhS7+U4gVvL8bLJYBy4ghx7kwCw5VbAteh
j+Wwe1V4BGeMA/FPP9k4e3Gend0xDCwqpL8TmWR2w9viRNKN73d+Y7rDCr0GkV2D5isef7B8uCi3
1jJW9boyUTZnu0PHttSHSQszTCYih2+a8G03D4kUG3IljnhWZd0PzgMxEdsY7Z5qbXSsWOCo6577
83A1t6mVhYvQc7QVcSJPPnpypCa/tkZ5EF2i9lCIzfefHOmadzjBYXFINo2gZyDCMRfwxDKgEHun
ylPsH1Ka/NU+8MVQNb/eHh5T9yooxdqdAu+z5BCfLRYfpplSg/nrxW9+hOrkPQHTXS40ha0Jt+zi
U9hyAXCKyidA/bGxbbe+59Y7TZFVCTT1683hHVv9VOCj2eGczShrMADxdBsA9YT6Ggw5vaZ97tAv
tcedh+Jt2RtFh/M0KZ77iAFL8eqFP6tYqfBgvV/PQcsNFCqAkoKjfyQ3RUbCpQpaVBhVGI7WcTPx
WthIkq5rmeqqHiq7FyzbI2TKsloFDRgc6VWpXv9OuWiQmv0tPotI8rCZJHN5kHikGel+r1m8KYtX
9srM28zp/sV2qSyEcO1EInG66rO04VqUQtrhDeVq3MI+ondqIjXHYcbT9TRE2j5x9Muvdo1gofmH
fo7ue09tGTxpPcQz7mbsyd4aMdLlFKF7rkXtTJpP2ieT1SBdGEuxWWnYQ/q98wVZ9dzT1W2CR3AD
vvPgYlXOuxKHS0ZPU1JqRTunUVIbxBsIChItSHJWnLNzC4WZUBB/ujSTlKhMhDJZ0NyOjcEwEuw1
js5jmfYBuK77Xsmiy8lHRNWDoOrX5SNboIFi/fwATojvYB7l82QX7rN4W1E66cMYyJGP2mTbnP8C
m24s9OgAiZ+ez/9BQNoUOvmTjkbU3W1c+4SuJQ9E7NqlDKPO11mqVdZa+B8cu/VPs88rg1n7bviH
CvknnHYTxWAu2MNuZy0BfgoqSvL3gmKY7lj2eU/LOS5PNEfA8nv/RUuGMPTuwaQlf7m/HySYn583
Krv+kYz8xGOAVoAwFiSx3c042P+OO9Nu3PjmQyC4k+cMjHt+eMe6eWzwvC/6Cy4verPluyhF3iB8
hTspW4KkbnEKNpuJ5C606kNMn0fn+0x8Me0kuu8q0c+3uoSEodgsrbrhcC1U3k2FvEw7se0JH8Hw
Ng8UEg1gXUuAXSfB1/d6Kxh2WTHIT97WE339y8JXfan6peXi6UuRlfkvcQY+BQK1RZKpQOBLi7Sd
eSbIE3K9W+eBKo+pD4vCVNSMN5Jw5Cf+aHzbAFwBAN7wL3ddDeADTphadabrskmpJxjy/C8iRRKz
7yv/22d0EBNxaKHPJf8ja4LFLFYd5zSmlk08rbr64PZQrmqSQGTlrDPa61n555oqWxang+81CgK7
mJgq6JituO3W5Q+dtzz75aglgxFuHMzvt0qf7WX/32H3QkBqPrVo0nAWKTVRr68vM5wL49nwZMo+
1eyJ/hXq3gMYSG/2lo/JWkoPgY/EK/kmexRxTzfJHX7h0RRuxJWozwexno3yQjuzPohKLwsvagUd
ubi2YZ7UBi+BEBkFdbxDsHMYfCjvEvjBHK6pRppGh1lfCdCWPl7YNI2ZeaabRf5TEtJRiZ2QCVxL
bE7akwCjCL2W/iuyghPYbUTuFF+7qgJtgJnVqL3XTmXXvbio/OvUGxodKkHIuRMnhsbgAmUPWmYj
7qiulTbqCTDcD4fb5HAfZdLaPWkTkx439xg/tCLF4YKvRliOqZhX/DSgRvT8SR6znLE6fIOAncK/
UiKGOYgO5+xJ8GT/qIqefln8YuNw3uDgzFjfeugBkXuvqKqF9+VhOtFoIlTnBpA2KcUfX0a1s8Gw
tI5SilpByvBeLmj0LxIZ5iksM2yuM7zZ0A6CzZ2+qx9Xs0cc8VIlr7tiKE65CVhFTbNaMezAWP4q
yO+QSCrr91zYWCkJ7MRaSkkELaIwmPXAXMo8JWBxZ16tDb3emq60fVfNibVNM8fIECkafc/R7tms
SOD3eUW+GLqnXQQCKAiPj1pVQoD7PxbKZAOuor6a34cLJfLTVEB/Bq9TzcDDogK7I0eDUL2G3ywy
6WXau7DrKf2BU30B9jIdQKhJPdljzT+RkuhWKXa5wRdPtxxaAIV+L3PwVxFI08781CoEZAUq23fE
U0Hc8vmBlVU3A6/cF97F/l6Yp+fuKOZ9cmtJ+Tiyxcm9e9z3Bc631PvDr6EDtgcYNV3trHzE/6pp
/X/tbmTbaQ2KlfOOXCPlWAQm/HH2X2OMxXtGFfELnnN0DU2oCyEYniZk4ZIXI0GWOdY/zB7wHyNW
Db1fOe/rajtwa+Iw1LpyVJ66mEJV2L6oHJGKajsH/z5FNnf+14jXMQ3enZjBsUIljBXW5M0m5YMw
QWGjlCmn5fr5EcBkpUKtctfsRsmZX1FnN5Gvv9bFPrKfACPKLzPAzvG1qOLDLpdaA7CfWMLtaeno
bwsR0QSueh4ErbmvuNcV2D588MD3SAYwSZKpu8+u+L9XqHc/7ATdHjhdIokGQnoKYbfNJKBLVd+Q
ZtrK1XyairgTeEIZLm/0c6eKOUT/2wLt93QiOQN3ioG5HMJ1JgcWqXOFiAymQVnecTrk3DbhYP7x
yZO+/WIU40Sk/D4zm51kb24fg3iE7Zt5sUB90ce0G3IT08tGcc6osdJ196sMK/OWGb30ijxBr8Xh
n6Z5xHYdjRY+1vhfgiLrzSXuoME73AOeROarNHlwfSVnPcdfzpkRs2xhNOnIgcTSF+nbiZddpIhN
WjyytBbt28/jJWIG3iBYaTrltfZarGCm7q2mXOvQb3s23F/nkXPYXth4XliBLYnixjFKT97S6X3b
Qe7MVFfx3vyVuc3XhbCa0xqE8bSqdimX9+wLTJM9iUsj/pyWPiL0n4UoLo3H+O9KZ7kDDmNeAQGd
kt6sym9Mwhp5ed/R9y77jBdvUEVsPfxtUecObXwdtcwq6jNgHc4qQPkhidQyacK5iRpH7mgN4aDB
dgip+9euDgbXu4GjmS2rA1GjjxFpoI3hdzwZuj47BlO7Qd6LQxqzSNzHGaDNDQ3llgiKl2W+S5jh
wlLyc1oWjDcGcRvI84i5xB55ql6p2ef+H6xFiZGac7N+kqz7omiOI6vr6Iy752x+NZXXFKQBovZE
doMuoTGaIacc6UuckkRAhlIAudBRfOKboF1jZQiK3JN4UGq+V3hkyvLLv5v1AxNht3cdHx+5Rt+u
orpwx+q5qmW0HJ1WsZmIYb/TAdc89T8Ef13j7FNsInMQl9XHAibkJ7h+7MCNGue00Lk1ODj/Iowx
0Cidje6XR39YWZ1kszkQTlNZERkEYGv5SClFu5t1wqxKcGGDV2z+3jqohitOf5JQ8pFhDWVq/lFI
nC63Q0rJ07ANQIrJ8q83g19BoGt7SvT0c3Y7+XWNEmydilT1Aw8HEHUf20Jl5eQR53FvK8tFM0nO
HqFohZJkY/4FlfT07WzuLCqv2pgWavSWvtX/iwMhkSjeXTai4smDKztxMrzLcKdOw++aa/cvOPpB
h6fkgLzbmUXC0qBFa9/st+Mq/lyxkIj8kvWwP6hWLjcaTpmktbh9PN/e1oZEceLKCrwdog7Gt1bl
/ktkepVUumpoLFh1gNNyFusUAxSVsy8sw1BaVLrUYuLendxqSRws2l2M9F1AmZvhDrSbOlf6s/ej
iJjbljA8Savt6bKr4BjhaGlT7K0NCD7+lri7F0u/xClVdlOrAhVfQrC8H5CAHuC2jAS6OQXaGCPi
lt6dPECxcBwJDcxOskjC5GWkFNC+p/2YLWySJVx3j0N5tS70E2VfDpchC5JzTUtN4BVL45DpQJc2
R4TFnWYm7QNjYOBr3COHhhy6p6uyh4KVsLXwjtE847vxqYJlpBE8jerZ2B3UqcJJhm9iAXl2PmSh
zdBydQWcVWGbKUI1bRfy9juBRuwby6cocsBgXNZv4w01wF72H95MH+qskcxPEH6IUN4L+M0u+P6f
zNynJEs0gnT3X81knZ3+F5l8ERCMdoTFQegsnz8tDgY/MJZWIe6Z4QKU+tN3IHa344r6B3eyQnze
/WZyG4yUA8+POP/e2rtDAZ0UnIYWWY35l6/qS9CESK0Ig53J7IMrgdT8B1YqpmCMkDJ0re1AbnTJ
ZTsAFRGGPx8VXmF858XUPdGPgoNscPFbFp2AFyps6jf53H8UGHjjChc0nP7tonKT7iAaAX1yJfq3
AK63g6gTTms6lWb11eivci0ps80IPpdB4r5oRXAfYFFzbxbDMLhvHDnrK18VmVUgrHlrdVdu7T+c
3gYMYRx9n17K1im/bmJ8LKheiubY4ceb9vADyrksE2cc/rBu/dtQIOxKsIN8WYMP13KzvY9dO0zw
9/jyuzetxMa83p+G9CbKzF+tjY2e0K8DAzFOCO4AbDVNydY4f+o7WU/ozlqwwOi8/cqpiEA7+qjl
BzdhPxxNm9YZV4OP556ByGryjOjAEGXTp0QUW2pD34DZDoxJzUHwjYB+tEyP9PMGtNcWdmuv7Ra7
OzgXsXr1XnWDHQxSGw6IJ5JDRBRonVJVPXQG/uK+34o0JZzBgK7tgBPBAqWdZuR5CIZ/AwddS0RT
WsalJThJbcwkZQzXMfJJLUnEstKC0do83Tysr+NRKJnPULzSOk3MWtVHKlb02PNzBL63sS2zeD0I
zC0LdlOFzZaThOTTrj4Pue2h9RZJHSkfLYTQlWBggM1Z4O2RFjZyb9jAUZHUytl0XUNr7sDak8Xi
X9HT0PNGbG+OpglL1IeE9jBM8kkhYeryvIgsqz9vZHE/2BZq9g//N9ptr9UUb9p2mmzuT7XbyiEf
aWq+ps32PGqzm90W1udR/083i+OuloahmAzSJb0VzKjjwcJyU1S7xc60e9D9zDh2kpoSdYhAX5v6
CKDetmylgA/MVhGX7KENWzEkLUhggW0Nlntl1FSSdpHukcnp2DwNhqgh9kp276vYG/Z7exs+LziU
mFyRH/HEb/aJwSwuc4VphRklkUULz8/cYp0mqBCtsHS8Om1aei58CcErnnhypZuyrEEa5Dohkh9f
Mz0ZFHbwGh3iQXPP7tQDdTgAPWvrQpZ6SPVkrUdEzGc7sjNYfbHAub5+FREcfqBwZ+qSBd3znpWQ
izSg6TJ2gmEKW+/N11qv0GirsEkk/BJO26DsWeeoHNxYgnwuZmXqbFEDO5hEMxuh4RbQg+gKB80x
9B5Wm9jxutFbS6tcv115ndpqInz28Q6EvI5jKe1ORnNprC94YjPkU46HHw9aRmE8J81gBMdOU1ru
85ae1ZVsjPhvAtX2yUvF0p8gSDdGfUXSlhLT159d1Qzv/EGHGB4k7rIRZQ8xgF5S2kmhexwa3Btn
0l+jGbh2ZRaj3j1GkoQhFWWIGPToZMlizUCpR0rYfUaZc1UUUwzgTq3XJQBCugZSmK9vyW5jwOrN
p6x7A7km7kZp8l+gUu9tHtCL3zJsh3TI0Li9TcLKt4jTzTQ+WslQz/HVdkeSef6ksTkCCxXnY9mJ
1U2b9UU31LzqFOCVL6JEG6OmJwoofhUWE0UY4iL50Txv5rc0mRdvyUK8GcV5rm1hsSURvGoqA/m7
eEKBywf5ezAYeaGcthnMaTlG2Sl2KCqOnGdUP0MTlzCyLdRyyUmmjTkoMI3JQDvPNmLWVdJp1lQ7
fPnA9UONA7PJpETEn7yeUgDpk90ag1tOVMv7AUYhO0qJmRmnLcoxxBdedVLNxRY95vpiOT3OcRAA
sOsaTsEtaGdU4uzuVKEq3/Y1GZsMWEWuJ8xVe/uWCi4wotXyQQVd58SMXif1GXPy3JlwRrqDa1uA
yJXlHmAsTV3THBbtDxSTRFTeMXK/wyBrh/TPmtCrfkiJTDlOOtKeL3KIVDm1syWyypNlpoRws5CT
sHVDThI6f4vOGI31MddG4WUA8H6T32JJJ8b8Nh5Mpn/GO/MBaLwpSQh5G912Lr6KRgVdt5yYwih0
2ZXRWPyyrmmS7IWNDk3JojzDTsolmZR64cDtK1/QdZn+laNcHn3fesb/WUgFoNZmz4a/grqeN+EB
6jk8HRh3eaVYTLT8NqDAxKY4u5z/rvlqvY9D8PwyBHUv97GGPsgLTcwqYclCiqFbC5W17cQ5Vee2
feXOa+1pO5vuZ3NKdUmk6tjQ2ZeWprV5iJgYiIC2MFQuyqALp77kdN3y2N+ICPRq03o+wEKcq2Z5
mmf1h49Ioi19LXuBIY1L/DOfERkgMoEs+RBKSdfWu9xiopbugoo4SUBmE9WI85ioxxt6feyrR5YL
WodIjdM+vM2t4SdNiKT7hVMI5L6lb40AMFVnhnaoZO7AOpmP6K+iPqwbr7PRSsaaJ8hNBfgwh9Jf
yGeHEbpSuzuNaqTqvUVDin/VK+tGsGEqYnNC1+gH29QQ5+kZVD7J76toYO9ONlwQe1YYyzBCLonk
o06cSZgPeWPfvXx4vw4RW5G7kc0EbBaHGWYJFrGpjygoyJG/xhIT12b/iNZhQxLcIqyPcnChw2QX
Rwnvewr7LkA3UlRIpfj+GL0L4WlHNL58TrLpcuTgCLu6qq8tlD1att6fdhjC16Vf7THVl5N+EJIq
QgaHZIDuS+ztbXHfMqMFQVmdyS2SQDdYLpYLI+ecrcUDPoEkZhjG4fXyu74TpFEabFg7Gk8Q/fta
FR5DndnBF8/IcaCBKHgsKlX1R0G3tFljngeaDmOCXMHIdV5ZyXBW73ph1xF2bOJr0R5tTIFOWhmV
aeIhW9EpVv2TaKsOlgRV6ezFBex8M9ZfNSTMp08UIfy1XDsHAYAHp8/7cBJMfgEJcHQN6bC3uJtn
M0wIyy+SH17Z7GIlhqWsAku1SsUh3Zkp4MbP30R22bsrbux57isnU4eE1Fe0bp2GGMZi93ahoo7O
iUbCCAujetxLcBnfTxa/4eXtQscrccLAEP3gZEGy6Qznpw7AdeVyTDHqa1PGNbYG+CqANXtyMtHf
/qgBlYUfDAbVtc36sJIlHXyOWKediQ9yj0hyZD4qbCS+7UCBlckatYSqSV+lOZEOBbta3ogUQoTj
5ngnRhE4Iu1MEchBkNyssCFsWA4NCUKLk3lGKJIQ9uHJ5GlSa1EVpBE+IODQG8dOYXAbKItN2J64
NFiodD7HnzZFuGri8MR0m18th9zZWv9GO3i156+cVsKUbtV85ZqN3Wo7MGn38nauLMqcu5BgJpVD
VXNlmqjmKoBWPagIpwPSBf4mQ+0xbO4U7g5J+1ECqsW3syJRPv2foZBWbaEd5jTQ17iXD0WDa9Tl
IfVkH0cmba4FxCTpgUU41Kywci72IhNk1jMHs1lpm08CBI+/mnGGK1fAHk2OXRHxC8mOyux6Tssx
AoG3fJ61uzvrL5q+bI1rBLUQE4/1gZnkpCJDad1t5yBt3Wz/+WvzeSed7eZv4/0FGH6xUTJeMDjr
80YoplOrUpU+bWXjQOatgCvG4pp9Af9n9SqPFiyqcTfuRUqOTGUldoTOZ3SjQ0LyO4JHnJEczCQb
zaoGAtMmoFUYnpd/N5oQ78l3GDIXa1aYyZjvbZs6u08nAN1KZGyOiBXnnqZHDLRbY70ZlAsfodHF
LIQEvP4UT1OGoVCMlp6PXPdWKcG86m+ahJp7awu/Y3r8kZolWQjAOSnyQxO+uC+PJRY+NzQ4azH/
3XfcFBzlQneNIj6bHimDrv76PWxkHxpxFdB9qaIy5aXe2JDFsTasi0LFspyz3fJTWqm7TYIb//OF
iDStZR283YNVUrEdqIjlqvrtg370LCQr2Hc3zt6oTcYQgBNQDq/QM0g2Rme6CCBg4a13FhtluBXg
tuGW3Oi/MU5bmd5tAG04Q8CgRhZTciS/BOBkEakWj5foewnAKVIf90j0/hxEXa46quCYS+ETDwCB
SGPKCgNzhhznYJoY0ZHL3q9x48T/FVDJnnTKYB0HF6VXsBuoq3PbFptkVZDcttqPCTLAFu6w8UU9
rA5k95YAybOSJTBeKJ5oDiLjQjU7PM0wufoHZ5zFJ6ksDb9Hl/qU3EHAwbOBptEiln55UNBAFn5j
VBke7C7acTj4c62cOdRFTCv8EnuFCZtruzOAbOPzNGzvLFIU6tZxU3fQsna5KaBpuUTwcNWjfFeA
iP0Dv6guc8v0Nx4HsszsPQowVQoI5P+lkqn0JUvzIHhtKo5u191gn6ZYZSw12YC6t3QeiK2y0l2m
DEC0GxCF8ucrsIqLY4gRE8lkt1N2LhXVlFGAZCtQLnRByIMb3FIgjD3XECe0jmq4cEcUpgBqHWKI
2q8r8ZHAlKYlAp9wve83uFF1bK4phFPMCmbNwqnTM4fYILg/XIDzCgTJ+OP0Jc+S5Kh++SyddksG
+yC+mZYyWop+c7VD+ksG1Sp0OfOQEyZ7B/nkuv1yS6Fp2e+RLL+em6gskXqHZLzC1m+y9pcbfga3
SQClZoXqfOMqei7W07ITeT0WSQhp5/QoiuCL9LGBWhLXaVcwGJ2TxxhU3g09DEUsb9RNHUwCtkZZ
ombIA7KYo4ATt82eg6vBzBr+LdBNQ7qbZZBCFGeM+vUkLELgVVZTwtXLwg7kr94wHR6KBPqa151k
vW2tdKsVLGbeOv4M2m6TztUE4ExldMLNWw1X4Rzv4w+wO0zgHa3Z/R2FLmVirN7O3ke3Fo9AExR6
B+zBMRSmmt9uxCYp9qs7A/iqVP6egBV3KzWFtGFAy5Y2J/xDos4EtNJtWwzZeXDTIpW5dFgKkUrM
8NKb8MF4MsCeQz6UFEfSRLCjxB50qjXh4Bwo6qbjkAKEexOjTVaW1LKXtm/4J/AwTmzZzBpYFqtW
whTVZCVYJHaRoMh6HkmN8hinPUiAwJi2a/oKTO8cG74MpRT9ZGzVSn8VdM1Kyt7JxCrSxrKFknd/
Y4vPLGojzXaBOoH+IucoqxuxA6WzWokKl0I6wy9DZG83LxAuRI+skDikLdxIU4NSpGwoRjEQDnVy
ooLRgtog8akdG82w/0lxLKIeI8oL3A/YDIwb7B06kEUZ2trqlCRhhmSpk71XKnnUy1/5HL/rSGBu
PmVI4gvxbGcwXODUKH15NmkdtMax7D8AhkImPUOLFy6lbupmFPHXJGSvFWJi3eiUppqOJT4oKS49
oiKQme65YEpeRUcz8VuuiR65hzTtoHI2mT+VJMpb7V2VNqdU4Z/+kjd8AK7JjiQHr5McmhnPn6F1
uB4Zwh8M4P5JFeda3h/+grVA3zwRjMv3JP89ZVXhKXkqoxbst+hauf/ppT8ni+7VVp4vM94Kx0bZ
mooL3Do1W2fqM8FrytszH70tyxOTiPkoaj6Rvvsh9Xv4UcSUR1VtvrOYxBMhsVarQ5GvpVn6KQnR
MKOfLMgONLuAYJP+1a7GpOWJnZcTTRKNxoz9WVH4nZCD/OTdxONd8DPkKPQY+nNWW+D2bfaD7L5m
3N649BTUEnCoMmZRIUFIlLRXT/Ppr8T6UXKX12wrmQ6QSeJ0zi7oQi4BgPTm2N73G7Np6qFQd8g6
NS8EndcwJltbHY1JT0wmS8jbultXTxln4njG0aKBcj94Eg+Blr2YNvsV5Y9D9JlUXYIDvdy174b8
f69X37tK4jpG/dTJcvqQXFUHX6pImQMEFiuCafUOWxboZUyWrwqaP3Yxfr0PR+e4RJyryCpw43DH
bO9Js/EzrR/Db23l7cQMUNnZ//IHlCMnXkQbqSJ+Bkpz+QN6I4zGmTtdURUnBBJG9t9PynABR2YU
FcsCU1BnsfyZkkUjCUNbCUCa5YH2Tyk31WtbDiJ6x971hd2X9vbT7tynULTVBmZz8EOPv8huveFt
7OJlDCqOWMiIL8VYkHIDpOh5dYarvb5YCEqnDKNfAlbvm0bkl92s2fXkeMnJ3sNEjJue14PvYWt8
EIr/jkvGIScE4TTV0ZlsLvNPJB1mbkGWuvfbMsXNqBG1DhZyZJEhjMlDgCXsHNTqNaXep+wg7Z7e
nXRsPZVld04JEGRhWcs4svPrTQj/YdItuahI6vCL+lQy7P3KhxbDQudfEI1FWMb+noYJAAt19gD/
QiSrBW0/FrJWkw/UR6EWbAPgtRzGvO23AGUM///cA9APyV9P4kPp13mU/3YqFnXxC+eh4fAedc+Z
HH8Lfl3uqIjqy9sLrEntnvFhqZaUgaHqI/T3jz2Sa4GDusCOZTqDhEYXnysfXMLZ7bdbAPe+2fqs
6Q4IsNi/lJJD0QwcILRbmK2RFNTJFr1sO6Vg6drtWQlUgfssz4tUunPdtP13qINk3Re+oKyIkXwn
tDJY6EUbIjcfBwtiW/XSpxZx/HF9/Ex8VuoGmqoIC7855GPVE5QgPaVL0krCOG+LObxjMIBGbhaq
cDcondnySFQfrLwJXXlftB3Ng5mRNXHqZ0FXuYIVlSylA1YvKINf4A/rYC991S7HKNNoHuVH2DZK
VR8RRAFZvgV4qoR1GfFaQdz7OQztz2CV9pSUub+8TOpCHwvAQGyRSfpoqqoCayuge8wcukgzA1tW
5afey8x28b3KefWZ6I0pkDESX8P9pL2AVq88b6YEuoARsG6cKrc+aNQGT0ibA+1nPdz9oTZWPMaA
pzB5j4+8+iGBUgBQW6bp55iepIw69rH9apT4iw1efe75frQ84ToAS8ubzX9hdVLc3jW20I9lAClF
YA20NWLBir9mhYrHK8Ahe7yzvgSIAZJpPhhpOVHqf5EM6CDhWswbXge5ZnMjg8sDxe5Dk0VILr+X
6GSRL43qBnvVcdI3Y+EQ655kWt7R157Q9zDKeLiNLYj1QaEeLQRNL69w7IT+L5Fwrq3YnQ8K3+T7
vM4RMlnG3byAGxphx3bdv7wVSRrpxApDW813rHgNhQywzhe7POmIjCeJ/Ezy8aVYE+to6CG46cCx
8xYu9KDFrRPTF1nnOKaediyygBAxmq1RYcyNfCZbfMC3d9Moku+LfaBTGWIunGZ6BjwFDT77VPOE
oNS7iNnX1VZ6FaWtNwpbwtA8WDBb7lYd5VdSr1GfXNx/A3xik17PzjcrRKMfXyxIdOzD2Bzh4Dvw
3qUTL43nxRT47j8VDTCNl+VyzjogdNyvnO7vIkckPqW7tMsVVy09OBQ1Ujznj6MeTuBExfEx40V+
Qah7FEJqexujBaVqTBO0850HCBLs9nwSbx9ryxOMvmIOM26wBb/EapPRpuLyFybw3kzjN0gTZWaz
LuhaAR79RscRomeg3D48apqawNnNQCf9qhLJkpP/JApOz1lkkxEC8QORLUJGYARQaSsJD1Ne5Bjq
OYUGuvTyqMlwSYb6mPjAenxlSkCjreuPbDltWA/q9LGZ4Zkft9gvLzCxjTAbVzSVqQyV8j05Rc1+
SR7EKxBWanLk56zUubgofWbeo9fsV8IFOz4NE7s1Lp0YVQdllmKYkmsPeK7Zxob/a1WjzG7RO+Li
1ebj3GvOZJ3uWjlqW3ai9mMnH8pZvSl19Go37MK9q2fsrnDoS/XcGSYAWDWhgg0+EoKNCudWvi+6
3LJYW2CUA/2p5i9+s3C3ix9lHhYdTE/LT9v4gt8koUHNksqxzpSbTM7YiA9SxJoJMbhiMjAuA+Oq
uRXHXimJ0F1QXW5/IufU3bp/DS8NTC92M0dNs+Sz+BN+BkKxzFF9bZ3SezZdrCn2LpqO0n7YncGF
VLia5KSozDTDELIl80mGEgUSuK5TgIUflkzzZrNT5udqo0QP9qswsBOhcq0wCUujOIEOKj47nq3O
qNvagtDP9/O3/sE9filik9Khr6IBlRiSzK+XpX3JWf3cn8qWOHvzFFo/mtu5Sz6PykzH1MsnAqvr
+AZo3YX2FcsJKHMjXJeNB+MAOCPyUSA5HNvBhln/fqFnRd67EF/mONPHag6qmslxwfLXeWYhNSgS
+0wr7/55WjPPeJJ+p42zxYkuNy34Rqj/of4JZ0gvifI8/g883G7mXmxtxloeTp4svHiSgz4fEoog
Ox0+P1X4OFkgSziXe4TrhDLe0yQbG+RmuB14TDech0sCdYaZFx8N0IRilAGjIVJeZ/oQi1tXlY9U
1WPbe7xVjrDZmbq/TCsEpdbG8o97VVbVA2m17Cq427xbx0G8MKFTod2l9qLjH80AtmgOlI711518
ktOsrxakjv6ENGZN38N1Mla7heAerOph0HwBYzoF2CQVOTSqrf5cwLqezRg7Cj8Js0krrsYvZW6Y
KIOsutbDZrDymiyIfD3Botv/D3XPLw2jEL6oNLPsDzkyrJAjRk2hGaczv09ixDTEfaxzHSygKxXa
lRA4AVVb6OrvJH6TxQmYDu27OjPmHSvWKYdsqlD6jX6Jrf4LUlqXfRjLVzTL+BTlYWq2PYiiIEca
VRzaiAF2XgL0gyjHgX4wyOXDTwh4wll7wC7TIag3XgoC8jxT0dqHW6u8FzBcD0HeFFyKhwH1/Av7
j67OE+kT3B9nBFlXEDdSfhBa9cUeCVVNeugxFUAdIJyvbAiCDZ13dLtSeaeYdiVlIl+qE3DhvQXs
Lwk8d020gdFbzTKKIaUJr3rT60tmJ/qB30mTTWO+zENndSb5V01xjDwC9ndbjeCjlG9Icb2yW2Da
7+VhZiYY+A+4gQZBsAil4kIVqcB7AnjSDj+JlJViB7lCcwgTCMuzvUN3P0oZITGpiAihRYnNtZay
5RkkBF9ahqN39V+a7kNc9TR1c+WUEo2Q426k2T8FV2e85xFr06Y0Ftt0i0a+mkYxYhQI40odF86A
dzUooBsHBxuTnwmXfy/u65sbXpD3wlRjUXCW/y1gH+Z82H1hesYuSUG/AqCwe/EQdfhyP1frnkSr
FzggljjK2YCjD7CTtb7Itwy+GEzLUjFCe2XRDsk0AL5DrzP5mH+g2TUcN9FeLE94N1h33WKfwPkn
XGH6tHFgJ8vIWqGy9a0S1iytfuJ6en5ki3xJKHcMiWAY3yBzlejlAzVEYzcr684mtZMYna5A4nEP
PtPIDEsJzVJbIxS4WWILq0nWRBBu2w+DGWSK5erJHpJI8Ik/C+KlN0I2DY5widSP7Ss6XMfC3UTw
Xs5IDVjT19mSxxKLK8Xq+e/S5lNSEQngDUEvtXBRdocRDcCda9Yo+XkKUdFmcmUtmySPpO3PJgal
WbM/rykV6CQnOlXbLa16epokhGpkLm8byxr+viSC0guuNGlny7monadq74MsW4MWnj/FYn9g+hEc
9tVUTTYA3la7InpeETdbzD3I1P9TFAN6+VL6yuQU2C4zbpQPQnsIBe5+AZUrvyByVY4KZmGQRPTC
jGjwRb7v0DgnvOq5Y0ud0hzM0rR8RF082z4+JoYNhc1Dcmsywk2oJXUNZ3hj6lkq//Q2xCVyfgTM
yMHjXziW3mW3GCxs3o5Zb8oQSTRX+XjRHpuZ1xP2l+X3fH+vHb2dQCTFGSuDjf/WK/UYxLbi9hYh
eUFNegXYfy3FHyYSWSmNtiQ31/XEP6nazMznJe+UCd8lu3XrpwDjIG05wdsTeDOkirhnFSgsYYf9
R+PUFFaMzKLrhe8Up3NG0zfeCEnMT8PkypykSv1zdK8kst7g6n23Z50ASQI+9K0vL3gpKzf7z4M1
9flUsPSwBMNpxvz69Uygp6PR0m9fc/2US8Td0U/YePrYSj2QXr0+tEC8uIoPvfsCCHfZyQKwiLrr
dQwDPIGcuNqCkqLSEQxRN4pBywti4wdYglEzYr+hgrkpbXHfAq5v9GMSqT9WjyTcaiGCYienKxb9
SEuhx+gxRzwpadDqh9XQPStzUkej6dvCkgmYShuvXwQRWVTZqJ0McXpMXK7prozZp1S8m21x2DWz
GGHZK6GcNROLvmEYAvePJeGiLbBw/Y/QgiYuwpGu6qGHN1kQFxkTtI/sDac/lej2lc1vmSgR4lXd
5z3BJ50Hb8gwA6HgZK2L2DyaxyS8J+U5APqsbsw6HylIc8Rr9wKp4H8wIeMVEUruiClM85ccCyT7
6e4W/4kB9j5C+1hnIF+5gasMsHpiZp8QlvDLg1lbwVwbgJcFG+2oy0j8qDQD++Qf+s4bNhqiA4Ce
FLm7h3GczFGMXE9MrOv2IgV7rg6HjhLXowdMQM46njOOe3v/h75AGKQMzCvEUtyaUlQqqT6I2LgA
zthVRF3b1ChxdJA2haylbcdlifxw2yoact2OLjpbiW/18yVmhBYqbZtSXBCxWqLVy8Lb6OY5+hjQ
1GM2sYdBqniSYWKb/5UUT6MW+QRc8lCexLPlAjcJK1k6DuFZSfCbdwbHCeg+w4PoKKaHTzDzkZN0
PKO0VY4rFc5fIQYFjBpFam2xpX2ZoCZRTLJoUmvP4ygq+VaHSYNMtQk0ZpuAUuJnIILhmxh4xl2Q
N1o9aztSnXkLT6Iu4SJc5rovXwy+NZDb3uoJOhR/am4mlrwch7vkCz8S9zsnai2DJrnuuevokup3
ewy8mwe1+X+Y3w+OjrR4Jr+bZzgek/unCqTo3r83w8LLhoZRU81utndlAefJLfdqojh0lgySW1ZE
jggh0gVldcnVVyP7v/6IMZpcKAZog5rcFRNpZ2qiHWVmm4/DuKPvHTiQak8S7jZkssNztgi1E8Fe
ysRBAdZ0p7nM2sffDF7QniAOgDzdGl22MV2b/59gkDPnFcxKqAMNQoaf/iAWeAb2O6jeHagZSPxS
0zlu8imJeL9atBTOgRjXtidUY26kOoNDtY3ldc/g33MsK22ge6mdzqwdyVEesUIJKOr/aWWX0bg4
fku9APSnPigRdoOMX3knZt2kV49tWG85M+at/3i+wqojPqYh7cW5F7mfxvZeqvn4WJ0Kb+9Fv/YH
QAqml/RDafLRNx5kI03LNInX4AH/Q1iqEzdaGrzflXvEJVlMryLreOq7he2499DfzKU5pgZJBVBV
yCp3tHIAYEKm4zr+BfrDmcFAfv8iQFtlcmUbclI3dcSlZVChnN/OqYeJWs+Jxg4p5jn7BW64UwRq
N1uTvFD9tj0jcf3cwuVgfcilzqmV5/K3eGY6yYMrTlu/QQyLFs3O2GKPfB5g29u7Rq1kZ/fqpnBS
imzjFfB8GBcuiLcJZdAQ46Hnxya0zYL+LiMw/g0XHw/EGqx8eg9FkfkGAoU+00Pi+JrfwHpPBY+c
4Izc7xgLGUJJUm6ieki+Hs0b3O5YbnSg/UYyXVPS5Hvx/vvOd99wrKakjwCaHVcD9PzhGYff5GE9
G6lyZzTFQyanhq9BbijmvKmsf8vRdBlJKBFE/58BDOWz8NgaPvtQtuajEnRi+s3sXb6cfj/SwxbX
EKBWua6GyfKkMJqkZSSJS1UmOjj8+XRP25MqJJqaOpbEm8Khluygv9QHUQJ//EeBU3Wy6RF9XlTu
tapZONimVXyVdKoyFGhc2ROJB4Ecv9FfMUHdVfYQIlHQq8IykcF7N90dNrBVHjw6fjMs5OzilvrH
2biJ+6XHv8M4wvglB854h2S5hfmSFUBTYnF9Hx+nDLLWWtYn1qXEYWteqpMZsFYRbrA6TB2ek9Ca
hrDeOOYl1bllIQbOs8j4eru/GKbWuj+hu3sg6heLvT6RVub+KZq8xV8ZXEEOTiurJU6kT0oggOMb
pfUbX4BDWO29tK7AnSCQwm5PAiqQbJswaI/LxUhkyop1Ng4Wb5/4GoqmES8zFsAOs/l+ZpO3Roww
go7DEm/waduObI+ycp6OJux4ggEcgOaxE8Np5aF+wRK+WJ4LKK0KwPLXk1kIXjOdL1yGZLy/lXsv
nVEZo8Nk6SsO7SOc2FI/IJXwKCM9wQvJpWv/CKaP3z3Mn2X4FmhSVjN8yDLhELBJEGbvz/vsOBcC
9ENR1ebBlMk4ypzLZAmwNXT+1fcvXMwBS4lpA8ZY8wrMLiP95zsWwWkRxClxhTQlCwZT2zAL8o/h
diHeZ68WLZZA7+21bn/F6HZZIUpwMr8cTHgsPoxy21NFhPm24WA64BfYpsrmxxbt5HkB3YsDC09v
MBF0Faq+gGtZU8aoFt4F2a26Ebh/BZM+3x/NhjUuY2uW5qmb9I7byhy+6nAiabqsYMoh6/PEeSzM
s0xP/FbRntBAesufBVNCYAIrRMZBKyFPSHlq/hsVm5v9vU8oiQOceVjuTg2mop4LSyk+ER/jpBID
38dyme6NCBulhar1t8uxSpuVPhot1lWpqvCX/vDjCDb/UvTyiU4OAb8cQqOki2SHaNMb0DDB32vm
cSZq2XZ/GJeCIo3Uem55usyrcxlUrtdz8HGoUxLu8BN5d5aiDTu0R2quNwsyTkH/cz0XdZ+6561n
vzZD6yriGxl4W7JW7rKZbqsH5rCKFe7fmGMloF/gUb37JZuZ0rTgoCfszunKoaDSUHU9aoqWGQL/
GWNgSog4d5eGYahJGJ8j1OgJ1OflonX6N9pH55B1yfe/ykyci+F1ZceJ9EChpm8YLVe99qT86qeT
fM5oAE/+GrAYrwPLlScnOIiQS6/XKes5T4oaau9EoRtMFTjc8PWsEazj3vDdOn8/9+H8SbivLXXL
7Xv5dZt0BBfG01zOaG3Q7X26dd/wfj9bi0qhZXREtbkbJr/TCehwvARjOZXFxwuKrC54LCL2xRK2
Q6sXbzrXX6gUeoF2yPDHYn+1DwWuLoJFtCneYQDxkbw7JM47hwaklCSm2f+GOP/ETDwSCH30nAtk
db6ShE6EDZtw6DKB/QbVcKJwmGOFYuVhIqquUthb16yj+WE+EgJexmt+61fCZikGzJ0f3Jn2PpvD
5hAv1uXqSypsiYaxJuFRL7kl8/Z20OjC19koC1dkCVywLUG5CoZfH+vT52M1xf/RY/Qm7KXWMlV+
2H301Ta46djvk5RxXqSrm3pCCfCwZQz4Mxae/Vky+BRJtz1OXtxSwklvAVzcWGfOtGZazJWnXylw
r5We/w7uYq0VKjoo6dmeA9iSg13KO5YnQp8pAxpTU5hmwohjz+AdbEgI3cTYJZZnAc5jJks5ciAA
l6LIid54l5j5dXUI5t+z25mvmgDnEU1pj29aegzLLqHhKbPBtM7WcxJtYjkMHKPCTTUaosWLBMfg
30ziixzY18YHSnQ4YL7s6w9J9PShZq4VVEWFwxMTBM7MWC005KmogaJUw8Af5H+KRnsalb0XCgBb
cMgFO41wJ3c27jfDiwY/smbHmx/ZNpPm5VO+BnNn4+lZJLfnjIMEHTNw83CiZcjO2/RjYjMCkiy9
P6wCz1cgYBQx8u7WeAee5hjuiyPJ0pto5GwljmY7qMna+smFBw4T2WUyqFR97F9LRrl8YKbJG0TM
Pqo72RTxBwGXG4wh5j2g7xnkvj6gewPOZrsPP1s6uABzt9G8k5ey0L6LU1SAo3nk76MeaFePeXTq
mqpSZmQuL+j/5YN5rhT2JW8g4yPHcOTQ3lwys5zAnW8phQVbxCAtfDtGr11ASIjjjfTmzMylQ+5F
78Tvzo9byGJ34Qg2bYgEJBdNSUVbjbzV46Lls/b8A6sLHB4tA+E8NQ2oSBfHW1G4NQD/Rzb8HoLx
e0k/YD4I9gJ0LmM9dmB2Y7xhyzSaGyGYc8iBPLERGPpOgXxqcElcKwejS9XURr28JVtniioCIbUy
4IYOvNHAxJr+MKQaZE72tVWZfme82WatEXZuTjUU758bltsEhPGW7A6h94nWMBpNcyeKhXszwwQG
8z8WKVueBiKyW+FKJbVY1D1W2akCdpGEi3pmY6aS7SzT+Jy9bBttlYzREph9+pQp5edSX5VBOCGG
eMV5Bbp4Y9qFliiJZtBxeohvE78ZjeHPgC45Nvq3JQ1eKC+Iq6rxwbV07oG2AwdotHoeBUeW4Tl6
3z8HyPekyd6bq2aHqFNoE8AQijsW4AcnHHnhqNxHa89HHQ1SRAf02+pxVPZ4o0zf58AuQY8Y5np1
dkJj/cynSTxYoPsb+UbYJ1oKbPps7GK6y9bZvCd2U8fRG/5bEYpDJ7mX7FPLkcdEWQ/GwF+wpRgm
9gAeV8SOn2DRIDiumdUiYOsvtzIjKBkehehmGC1VefI8XAwnhwNhITm3F2oAe/PPVLDTp1uWwXFF
/CVzzsiyUhSe51LEQHGlso4jHD7xSU61pxEsnDJfPe53y6GFNsjDO5XDtyrkJaxMVNDu/2KwyIbw
u7JMUu9NB/9bmBssY7KRH/NRpQIVwVZNy4/UQA3w3AcBWLh/XXXzIdZmzWKsl7kLJEjxnohp+qGg
ruAG+6ZqKQgVLoJzC+hpYVh8HfbTSxYu6U3Obs9rNScCXjeTB4J3W4pbEZyYL2tlSUylC/1ovZHp
H595n+VGg2ELva5o4N3rMdb4+0E9rOhYI7JYFRSsuyCorUmhES9Ggokqnj9kBDVZlh/njWw88aKr
qfxPH20TX0RFoZJpBzed1vRThewhYr+k+MFlTbvy3aLcVZwNf0MMkKSaS2Sho7HI2J24bL3rcLIw
E/pFWE333jxa14n12RPoEN0nfP8shCjxQb1dfkCwqosXiZV22zhKvGgixpIHexZ3s/+NhDBcZOD2
kXlqiOWSgbz98x812yx3AZtB3f4kAeZQJkDRjuqdUJ/uGYPm5yHe82Ubr8UYOR8Vwbza7cFA6L6j
J0xCRHBnJRSFt0UXj6Ad0AxsSSz3zpf6U6l34MfH7diteptX1xVoRQFx22U2SCHhnwlGMLRahR2T
slFDmQy7yWht2/7iUcq5EfR/jy2/fmcMVTFC4RvYO26oOgk5Gw4H7xOMJnZnB/KQo4Rb//P6Soka
XbnvU7lAKl0KJ1oYdJF/LbvkwQw6AMTpNEJpLRYwXKwbb9ndPEiqF2lyJoz9hEv+vxfQejE/iH6a
2TiyBCm3Hqu6OHaRdadRUMPGZ5eMH4fM3SzBl/V7ANAJjoSESmxHS32bF5Ck22iYodPl38y6BYnG
CJBNpBoopUrfW6LvD/2fIx44RXR1dR0d58coSO8F7QHLnLjCW+jfxm0SmLu6xsg5SNuMtgRl0m1p
siZdsbx0yRoRrbugcfDEdRgW0dVcd99RaQ8lbvgCBNub7YlYFMU1t7SlNUIY5YdTXBDoTFeSo673
L2vRDoKGqjtP6SzCnAoqQXDufymuD4Q7HrmO04JPJjqQdigB9nuGAWDsH0dbIffi+JWdK4cnhcub
CtDsWl4Ces7p4mJ3WvW+ka5dEWe5KB59U4nulamei0ugmxQeL8q467ViEyhlcvl+oKz/c1BdVmSV
5gRarEgPBYHWGVWOLLrzTg6nw7SY6g64qGD9tSFsyyMmE7fPNcp9m0ptO3MjQaCmuHYVf1casiZn
3M7fPflSTtMA5kPuFX1rC5cdTwSfTjNVh7zJa6dSQXO2RXrTHJmimWZLs9u2+GKWYiPbd7liVv3E
YyPGVo3Ggx6gf/402t+604RhXrIMC8XVy931idGpDcdCnTGJeXjY22EBu+E5/DRVxvsdjm3WqnUM
c6eyFJEyJw5zmycP0PEIaPSmX8yukObBmFYGBqlt5yg1pFLOukNv/R5fUFCjmZ1hhxkWZBO4GscS
xRP1aXVIv4SWfC3RILcwvtzrrIPtRx5AUlGwW4VglG58E6WIMv+kLbuGFmAbncRx7y4IubTD1ArJ
w6v5eWtBSe3jBLjMPjJ4VfQN2InVJxPLv6ZCWtYWXuENPrzH372YieTMYuoA7PYiJ7wspcxdXHTE
AGf6thDO1PapoHdnJsRFrkLyRGkhoqoTlokX0Gh0dDKnzRQeyGz5X/j3FWHUZiS8ntYFmbzuBtVn
SBtLI/OzYOQ/gR6tQWAzk5oAAxaWfLxNKbvGBIJgusmfuWcY1gqPFxT//tAvXCH3lO+H0TYlr9uI
5B0HwnxvrYJo7iqkiGulXZNtKOy4EEh36K3rGjH+4Re08aRjYS7xlymQMwvhMJFr23rjrse8jOVY
1IdJqEA5l7gxhflSjWC/zrls0OUbPBTm5ufL8UWcEcHUXsiFTxW0+fgpGbm/gfc/o4MmTj/nTRpk
5lYAt9MtVPll2XiC5x4+xcr+R58vFvGr+9eQDCffAxvxIBnX2qmY8uOw4DR7mjbUFkJ2xXo6NQ/y
S0B9F878G1v9EB9nHTi+kqwtE0yJ0b+tjL+SG8lhcYJ9K0PgLGk40ErW0Bz91/k2/NKnILhrMsO/
dV7K60+2O4tbmpGvwd+IKwEHgLUPJtVSOXZIxgq173bxZwXaS90QjmhjdbiZdmAebuAh9n7zpfWs
Stznpg/hI+V7oi35FtIYAZ/MAYfeoreZiXfrHlVlhE22tVkH4ubaU3Xeruk/kLgQHNjOJZw/ph0K
XKfC/migVDakK0UGvH37O/2WTfVERQ0bSs4giNs0VjArB51Z+lLZOjbCIbeFhJrYbyrki64RPlSr
OpyKLZyplbHogOPuy0MVYaWNeialCBL78gnlPC+30l10smHJMmwdf2UMKiSdPWryxbLH2uM4WOvF
4peRN18FuNj5GGtoE2yh3OVzbHu9uRr1xZxPGH71GNi3qa89q0KH0Q0GgvpcFRs4aCxwp5cKi9tK
0Xldl0aa7ew/bji+x9TkbgAmfP5vhtRzfUO6pO0NivXn9cPWB07au+nEhsByQxtWJ/jiDYBihDTK
rWVFzJ4AJVPyvIgLyf6OS7r52N2+pDWat7RyC3Ih0YaAfD4II0MW3gGlsAGFQtoAuteSlAVh7mbD
Tci9/RfEP1ddMmv7KeMKYYy7HqS/Lv50x2xcct1lTAuHsTMav0B+4MdOb8NO/T0d1pYGI9OUB/bQ
asKAulbu3u17f+VN9K2PkX5FmVnpZcxtbqYxp6S40ZqSYXEC9AUSlsoVNxYhXQGZgg9EDoepO0St
7OC8cMrQqVmEln/fwh/1usbZ4Fnohxy7c58OnaErFPBHdY8uKkYCYupq0My5xotDElac+mndKC8+
c0bF2nxy9flFb5CP/6MwW48SyMZObnqHzKOcv9/CfbCcgYqkG+XAzfNy//BcSIcQK35o9739KO0j
ZRpiUDikWUbWY/ee7QoR3GsLHgOSiQgxrF7Xrkbi4CmoDILaQ/DYWwCzLAS7pdKrRRF52eZ/NB5a
6YgMLpvSmaPTJEp9a8LlH5x+we6Yc0t7JPltUdRMiZaKS630hzn8kSTkpcFo4ofUwos1Hi7gt2yF
SknBFG09KvQlRHx+y0ZghWxr0/re0HYg2sbsMZF2nTYc5F16fBW3tMYWDjqvAWGI2C7yO2xYKun7
GxhWhN3Dk+kMRwLtSzX0dg2q2cnPb+vFdULIcP+QP6nLiMuNf/pb9nwleXFtUe/1Bdy2LMG/FBSN
X7ii+hcwHC9EQ+jlhGhudqC0J/ytfSU/7gHdo6Ov2aU5ORvAH+DWmh7VHAIOXB4gDjGCfTAICwlc
hhJPyI0iwzopCx1V1Uh0k97NCKs0t3jqiceywFetQiLLYG7uYz0ZWI6dv1Ddsj3Hr+X2auKufgMt
S3TSMWw0csxDAh0lQhM89HFA3jFcbBVYlo65viT7Kmy7AO3pJELmQnbQ49fwPldYnQCiS7zg6iph
0caxMspN8WLC9Pweu4Lnu8KtZ/bwP/dhFdTUM04rL9n/+6PAYfjJyA0kFO7jYVZbg7/FbT1bAwx0
UHVacuQvdOQiJ0tlScmOacxADobD6Yg0UHjbtKJWAEKUTcxFKdNihGu4oYeTtWepDH1rD99ynCgN
yYnr9c3J9ldOMkL0f5i4A+o0sgHwrWNfawTF7nDmyJnN+MFOsD4zboiIeYAGBzi0uBqS/1T8rMZs
WXBuYOqyrV4+UyBwuGQaGrtdubDbYwtpZNyo2j1wHIwQI2ONom+cfh1JXILa8cvejO8oObqZCi9P
DrtrDFkhdEuCvl1FGL/mpfmenyELwn7HQN0QU19U2Oc50DkAetGYO4OTsrsDuyX1iVL7+1G9BEYc
bLTQK5j5q2g94zpyaz8VdN71UHEPsRbOL22FY+31F5SM2elZa8lstHrwICY5u5YBqgpAwURhLkLy
tdOE4CXssAt152EzXE4tHGRjA+ZTW/DHQVsJX/iMflYIyNsoTifUaJHt02VIkmF9WXrDSYWhdWuV
Radwr+8gAlunlW74Qi5VfuLJT/Iyci5iwSESfSXR/W8AeYGHftwa1EYIqGY5R6/1etkBNimCU0v6
QsScOyZSu3Ixg2+ylz4UiMktlzGyqbaRhiRYuqHkxpA7T2c6GHK41bi/oRCIeLyYTBqmB8cdEJ79
61qOozQVMniKMvrIk5CwdTrPxird1XxafStYI82tB87LKf8a5McFCbsPm3AyglwtTzc/M5Vn4Vsp
p9OuxhR4UPlbngSjvb5YpsOfjVj9vJcEBOsME2cGEl2oYUZP1fWhTBVSECFByKjS7LWFIg1UaCeq
I4Mcj1UKUy2Pz0YhTG3XvxjtzW3Is4G0uOoFg7zKWlBJeAz7lesARJrpBmBSs1QvLx12FIydWk1G
4aBXbbiwIa1Aw4NtQqG0DpGVXCXaAVz/cOYYSvyTMn3xlPb0iMqlm4kMeD0D+AlCI11jL8PlpOPg
2IaVWyql9Q36sBHJ22HQfWDJffbHO3Xx5gKLuHDtrrFPBqxTCfe5Zu/a2pdAqbbRn5+Tv0JGU6v1
yxhhzdqQTAhELexwPCIN7uGLGHtAAUQy4xvR44/+bRqTlHpORcYkIYk/RRpidxoAR0NHdx3JfJ8O
/l8XCqQnaYrv/n+eJY3FqK8XnBbkjs3+hXNlMFZKtgbUDGd4pdNLhJLGytn9WC0SvPck1Ra27NQm
rGBlbReSTrmfGvjtafgw763kpomgQeZ2dOobrLfkVLywKWzurJYfXz7M+w4BUyC+0ygFkCyD3hHo
tRDIti0BymEZCId75GmJv0sKj+tmRf3zs6BrVMPhFtkPFwBZBkqgysuyKyJjJ4Rzkv9HlQn21zeO
YuK+WM97QrkOsJwJyhsh6ZUusB3wgHGmoCsEA77judVCv+AbTFsR3+FMTDLAhE6Ovfh/wHleiwkF
qiGojBiwTjqjhwKv/KeJIDiZAqerXliHfBZSUs1orZfveRE+Vwix+oPx70wNB4yc3I4qjbqArFi4
U8MBY+kQ6G1SFpVz93QsfOd7pjXJwEX5lr7ibzPTgVmIKDevVEJwtcxuufwFUbBqteu9togr6W9/
zp1qvfKbhZNad2x8hJ26+n9iyr43xUh9whhsrrt/TYNSiRK+fbu2+Mog/uC9mau22LlRviVtLx0i
28nk2y2rLnmqXggYoPnk1yUNb/bZIhcBciz+N5yNfqBcap132q8hpldripdH1EynSbKArbBybyiu
18B96BzuyIr0WjnqAI2aN6EPJVLinVJwpm7jCm1ZSVS/bJjuEki3OQaDnfH+PBfsYvCiJ8ODkE2Q
FK/F4B2RRCy0NQp+8nW6YAQjWqAsa29HNkJ+YUIMjN6T8Jz6oo2wjJGjXgSosPHNrQh05bvSq8UO
97FfDm9m+mgbyJXn70BH6GjQgKlXDfIQu0iQYlmkoY5jxRTWBVv7yf8h67VskHHJDzpOho+vF7qo
2mCZ7JPRiNnR7DMmBAOdz84Pl9yDNSeUvo75eXg/a+5x7Bare37Drqe+qY3rrmDKPHxK3/Emx8fK
WkjwufT7FqA6kuvyMWNoSPD7esbF8seWTlK7rDhTgoqmRDfI6rENsON7HGBUe17NOk1uVT5bJ1Td
ogLnXAWsfrNtoJjivsN7y9K3i6d0BwOEcLiBXzolj1p7UnD0+kmbFS2wKVccjNL4ktxGzqQf5kXR
XXFepZmugmzI1mVyeGX4PgX9XmkkRQGAlSBJV1Dp66xhbRHOM8YtYTcsggKdECKopwDuxemD3AeL
ILi+RO0rjuEGgufKSf6amWPHFwQEOG8LID3x9lsBmO4Xt14bSPNNqzg9s2a/GMh2HoyT65Qmm59O
Vvg1VQ3/TEqA/W+SdTknA1kJbYSNhyFh90fUIc4obPzclpW6OxQWKBQiH2taofeQm7q2gW2A8ANa
wUAxDnzFYa/4iqS2j0hFQTBr0OIHQ1MVPKG5zCI03AV0PARjXVs1AqKvxeIdl4JVpsJB2Uq+/d/G
K6DWx4Stjou8VpMGAIrP3A/xOaw74o9QvPL5eFlF8AlDJZqw9j/dOmC879fiWtxDPTz3+1jodmU/
hvNXM3RVhd1kd/MqYncf2/fkKRJP4dRyRzR7BxBX8fp/6rz2nDfqxye1l1LmlL/3yezae4N2quSX
DXW8jAPt/IAUuZTsXrTj/74J6f/gvgAQBhkNSttnGjNMQ8assU+cdYBbffAr+T1cBolVUJcfL9QL
I6tAb/IfPLwQOMGuZPlZdVASQLLpMs3iofCAotMEEaRuFf1/Y5d6m2YSOCIlFujX/mqKcqyFfTWz
lKc0PEJjx9PT3MuOYASj+gmqONGXdtZialBJnbmq8ehFBf4t9tcE07Wo8kEhOESYQbuq+6xSGjP4
LL0TfMVq/sZ5H1KBU0bz+K0sAG9YOfAuGxfntxhbNryx3/NPLMSRzVz0qL00Hvmh8Ms7AWnAcv/r
Y9tQzc6e6F0LVfomZ0JkZHktM7BqQfmq4VIS9EG5BQRMi0vFD3/0oASDrAPypGZ5EPecw6l3Kj4r
CAgxpYGWHpHC1Y4af/8QW2kM+lPuG1DcPFSxrf+MsqGQA+AOYsF7IvLzBpMQhuIarJlHaM//C2RM
P2m2W+Z4LOoSU2LAg5WhYhv1jP/bxSNXLFr9a2slPW5iFsNvm7BUSRCnMfY9ebEGHu9Dwv8pJwxo
QnfxtjHJW4cN+zFHrFu9sUSuhotPu80N1pIujUnfZjJFzfgJQMWLGNrk2vo6N1hR1po23nGIEiz0
QE+2fEshH/BEiwM/AwIzSUsb4DQzdhThDk5DNgq4f4GiVUR0jOrWECIWf+cBc49S+RcDvkE9F/0o
LeGott11+jQxvJNX9u9+otSrKpKvJ56Rp9xHOwnTKCwBHcHX0YZlH3BXPD5fJ0IcOByk2GuzJYra
r+LzSlQwARnZiJ0cvunBqAHaLsk3e16UTSLX3/noHBt9m0SRjAt1BtlbxNVtxGl8K7oLv2sR/wI5
MR/i55G5dBob7lwfulhvanR9TCS1Y1L7Prv5gMEL15eyZeC6zVeE+On8YMN/fJtNHxDe5/HisoUl
7mhnqPoxjTMJmbA/a2KIC8dUuSIoSYS0xMxMBlEKhnX33R7S3VCYCsoABF4XNE5N7paFTvPG7taJ
OVykoEzIrR4uhtxlfIzjrg8Hwqggqdq3ZJ+tJLov2qBg1OxkW5BtLkNq7ktnI/LP7nP2cYDQKJQU
V1oLhSTWc5ly/xTrzd9yW3MPcwgvWIvSLIIq9RdZwR6ONf/XLg9SJgZGCl2uwPRMCGCnM0VyfOy3
VwmBr3SIB+LgraxzjQ9+HoF0kuMJvIdKGjL58bs7fGFhCZjjFhgXMJC400ip6g6+rH37FOG+LbYA
CX1/FS8xc8Nm/NkWbgG/SW8ptBBiEUuFB4fIZomIf1E5GUPZAKaAlf9p51Q9uUfORzHB4SgRs5F7
2yK2gdGEia1grSrZxqvPZtH4SZahQGVKH/2yyhrZMIYMaljbyodfbEfmYMd/mhOKCuWHaU2+W7ty
YkAQ+y339XosF1veqt8BatMOQDsAPySMegcWjLCAmKq6d2GGk3rlPWGWpi8mt+4whP/hxkH99D8n
aousPl7UReukqlm54LMhvIVPx1hlKL/3kWclO/GRt6CvwyaLXgPkkIxIGyKUYn5yoIM2Yc37vOj3
ulP6g3bdYaPfSBy3mBzzL/nBmxR2YY5K2mujgKHwIP+dJGEB4rtWqub5vW2zSJbuvSRFamiOQBOD
cNK4/iNWX0NST9bPtu5m7gIoZKj/7l9KwZYL6ji6BHPwvNG59fZZmkIygcvXto8FNkg8y+DtPKtR
Ej+6IVFz5KL4SXc9F8OSJvFBby3DfDupLPZ4TFCALD4TlIj8k3pZVCYuszfYeu4EK6Jdl2Kr2B69
8u5mdwKYTXXbsJwiFb/pivQaAzXI+pr57REhgAuTLicBPOWSL9JK1vIuwaMBAZ+lWKmt79FEOh+v
eqg27iUHX63SKrKV+sSPeCWQEGbnHbtufBcNeQ5gaAbzmbrzb3zm2Infxi5QLqKGiq2PDScqGnZ1
4/NjvAx8IhTVEk894PPGDXpYiR/+x/3ahbR7SxjfZwU/yMPr9cT55fdPrTvXOsQvKI0yYWFZ/qrC
rytpJt5UUPZTUYlwv657JQmL2j+T1I/fa6W9fcruM1s0GPDNFCLKlsKYIAGNxRqEGJdY1soXdTcb
zUZE19L0zuhQvAPgFxidUkvybn7KqewqxzHv0vCvTIOQoD+a3ofUo8y66lR+iK96zQnvaDFcypDT
8Gpo5i0G5Zk2lDkrPeR/uq1j6bzDDIYvDEFQtaA/KrKs+XedzxFUYJlxHKfJl39W5495VM/cLSU5
NxCibJj51B5FCu6UgNOYNeyNBFF+ryTfRSF/2MScsDevzKg8HYZj7kMfJL+mo5MGzFg2xZ2OYFQS
KjL0jjKbR1Wwvh8So/4Lbu7imQwxRHX+4QpAcOREIhh8xRhCBCHyU4eWZ28li25TfgfEPzIHngdH
lky0hyyXZKnnjYinnVPIvGb2EFUhhjk1jVzZu9FeVbdmzBfQy4NCxtqoVXzRnpBCEmIw+iU/++KN
DzLW91LTFYTgF5LSqmhsgxKVR5i5vpHppnP/7nWESXshAQDQuPqOHJbnpaEeJ4iubFB8YX1SI+iD
Lh6m4s2qQ8tHNhigdl+lnr2SSTpXJm7s7vIip58YkfpqBeQbTOmxJJn4mR2l6CxLNIuWnAnV3VL/
3hy+CFca1XWyTF91OZty1dBaGY2GEC135YxGNRWYHsdjkIXZcnxe4dTHeeGk1IoGqEZ7BDJycPUY
HEz9lJG2oq4LbLIAMPCKpTOotTVLBxAeY5eJaduE1UK2ipv2Fb8IJhtTUNFMH0NNTouSRPSaSx/n
IufrmPRZD/sAFCP7ACniheUHWTBMu/QW1GlwSSfYEzLdvr98J44dgnV/n/AuONLnEmqoH5SKAX6O
lbI4j/ys8sES8dfvwqGSdE4dPLiu7pOQEkOlInHSHPpnetRJpQDcoloGOfwMhLCcyVL97X0hpUDa
714cJS44Mf3ytAkwqfLBGKfsu8SuXnzeEWSIQUtjijSwKE2uVhyou180Ti/YzkiYZ3bp7/nc1Cud
n/IALubYmweV8cWETz1wt6ffWx0t6k+Wd52ChA6JrKCmRvjpclNCQXfzXniT9kHxfTymUTuhkV+B
JXLPDNH+yskGtLhCPqgqH9gtXU0Z8GJw0Y8pTMb1lubK8h53ilsZCbqJaRIgXF7L/NQA1zEHvH38
rIDUvzj1u7atnojknZ0TLL2ijOQwZIJq9AA52IoFIkrkOmcZsx7NxxLTQfIPEOBGg/XFkLVAz5nf
WMR14bcs/Bc5E2Q1j4XXjG5vqWuytQyuf1dXZO0QKB6RvJdRKexxn7nY7+xJ/kOapDBT/dPSiwri
OSNXmdX0bqEJfoX0F4GOoaH+iIp993pl/auZI4iNuAYyCtOa0APBl6pswpXTpwF8o9XdtRYUiwrJ
rgCDPDq5rGuanmbcUz5jkR8cL20rS3ZbfquTYlyv876DwJpYvFCR57RBfVgTYKCp6c5uO8/dbTjc
Csu6g370LJE/6HLFB64OZ076JqCsNT/wRahfqI1vmirflAZioudbZzIwHmrGEpXxEyLiFm07kNf6
jlJesrFTB2tK0GBzlPfUaFZ0NGjG38ergMcuH9e7sUTk4KjYKCTiWJjh5fgHgTP0yRJfOiX3/ho0
j/RdMMXBejxROvJluQ/V7P5fzwNgathOYU15TG4OEUvcd2a6MFrMdFZGok1IC+aeC+eH1qSx7Y7+
utznN7DcgUcri8dbOeFO1vO+kd7nDWlKQ3Eoq+MHEd9lz92AXbaK9QUZW58lT2d4NZb36Y+MSC4K
u+6eYCRPyNboo1E3O3Q9mvAK5Mc7vagSNb2cT1WVvQ0Twbr11aOQWs7e1pokjMVg75oa1uMu44jV
EpgjVOgi7/m26yLBj1H27OW3PrCc9Ookjn9iYL4AnMbc+vW3U4thSm89Wdj3weDT/TTQ1NfkhzPr
jNAk+hu4h27IpgRaVSDgEsJEFMbTgabvQdePJ0AH8jy0HUUfIAVWd+s7OywJ1WtrvA8KqkWQ65x3
N4w1Vb/qjkKMLGaoq5k8H/N7VHDvIUia1eUXjaCT7J9e061r/aHpmgP/XYWsT3gqHB2htTpMWtDu
42vA6W+uAmCukG4tSWggulZqqgWWyqGV11PinGmeqNjKvMnSyrJ0GWa5SX2m0EO0pd3jfCIpc8EN
b4+AitDAYlqLa15BI+2qP5lO2nTK1NT34HsgrLmUOTqYAxWPwVo2abxXOqPaALNxLf8IOM5Psm7R
dpwqBbkpDzmDZgbcgUpxhzBxyBwkRLg1Ea7Z1APnUHG4NmRLRqISVY/DYoCax9rM0o8LtcCLJyWm
kSuylX5zxOU9RRx5Q+d+dJHG2BLHBDPLeUgK71eJQoYvhgv6jfrIZlZtM/dPYO2mXQ+ZwEF54DKC
T7qetmCJZZrdNs120O4yzLbjLscuknNNzRjnpW/bYCyi8/ySUf+gNoMFhBlKwqiLRhzMFs/zRx/F
DhWmpkNDceIDUmbwIeAJiGQ7eTzQfSPcdvzYZ7epIyME0IRKds5tpyL/6bGgDvv5+r3im9ft2ddw
Uz3g91+0n/QiDvGhGGkxKD1a0FlR91Nzj0teTBbEOEuLsrJwjVrfF7A9KstYr6niGasvz9KBBTNQ
d1wa6zGRQMTLllMyauuwg8DL9CHh1ESd+909t9PVZURV8Q/TBsdDBFG6s70KHmonx9dIHQDnjine
rXtFkQBYZVnM2y7CEuFoskLpG2lzkli8wDl+1B2s9xvMa/Vmu6iwe9hD8gSdjIDohFnPh59MgjvK
ZvdJ7PZl4JS01uCgjsmcRaYcsBvAEbJt/JGDUWvtVDhyyBFIDUDuUQVr7lcy6zGxV2kN8bXtaMwu
dd5AEq+48gZtpFEjVNCgeTmoFgZi1AdotC+C7m+SaUD4M1oYzdwaV4kFGF8jg+/jZmF8kDzx+5tp
il3B7q6dPVhnN090IbwE2QrhTiqNWnTcpEftHyfRGMeP4H2dsmKJo8iwQd07i7LiqUGuBLrX2Urq
zdCJq3kUOIkL4V0Yzzq+t7Ftsf8DzV9VIXpto/eadv2vW/M5vH3AsbZIEcW+yr5xex5YQSruTzmM
aThMMLg5ESqD6cbKZLb5bONN3bb2sxwwtV1nhJaOSF3olLl4fT1kULjSZNaUwxNJwHhyJnomRzam
bflbAD0/U86p0sIu7zlS7L2/TSm+lAHMjA0GxF+ahiklIpQ7TxwuKEQaDokFypKoK6hAzD53tL+E
NOzZVg7BNPeO6X9XSrGO7NrwdBwgiwqW6rKB7VRhUo30QUIU8+wOLQ4YOC9tvGdbB4sC/DS5Pkps
TjXiOg+r5RY1NSgogHEXDbQ+qMlqh43bxupotVnkSsacH4AfqI47FayJagxJj1zZjTJyn1e9FYK6
HWCwtQCaNZxWPIizmdrG+dm98QPM4iKG6Pq23S7J4kS3GcCpMs3PWvnZV/DaOLklr5kPn/EOq8Zs
gbEuSc8VDbdJ0XFGothbScx21VtfckhxdAHZyiA4ZiNVpWbD6jGcuEDnFmKeE8lKLuIpdptiHlfB
0/FjAxPt5QADolv+i9d0PbR7DL79wqn68RDCiVqOL3aFEC1pWTdReTDOT1wHDvogg0xTM9iqpxKe
yHQ6rI6C7OK0y3GJnzBC9DjaGnDsebxzWuFiri8sRYwRdu0kReqaPaUqlb2DmmcbLHIxA+Xru1/t
PJ5qLS2DHD336gGJpJwl35BMOH+3FLxobP4slq/cJxsMBRICwToqi1D+NW6d8WlLX2YAlc4d9cPN
AdRAQ46Rf7BbsGLDG7HnwrlVdmuUelUDnd7bRyL17O7skhk5Ia687XRARjRXaYPss4qRAmEAtN2S
J6mnTYtByxVyYwEApXi3vVLthoQPOYNn+fTYTZzqluN61vPQAQdwM2Rz3GsG7jGxB7InNeh7z7B2
IKkrUPLzxwnQbyNAg5f+hL70y8T1Yj1g28hJH/FdNCkDFnaFwO1KiOQ6J1Fug6xdao8lUmMSi6yO
VwjhzJBhzbACwwTJQ8fkWisAcjwgPVpFMBSRBRCsWcmTBrAheK4d9Y5qbpe3Pp24ycx3Pk0z69xn
k1KsZ1cErnyoEItt5y1fN8oq089MAjDDLm7vJSUyZofE+N2hYx1YDecwHRPHzfsGI9/vKNsDiX4B
FrZkelDUNTLlx7MRVBMbHWnkFMc8Tp8RtDj8hX1jySWwRwvBxNV4MjvLIAFS13Klc7vmR4mwf4VE
kiCiBQ3Gu8JnZN44NZwXbGVRpqzd5aMjNJqFKBp2NmzDMNul99qXYlB30WpZ2rfNtn+UAfZEQaDG
sl5vGK2a0+9ZtS+CahPiN5gcLHUDLPqirIGeZR0y2SC7mVvd6nBrGrl7o6uk0JBfxS62HkhCjtox
eXsSzrIBFBhUE6rQ1bRXtCIJMqhrZA4cF60x2PAW2kLQSI2l/DslVu/+IG2Bprpkhli5KQKzdj9p
i3IHasD1V0Karo9B0mt7QYEGON/dmQ1XrLdNKQn4Cd0U+HWuS9iHDVn0BAdLoYNzrAYTdIqfaeQH
8nVhwNygGo8ghEEzN/AQN7j0lToJ+Bat/QJOr9/ocib1pmrlMzn/nu4HIpNLxrgMk27r5IeFYU3q
fSaO8d1emh64S6vIseX8evnFq1qdfNpGnO0i+g4upSt4kdUz2G5fKVIA/Vtyj2ZEjDGldW5kHWkN
qfl+ZffQ3HR7SI88sUcDj1PYHAeGPcyxNKjsSbyKokNpOBOXTPFoQVleWBnGEYzNm5a3PUJ4+unU
ZrIQDkw4Q368a92JRu/lcxJdQe687nB9j6QI0bVC8iOH4NWxXttlOr63uqAuT8yaIkxRecXji9dR
FSMXG60yxg7WBdbNOPYyAwTu/NEpAc3wMhXX+5IOL/33xyr4WgcLYKrjmwyoKp+ZF0KQCBRTPmJi
Y6j1QXICk0WhhP7IwNVbfN8b7xFBl2xAgCkkGphmcUAIQjW1YgqzosXT+cZ23jB7O/K8ALBWRR8D
uBwFypjJ9KArHVpBzpDeWHXfrNTVdlG4jHX9RYsJMY2OTNmOqV0AFZfnTh2W/HoQAEu4wC52PoZ1
9DOTem5mnfz28jh3cBiXrts7sC1LBgkOJL8Rn9/K4uICttm9T7IJXxBDW5P+ElQ4T7oiswHI5q/6
OuGKButoMtG3n7NWy3laKTj//noc9Mf+ZmM/RmCVy01QQylZuP+C61gHUkuSCqRwJLLp18UcyHb5
5xt1CKLsIK3hpvxsgK6yJi3OsoVEmbGm26eIC/LTF4fvcFljqzyD4ngOBzetPjYc3GojCXsuRFoR
e1HSOPAAK6g3LS81QsDhVhor6A5pP/jGdobYNcMx2EixOypsYLUC5qmWr+u4RXQ3HwLSuwWN7j1E
CQIRfHFPwHUl3qgvUn8t7ZE7N9Lpn0Nx76L3xOM4b4PTSzY2QV1jjcdMVJNofO6ivcB4U77jSOAj
u5VL4hvha6Ga1jcOWaXs8sJ1y/kZAI6uBObPtX0RQryMGGfcxkPbcb2oCBdtW5mlGRZ1wZtqn76k
Syi+1+wn+bjcAPXy2rybzZ//5vpBIM75Krd+n2npxt6hTFoZk5UJc4JTMOYZTnevi/iF1+j4le40
b6z9HtlKsqDPQfW15/+hhBZMcYvWmEXF3zqAo4oLBZB1sEbmg58TnCGeOB6xx/o+ujmElxLw4xNZ
ND7BHxo/0+9UKH1nczHk7mBAvOg5QkKlVoM6ooUYtieoOCAEmhbYtlozM87KajJTHPJfzJsGlRM4
MAob37XWDvtCpANIb22Ll6BnQQNP5/GL1B9DczOHR6H4AkZ1MHF+mPv6+jeN6yI4yWrh2Cywb04S
N0gvyrSKtri4NPF4mJCPLFZGefal6AyxVxIj05fa6ZwPnuwscRMeptuYjEtp1oD6uW3RP9rPxVBO
21bi5o9AyXxqXLjHoRjJo+JBlSJOcj692zeBDZy6dklVlbjZz/c8oSWZfL7gGtE9jcBRM7vKtZCN
JEg0GjZ5aL/sB0lbtFcsCjRthE69C29L9zczgFcBT5QG2cqnXZ5kSL0kgoW5sU14swMoVqXwEDDk
nWAEO6mfM3M0eWIFrJpf3ECjI8N+UTXliNSguCmvdYVvhPofUvWMh0kZOm0MXgBs0mx59SKioJ0y
RRgbKBGkQPOEk6cnRcCBZafGqq1+Ts4aTIsTVJmc/q1ytxsCC1/N546Jgp5Yp6Vrnhyq9HUnIIbI
+ToDWz3A/2wZiwyDwqkc3UdYO2M1r0GJeKjFuDmJW7RPtCmv0O0lG52EgsV6RsawiofPBwmGC+Es
zRnBGR2ZSivc0kWfgC8OSgR58dAolANVhZ1pYUZsEh2PaNNRbgmYWbpjAx/iRh7tsx6sI3bTGzwV
QPphp/un8Bt6ylLZuUwx/Occ3u4YyKH1760/BYL8XLoPVulFBRjz79qxq6rTgKL3AURtMfJqr7mE
cAms9RHiebG9NwasNeYMej3K3npXFIgrb9Ri8nk5aJiYwPX4IpQCAfEfOou1BQwvbUnX2nCWG4v5
h5JbU3H0gOBJoGzDAeinSMSuQ+P+KtZZj3zm9PY6Y2apAwjQogqUkeqWOf9P+KMB5MXXvY1EijO5
qdweRua0EjvBSyXBy7YU4zpTReYyMnD6E2+CcscRW+aeNPvtpA/E41czhvIKm92ds1REHzhE2gmA
zoQgnnB45df1Ja+v+iolRR1dc6AGI/M7Gjj7spwJePIPX7+Xf3C3igUuabHwff7RULOm8z9B7P0c
+qBoJumUFQMw/uHJ7HnZI4dbcyM3kLLVy8Cd3UM+mmey6qL0Ph0vrY7/UTXT/HnVT+94qdNnynrf
XgI7STYCMszmiuop+aoeNZa3GEiAx4l4Lil4oB/+UVOFV8TTQlTtEvPobP2BOgZrzpip0F8d+zvO
LchmVVIG8YCPAO8JtM6ML0hPccfvzUTJNbCxwLVmjdfv2/ZgVG6JaW0H05ozLbvhj4TyqrnEufJ+
65i5r7Nnl8brY5btu1dgat9rWk5NuNLq7wJwId2Odv+5eQQ2+JhNnvj/QbfyvjvNd6BB4hGb/RVy
PWbBEkOONQ/+kOdKxUFq+1WctGJCBISMFTZ5cUid58IrbUI9tvWe8ftknoyJTqao8CSyXMBFFo4I
ec2X4hPZrstf15dZtTjdGP6xLlcaKgxcpTiharn40YD/edphjuG2BwSz6cgBgQWoPcFYeiRc2BVp
fOGpi8P7p0WVRweGdO8Vduww6die0TiU21u5JOvHgzDXFCHSpsJM6uT1PZpwWXQmcC6MA38v027T
KiWkxsIVisPh1jWi8oYh/hdxUgrnBLy068iHtxq/APCoWrborKNXlefCvOk+QdBXb6XSAUQPKoAr
9ID98Vqs6adVO1Q8vemptoTao0jk5eeAM47AHqimAB6E2s2aN5MncJiFt9w6jP5SSw+hxywJV5Fq
gQIWQSFcc/Bth2B5njQ5DfAoCKnXA19TtFcwf8isykPs4eJjpIOsdxdvg05UnGuL6TosgwEusVjW
yjrBMfQTwvfQDzIdhhNBeyl/+8tX9EwIuAnK1aL8EEiXx7bOuOEqATih9KdtYg+ABB+cb0I4WRyz
XjYkjJtA3Fpvb1juLuBiMqNTniZiWiyxxJSFVqfhHllSJUskVS5lGePpeL4avVY/0/kLEptrm60B
nQzZ+MN07gOiwBAnnspkKbmZj+uiJVgdV7Fjs3QlF9rvZXlPBsSgG2cTcilS2stOTmLPHeHY55hF
vKSg6wsJpChmllklRhLNRCTRBh39fcfL3B8Ey8ZnaeFIqS1by3Gwinjj/dBXHHTxoLo3mMTf2+hN
NbRazHgJs3EZHfxi4rBDjbHUTZJaknDn/trKniuV9Noq+q2klzktjiZtfHKOZC3FObZdH8iUbkwp
d82cXS/c6+P/9a2jMnTzNz7pzg91OCBelh1HP/5s0yWNnycbYK+udyy9kqZJEn+KfjVAKiFOPhSV
7i+8WrXTfCwhxcGiHxazsJt+OFnO5hF/6nAaS51IUPx8Vd9sOlFg7/P8B7aotuJMRY7ENsX8RyRa
8aCsw+iKqmMrbO9AaJl7gtZdXQR+m/9a9zoNWEpsLiSv4ZC8L+PFIevbZol7+gxJ1Dd+9arx494x
rPYYVy3z3Kq2G4lG55SW2/turQ7j1m8b78t3r+7ZzIGVK7mNNz3C7nntV7NtT7pIHorUKF3H/rQC
8KSVAJ3rKWVNI0BpKdpqPsleObN70rruXN++d/v1WVTg8wCf6EeE1KoM9Qk6GjGss3mUmsDWpO1J
6wyKmDMR6fAUIMb4d9vlLfiT0i7Qn/zRHpeYuMpdo8QobnBsAPJTK7cwlJHx27PCUJ1QJNHtQbvh
APzYnP6aQZbTsir5lIJXcWQN2Xub2eS3hLRkvqRsEhYgZ1wiHbxn1/g0kL9d2S5dZDwY3wnOGcOU
GuCa+18PXQGEwesW505RmlSKIGkgnMegXfCHBTGnm+54NseY5gInybWM53Z4wRPGvduL/rmcmbX9
lEZdd0+snp/B80yHs3/xsVbRU6i6BiYF358pcGEAlebHoltHX2XAbSbzqWaT1ev9KpL8UWscCjrb
kJTTVAyOjn504fU9xIMN81Z16ore4rWb0OAfTMiJq+9rWPsayT79woKCmHDfTlfs4GlVVKijplE3
kivpfZMNaCxcMmwHfMnfCDh0aMjgPNMH7+STFFlOVC/UuL30/0krdRF8b8ZhP7avfYBbhiWkvNEH
b5dLNzXu2ax5rhyrC5jPwaihHSE6t2X4Us6wIMthfBFI2cqnXXQ8jhIM240YaiGloeRQoCcxdMdk
Iia4vYoNbalyp98984V3hoHla+8lmpTtDQqQ4F2z4/GAvQ5BbiE0TJ7VUUBlO8t5PL1TMPs3XNam
joqAASyxuZZRbjmYDtTlPlhoosO46iglQsHrW7S3eW33pajl5RL21xka+/idPwqJrooaB4mYd0Ir
ydQ73t6kLY1lWoTazB03ScMpD4w1+S+tZh523BclVUicYzoBaDrpn6LEvyhLoiGnxCAXIbyjlzgt
Uvd4LDbz7VzoYazzqKgCMLWblQkxgqDGMgoMT94fQ6UQtV8H9dxiLxJgNbgSBk6GeWQekQarsYGM
7xOlGJGVLSyBlShvLVE1TcJJgZZzvt9lTiNAMKJAL75XL1iNdq3ls1nfZvmLx0JAGDT8KwWEU4nR
jpLNSJo/ClAxUzQlpAbef7LlW918lJ/RGrWB2hxuTUJGT9jCcOAxCNiO+JawZu0Ave6cZy+pWB/R
hHd97GQ3ldWpcb6i9pbhkhoqVhx/N2ZJ55wdNHVRs54Q+J2eAz2wUpiIuCHmBH7yeXFoQmwxmgu4
T6KzbivQWVUjc5N4+VYJENzEpCKQe3S0ebTO+o5AKBQw09PHU+dEO9QuSw/m1nUzYvtuhbdDtNux
gqSu/nqjv61FzHHlQLsTsFfAi+gZj6tQz2M+Kz4JPxNI+2DSyIDYDsB2m0M6F6Uenqk5AUABHN7B
89oSZEBSZSUTecQbTSPSfr4GRVFP5B/nEARVM5UxBVmE5O+N3iteOJWqy/TM7lrpXlvjH85wBFWZ
dtyYV9EDjKOl7eKWrTDzJJbOAmsNPG+3ES9X62NOYf0djLgQSP7+d7cBMzbFAweYjkxjfltEHMrb
pDgL9XfISpZLWCWDhb+BhYgAEOwD2D+6jrVfBWOy8DgmzG/klp3T6DzOJ00xLjpN+rwJ3w+yrizv
vIg6I+MwmykgwC03JDY9nKb0E0LO4Z9MpO1TauRv+E5XZM5Iou2mPF1inzfCDiNwcV5dC0NBKfsz
PgogiIxIbrG4f84hLiUbOGfEcxC55cmBshdl3f3fSH5uK+zySCjaAEVUMUzbDmSDn+5SKEUEZPwX
C7xOcFQlApbs4AD1gD9b2mtUh9vXnjLvy8ZUzjnJCmeZcjEKeeLRZUOaGytrVE3vSVYoNy/TskY4
EauPSq5n0Sz6FL5xKYyqJGcarGI+yq0fHzC1YU5GHpAVIrKXglqnndFlVCAAWEXdTnm6MBXfhT5H
QDvoIQtJB5AleNzExz9vumEIzvlaXnuCUDRqzV4PAc9m027CyM13e1htKfCtQrD7JQ/7+5fmuTTF
r/G3tYc3Is/MuUIxhB205a2c771Lf60MhmZzmpS6MvNfaqobmSvdV7yINySyXjY5xQGkQmVkiqBz
Avln/513jEnfTfMGksO4w8uGCV/u7OgWXuDQnURVpnDA/6FdGxjEYIRe5xRAYDqTkOR4bcod/DyG
je93/evadGt1VPHxWxgwJWgJP3F9HbH4W9xhhKGMkuFHXVMUiYrYmHS+xG1yugaL2IwxP6eLsYry
0Vg/xkYDgk7mKjjODJ9oQ7B+80XHpI9e+A5vbu7pD/4SzlQgeCb6kTeqUrrf9xAFJnq1wbfNqSEe
Q3juaHaRR3Vnm2He9jPIim7Af8OAjhFSQlJSW4mtxspBRObKUr12iT6OijlIweMw63ktdBBrs1rL
ltT4HuPtyiNDFqOBlx0xqT0mwFnh3xtPH8VS6a1k7xtwV0sTHesBcYFKGAIV3/cu8DA+WhoqvW+I
B8bh2p6wztDr3qeE+ckXqn8WTm6gpqhkFn9F6D/N+68PCUgaGP0+bwfr7RTbcRTGOkM8NliLP5z5
IR5OLISW1BQ0CXlDXLqHw2ffbBoW0GFfABv/jBmjDJx5UvBR6Xx+BBNPXFZncmBQrf6drBuJBJUj
4P0QFCIApN4XuCBI5H6sy5PWXObUTdB19Kx4i4vzfFnt6FlEn0OKAZdBWLRSvYHcrMRgXvIb4lp6
zl0BvCV4JV9PWEuhahFJmxo1XpAJTbSXH78TfKSw+r9oiBzjiD7iSHiLd4RpnLdsbFAknwS6t+8H
f8DMonBawd2JRju6IQEYzhjlfcb8OxBKR5JygcdSY4KkAS1ii9eeUp5moty+BJ5WBQmo3gSeQGI8
4XathYY4+XTcICQdxqdm2BT6c4T7HFV+JvuLnRFBEtyLP3k6MHpu4cHldFErQuokEQBFn53t1G8V
qkli32+JCi/2I4+mhDkbGD86Z/eR4yMAB0RB1MgUuvjnu+AKx2JdtyeZK/NFmycm/S0EK/sDpYuP
IWoiLd+DTwBjDUtw3GnwAbrvLez2gCJlFywqeO5Y73dNWQtBWcXZErkSp/RxgVfVyb40iwLj7Uc8
0/zoxtLmcynFNOscqPb+ETFryYharEz2r0FeC51s5mVh1kfrhv8zJmiDUezc+cwshqfZfkQFw78d
//ACpMlzbx+A+3hvSuuxPKFP1Lr/KQghWAUu9QERcC0fJxZBC4YdxAnH432vax8bqh6CElAv1vbW
r063WsEEFxgUKOMFuS8aGcrnBXtwtv4AhEaPj+93Og2CLv0hcL7VtYCFwZ0ujQqKhYecumdg92Az
BxZ9EmYv8XaisfbYBWX8Qz0tU+ovZ/X9GOu9IQ/mAFLJ1aoRaAlLhlYmtQYDYJCNTDcoEd+lRh+N
+r1xROJ2nkowzkSgyoD4/O2KrO4Bshf/rbo8nI8sNJvFYWqtzGkNsfX96by+Ab8NcBgxqFG6wsws
QxRFPY2ebzQnIKXKU5/5x53G2vXhoNFXzK8w9OB++tW4UDOwUQm3psOB91475VrHT6OBn1UogGAd
PShI/bRsNXB+pZ/LzlXMIgCEfffti4Q4bJiKoaWg3f1rPxM5TXuxnhSyI7D16964d53mcuw5BRef
2pvC291XyRZo5h+VfJqqG9WeV2XRWemEfFcVmwIU0cckuu6sP9V33ckB3oY5Yvve6Uu1HaI13yX6
LETNHQuYU36VpiaAvxYm0Hndw2Rn7qfwOZzOFfpPrOTIWZOyQAEIt5gLMDfojNneeWvAKWuXoi7v
KxQDak6Y2LRuCMx2V3ym5fHL74ZZgzIQuQzspOqGXiSYn+8s4aD1ib/PFUB26oJgQZI8HLrI0MCd
O9fGZ5zv4RbuSbr0qA==
`protect end_protected

